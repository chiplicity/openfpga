* NGSPICE file created from grid_io_left_left.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A Y VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_4 abstract view
.subckt sky130_fd_sc_hd__ebufn_4 A TE_B Z VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 D Q CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N X VGND VNB VPB VPWR
.ends

.subckt grid_io_left_left IO_ISOL_N ccff_head ccff_tail gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT prog_clk right_width_0_height_0__pin_0_
+ right_width_0_height_0__pin_1_lower right_width_0_height_0__pin_1_upper VPWR VGND
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
+ logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__inv_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN
+ logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y right_width_0_height_0__pin_1_lower
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__ebufn_4
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE right_width_0_height_0__pin_0_
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR gfpga_pad_EMBEDDED_IO_HD_SOC_OUT VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__ebufn_4
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0_ right_width_0_height_0__pin_1_lower right_width_0_height_0__pin_1_upper VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ ccff_head ccff_tail prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE ccff_tail
+ IO_ISOL_N gfpga_pad_EMBEDDED_IO_HD_SOC_DIR VGND VGND VPWR VPWR sky130_fd_sc_hd__or2b_4
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
.ends

