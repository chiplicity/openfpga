VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_1__0_
  CLASS BLOCK ;
  FOREIGN sb_1__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 120.000 BY 120.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 2.400 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 2.760 120.000 3.360 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 8.880 120.000 9.480 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 2.400 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 15.000 120.000 15.600 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 21.120 120.000 21.720 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 2.400 ;
    END
  END address[6]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.310 117.600 3.590 120.000 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 27.920 120.000 28.520 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 34.040 120.000 34.640 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.750 117.600 10.030 120.000 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 2.400 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 2.400 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 2.400 4.040 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 2.400 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 117.600 16.930 120.000 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 2.400 10.840 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 2.400 17.640 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 2.400 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 2.400 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 2.400 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 2.400 25.120 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 40.160 120.000 40.760 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 23.090 117.600 23.370 120.000 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 2.400 ;
    END
  END chanx_left_out[8]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.990 117.600 30.270 120.000 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 46.280 120.000 46.880 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.430 117.600 36.710 120.000 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 2.400 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 2.400 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 2.400 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 2.400 31.920 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 2.400 38.720 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.330 117.600 43.610 120.000 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 2.400 46.200 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 49.770 117.600 50.050 120.000 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 53.080 120.000 53.680 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 2.400 53.000 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 59.200 120.000 59.800 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 2.400 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 56.670 117.600 56.950 120.000 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 2.400 59.800 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 2.400 67.280 ;
    END
  END chanx_right_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.110 117.600 63.390 120.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 65.320 120.000 65.920 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 2.400 74.080 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.010 117.600 70.290 120.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 2.400 80.880 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 2.400 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 2.400 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 2.400 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 2.400 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 2.400 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 2.400 88.360 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 2.400 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 2.400 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 71.440 120.000 72.040 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 78.240 120.000 78.840 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 84.360 120.000 84.960 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.560 2.400 95.160 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 90.480 120.000 91.080 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 2.400 ;
    END
  END enable
  PIN left_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 83.350 117.600 83.630 120.000 ;
    END
  END left_bottom_grid_pin_11_
  PIN left_bottom_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 2.400 ;
    END
  END left_bottom_grid_pin_13_
  PIN left_bottom_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 109.520 120.000 110.120 ;
    END
  END left_bottom_grid_pin_15_
  PIN left_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 96.600 120.000 97.200 ;
    END
  END left_bottom_grid_pin_1_
  PIN left_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 103.400 120.000 104.000 ;
    END
  END left_bottom_grid_pin_3_
  PIN left_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.450 117.600 76.730 120.000 ;
    END
  END left_bottom_grid_pin_5_
  PIN left_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 2.400 ;
    END
  END left_bottom_grid_pin_7_
  PIN left_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 2.400 101.960 ;
    END
  END left_bottom_grid_pin_9_
  PIN left_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 2.400 ;
    END
  END left_top_grid_pin_10_
  PIN right_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.690 117.600 96.970 120.000 ;
    END
  END right_bottom_grid_pin_11_
  PIN right_bottom_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.130 117.600 103.410 120.000 ;
    END
  END right_bottom_grid_pin_13_
  PIN right_bottom_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.030 117.600 110.310 120.000 ;
    END
  END right_bottom_grid_pin_15_
  PIN right_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 2.400 109.440 ;
    END
  END right_bottom_grid_pin_1_
  PIN right_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 2.400 116.240 ;
    END
  END right_bottom_grid_pin_3_
  PIN right_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 2.400 ;
    END
  END right_bottom_grid_pin_5_
  PIN right_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 89.790 117.600 90.070 120.000 ;
    END
  END right_bottom_grid_pin_7_
  PIN right_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 115.640 120.000 116.240 ;
    END
  END right_bottom_grid_pin_9_
  PIN right_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 116.470 117.600 116.750 120.000 ;
    END
  END right_top_grid_pin_10_
  PIN top_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 2.400 ;
    END
  END top_left_grid_pin_13_
  PIN top_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 2.400 ;
    END
  END top_right_grid_pin_11_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 24.720 10.640 26.320 109.040 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 44.720 10.640 46.320 109.040 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 114.080 108.885 ;
      LAYER met1 ;
        RECT 0.530 0.380 118.150 117.940 ;
      LAYER met2 ;
        RECT 0.550 117.320 3.030 118.050 ;
        RECT 3.870 117.320 9.470 118.050 ;
        RECT 10.310 117.320 16.370 118.050 ;
        RECT 17.210 117.320 22.810 118.050 ;
        RECT 23.650 117.320 29.710 118.050 ;
        RECT 30.550 117.320 36.150 118.050 ;
        RECT 36.990 117.320 43.050 118.050 ;
        RECT 43.890 117.320 49.490 118.050 ;
        RECT 50.330 117.320 56.390 118.050 ;
        RECT 57.230 117.320 62.830 118.050 ;
        RECT 63.670 117.320 69.730 118.050 ;
        RECT 70.570 117.320 76.170 118.050 ;
        RECT 77.010 117.320 83.070 118.050 ;
        RECT 83.910 117.320 89.510 118.050 ;
        RECT 90.350 117.320 96.410 118.050 ;
        RECT 97.250 117.320 102.850 118.050 ;
        RECT 103.690 117.320 109.750 118.050 ;
        RECT 110.590 117.320 116.190 118.050 ;
        RECT 117.030 117.320 118.130 118.050 ;
        RECT 0.550 2.680 118.130 117.320 ;
        RECT 0.550 0.270 1.650 2.680 ;
        RECT 2.490 0.270 5.790 2.680 ;
        RECT 6.630 0.270 9.930 2.680 ;
        RECT 10.770 0.270 14.070 2.680 ;
        RECT 14.910 0.270 18.210 2.680 ;
        RECT 19.050 0.270 22.350 2.680 ;
        RECT 23.190 0.270 26.490 2.680 ;
        RECT 27.330 0.270 30.630 2.680 ;
        RECT 31.470 0.270 34.770 2.680 ;
        RECT 35.610 0.270 38.910 2.680 ;
        RECT 39.750 0.270 43.050 2.680 ;
        RECT 43.890 0.270 47.190 2.680 ;
        RECT 48.030 0.270 51.330 2.680 ;
        RECT 52.170 0.270 55.470 2.680 ;
        RECT 56.310 0.270 59.610 2.680 ;
        RECT 60.450 0.270 63.750 2.680 ;
        RECT 64.590 0.270 67.890 2.680 ;
        RECT 68.730 0.270 72.030 2.680 ;
        RECT 72.870 0.270 76.170 2.680 ;
        RECT 77.010 0.270 80.310 2.680 ;
        RECT 81.150 0.270 84.450 2.680 ;
        RECT 85.290 0.270 88.590 2.680 ;
        RECT 89.430 0.270 92.730 2.680 ;
        RECT 93.570 0.270 96.870 2.680 ;
        RECT 97.710 0.270 101.010 2.680 ;
        RECT 101.850 0.270 105.150 2.680 ;
        RECT 105.990 0.270 109.290 2.680 ;
        RECT 110.130 0.270 113.430 2.680 ;
        RECT 114.270 0.270 117.570 2.680 ;
      LAYER met3 ;
        RECT 2.800 115.240 117.200 115.640 ;
        RECT 0.270 110.520 118.370 115.240 ;
        RECT 0.270 109.840 117.200 110.520 ;
        RECT 2.800 109.120 117.200 109.840 ;
        RECT 2.800 108.440 118.370 109.120 ;
        RECT 0.270 104.400 118.370 108.440 ;
        RECT 0.270 103.000 117.200 104.400 ;
        RECT 0.270 102.360 118.370 103.000 ;
        RECT 2.800 100.960 118.370 102.360 ;
        RECT 0.270 97.600 118.370 100.960 ;
        RECT 0.270 96.200 117.200 97.600 ;
        RECT 0.270 95.560 118.370 96.200 ;
        RECT 2.800 94.160 118.370 95.560 ;
        RECT 0.270 91.480 118.370 94.160 ;
        RECT 0.270 90.080 117.200 91.480 ;
        RECT 0.270 88.760 118.370 90.080 ;
        RECT 2.800 87.360 118.370 88.760 ;
        RECT 0.270 85.360 118.370 87.360 ;
        RECT 0.270 83.960 117.200 85.360 ;
        RECT 0.270 81.280 118.370 83.960 ;
        RECT 2.800 79.880 118.370 81.280 ;
        RECT 0.270 79.240 118.370 79.880 ;
        RECT 0.270 77.840 117.200 79.240 ;
        RECT 0.270 74.480 118.370 77.840 ;
        RECT 2.800 73.080 118.370 74.480 ;
        RECT 0.270 72.440 118.370 73.080 ;
        RECT 0.270 71.040 117.200 72.440 ;
        RECT 0.270 67.680 118.370 71.040 ;
        RECT 2.800 66.320 118.370 67.680 ;
        RECT 2.800 66.280 117.200 66.320 ;
        RECT 0.270 64.920 117.200 66.280 ;
        RECT 0.270 60.200 118.370 64.920 ;
        RECT 2.800 58.800 117.200 60.200 ;
        RECT 0.270 54.080 118.370 58.800 ;
        RECT 0.270 53.400 117.200 54.080 ;
        RECT 2.800 52.680 117.200 53.400 ;
        RECT 2.800 52.000 118.370 52.680 ;
        RECT 0.270 47.280 118.370 52.000 ;
        RECT 0.270 46.600 117.200 47.280 ;
        RECT 2.800 45.880 117.200 46.600 ;
        RECT 2.800 45.200 118.370 45.880 ;
        RECT 0.270 41.160 118.370 45.200 ;
        RECT 0.270 39.760 117.200 41.160 ;
        RECT 0.270 39.120 118.370 39.760 ;
        RECT 2.800 37.720 118.370 39.120 ;
        RECT 0.270 35.040 118.370 37.720 ;
        RECT 0.270 33.640 117.200 35.040 ;
        RECT 0.270 32.320 118.370 33.640 ;
        RECT 2.800 30.920 118.370 32.320 ;
        RECT 0.270 28.920 118.370 30.920 ;
        RECT 0.270 27.520 117.200 28.920 ;
        RECT 0.270 25.520 118.370 27.520 ;
        RECT 2.800 24.120 118.370 25.520 ;
        RECT 0.270 22.120 118.370 24.120 ;
        RECT 0.270 20.720 117.200 22.120 ;
        RECT 0.270 18.040 118.370 20.720 ;
        RECT 2.800 16.640 118.370 18.040 ;
        RECT 0.270 16.000 118.370 16.640 ;
        RECT 0.270 14.600 117.200 16.000 ;
        RECT 0.270 11.240 118.370 14.600 ;
        RECT 2.800 9.880 118.370 11.240 ;
        RECT 2.800 9.840 117.200 9.880 ;
        RECT 0.270 8.480 117.200 9.840 ;
        RECT 0.270 4.440 118.370 8.480 ;
        RECT 2.800 3.760 118.370 4.440 ;
        RECT 2.800 3.040 117.200 3.760 ;
        RECT 0.270 2.895 117.200 3.040 ;
      LAYER met4 ;
        RECT 0.295 10.640 24.320 109.040 ;
        RECT 26.720 10.640 44.320 109.040 ;
        RECT 46.720 10.640 106.320 109.040 ;
  END
END sb_1__0_
END LIBRARY

