magic
tech EFS8A
magscale 1 2
timestamp 1602095374
<< locali >>
rect 15887 19873 16014 19907
rect 13783 19465 13921 19499
rect 13093 18207 13127 18309
rect 14013 18071 14047 18241
rect 6503 17697 6630 17731
rect 10327 16745 10333 16779
rect 17319 16745 17325 16779
rect 10327 16677 10361 16745
rect 17319 16677 17353 16745
rect 15703 15521 15830 15555
rect 18371 15521 18406 15555
rect 10327 14807 10361 14875
rect 10327 14773 10333 14807
rect 15663 14569 15669 14603
rect 15663 14501 15697 14569
rect 2179 13753 2224 13787
rect 8395 13719 8429 13787
rect 8395 13685 8401 13719
rect 9972 13413 10044 13447
rect 7757 11543 7791 11713
rect 6647 11305 6653 11339
rect 16031 11305 16037 11339
rect 6647 11237 6681 11305
rect 16031 11237 16065 11305
rect 18423 10455 18457 10523
rect 18423 10421 18429 10455
rect 3927 10081 4146 10115
rect 16899 10081 16934 10115
rect 6101 9367 6135 9605
rect 10051 9129 10057 9163
rect 10051 9061 10085 9129
rect 21223 8381 21350 8415
rect 2139 8041 2145 8075
rect 2139 7973 2173 8041
rect 19751 6817 19878 6851
rect 17727 5797 17772 5831
rect 16439 5729 16474 5763
rect 6377 5015 6411 5321
rect 7665 5151 7699 5321
rect 7757 5083 7791 5321
rect 7573 5049 7791 5083
rect 8159 4641 8286 4675
rect 3617 3995 3651 4165
rect 9999 3621 10044 3655
rect 5767 3553 5802 3587
rect 19211 3145 19349 3179
rect 14467 2839 14501 2907
rect 14467 2805 14473 2839
rect 14139 2465 14219 2499
<< viali >>
rect 20085 21641 20119 21675
rect 8560 21437 8594 21471
rect 19600 21437 19634 21471
rect 8631 21301 8665 21335
rect 9045 21301 9079 21335
rect 19671 21301 19705 21335
rect 8585 21097 8619 21131
rect 12541 21097 12575 21131
rect 18245 21097 18279 21131
rect 12357 20961 12391 20995
rect 18061 20961 18095 20995
rect 19876 20961 19910 20995
rect 19947 20757 19981 20791
rect 2697 20553 2731 20587
rect 4537 20553 4571 20587
rect 7941 20553 7975 20587
rect 8401 20553 8435 20587
rect 14197 20553 14231 20587
rect 17233 20553 17267 20587
rect 19165 20553 19199 20587
rect 21097 20553 21131 20587
rect 19993 20485 20027 20519
rect 12817 20417 12851 20451
rect 2212 20349 2246 20383
rect 4144 20349 4178 20383
rect 7757 20349 7791 20383
rect 14013 20349 14047 20383
rect 14565 20349 14599 20383
rect 16748 20349 16782 20383
rect 18981 20349 19015 20383
rect 19533 20349 19567 20383
rect 20913 20349 20947 20383
rect 21465 20349 21499 20383
rect 9413 20281 9447 20315
rect 9505 20281 9539 20315
rect 10057 20281 10091 20315
rect 11897 20281 11931 20315
rect 12541 20281 12575 20315
rect 12633 20281 12667 20315
rect 18245 20281 18279 20315
rect 2283 20213 2317 20247
rect 4215 20213 4249 20247
rect 9229 20213 9263 20247
rect 11345 20213 11379 20247
rect 12265 20213 12299 20247
rect 16819 20213 16853 20247
rect 8769 19941 8803 19975
rect 9873 19941 9907 19975
rect 11713 19941 11747 19975
rect 12541 19941 12575 19975
rect 13277 19941 13311 19975
rect 17325 19941 17359 19975
rect 19349 19941 19383 19975
rect 19441 19941 19475 19975
rect 1476 19873 1510 19907
rect 8125 19873 8159 19907
rect 15853 19873 15887 19907
rect 20980 19873 21014 19907
rect 9781 19805 9815 19839
rect 10057 19805 10091 19839
rect 11621 19805 11655 19839
rect 13185 19805 13219 19839
rect 17233 19805 17267 19839
rect 17877 19805 17911 19839
rect 19993 19805 20027 19839
rect 12173 19737 12207 19771
rect 13737 19737 13771 19771
rect 1547 19669 1581 19703
rect 9413 19669 9447 19703
rect 16083 19669 16117 19703
rect 16497 19669 16531 19703
rect 21051 19669 21085 19703
rect 1593 19465 1627 19499
rect 8033 19465 8067 19499
rect 9413 19465 9447 19499
rect 9781 19465 9815 19499
rect 10149 19465 10183 19499
rect 12173 19465 12207 19499
rect 13369 19465 13403 19499
rect 13921 19465 13955 19499
rect 18429 19465 18463 19499
rect 20913 19465 20947 19499
rect 21649 19465 21683 19499
rect 20177 19397 20211 19431
rect 11529 19329 11563 19363
rect 11805 19329 11839 19363
rect 17785 19329 17819 19363
rect 19625 19329 19659 19363
rect 8493 19261 8527 19295
rect 10701 19261 10735 19295
rect 11437 19261 11471 19295
rect 12500 19261 12534 19295
rect 13712 19261 13746 19295
rect 14105 19261 14139 19295
rect 15301 19261 15335 19295
rect 15428 19261 15462 19295
rect 17141 19261 17175 19295
rect 21148 19261 21182 19295
rect 8401 19193 8435 19227
rect 8855 19193 8889 19227
rect 12587 19193 12621 19227
rect 15531 19193 15565 19227
rect 16497 19193 16531 19227
rect 16589 19193 16623 19227
rect 17509 19193 17543 19227
rect 19441 19193 19475 19227
rect 19717 19193 19751 19227
rect 20637 19193 20671 19227
rect 21235 19193 21269 19227
rect 12909 19125 12943 19159
rect 16037 19125 16071 19159
rect 18521 19125 18555 19159
rect 18981 19125 19015 19159
rect 10701 18921 10735 18955
rect 13553 18921 13587 18955
rect 14335 18921 14369 18955
rect 16497 18921 16531 18955
rect 10102 18853 10136 18887
rect 11713 18853 11747 18887
rect 12265 18853 12299 18887
rect 15622 18853 15656 18887
rect 17141 18853 17175 18887
rect 17233 18853 17267 18887
rect 18889 18853 18923 18887
rect 1444 18785 1478 18819
rect 13128 18785 13162 18819
rect 14232 18785 14266 18819
rect 9781 18717 9815 18751
rect 11621 18717 11655 18751
rect 13231 18717 13265 18751
rect 15301 18717 15335 18751
rect 18797 18717 18831 18751
rect 19073 18717 19107 18751
rect 16221 18649 16255 18683
rect 17693 18649 17727 18683
rect 1547 18581 1581 18615
rect 8585 18581 8619 18615
rect 19717 18581 19751 18615
rect 1869 18377 1903 18411
rect 7665 18377 7699 18411
rect 9321 18377 9355 18411
rect 11253 18377 11287 18411
rect 12173 18377 12207 18411
rect 15209 18377 15243 18411
rect 17693 18377 17727 18411
rect 19257 18377 19291 18411
rect 21189 18377 21223 18411
rect 8125 18309 8159 18343
rect 13093 18309 13127 18343
rect 17417 18309 17451 18343
rect 8309 18241 8343 18275
rect 8953 18241 8987 18275
rect 10149 18241 10183 18275
rect 1476 18173 1510 18207
rect 2237 18173 2271 18207
rect 11412 18173 11446 18207
rect 12516 18173 12550 18207
rect 13093 18173 13127 18207
rect 14013 18241 14047 18275
rect 18245 18241 18279 18275
rect 19533 18241 19567 18275
rect 19993 18241 20027 18275
rect 8401 18105 8435 18139
rect 9873 18105 9907 18139
rect 9965 18105 9999 18139
rect 13001 18105 13035 18139
rect 14289 18173 14323 18207
rect 16532 18173 16566 18207
rect 16957 18173 16991 18207
rect 18496 18173 18530 18207
rect 21005 18173 21039 18207
rect 14610 18105 14644 18139
rect 15485 18105 15519 18139
rect 19625 18105 19659 18139
rect 1547 18037 1581 18071
rect 9689 18037 9723 18071
rect 10793 18037 10827 18071
rect 11483 18037 11517 18071
rect 11897 18037 11931 18071
rect 12587 18037 12621 18071
rect 13277 18037 13311 18071
rect 13737 18037 13771 18071
rect 14013 18037 14047 18071
rect 14197 18037 14231 18071
rect 15853 18037 15887 18071
rect 16635 18037 16669 18071
rect 18567 18037 18601 18071
rect 18981 18037 19015 18071
rect 21557 18037 21591 18071
rect 2237 17833 2271 17867
rect 19901 17833 19935 17867
rect 21097 17833 21131 17867
rect 9965 17765 9999 17799
rect 11713 17765 11747 17799
rect 14381 17765 14415 17799
rect 16865 17765 16899 17799
rect 16957 17765 16991 17799
rect 18981 17765 19015 17799
rect 19073 17765 19107 17799
rect 4905 17697 4939 17731
rect 5365 17697 5399 17731
rect 6469 17697 6503 17731
rect 10333 17697 10367 17731
rect 13645 17697 13679 17731
rect 14105 17697 14139 17731
rect 15336 17697 15370 17731
rect 20913 17697 20947 17731
rect 5457 17629 5491 17663
rect 8585 17629 8619 17663
rect 10885 17629 10919 17663
rect 11621 17629 11655 17663
rect 11897 17629 11931 17663
rect 18337 17629 18371 17663
rect 19257 17629 19291 17663
rect 10517 17561 10551 17595
rect 17417 17561 17451 17595
rect 6699 17493 6733 17527
rect 8493 17493 8527 17527
rect 12541 17493 12575 17527
rect 13553 17493 13587 17527
rect 14657 17493 14691 17527
rect 15439 17493 15473 17527
rect 15761 17493 15795 17527
rect 5089 17289 5123 17323
rect 10333 17289 10367 17323
rect 12173 17289 12207 17323
rect 14841 17289 14875 17323
rect 15209 17289 15243 17323
rect 17141 17289 17175 17323
rect 19625 17289 19659 17323
rect 21465 17289 21499 17323
rect 21741 17289 21775 17323
rect 8217 17221 8251 17255
rect 13277 17221 13311 17255
rect 16221 17221 16255 17255
rect 19257 17221 19291 17255
rect 2329 17153 2363 17187
rect 2605 17153 2639 17187
rect 4629 17153 4663 17187
rect 6285 17153 6319 17187
rect 6929 17153 6963 17187
rect 10793 17153 10827 17187
rect 11437 17153 11471 17187
rect 14197 17153 14231 17187
rect 15301 17153 15335 17187
rect 16865 17153 16899 17187
rect 18337 17153 18371 17187
rect 8401 17085 8435 17119
rect 8861 17085 8895 17119
rect 12484 17085 12518 17119
rect 13461 17085 13495 17119
rect 13921 17085 13955 17119
rect 20980 17085 21014 17119
rect 2421 17017 2455 17051
rect 3617 17017 3651 17051
rect 4169 17017 4203 17051
rect 4261 17017 4295 17051
rect 7021 17017 7055 17051
rect 7573 17017 7607 17051
rect 10885 17017 10919 17051
rect 13001 17017 13035 17051
rect 15622 17017 15656 17051
rect 18429 17017 18463 17051
rect 18981 17017 19015 17051
rect 2145 16949 2179 16983
rect 3893 16949 3927 16983
rect 5549 16949 5583 16983
rect 6653 16949 6687 16983
rect 8493 16949 8527 16983
rect 9965 16949 9999 16983
rect 11713 16949 11747 16983
rect 12587 16949 12621 16983
rect 17877 16949 17911 16983
rect 21051 16949 21085 16983
rect 8769 16745 8803 16779
rect 10333 16745 10367 16779
rect 10885 16745 10919 16779
rect 15577 16745 15611 16779
rect 17325 16745 17359 16779
rect 17877 16745 17911 16779
rect 21097 16745 21131 16779
rect 4215 16677 4249 16711
rect 5819 16677 5853 16711
rect 8211 16677 8245 16711
rect 11897 16677 11931 16711
rect 18337 16677 18371 16711
rect 18889 16677 18923 16711
rect 4123 16609 4157 16643
rect 5457 16609 5491 16643
rect 13645 16609 13679 16643
rect 14105 16609 14139 16643
rect 15301 16609 15335 16643
rect 15761 16609 15795 16643
rect 20913 16609 20947 16643
rect 7849 16541 7883 16575
rect 9965 16541 9999 16575
rect 11805 16541 11839 16575
rect 12173 16541 12207 16575
rect 14381 16541 14415 16575
rect 16957 16541 16991 16575
rect 18797 16541 18831 16575
rect 19073 16541 19107 16575
rect 2605 16405 2639 16439
rect 6377 16405 6411 16439
rect 6837 16405 6871 16439
rect 13461 16405 13495 16439
rect 5825 16201 5859 16235
rect 7941 16201 7975 16235
rect 8309 16201 8343 16235
rect 10149 16201 10183 16235
rect 11897 16201 11931 16235
rect 13369 16201 13403 16235
rect 15301 16201 15335 16235
rect 16037 16201 16071 16235
rect 17141 16201 17175 16235
rect 19533 16201 19567 16235
rect 21189 16201 21223 16235
rect 1593 16133 1627 16167
rect 11437 16133 11471 16167
rect 12173 16133 12207 16167
rect 17785 16133 17819 16167
rect 3985 16065 4019 16099
rect 5549 16065 5583 16099
rect 6285 16065 6319 16099
rect 6929 16065 6963 16099
rect 7205 16065 7239 16099
rect 10885 16065 10919 16099
rect 14933 16065 14967 16099
rect 18337 16065 18371 16099
rect 20177 16065 20211 16099
rect 20453 16065 20487 16099
rect 1409 15997 1443 16031
rect 1961 15997 1995 16031
rect 2421 15997 2455 16031
rect 2789 15997 2823 16031
rect 3065 15997 3099 16031
rect 3249 15997 3283 16031
rect 4077 15997 4111 16031
rect 8953 15997 8987 16031
rect 9321 15997 9355 16031
rect 9505 15997 9539 16031
rect 14197 15997 14231 16031
rect 14657 15997 14691 16031
rect 15669 15997 15703 16031
rect 16221 15997 16255 16031
rect 19257 15997 19291 16031
rect 19901 15997 19935 16031
rect 3617 15929 3651 15963
rect 4439 15929 4473 15963
rect 7021 15929 7055 15963
rect 9781 15929 9815 15963
rect 10701 15929 10735 15963
rect 10977 15929 11011 15963
rect 16542 15929 16576 15963
rect 17417 15929 17451 15963
rect 18658 15929 18692 15963
rect 20269 15929 20303 15963
rect 4997 15861 5031 15895
rect 6561 15861 6595 15895
rect 13645 15861 13679 15895
rect 14013 15861 14047 15895
rect 4261 15657 4295 15691
rect 8401 15657 8435 15691
rect 9045 15657 9079 15691
rect 10701 15657 10735 15691
rect 11161 15657 11195 15691
rect 16589 15657 16623 15691
rect 17785 15657 17819 15691
rect 18797 15657 18831 15691
rect 20085 15657 20119 15691
rect 2605 15589 2639 15623
rect 4721 15589 4755 15623
rect 6561 15589 6595 15623
rect 11621 15589 11655 15623
rect 14381 15589 14415 15623
rect 16221 15589 16255 15623
rect 16957 15589 16991 15623
rect 1476 15521 1510 15555
rect 9689 15521 9723 15555
rect 10149 15521 10183 15555
rect 13645 15521 13679 15555
rect 14197 15521 14231 15555
rect 14657 15521 14691 15555
rect 15669 15521 15703 15555
rect 18337 15521 18371 15555
rect 19384 15521 19418 15555
rect 2513 15453 2547 15487
rect 4629 15453 4663 15487
rect 4905 15453 4939 15487
rect 6469 15453 6503 15487
rect 7941 15453 7975 15487
rect 10425 15453 10459 15487
rect 11529 15453 11563 15487
rect 12173 15453 12207 15487
rect 16854 15453 16888 15487
rect 17325 15453 17359 15487
rect 2329 15385 2363 15419
rect 3065 15385 3099 15419
rect 7021 15385 7055 15419
rect 1547 15317 1581 15351
rect 1869 15317 1903 15351
rect 12541 15317 12575 15351
rect 15899 15317 15933 15351
rect 18475 15317 18509 15351
rect 19487 15317 19521 15351
rect 2697 15113 2731 15147
rect 2973 15113 3007 15147
rect 4077 15113 4111 15147
rect 6469 15113 6503 15147
rect 9873 15113 9907 15147
rect 10885 15113 10919 15147
rect 11529 15113 11563 15147
rect 11805 15113 11839 15147
rect 15025 15113 15059 15147
rect 15761 15113 15795 15147
rect 18337 15113 18371 15147
rect 19533 15113 19567 15147
rect 21465 15113 21499 15147
rect 3341 15045 3375 15079
rect 7481 15045 7515 15079
rect 1777 14977 1811 15011
rect 4629 14977 4663 15011
rect 4905 14977 4939 15011
rect 6929 14977 6963 15011
rect 7849 14977 7883 15011
rect 12817 14977 12851 15011
rect 16681 14977 16715 15011
rect 8401 14909 8435 14943
rect 8861 14909 8895 14943
rect 9137 14909 9171 14943
rect 9965 14909 9999 14943
rect 14289 14909 14323 14943
rect 14473 14909 14507 14943
rect 20980 14909 21014 14943
rect 1685 14841 1719 14875
rect 2098 14841 2132 14875
rect 4721 14841 4755 14875
rect 6101 14841 6135 14875
rect 7021 14841 7055 14875
rect 8217 14841 8251 14875
rect 12541 14841 12575 14875
rect 12633 14841 12667 14875
rect 14749 14841 14783 14875
rect 16405 14841 16439 14875
rect 16497 14841 16531 14875
rect 4445 14773 4479 14807
rect 5641 14773 5675 14807
rect 9413 14773 9447 14807
rect 10333 14773 10367 14807
rect 12173 14773 12207 14807
rect 13645 14773 13679 14807
rect 16221 14773 16255 14807
rect 17325 14773 17359 14807
rect 19073 14773 19107 14807
rect 21051 14773 21085 14807
rect 1961 14569 1995 14603
rect 4997 14569 5031 14603
rect 8033 14569 8067 14603
rect 9873 14569 9907 14603
rect 10241 14569 10275 14603
rect 11437 14569 11471 14603
rect 14381 14569 14415 14603
rect 15669 14569 15703 14603
rect 16221 14569 16255 14603
rect 16865 14569 16899 14603
rect 4398 14501 4432 14535
rect 5273 14501 5307 14535
rect 6285 14501 6319 14535
rect 10838 14501 10872 14535
rect 17233 14501 17267 14535
rect 19257 14501 19291 14535
rect 19349 14501 19383 14535
rect 1961 14433 1995 14467
rect 2237 14433 2271 14467
rect 8033 14433 8067 14467
rect 8309 14433 8343 14467
rect 10517 14433 10551 14467
rect 13369 14433 13403 14467
rect 13921 14433 13955 14467
rect 15301 14433 15335 14467
rect 4077 14365 4111 14399
rect 6193 14365 6227 14399
rect 6837 14365 6871 14399
rect 14105 14365 14139 14399
rect 17141 14365 17175 14399
rect 17785 14365 17819 14399
rect 19533 14365 19567 14399
rect 2697 14229 2731 14263
rect 3893 14229 3927 14263
rect 5917 14229 5951 14263
rect 7113 14229 7147 14263
rect 12541 14229 12575 14263
rect 14749 14229 14783 14263
rect 1777 14025 1811 14059
rect 3801 14025 3835 14059
rect 5365 14025 5399 14059
rect 6377 14025 6411 14059
rect 10241 14025 10275 14059
rect 12173 14025 12207 14059
rect 15669 14025 15703 14059
rect 16221 14025 16255 14059
rect 17417 14025 17451 14059
rect 17785 14025 17819 14059
rect 19165 14025 19199 14059
rect 5687 13957 5721 13991
rect 8953 13957 8987 13991
rect 9873 13957 9907 13991
rect 11069 13957 11103 13991
rect 13461 13957 13495 13991
rect 15025 13957 15059 13991
rect 1869 13889 1903 13923
rect 4066 13889 4100 13923
rect 4721 13889 4755 13923
rect 8033 13889 8067 13923
rect 9229 13889 9263 13923
rect 10517 13889 10551 13923
rect 11437 13889 11471 13923
rect 12817 13889 12851 13923
rect 14105 13889 14139 13923
rect 17141 13889 17175 13923
rect 2789 13821 2823 13855
rect 5600 13821 5634 13855
rect 6888 13821 6922 13855
rect 7297 13821 7331 13855
rect 18372 13821 18406 13855
rect 18475 13821 18509 13855
rect 20980 13821 21014 13855
rect 2145 13753 2179 13787
rect 4169 13753 4203 13787
rect 4997 13753 5031 13787
rect 10609 13753 10643 13787
rect 12541 13753 12575 13787
rect 12633 13753 12667 13787
rect 14013 13753 14047 13787
rect 14467 13753 14501 13787
rect 16497 13753 16531 13787
rect 16589 13753 16623 13787
rect 18889 13753 18923 13787
rect 19441 13753 19475 13787
rect 19533 13753 19567 13787
rect 20085 13753 20119 13787
rect 21465 13753 21499 13787
rect 3157 13685 3191 13719
rect 3525 13685 3559 13719
rect 6009 13685 6043 13719
rect 6975 13685 7009 13719
rect 7941 13685 7975 13719
rect 8401 13685 8435 13719
rect 15301 13685 15335 13719
rect 20361 13685 20395 13719
rect 21051 13685 21085 13719
rect 4169 13481 4203 13515
rect 6837 13481 6871 13515
rect 7113 13481 7147 13515
rect 7849 13481 7883 13515
rect 10609 13481 10643 13515
rect 10885 13481 10919 13515
rect 14105 13481 14139 13515
rect 18061 13481 18095 13515
rect 19625 13481 19659 13515
rect 2237 13413 2271 13447
rect 6279 13413 6313 13447
rect 9938 13413 9972 13447
rect 11713 13413 11747 13447
rect 12265 13413 12299 13447
rect 16865 13413 16899 13447
rect 18705 13413 18739 13447
rect 19257 13413 19291 13447
rect 21097 13413 21131 13447
rect 21649 13413 21683 13447
rect 1777 13345 1811 13379
rect 2053 13345 2087 13379
rect 4169 13345 4203 13379
rect 4629 13345 4663 13379
rect 8620 13345 8654 13379
rect 8723 13345 8757 13379
rect 15704 13345 15738 13379
rect 5917 13277 5951 13311
rect 9689 13277 9723 13311
rect 11621 13277 11655 13311
rect 16773 13277 16807 13311
rect 17417 13277 17451 13311
rect 18613 13277 18647 13311
rect 21005 13277 21039 13311
rect 2881 13209 2915 13243
rect 15807 13209 15841 13243
rect 2513 13141 2547 13175
rect 3801 13141 3835 13175
rect 5733 13141 5767 13175
rect 8217 13141 8251 13175
rect 9137 13141 9171 13175
rect 13461 13141 13495 13175
rect 13829 13141 13863 13175
rect 16497 13141 16531 13175
rect 19993 13141 20027 13175
rect 3157 12937 3191 12971
rect 5779 12937 5813 12971
rect 8217 12937 8251 12971
rect 8585 12937 8619 12971
rect 10609 12937 10643 12971
rect 12173 12937 12207 12971
rect 12587 12937 12621 12971
rect 13461 12937 13495 12971
rect 16773 12937 16807 12971
rect 17417 12937 17451 12971
rect 19533 12937 19567 12971
rect 20913 12937 20947 12971
rect 22109 12937 22143 12971
rect 1777 12869 1811 12903
rect 6561 12869 6595 12903
rect 7481 12869 7515 12903
rect 11805 12869 11839 12903
rect 16037 12869 16071 12903
rect 17785 12869 17819 12903
rect 20269 12869 20303 12903
rect 21373 12869 21407 12903
rect 4537 12801 4571 12835
rect 6929 12801 6963 12835
rect 7849 12801 7883 12835
rect 9597 12801 9631 12835
rect 10241 12801 10275 12835
rect 11529 12801 11563 12835
rect 18153 12801 18187 12835
rect 18429 12801 18463 12835
rect 19717 12801 19751 12835
rect 1685 12733 1719 12767
rect 1961 12733 1995 12767
rect 3801 12733 3835 12767
rect 3893 12733 3927 12767
rect 4077 12733 4111 12767
rect 5708 12733 5742 12767
rect 8861 12733 8895 12767
rect 9413 12733 9447 12767
rect 12516 12733 12550 12767
rect 13001 12733 13035 12767
rect 13553 12733 13587 12767
rect 14105 12733 14139 12767
rect 14289 12733 14323 12767
rect 14657 12733 14691 12767
rect 15117 12733 15151 12767
rect 16932 12733 16966 12767
rect 19165 12733 19199 12767
rect 21189 12733 21223 12767
rect 21741 12733 21775 12767
rect 2421 12665 2455 12699
rect 7021 12665 7055 12699
rect 10885 12665 10919 12699
rect 10977 12665 11011 12699
rect 15025 12665 15059 12699
rect 15479 12665 15513 12699
rect 18245 12665 18279 12699
rect 19809 12665 19843 12699
rect 2697 12597 2731 12631
rect 3709 12597 3743 12631
rect 4905 12597 4939 12631
rect 5273 12597 5307 12631
rect 6101 12597 6135 12631
rect 9965 12597 9999 12631
rect 16313 12597 16347 12631
rect 17003 12597 17037 12631
rect 3801 12393 3835 12427
rect 5733 12393 5767 12427
rect 8125 12393 8159 12427
rect 10287 12393 10321 12427
rect 10885 12393 10919 12427
rect 16313 12393 16347 12427
rect 17049 12393 17083 12427
rect 18797 12393 18831 12427
rect 20361 12393 20395 12427
rect 2881 12325 2915 12359
rect 15755 12325 15789 12359
rect 17963 12325 17997 12359
rect 21005 12325 21039 12359
rect 21097 12325 21131 12359
rect 1777 12257 1811 12291
rect 1869 12257 1903 12291
rect 2053 12257 2087 12291
rect 2513 12257 2547 12291
rect 4169 12257 4203 12291
rect 5917 12257 5951 12291
rect 6193 12257 6227 12291
rect 6929 12257 6963 12291
rect 7665 12257 7699 12291
rect 7941 12257 7975 12291
rect 10216 12257 10250 12291
rect 11897 12257 11931 12291
rect 12081 12257 12115 12291
rect 13645 12257 13679 12291
rect 14197 12257 14231 12291
rect 18521 12257 18555 12291
rect 19717 12257 19751 12291
rect 1685 12189 1719 12223
rect 4813 12189 4847 12223
rect 12173 12189 12207 12223
rect 12725 12189 12759 12223
rect 14381 12189 14415 12223
rect 15393 12189 15427 12223
rect 17601 12189 17635 12223
rect 21649 12189 21683 12223
rect 7757 12121 7791 12155
rect 8769 12121 8803 12155
rect 19901 12121 19935 12155
rect 7205 12053 7239 12087
rect 9137 12053 9171 12087
rect 13001 12053 13035 12087
rect 16589 12053 16623 12087
rect 3065 11849 3099 11883
rect 3709 11849 3743 11883
rect 4905 11849 4939 11883
rect 5733 11849 5767 11883
rect 12173 11849 12207 11883
rect 13645 11849 13679 11883
rect 15761 11849 15795 11883
rect 19717 11849 19751 11883
rect 21373 11849 21407 11883
rect 3433 11781 3467 11815
rect 3985 11781 4019 11815
rect 6929 11781 6963 11815
rect 11253 11781 11287 11815
rect 15485 11781 15519 11815
rect 18245 11781 18279 11815
rect 21097 11781 21131 11815
rect 2697 11713 2731 11747
rect 7757 11713 7791 11747
rect 8585 11713 8619 11747
rect 11483 11713 11517 11747
rect 12541 11713 12575 11747
rect 12817 11713 12851 11747
rect 14749 11713 14783 11747
rect 17141 11713 17175 11747
rect 2237 11645 2271 11679
rect 3893 11645 3927 11679
rect 4169 11645 4203 11679
rect 6561 11645 6595 11679
rect 6837 11645 6871 11679
rect 7113 11645 7147 11679
rect 7573 11645 7607 11679
rect 2329 11577 2363 11611
rect 6101 11577 6135 11611
rect 8769 11645 8803 11679
rect 9229 11645 9263 11679
rect 9597 11645 9631 11679
rect 9965 11645 9999 11679
rect 11396 11645 11430 11679
rect 14013 11645 14047 11679
rect 14473 11645 14507 11679
rect 21592 11645 21626 11679
rect 22017 11645 22051 11679
rect 12633 11577 12667 11611
rect 16497 11577 16531 11611
rect 16589 11577 16623 11611
rect 20085 11577 20119 11611
rect 20177 11577 20211 11611
rect 20729 11577 20763 11611
rect 4353 11509 4387 11543
rect 7757 11509 7791 11543
rect 7941 11509 7975 11543
rect 8217 11509 8251 11543
rect 9045 11509 9079 11543
rect 10609 11509 10643 11543
rect 11897 11509 11931 11543
rect 16313 11509 16347 11543
rect 17693 11509 17727 11543
rect 18981 11509 19015 11543
rect 21695 11509 21729 11543
rect 1777 11305 1811 11339
rect 2881 11305 2915 11339
rect 6653 11305 6687 11339
rect 9137 11305 9171 11339
rect 11345 11305 11379 11339
rect 14013 11305 14047 11339
rect 16037 11305 16071 11339
rect 16589 11305 16623 11339
rect 8769 11237 8803 11271
rect 10787 11237 10821 11271
rect 12494 11237 12528 11271
rect 20361 11237 20395 11271
rect 21097 11237 21131 11271
rect 21649 11237 21683 11271
rect 1777 11169 1811 11203
rect 2053 11169 2087 11203
rect 4721 11169 4755 11203
rect 5181 11169 5215 11203
rect 8033 11169 8067 11203
rect 8309 11169 8343 11203
rect 12173 11169 12207 11203
rect 18280 11169 18314 11203
rect 19901 11169 19935 11203
rect 19993 11169 20027 11203
rect 2513 11101 2547 11135
rect 5457 11101 5491 11135
rect 6285 11101 6319 11135
rect 10425 11101 10459 11135
rect 15669 11101 15703 11135
rect 21005 11101 21039 11135
rect 8125 11033 8159 11067
rect 13737 11033 13771 11067
rect 14473 11033 14507 11067
rect 4353 10965 4387 10999
rect 7205 10965 7239 10999
rect 7757 10965 7791 10999
rect 13093 10965 13127 10999
rect 15577 10965 15611 10999
rect 18153 10965 18187 10999
rect 18383 10965 18417 10999
rect 20637 10965 20671 10999
rect 1593 10761 1627 10795
rect 2421 10761 2455 10795
rect 4445 10761 4479 10795
rect 5917 10761 5951 10795
rect 6377 10761 6411 10795
rect 10425 10761 10459 10795
rect 11897 10761 11931 10795
rect 18981 10761 19015 10795
rect 19349 10761 19383 10795
rect 21281 10761 21315 10795
rect 21557 10761 21591 10795
rect 2053 10693 2087 10727
rect 14933 10693 14967 10727
rect 19993 10693 20027 10727
rect 2697 10625 2731 10659
rect 2973 10625 3007 10659
rect 7251 10625 7285 10659
rect 20269 10625 20303 10659
rect 20729 10625 20763 10659
rect 1409 10557 1443 10591
rect 4629 10557 4663 10591
rect 5089 10557 5123 10591
rect 7164 10557 7198 10591
rect 8125 10557 8159 10591
rect 8585 10557 8619 10591
rect 8953 10557 8987 10591
rect 9321 10557 9355 10591
rect 10517 10557 10551 10591
rect 11069 10557 11103 10591
rect 14289 10557 14323 10591
rect 15117 10557 15151 10591
rect 15577 10557 15611 10591
rect 15945 10557 15979 10591
rect 16313 10557 16347 10591
rect 16589 10557 16623 10591
rect 17417 10557 17451 10591
rect 18061 10557 18095 10591
rect 2789 10489 2823 10523
rect 5365 10489 5399 10523
rect 7665 10489 7699 10523
rect 10057 10489 10091 10523
rect 12817 10489 12851 10523
rect 12909 10489 12943 10523
rect 13461 10489 13495 10523
rect 14565 10489 14599 10523
rect 16865 10489 16899 10523
rect 17877 10489 17911 10523
rect 20361 10489 20395 10523
rect 3801 10421 3835 10455
rect 4077 10421 4111 10455
rect 8033 10421 8067 10455
rect 8401 10421 8435 10455
rect 10793 10421 10827 10455
rect 12265 10421 12299 10455
rect 18429 10421 18463 10455
rect 2605 10217 2639 10251
rect 4721 10217 4755 10251
rect 8677 10217 8711 10251
rect 10517 10217 10551 10251
rect 10885 10217 10919 10251
rect 12817 10217 12851 10251
rect 15577 10217 15611 10251
rect 16405 10217 16439 10251
rect 19855 10217 19889 10251
rect 21097 10217 21131 10251
rect 2047 10149 2081 10183
rect 2973 10149 3007 10183
rect 5089 10149 5123 10183
rect 5819 10149 5853 10183
rect 7389 10149 7423 10183
rect 11437 10149 11471 10183
rect 14013 10149 14047 10183
rect 18061 10149 18095 10183
rect 20269 10149 20303 10183
rect 1685 10081 1719 10115
rect 3249 10081 3283 10115
rect 3893 10081 3927 10115
rect 6377 10081 6411 10115
rect 13277 10081 13311 10115
rect 13553 10081 13587 10115
rect 15485 10081 15519 10115
rect 15853 10081 15887 10115
rect 16865 10081 16899 10115
rect 19752 10081 19786 10115
rect 20913 10081 20947 10115
rect 5457 10013 5491 10047
rect 7297 10013 7331 10047
rect 7573 10013 7607 10047
rect 11345 10013 11379 10047
rect 11621 10013 11655 10047
rect 13093 10013 13127 10047
rect 17969 10013 18003 10047
rect 18613 10013 18647 10047
rect 4215 9945 4249 9979
rect 6745 9945 6779 9979
rect 13369 9945 13403 9979
rect 3617 9877 3651 9911
rect 7113 9877 7147 9911
rect 8217 9877 8251 9911
rect 9045 9877 9079 9911
rect 15025 9877 15059 9911
rect 17003 9877 17037 9911
rect 18889 9877 18923 9911
rect 2053 9673 2087 9707
rect 5825 9673 5859 9707
rect 6653 9673 6687 9707
rect 8125 9673 8159 9707
rect 11621 9673 11655 9707
rect 16865 9673 16899 9707
rect 21557 9673 21591 9707
rect 6101 9605 6135 9639
rect 13461 9605 13495 9639
rect 14565 9605 14599 9639
rect 19073 9605 19107 9639
rect 2881 9537 2915 9571
rect 1409 9469 1443 9503
rect 4077 9469 4111 9503
rect 2973 9401 3007 9435
rect 3525 9401 3559 9435
rect 4445 9401 4479 9435
rect 4537 9401 4571 9435
rect 5089 9401 5123 9435
rect 11345 9537 11379 9571
rect 18153 9537 18187 9571
rect 20637 9537 20671 9571
rect 8861 9469 8895 9503
rect 8953 9469 8987 9503
rect 9505 9469 9539 9503
rect 12265 9469 12299 9503
rect 12449 9469 12483 9503
rect 12909 9469 12943 9503
rect 14064 9469 14098 9503
rect 15025 9469 15059 9503
rect 15485 9469 15519 9503
rect 15853 9469 15887 9503
rect 16221 9469 16255 9503
rect 6929 9401 6963 9435
rect 7021 9401 7055 9435
rect 7573 9401 7607 9435
rect 9689 9401 9723 9435
rect 10149 9401 10183 9435
rect 10701 9401 10735 9435
rect 10793 9401 10827 9435
rect 14151 9401 14185 9435
rect 14841 9401 14875 9435
rect 18245 9401 18279 9435
rect 18797 9401 18831 9435
rect 20453 9401 20487 9435
rect 20729 9401 20763 9435
rect 21281 9401 21315 9435
rect 1593 9333 1627 9367
rect 2329 9333 2363 9367
rect 5549 9333 5583 9367
rect 6101 9333 6135 9367
rect 6285 9333 6319 9367
rect 8493 9333 8527 9367
rect 10425 9333 10459 9367
rect 12725 9333 12759 9367
rect 13829 9333 13863 9367
rect 16221 9333 16255 9367
rect 17509 9333 17543 9367
rect 17877 9333 17911 9367
rect 19717 9333 19751 9367
rect 3157 9129 3191 9163
rect 3525 9129 3559 9163
rect 3893 9129 3927 9163
rect 4215 9129 4249 9163
rect 6929 9129 6963 9163
rect 9045 9129 9079 9163
rect 10057 9129 10091 9163
rect 11575 9129 11609 9163
rect 14749 9129 14783 9163
rect 15485 9129 15519 9163
rect 20637 9129 20671 9163
rect 5727 9061 5761 9095
rect 7297 9061 7331 9095
rect 11345 9061 11379 9095
rect 13046 9061 13080 9095
rect 16358 9061 16392 9095
rect 18521 9061 18555 9095
rect 18613 9061 18647 9095
rect 21005 9061 21039 9095
rect 21097 9061 21131 9095
rect 2053 8993 2087 9027
rect 2329 8993 2363 9027
rect 2789 8993 2823 9027
rect 4144 8993 4178 9027
rect 6285 8993 6319 9027
rect 9689 8993 9723 9027
rect 11472 8993 11506 9027
rect 12725 8993 12759 9027
rect 2145 8925 2179 8959
rect 5365 8925 5399 8959
rect 7205 8925 7239 8959
rect 7573 8925 7607 8959
rect 12449 8925 12483 8959
rect 13921 8925 13955 8959
rect 15025 8925 15059 8959
rect 16037 8925 16071 8959
rect 18981 8925 19015 8959
rect 21281 8925 21315 8959
rect 16957 8857 16991 8891
rect 1685 8789 1719 8823
rect 4721 8789 4755 8823
rect 4997 8789 5031 8823
rect 10609 8789 10643 8823
rect 13645 8789 13679 8823
rect 15853 8789 15887 8823
rect 18245 8789 18279 8823
rect 2881 8585 2915 8619
rect 4077 8585 4111 8619
rect 6653 8585 6687 8619
rect 10517 8585 10551 8619
rect 11897 8585 11931 8619
rect 15485 8585 15519 8619
rect 15853 8585 15887 8619
rect 17233 8585 17267 8619
rect 20913 8585 20947 8619
rect 21741 8585 21775 8619
rect 3249 8517 3283 8551
rect 7849 8517 7883 8551
rect 16957 8517 16991 8551
rect 2513 8449 2547 8483
rect 5365 8449 5399 8483
rect 6009 8449 6043 8483
rect 11437 8449 11471 8483
rect 12725 8449 12759 8483
rect 13185 8449 13219 8483
rect 13461 8449 13495 8483
rect 18245 8449 18279 8483
rect 1685 8381 1719 8415
rect 1961 8381 1995 8415
rect 3592 8381 3626 8415
rect 4721 8381 4755 8415
rect 5089 8381 5123 8415
rect 5733 8381 5767 8415
rect 6904 8381 6938 8415
rect 8033 8381 8067 8415
rect 8585 8381 8619 8415
rect 8769 8381 8803 8415
rect 9597 8381 9631 8415
rect 10793 8381 10827 8415
rect 16037 8381 16071 8415
rect 19257 8381 19291 8415
rect 19533 8381 19567 8415
rect 19809 8381 19843 8415
rect 21189 8381 21223 8415
rect 22109 8381 22143 8415
rect 9959 8313 9993 8347
rect 12265 8313 12299 8347
rect 13277 8313 13311 8347
rect 16358 8313 16392 8347
rect 17877 8313 17911 8347
rect 18337 8313 18371 8347
rect 18889 8313 18923 8347
rect 19717 8313 19751 8347
rect 1777 8245 1811 8279
rect 3663 8245 3697 8279
rect 4445 8245 4479 8279
rect 6975 8245 7009 8279
rect 7389 8245 7423 8279
rect 9137 8245 9171 8279
rect 9505 8245 9539 8279
rect 15209 8245 15243 8279
rect 21419 8245 21453 8279
rect 1685 8041 1719 8075
rect 2145 8041 2179 8075
rect 2697 8041 2731 8075
rect 7665 8041 7699 8075
rect 8125 8041 8159 8075
rect 9505 8041 9539 8075
rect 15393 8041 15427 8075
rect 19073 8041 19107 8075
rect 19625 8041 19659 8075
rect 4169 7973 4203 8007
rect 4261 7973 4295 8007
rect 6561 7973 6595 8007
rect 6745 7973 6779 8007
rect 6837 7973 6871 8007
rect 12678 7973 12712 8007
rect 18245 7973 18279 8007
rect 20913 7973 20947 8007
rect 5708 7905 5742 7939
rect 10977 7905 11011 7939
rect 11253 7905 11287 7939
rect 15301 7905 15335 7939
rect 15761 7905 15795 7939
rect 16129 7905 16163 7939
rect 16497 7905 16531 7939
rect 21005 7905 21039 7939
rect 1777 7837 1811 7871
rect 4445 7837 4479 7871
rect 7021 7837 7055 7871
rect 9781 7837 9815 7871
rect 10425 7837 10459 7871
rect 11529 7837 11563 7871
rect 12357 7837 12391 7871
rect 18153 7837 18187 7871
rect 13277 7769 13311 7803
rect 18705 7769 18739 7803
rect 5779 7701 5813 7735
rect 8861 7701 8895 7735
rect 13553 7701 13587 7735
rect 2881 7497 2915 7531
rect 6285 7497 6319 7531
rect 8677 7497 8711 7531
rect 10333 7497 10367 7531
rect 11437 7497 11471 7531
rect 11805 7497 11839 7531
rect 12633 7497 12667 7531
rect 16037 7497 16071 7531
rect 17095 7497 17129 7531
rect 21097 7497 21131 7531
rect 13461 7429 13495 7463
rect 15393 7429 15427 7463
rect 19257 7429 19291 7463
rect 21465 7429 21499 7463
rect 1777 7361 1811 7395
rect 2605 7361 2639 7395
rect 4169 7361 4203 7395
rect 6929 7361 6963 7395
rect 7389 7361 7423 7395
rect 9505 7361 9539 7395
rect 10517 7361 10551 7395
rect 10977 7361 11011 7395
rect 12265 7361 12299 7395
rect 18337 7361 18371 7395
rect 19625 7361 19659 7395
rect 4537 7293 4571 7327
rect 4997 7293 5031 7327
rect 5917 7293 5951 7327
rect 8769 7293 8803 7327
rect 8861 7293 8895 7327
rect 9045 7293 9079 7327
rect 9965 7293 9999 7327
rect 14933 7293 14967 7327
rect 15669 7293 15703 7327
rect 16992 7293 17026 7327
rect 17417 7293 17451 7327
rect 19947 7293 19981 7327
rect 20913 7293 20947 7327
rect 1961 7225 1995 7259
rect 2053 7225 2087 7259
rect 3525 7225 3559 7259
rect 3617 7225 3651 7259
rect 4905 7225 4939 7259
rect 5359 7225 5393 7259
rect 7021 7225 7055 7259
rect 8309 7225 8343 7259
rect 10609 7225 10643 7259
rect 12909 7225 12943 7259
rect 13001 7225 13035 7259
rect 18429 7225 18463 7259
rect 18981 7225 19015 7259
rect 20039 7225 20073 7259
rect 20729 7225 20763 7259
rect 3341 7157 3375 7191
rect 6653 7157 6687 7191
rect 7849 7157 7883 7191
rect 17877 7157 17911 7191
rect 20453 7157 20487 7191
rect 1593 6953 1627 6987
rect 1961 6953 1995 6987
rect 2513 6953 2547 6987
rect 3893 6953 3927 6987
rect 4261 6953 4295 6987
rect 4721 6953 4755 6987
rect 7573 6953 7607 6987
rect 14657 6953 14691 6987
rect 18521 6953 18555 6987
rect 18797 6953 18831 6987
rect 2421 6885 2455 6919
rect 6469 6885 6503 6919
rect 6745 6885 6779 6919
rect 10333 6885 10367 6919
rect 12357 6885 12391 6919
rect 17922 6885 17956 6919
rect 21005 6885 21039 6919
rect 21097 6885 21131 6919
rect 1409 6817 1443 6851
rect 4537 6817 4571 6851
rect 4997 6817 5031 6851
rect 8620 6817 8654 6851
rect 13788 6817 13822 6851
rect 15301 6817 15335 6851
rect 15853 6817 15887 6851
rect 16129 6817 16163 6851
rect 16497 6817 16531 6851
rect 19717 6817 19751 6851
rect 6101 6749 6135 6783
rect 6653 6749 6687 6783
rect 7021 6749 7055 6783
rect 8723 6749 8757 6783
rect 10241 6749 10275 6783
rect 12265 6749 12299 6783
rect 13875 6749 13909 6783
rect 16773 6749 16807 6783
rect 17601 6749 17635 6783
rect 21281 6749 21315 6783
rect 10793 6681 10827 6715
rect 12817 6681 12851 6715
rect 13185 6681 13219 6715
rect 3525 6613 3559 6647
rect 5457 6613 5491 6647
rect 14197 6613 14231 6647
rect 19947 6613 19981 6647
rect 3111 6409 3145 6443
rect 4353 6409 4387 6443
rect 7941 6409 7975 6443
rect 8677 6409 8711 6443
rect 9413 6409 9447 6443
rect 9965 6409 9999 6443
rect 11069 6409 11103 6443
rect 11897 6409 11931 6443
rect 12265 6409 12299 6443
rect 13645 6409 13679 6443
rect 16405 6409 16439 6443
rect 16773 6409 16807 6443
rect 17785 6409 17819 6443
rect 18337 6409 18371 6443
rect 19073 6409 19107 6443
rect 21833 6409 21867 6443
rect 3985 6341 4019 6375
rect 5089 6341 5123 6375
rect 5273 6341 5307 6375
rect 6929 6341 6963 6375
rect 14197 6341 14231 6375
rect 16129 6341 16163 6375
rect 19901 6341 19935 6375
rect 21465 6341 21499 6375
rect 2881 6273 2915 6307
rect 7297 6273 7331 6307
rect 10793 6273 10827 6307
rect 12909 6273 12943 6307
rect 15761 6273 15795 6307
rect 20545 6273 20579 6307
rect 2053 6205 2087 6239
rect 3040 6205 3074 6239
rect 3433 6205 3467 6239
rect 5181 6205 5215 6239
rect 5457 6205 5491 6239
rect 6285 6205 6319 6239
rect 6837 6205 6871 6239
rect 7113 6205 7147 6239
rect 8493 6205 8527 6239
rect 14105 6205 14139 6239
rect 14381 6205 14415 6239
rect 14841 6205 14875 6239
rect 17024 6205 17058 6239
rect 18705 6205 18739 6239
rect 5917 6137 5951 6171
rect 10149 6137 10183 6171
rect 10241 6137 10275 6171
rect 12633 6137 12667 6171
rect 12725 6137 12759 6171
rect 17509 6137 17543 6171
rect 20361 6137 20395 6171
rect 20637 6137 20671 6171
rect 21189 6137 21223 6171
rect 1685 6069 1719 6103
rect 2421 6069 2455 6103
rect 4721 6069 4755 6103
rect 6561 6069 6595 6103
rect 8217 6069 8251 6103
rect 11437 6069 11471 6103
rect 14013 6069 14047 6103
rect 15301 6069 15335 6103
rect 17095 6069 17129 6103
rect 2789 5865 2823 5899
rect 4169 5865 4203 5899
rect 6285 5865 6319 5899
rect 10149 5865 10183 5899
rect 12265 5865 12299 5899
rect 19073 5865 19107 5899
rect 20545 5865 20579 5899
rect 1863 5797 1897 5831
rect 3433 5797 3467 5831
rect 10425 5797 10459 5831
rect 10977 5797 11011 5831
rect 17693 5797 17727 5831
rect 19349 5797 19383 5831
rect 19441 5797 19475 5831
rect 21097 5797 21131 5831
rect 1501 5729 1535 5763
rect 2421 5729 2455 5763
rect 4077 5729 4111 5763
rect 4721 5729 4755 5763
rect 5089 5729 5123 5763
rect 5457 5729 5491 5763
rect 6469 5729 6503 5763
rect 6745 5729 6779 5763
rect 8033 5729 8067 5763
rect 8125 5729 8159 5763
rect 14264 5729 14298 5763
rect 16405 5729 16439 5763
rect 3801 5661 3835 5695
rect 7205 5661 7239 5695
rect 10333 5661 10367 5695
rect 17417 5661 17451 5695
rect 21005 5661 21039 5695
rect 21281 5661 21315 5695
rect 6561 5593 6595 5627
rect 15945 5593 15979 5627
rect 18337 5593 18371 5627
rect 19901 5593 19935 5627
rect 7573 5525 7607 5559
rect 12633 5525 12667 5559
rect 14335 5525 14369 5559
rect 15669 5525 15703 5559
rect 16543 5525 16577 5559
rect 17325 5525 17359 5559
rect 2881 5321 2915 5355
rect 6101 5321 6135 5355
rect 6377 5321 6411 5355
rect 6561 5321 6595 5355
rect 7665 5321 7699 5355
rect 2145 5185 2179 5219
rect 5549 5185 5583 5219
rect 3249 5117 3283 5151
rect 3709 5117 3743 5151
rect 4445 5117 4479 5151
rect 4721 5117 4755 5151
rect 5089 5117 5123 5151
rect 1501 5049 1535 5083
rect 1593 5049 1627 5083
rect 3525 5049 3559 5083
rect 6929 5185 6963 5219
rect 6837 5117 6871 5151
rect 7113 5117 7147 5151
rect 7665 5117 7699 5151
rect 7757 5321 7791 5355
rect 10241 5321 10275 5355
rect 10609 5321 10643 5355
rect 17785 5321 17819 5355
rect 20913 5321 20947 5355
rect 22201 5321 22235 5355
rect 18981 5253 19015 5287
rect 21189 5253 21223 5287
rect 21925 5253 21959 5287
rect 8401 5185 8435 5219
rect 14749 5185 14783 5219
rect 20545 5185 20579 5219
rect 8309 5117 8343 5151
rect 8493 5117 8527 5151
rect 10885 5117 10919 5151
rect 12265 5117 12299 5151
rect 12725 5117 12759 5151
rect 13921 5117 13955 5151
rect 14657 5117 14691 5151
rect 15485 5117 15519 5151
rect 15577 5117 15611 5151
rect 16037 5117 16071 5151
rect 16405 5117 16439 5151
rect 16865 5117 16899 5151
rect 17049 5117 17083 5151
rect 18061 5117 18095 5151
rect 21440 5117 21474 5151
rect 9873 5049 9907 5083
rect 10793 5049 10827 5083
rect 12449 5049 12483 5083
rect 17417 5049 17451 5083
rect 18382 5049 18416 5083
rect 19901 5049 19935 5083
rect 19993 5049 20027 5083
rect 2421 4981 2455 5015
rect 3801 4981 3835 5015
rect 6377 4981 6411 5015
rect 7849 4981 7883 5015
rect 15117 4981 15151 5015
rect 19349 4981 19383 5015
rect 19717 4981 19751 5015
rect 21511 4981 21545 5015
rect 1685 4777 1719 4811
rect 3433 4777 3467 4811
rect 6193 4777 6227 4811
rect 9781 4777 9815 4811
rect 12081 4777 12115 4811
rect 14197 4777 14231 4811
rect 17509 4777 17543 4811
rect 18337 4777 18371 4811
rect 1961 4709 1995 4743
rect 4445 4709 4479 4743
rect 6561 4709 6595 4743
rect 17049 4709 17083 4743
rect 19349 4709 19383 4743
rect 19901 4709 19935 4743
rect 20913 4709 20947 4743
rect 6653 4641 6687 4675
rect 6929 4641 6963 4675
rect 8125 4641 8159 4675
rect 8769 4641 8803 4675
rect 9965 4641 9999 4675
rect 10425 4641 10459 4675
rect 10701 4641 10735 4675
rect 10885 4641 10919 4675
rect 11805 4641 11839 4675
rect 12265 4641 12299 4675
rect 12725 4641 12759 4675
rect 12817 4641 12851 4675
rect 13185 4641 13219 4675
rect 15025 4641 15059 4675
rect 15853 4641 15887 4675
rect 16037 4641 16071 4675
rect 16405 4641 16439 4675
rect 16773 4641 16807 4675
rect 17944 4641 17978 4675
rect 21005 4641 21039 4675
rect 1869 4573 1903 4607
rect 2145 4573 2179 4607
rect 4353 4573 4387 4607
rect 4721 4573 4755 4607
rect 6745 4573 6779 4607
rect 7389 4573 7423 4607
rect 13737 4573 13771 4607
rect 19257 4573 19291 4607
rect 8033 4505 8067 4539
rect 3709 4437 3743 4471
rect 8355 4437 8389 4471
rect 18015 4437 18049 4471
rect 2329 4233 2363 4267
rect 5457 4233 5491 4267
rect 5779 4233 5813 4267
rect 6653 4233 6687 4267
rect 7481 4233 7515 4267
rect 11253 4233 11287 4267
rect 17233 4233 17267 4267
rect 18337 4233 18371 4267
rect 18889 4233 18923 4267
rect 20913 4233 20947 4267
rect 3617 4165 3651 4199
rect 3709 4165 3743 4199
rect 7757 4165 7791 4199
rect 10149 4165 10183 4199
rect 15669 4165 15703 4199
rect 2605 4097 2639 4131
rect 3433 4029 3467 4063
rect 11621 4097 11655 4131
rect 13461 4097 13495 4131
rect 15945 4097 15979 4131
rect 17601 4097 17635 4131
rect 3893 4029 3927 4063
rect 5676 4029 5710 4063
rect 6101 4029 6135 4063
rect 6996 4029 7030 4063
rect 8125 4029 8159 4063
rect 8401 4029 8435 4063
rect 8769 4029 8803 4063
rect 9321 4029 9355 4063
rect 10609 4029 10643 4063
rect 12516 4029 12550 4063
rect 13829 4029 13863 4063
rect 14197 4029 14231 4063
rect 14381 4029 14415 4063
rect 14933 4029 14967 4063
rect 19073 4029 19107 4063
rect 1409 3961 1443 3995
rect 1869 3961 1903 3995
rect 3617 3961 3651 3995
rect 4214 3961 4248 3995
rect 10241 3961 10275 3995
rect 13001 3961 13035 3995
rect 16037 3961 16071 3995
rect 16589 3961 16623 3995
rect 19717 3961 19751 3995
rect 19993 3961 20027 3995
rect 4813 3893 4847 3927
rect 5089 3893 5123 3927
rect 7067 3893 7101 3927
rect 8033 3893 8067 3927
rect 9689 3893 9723 3927
rect 11989 3893 12023 3927
rect 12587 3893 12621 3927
rect 14749 3893 14783 3927
rect 16957 3893 16991 3927
rect 6745 3689 6779 3723
rect 8677 3689 8711 3723
rect 9413 3689 9447 3723
rect 11713 3689 11747 3723
rect 12725 3689 12759 3723
rect 13369 3689 13403 3723
rect 14749 3689 14783 3723
rect 15025 3689 15059 3723
rect 16313 3689 16347 3723
rect 16681 3689 16715 3723
rect 18107 3689 18141 3723
rect 19257 3689 19291 3723
rect 19441 3689 19475 3723
rect 21051 3689 21085 3723
rect 7389 3621 7423 3655
rect 9965 3621 9999 3655
rect 12126 3621 12160 3655
rect 15393 3621 15427 3655
rect 15485 3621 15519 3655
rect 4813 3553 4847 3587
rect 5733 3553 5767 3587
rect 8309 3553 8343 3587
rect 14289 3553 14323 3587
rect 16865 3553 16899 3587
rect 18036 3553 18070 3587
rect 20980 3553 21014 3587
rect 7297 3485 7331 3519
rect 9689 3485 9723 3519
rect 11805 3485 11839 3519
rect 14381 3485 14415 3519
rect 7849 3417 7883 3451
rect 13093 3417 13127 3451
rect 15945 3417 15979 3451
rect 17049 3417 17083 3451
rect 4445 3349 4479 3383
rect 5273 3349 5307 3383
rect 5871 3349 5905 3383
rect 7021 3349 7055 3383
rect 10609 3349 10643 3383
rect 10885 3349 10919 3383
rect 11253 3349 11287 3383
rect 1593 3145 1627 3179
rect 3341 3145 3375 3179
rect 4353 3145 4387 3179
rect 6561 3145 6595 3179
rect 8401 3145 8435 3179
rect 10977 3145 11011 3179
rect 13645 3145 13679 3179
rect 15025 3145 15059 3179
rect 15393 3145 15427 3179
rect 15669 3145 15703 3179
rect 16865 3145 16899 3179
rect 19349 3145 19383 3179
rect 21051 3145 21085 3179
rect 21465 3145 21499 3179
rect 3571 3077 3605 3111
rect 11345 3077 11379 3111
rect 14013 3077 14047 3111
rect 4537 3009 4571 3043
rect 4813 3009 4847 3043
rect 6285 3009 6319 3043
rect 6837 3009 6871 3043
rect 8585 3009 8619 3043
rect 9689 3009 9723 3043
rect 10609 3009 10643 3043
rect 12633 3009 12667 3043
rect 13277 3009 13311 3043
rect 14105 3009 14139 3043
rect 16221 3009 16255 3043
rect 1409 2941 1443 2975
rect 3500 2941 3534 2975
rect 3893 2941 3927 2975
rect 7757 2941 7791 2975
rect 8125 2941 8159 2975
rect 11161 2941 11195 2975
rect 19140 2941 19174 2975
rect 19533 2941 19567 2975
rect 20980 2941 21014 2975
rect 4629 2873 4663 2907
rect 7158 2873 7192 2907
rect 9137 2873 9171 2907
rect 9781 2873 9815 2907
rect 10333 2873 10367 2907
rect 12265 2873 12299 2907
rect 12725 2873 12759 2907
rect 15945 2873 15979 2907
rect 16037 2873 16071 2907
rect 2053 2805 2087 2839
rect 5825 2805 5859 2839
rect 9413 2805 9447 2839
rect 11805 2805 11839 2839
rect 14473 2805 14507 2839
rect 18061 2805 18095 2839
rect 18613 2805 18647 2839
rect 21833 2805 21867 2839
rect 1547 2601 1581 2635
rect 4215 2601 4249 2635
rect 8815 2601 8849 2635
rect 11897 2601 11931 2635
rect 12449 2601 12483 2635
rect 14381 2601 14415 2635
rect 16497 2601 16531 2635
rect 20085 2601 20119 2635
rect 3157 2533 3191 2567
rect 7297 2533 7331 2567
rect 7849 2533 7883 2567
rect 9137 2533 9171 2567
rect 9597 2533 9631 2567
rect 9965 2533 9999 2567
rect 11253 2533 11287 2567
rect 12817 2533 12851 2567
rect 13369 2533 13403 2567
rect 15301 2533 15335 2567
rect 15646 2533 15680 2567
rect 1444 2465 1478 2499
rect 1869 2465 1903 2499
rect 2513 2465 2547 2499
rect 4144 2465 4178 2499
rect 5181 2465 5215 2499
rect 5365 2465 5399 2499
rect 8712 2465 8746 2499
rect 11345 2465 11379 2499
rect 14105 2465 14139 2499
rect 17049 2465 17083 2499
rect 17601 2465 17635 2499
rect 18337 2465 18371 2499
rect 19533 2465 19567 2499
rect 21256 2465 21290 2499
rect 6009 2397 6043 2431
rect 6653 2397 6687 2431
rect 7205 2397 7239 2431
rect 9873 2397 9907 2431
rect 10333 2397 10367 2431
rect 12725 2397 12759 2431
rect 13645 2397 13679 2431
rect 14933 2397 14967 2431
rect 15577 2397 15611 2431
rect 18981 2397 19015 2431
rect 6377 2329 6411 2363
rect 8585 2329 8619 2363
rect 11529 2329 11563 2363
rect 16129 2329 16163 2363
rect 19717 2329 19751 2363
rect 2237 2261 2271 2295
rect 4629 2261 4663 2295
rect 17233 2261 17267 2295
rect 18521 2261 18555 2295
rect 21327 2261 21361 2295
rect 21741 2261 21775 2295
<< metal1 >>
rect 14 23536 20 23588
rect 72 23576 78 23588
rect 566 23576 572 23588
rect 72 23548 572 23576
rect 72 23536 78 23548
rect 566 23536 572 23548
rect 624 23536 630 23588
rect 1104 21786 22816 21808
rect 1104 21734 4982 21786
rect 5034 21734 5046 21786
rect 5098 21734 5110 21786
rect 5162 21734 5174 21786
rect 5226 21734 12982 21786
rect 13034 21734 13046 21786
rect 13098 21734 13110 21786
rect 13162 21734 13174 21786
rect 13226 21734 20982 21786
rect 21034 21734 21046 21786
rect 21098 21734 21110 21786
rect 21162 21734 21174 21786
rect 21226 21734 22816 21786
rect 1104 21712 22816 21734
rect 20070 21672 20076 21684
rect 20031 21644 20076 21672
rect 20070 21632 20076 21644
rect 20128 21632 20134 21684
rect 8548 21471 8606 21477
rect 8548 21437 8560 21471
rect 8594 21468 8606 21471
rect 19588 21471 19646 21477
rect 8594 21440 9076 21468
rect 8594 21437 8606 21440
rect 8548 21431 8606 21437
rect 8386 21292 8392 21344
rect 8444 21332 8450 21344
rect 9048 21341 9076 21440
rect 19588 21437 19600 21471
rect 19634 21468 19646 21471
rect 20070 21468 20076 21480
rect 19634 21440 20076 21468
rect 19634 21437 19646 21440
rect 19588 21431 19646 21437
rect 20070 21428 20076 21440
rect 20128 21428 20134 21480
rect 8619 21335 8677 21341
rect 8619 21332 8631 21335
rect 8444 21304 8631 21332
rect 8444 21292 8450 21304
rect 8619 21301 8631 21304
rect 8665 21301 8677 21335
rect 8619 21295 8677 21301
rect 9033 21335 9091 21341
rect 9033 21301 9045 21335
rect 9079 21332 9091 21335
rect 10042 21332 10048 21344
rect 9079 21304 10048 21332
rect 9079 21301 9091 21304
rect 9033 21295 9091 21301
rect 10042 21292 10048 21304
rect 10100 21292 10106 21344
rect 19334 21292 19340 21344
rect 19392 21332 19398 21344
rect 19659 21335 19717 21341
rect 19659 21332 19671 21335
rect 19392 21304 19671 21332
rect 19392 21292 19398 21304
rect 19659 21301 19671 21304
rect 19705 21301 19717 21335
rect 19659 21295 19717 21301
rect 1104 21242 22816 21264
rect 1104 21190 8982 21242
rect 9034 21190 9046 21242
rect 9098 21190 9110 21242
rect 9162 21190 9174 21242
rect 9226 21190 16982 21242
rect 17034 21190 17046 21242
rect 17098 21190 17110 21242
rect 17162 21190 17174 21242
rect 17226 21190 22816 21242
rect 1104 21168 22816 21190
rect 8573 21131 8631 21137
rect 8573 21097 8585 21131
rect 8619 21128 8631 21131
rect 9306 21128 9312 21140
rect 8619 21100 9312 21128
rect 8619 21097 8631 21100
rect 8573 21091 8631 21097
rect 9306 21088 9312 21100
rect 9364 21088 9370 21140
rect 12529 21131 12587 21137
rect 12529 21097 12541 21131
rect 12575 21128 12587 21131
rect 13262 21128 13268 21140
rect 12575 21100 13268 21128
rect 12575 21097 12587 21100
rect 12529 21091 12587 21097
rect 13262 21088 13268 21100
rect 13320 21088 13326 21140
rect 18233 21131 18291 21137
rect 18233 21097 18245 21131
rect 18279 21128 18291 21131
rect 19242 21128 19248 21140
rect 18279 21100 19248 21128
rect 18279 21097 18291 21100
rect 18233 21091 18291 21097
rect 19242 21088 19248 21100
rect 19300 21088 19306 21140
rect 12342 20992 12348 21004
rect 12303 20964 12348 20992
rect 12342 20952 12348 20964
rect 12400 20952 12406 21004
rect 18046 20992 18052 21004
rect 18007 20964 18052 20992
rect 18046 20952 18052 20964
rect 18104 20952 18110 21004
rect 19864 20995 19922 21001
rect 19864 20961 19876 20995
rect 19910 20992 19922 20995
rect 19978 20992 19984 21004
rect 19910 20964 19984 20992
rect 19910 20961 19922 20964
rect 19864 20955 19922 20961
rect 19978 20952 19984 20964
rect 20036 20952 20042 21004
rect 19518 20748 19524 20800
rect 19576 20788 19582 20800
rect 19935 20791 19993 20797
rect 19935 20788 19947 20791
rect 19576 20760 19947 20788
rect 19576 20748 19582 20760
rect 19935 20757 19947 20760
rect 19981 20757 19993 20791
rect 19935 20751 19993 20757
rect 1104 20698 22816 20720
rect 1104 20646 4982 20698
rect 5034 20646 5046 20698
rect 5098 20646 5110 20698
rect 5162 20646 5174 20698
rect 5226 20646 12982 20698
rect 13034 20646 13046 20698
rect 13098 20646 13110 20698
rect 13162 20646 13174 20698
rect 13226 20646 20982 20698
rect 21034 20646 21046 20698
rect 21098 20646 21110 20698
rect 21162 20646 21174 20698
rect 21226 20646 22816 20698
rect 1104 20624 22816 20646
rect 2685 20587 2743 20593
rect 2685 20553 2697 20587
rect 2731 20584 2743 20587
rect 2774 20584 2780 20596
rect 2731 20556 2780 20584
rect 2731 20553 2743 20556
rect 2685 20547 2743 20553
rect 2200 20383 2258 20389
rect 2200 20349 2212 20383
rect 2246 20380 2258 20383
rect 2700 20380 2728 20547
rect 2774 20544 2780 20556
rect 2832 20544 2838 20596
rect 4522 20584 4528 20596
rect 4483 20556 4528 20584
rect 4522 20544 4528 20556
rect 4580 20544 4586 20596
rect 7926 20584 7932 20596
rect 7887 20556 7932 20584
rect 7926 20544 7932 20556
rect 7984 20544 7990 20596
rect 8386 20584 8392 20596
rect 8347 20556 8392 20584
rect 8386 20544 8392 20556
rect 8444 20544 8450 20596
rect 14182 20584 14188 20596
rect 14143 20556 14188 20584
rect 14182 20544 14188 20556
rect 14240 20544 14246 20596
rect 17221 20587 17279 20593
rect 17221 20553 17233 20587
rect 17267 20584 17279 20587
rect 17862 20584 17868 20596
rect 17267 20556 17868 20584
rect 17267 20553 17279 20556
rect 17221 20547 17279 20553
rect 12250 20408 12256 20460
rect 12308 20448 12314 20460
rect 12805 20451 12863 20457
rect 12805 20448 12817 20451
rect 12308 20420 12817 20448
rect 12308 20408 12314 20420
rect 12805 20417 12817 20420
rect 12851 20417 12863 20451
rect 12805 20411 12863 20417
rect 2246 20352 2728 20380
rect 4132 20383 4190 20389
rect 2246 20349 2258 20352
rect 2200 20343 2258 20349
rect 4132 20349 4144 20383
rect 4178 20380 4190 20383
rect 4522 20380 4528 20392
rect 4178 20352 4528 20380
rect 4178 20349 4190 20352
rect 4132 20343 4190 20349
rect 4522 20340 4528 20352
rect 4580 20340 4586 20392
rect 7745 20383 7803 20389
rect 7745 20349 7757 20383
rect 7791 20380 7803 20383
rect 8386 20380 8392 20392
rect 7791 20352 8392 20380
rect 7791 20349 7803 20352
rect 7745 20343 7803 20349
rect 8386 20340 8392 20352
rect 8444 20340 8450 20392
rect 13906 20340 13912 20392
rect 13964 20380 13970 20392
rect 14001 20383 14059 20389
rect 14001 20380 14013 20383
rect 13964 20352 14013 20380
rect 13964 20340 13970 20352
rect 14001 20349 14013 20352
rect 14047 20380 14059 20383
rect 14553 20383 14611 20389
rect 14553 20380 14565 20383
rect 14047 20352 14565 20380
rect 14047 20349 14059 20352
rect 14001 20343 14059 20349
rect 14553 20349 14565 20352
rect 14599 20349 14611 20383
rect 14553 20343 14611 20349
rect 16736 20383 16794 20389
rect 16736 20349 16748 20383
rect 16782 20380 16794 20383
rect 17236 20380 17264 20547
rect 17862 20544 17868 20556
rect 17920 20544 17926 20596
rect 19153 20587 19211 20593
rect 19153 20553 19165 20587
rect 19199 20584 19211 20587
rect 20438 20584 20444 20596
rect 19199 20556 20444 20584
rect 19199 20553 19211 20556
rect 19153 20547 19211 20553
rect 20438 20544 20444 20556
rect 20496 20544 20502 20596
rect 21085 20587 21143 20593
rect 21085 20553 21097 20587
rect 21131 20584 21143 20587
rect 21726 20584 21732 20596
rect 21131 20556 21732 20584
rect 21131 20553 21143 20556
rect 21085 20547 21143 20553
rect 21726 20544 21732 20556
rect 21784 20544 21790 20596
rect 19978 20516 19984 20528
rect 19939 20488 19984 20516
rect 19978 20476 19984 20488
rect 20036 20476 20042 20528
rect 18966 20380 18972 20392
rect 16782 20352 17264 20380
rect 18927 20352 18972 20380
rect 16782 20349 16794 20352
rect 16736 20343 16794 20349
rect 18966 20340 18972 20352
rect 19024 20380 19030 20392
rect 19521 20383 19579 20389
rect 19521 20380 19533 20383
rect 19024 20352 19533 20380
rect 19024 20340 19030 20352
rect 19521 20349 19533 20352
rect 19567 20349 19579 20383
rect 19521 20343 19579 20349
rect 19886 20340 19892 20392
rect 19944 20380 19950 20392
rect 20901 20383 20959 20389
rect 20901 20380 20913 20383
rect 19944 20352 20913 20380
rect 19944 20340 19950 20352
rect 20901 20349 20913 20352
rect 20947 20380 20959 20383
rect 21453 20383 21511 20389
rect 21453 20380 21465 20383
rect 20947 20352 21465 20380
rect 20947 20349 20959 20352
rect 20901 20343 20959 20349
rect 21453 20349 21465 20352
rect 21499 20349 21511 20383
rect 21453 20343 21511 20349
rect 9398 20312 9404 20324
rect 9359 20284 9404 20312
rect 9398 20272 9404 20284
rect 9456 20272 9462 20324
rect 9493 20315 9551 20321
rect 9493 20281 9505 20315
rect 9539 20281 9551 20315
rect 10042 20312 10048 20324
rect 10003 20284 10048 20312
rect 9493 20275 9551 20281
rect 2271 20247 2329 20253
rect 2271 20213 2283 20247
rect 2317 20244 2329 20247
rect 2406 20244 2412 20256
rect 2317 20216 2412 20244
rect 2317 20213 2329 20216
rect 2271 20207 2329 20213
rect 2406 20204 2412 20216
rect 2464 20204 2470 20256
rect 4203 20247 4261 20253
rect 4203 20213 4215 20247
rect 4249 20244 4261 20247
rect 8846 20244 8852 20256
rect 4249 20216 8852 20244
rect 4249 20213 4261 20216
rect 4203 20207 4261 20213
rect 8846 20204 8852 20216
rect 8904 20204 8910 20256
rect 9217 20247 9275 20253
rect 9217 20213 9229 20247
rect 9263 20244 9275 20247
rect 9306 20244 9312 20256
rect 9263 20216 9312 20244
rect 9263 20213 9275 20216
rect 9217 20207 9275 20213
rect 9306 20204 9312 20216
rect 9364 20244 9370 20256
rect 9508 20244 9536 20275
rect 10042 20272 10048 20284
rect 10100 20272 10106 20324
rect 11885 20315 11943 20321
rect 11885 20281 11897 20315
rect 11931 20312 11943 20315
rect 12526 20312 12532 20324
rect 11931 20284 12532 20312
rect 11931 20281 11943 20284
rect 11885 20275 11943 20281
rect 12526 20272 12532 20284
rect 12584 20272 12590 20324
rect 12618 20272 12624 20324
rect 12676 20312 12682 20324
rect 12676 20284 12721 20312
rect 12676 20272 12682 20284
rect 16390 20272 16396 20324
rect 16448 20312 16454 20324
rect 18046 20312 18052 20324
rect 16448 20284 18052 20312
rect 16448 20272 16454 20284
rect 18046 20272 18052 20284
rect 18104 20312 18110 20324
rect 18233 20315 18291 20321
rect 18233 20312 18245 20315
rect 18104 20284 18245 20312
rect 18104 20272 18110 20284
rect 18233 20281 18245 20284
rect 18279 20281 18291 20315
rect 18233 20275 18291 20281
rect 9364 20216 9536 20244
rect 11333 20247 11391 20253
rect 9364 20204 9370 20216
rect 11333 20213 11345 20247
rect 11379 20244 11391 20247
rect 11606 20244 11612 20256
rect 11379 20216 11612 20244
rect 11379 20213 11391 20216
rect 11333 20207 11391 20213
rect 11606 20204 11612 20216
rect 11664 20204 11670 20256
rect 12253 20247 12311 20253
rect 12253 20213 12265 20247
rect 12299 20244 12311 20247
rect 12342 20244 12348 20256
rect 12299 20216 12348 20244
rect 12299 20213 12311 20216
rect 12253 20207 12311 20213
rect 12342 20204 12348 20216
rect 12400 20204 12406 20256
rect 14734 20204 14740 20256
rect 14792 20244 14798 20256
rect 16807 20247 16865 20253
rect 16807 20244 16819 20247
rect 14792 20216 16819 20244
rect 14792 20204 14798 20216
rect 16807 20213 16819 20216
rect 16853 20213 16865 20247
rect 16807 20207 16865 20213
rect 1104 20154 22816 20176
rect 1104 20102 8982 20154
rect 9034 20102 9046 20154
rect 9098 20102 9110 20154
rect 9162 20102 9174 20154
rect 9226 20102 16982 20154
rect 17034 20102 17046 20154
rect 17098 20102 17110 20154
rect 17162 20102 17174 20154
rect 17226 20102 22816 20154
rect 1104 20080 22816 20102
rect 18874 20000 18880 20052
rect 18932 20040 18938 20052
rect 18932 20012 19472 20040
rect 18932 20000 18938 20012
rect 8757 19975 8815 19981
rect 8757 19941 8769 19975
rect 8803 19972 8815 19975
rect 9766 19972 9772 19984
rect 8803 19944 9772 19972
rect 8803 19941 8815 19944
rect 8757 19935 8815 19941
rect 9766 19932 9772 19944
rect 9824 19972 9830 19984
rect 9861 19975 9919 19981
rect 9861 19972 9873 19975
rect 9824 19944 9873 19972
rect 9824 19932 9830 19944
rect 9861 19941 9873 19944
rect 9907 19941 9919 19975
rect 11698 19972 11704 19984
rect 11659 19944 11704 19972
rect 9861 19935 9919 19941
rect 11698 19932 11704 19944
rect 11756 19972 11762 19984
rect 12529 19975 12587 19981
rect 12529 19972 12541 19975
rect 11756 19944 12541 19972
rect 11756 19932 11762 19944
rect 12529 19941 12541 19944
rect 12575 19972 12587 19975
rect 12618 19972 12624 19984
rect 12575 19944 12624 19972
rect 12575 19941 12587 19944
rect 12529 19935 12587 19941
rect 12618 19932 12624 19944
rect 12676 19932 12682 19984
rect 13265 19975 13323 19981
rect 13265 19941 13277 19975
rect 13311 19972 13323 19975
rect 13354 19972 13360 19984
rect 13311 19944 13360 19972
rect 13311 19941 13323 19944
rect 13265 19935 13323 19941
rect 13354 19932 13360 19944
rect 13412 19932 13418 19984
rect 17313 19975 17371 19981
rect 17313 19941 17325 19975
rect 17359 19972 17371 19975
rect 17494 19972 17500 19984
rect 17359 19944 17500 19972
rect 17359 19941 17371 19944
rect 17313 19935 17371 19941
rect 17494 19932 17500 19944
rect 17552 19932 17558 19984
rect 19334 19972 19340 19984
rect 19295 19944 19340 19972
rect 19334 19932 19340 19944
rect 19392 19932 19398 19984
rect 19444 19981 19472 20012
rect 19429 19975 19487 19981
rect 19429 19941 19441 19975
rect 19475 19941 19487 19975
rect 19429 19935 19487 19941
rect 1464 19907 1522 19913
rect 1464 19873 1476 19907
rect 1510 19904 1522 19907
rect 1578 19904 1584 19916
rect 1510 19876 1584 19904
rect 1510 19873 1522 19876
rect 1464 19867 1522 19873
rect 1578 19864 1584 19876
rect 1636 19864 1642 19916
rect 8018 19864 8024 19916
rect 8076 19904 8082 19916
rect 8113 19907 8171 19913
rect 8113 19904 8125 19907
rect 8076 19876 8125 19904
rect 8076 19864 8082 19876
rect 8113 19873 8125 19876
rect 8159 19873 8171 19907
rect 15838 19904 15844 19916
rect 15799 19876 15844 19904
rect 8113 19867 8171 19873
rect 15838 19864 15844 19876
rect 15896 19864 15902 19916
rect 20806 19864 20812 19916
rect 20864 19904 20870 19916
rect 20968 19907 21026 19913
rect 20968 19904 20980 19907
rect 20864 19876 20980 19904
rect 20864 19864 20870 19876
rect 20968 19873 20980 19876
rect 21014 19904 21026 19907
rect 23014 19904 23020 19916
rect 21014 19876 23020 19904
rect 21014 19873 21026 19876
rect 20968 19867 21026 19873
rect 23014 19864 23020 19876
rect 23072 19864 23078 19916
rect 9769 19839 9827 19845
rect 9769 19805 9781 19839
rect 9815 19805 9827 19839
rect 10042 19836 10048 19848
rect 10003 19808 10048 19836
rect 9769 19799 9827 19805
rect 9784 19768 9812 19799
rect 10042 19796 10048 19808
rect 10100 19796 10106 19848
rect 11606 19836 11612 19848
rect 11567 19808 11612 19836
rect 11606 19796 11612 19808
rect 11664 19796 11670 19848
rect 13173 19839 13231 19845
rect 13173 19805 13185 19839
rect 13219 19836 13231 19839
rect 13538 19836 13544 19848
rect 13219 19808 13544 19836
rect 13219 19805 13231 19808
rect 13173 19799 13231 19805
rect 13538 19796 13544 19808
rect 13596 19796 13602 19848
rect 17218 19836 17224 19848
rect 17179 19808 17224 19836
rect 17218 19796 17224 19808
rect 17276 19796 17282 19848
rect 17865 19839 17923 19845
rect 17865 19805 17877 19839
rect 17911 19836 17923 19839
rect 19058 19836 19064 19848
rect 17911 19808 19064 19836
rect 17911 19805 17923 19808
rect 17865 19799 17923 19805
rect 19058 19796 19064 19808
rect 19116 19796 19122 19848
rect 19978 19836 19984 19848
rect 19939 19808 19984 19836
rect 19978 19796 19984 19808
rect 20036 19796 20042 19848
rect 10134 19768 10140 19780
rect 9784 19740 10140 19768
rect 10134 19728 10140 19740
rect 10192 19768 10198 19780
rect 12161 19771 12219 19777
rect 12161 19768 12173 19771
rect 10192 19740 12173 19768
rect 10192 19728 10198 19740
rect 12161 19737 12173 19740
rect 12207 19768 12219 19771
rect 13725 19771 13783 19777
rect 13725 19768 13737 19771
rect 12207 19740 13737 19768
rect 12207 19737 12219 19740
rect 12161 19731 12219 19737
rect 13725 19737 13737 19740
rect 13771 19737 13783 19771
rect 13725 19731 13783 19737
rect 1535 19703 1593 19709
rect 1535 19669 1547 19703
rect 1581 19700 1593 19703
rect 2866 19700 2872 19712
rect 1581 19672 2872 19700
rect 1581 19669 1593 19672
rect 1535 19663 1593 19669
rect 2866 19660 2872 19672
rect 2924 19660 2930 19712
rect 9398 19700 9404 19712
rect 9311 19672 9404 19700
rect 9398 19660 9404 19672
rect 9456 19700 9462 19712
rect 12250 19700 12256 19712
rect 9456 19672 12256 19700
rect 9456 19660 9462 19672
rect 12250 19660 12256 19672
rect 12308 19660 12314 19712
rect 16071 19703 16129 19709
rect 16071 19669 16083 19703
rect 16117 19700 16129 19703
rect 16298 19700 16304 19712
rect 16117 19672 16304 19700
rect 16117 19669 16129 19672
rect 16071 19663 16129 19669
rect 16298 19660 16304 19672
rect 16356 19660 16362 19712
rect 16485 19703 16543 19709
rect 16485 19669 16497 19703
rect 16531 19700 16543 19703
rect 16574 19700 16580 19712
rect 16531 19672 16580 19700
rect 16531 19669 16543 19672
rect 16485 19663 16543 19669
rect 16574 19660 16580 19672
rect 16632 19660 16638 19712
rect 20714 19660 20720 19712
rect 20772 19700 20778 19712
rect 21039 19703 21097 19709
rect 21039 19700 21051 19703
rect 20772 19672 21051 19700
rect 20772 19660 20778 19672
rect 21039 19669 21051 19672
rect 21085 19669 21097 19703
rect 21039 19663 21097 19669
rect 1104 19610 22816 19632
rect 1104 19558 4982 19610
rect 5034 19558 5046 19610
rect 5098 19558 5110 19610
rect 5162 19558 5174 19610
rect 5226 19558 12982 19610
rect 13034 19558 13046 19610
rect 13098 19558 13110 19610
rect 13162 19558 13174 19610
rect 13226 19558 20982 19610
rect 21034 19558 21046 19610
rect 21098 19558 21110 19610
rect 21162 19558 21174 19610
rect 21226 19558 22816 19610
rect 1104 19536 22816 19558
rect 1578 19496 1584 19508
rect 1539 19468 1584 19496
rect 1578 19456 1584 19468
rect 1636 19456 1642 19508
rect 8018 19496 8024 19508
rect 7979 19468 8024 19496
rect 8018 19456 8024 19468
rect 8076 19496 8082 19508
rect 9306 19496 9312 19508
rect 8076 19468 9312 19496
rect 8076 19456 8082 19468
rect 9306 19456 9312 19468
rect 9364 19496 9370 19508
rect 9401 19499 9459 19505
rect 9401 19496 9413 19499
rect 9364 19468 9413 19496
rect 9364 19456 9370 19468
rect 9401 19465 9413 19468
rect 9447 19465 9459 19499
rect 9766 19496 9772 19508
rect 9727 19468 9772 19496
rect 9401 19459 9459 19465
rect 9766 19456 9772 19468
rect 9824 19456 9830 19508
rect 10134 19496 10140 19508
rect 10095 19468 10140 19496
rect 10134 19456 10140 19468
rect 10192 19456 10198 19508
rect 11606 19456 11612 19508
rect 11664 19496 11670 19508
rect 12161 19499 12219 19505
rect 12161 19496 12173 19499
rect 11664 19468 12173 19496
rect 11664 19456 11670 19468
rect 12161 19465 12173 19468
rect 12207 19465 12219 19499
rect 13354 19496 13360 19508
rect 12161 19459 12219 19465
rect 12268 19468 13360 19496
rect 11517 19363 11575 19369
rect 11517 19329 11529 19363
rect 11563 19360 11575 19363
rect 11698 19360 11704 19372
rect 11563 19332 11704 19360
rect 11563 19329 11575 19332
rect 11517 19323 11575 19329
rect 11698 19320 11704 19332
rect 11756 19360 11762 19372
rect 11793 19363 11851 19369
rect 11793 19360 11805 19363
rect 11756 19332 11805 19360
rect 11756 19320 11762 19332
rect 11793 19329 11805 19332
rect 11839 19329 11851 19363
rect 11793 19323 11851 19329
rect 8481 19295 8539 19301
rect 8481 19261 8493 19295
rect 8527 19292 8539 19295
rect 8570 19292 8576 19304
rect 8527 19264 8576 19292
rect 8527 19261 8539 19264
rect 8481 19255 8539 19261
rect 8570 19252 8576 19264
rect 8628 19252 8634 19304
rect 10686 19292 10692 19304
rect 10599 19264 10692 19292
rect 10686 19252 10692 19264
rect 10744 19292 10750 19304
rect 11425 19295 11483 19301
rect 11425 19292 11437 19295
rect 10744 19264 11437 19292
rect 10744 19252 10750 19264
rect 11425 19261 11437 19264
rect 11471 19292 11483 19295
rect 11606 19292 11612 19304
rect 11471 19264 11612 19292
rect 11471 19261 11483 19264
rect 11425 19255 11483 19261
rect 11606 19252 11612 19264
rect 11664 19292 11670 19304
rect 12268 19292 12296 19468
rect 13354 19456 13360 19468
rect 13412 19456 13418 19508
rect 13906 19496 13912 19508
rect 13867 19468 13912 19496
rect 13906 19456 13912 19468
rect 13964 19456 13970 19508
rect 18417 19499 18475 19505
rect 18417 19465 18429 19499
rect 18463 19496 18475 19499
rect 19334 19496 19340 19508
rect 18463 19468 19340 19496
rect 18463 19465 18475 19468
rect 18417 19459 18475 19465
rect 19334 19456 19340 19468
rect 19392 19456 19398 19508
rect 20806 19456 20812 19508
rect 20864 19496 20870 19508
rect 20901 19499 20959 19505
rect 20901 19496 20913 19499
rect 20864 19468 20913 19496
rect 20864 19456 20870 19468
rect 20901 19465 20913 19468
rect 20947 19465 20959 19499
rect 21634 19496 21640 19508
rect 21595 19468 21640 19496
rect 20901 19459 20959 19465
rect 21634 19456 21640 19468
rect 21692 19456 21698 19508
rect 12526 19388 12532 19440
rect 12584 19428 12590 19440
rect 14734 19428 14740 19440
rect 12584 19400 14740 19428
rect 12584 19388 12590 19400
rect 14734 19388 14740 19400
rect 14792 19388 14798 19440
rect 19978 19388 19984 19440
rect 20036 19428 20042 19440
rect 20165 19431 20223 19437
rect 20165 19428 20177 19431
rect 20036 19400 20177 19428
rect 20036 19388 20042 19400
rect 20165 19397 20177 19400
rect 20211 19397 20223 19431
rect 20165 19391 20223 19397
rect 16206 19320 16212 19372
rect 16264 19360 16270 19372
rect 17218 19360 17224 19372
rect 16264 19332 17224 19360
rect 16264 19320 16270 19332
rect 17218 19320 17224 19332
rect 17276 19360 17282 19372
rect 17773 19363 17831 19369
rect 17773 19360 17785 19363
rect 17276 19332 17785 19360
rect 17276 19320 17282 19332
rect 17773 19329 17785 19332
rect 17819 19329 17831 19363
rect 17773 19323 17831 19329
rect 19613 19363 19671 19369
rect 19613 19329 19625 19363
rect 19659 19360 19671 19363
rect 19659 19332 20668 19360
rect 19659 19329 19671 19332
rect 19613 19323 19671 19329
rect 11664 19264 12296 19292
rect 12488 19295 12546 19301
rect 11664 19252 11670 19264
rect 12488 19261 12500 19295
rect 12534 19292 12546 19295
rect 13700 19295 13758 19301
rect 12534 19261 12547 19292
rect 12488 19255 12547 19261
rect 13700 19261 13712 19295
rect 13746 19292 13758 19295
rect 13998 19292 14004 19304
rect 13746 19264 14004 19292
rect 13746 19261 13758 19264
rect 13700 19255 13758 19261
rect 8389 19227 8447 19233
rect 8389 19193 8401 19227
rect 8435 19224 8447 19227
rect 8843 19227 8901 19233
rect 8843 19224 8855 19227
rect 8435 19196 8855 19224
rect 8435 19193 8447 19196
rect 8389 19187 8447 19193
rect 8843 19193 8855 19196
rect 8889 19224 8901 19227
rect 9674 19224 9680 19236
rect 8889 19196 9680 19224
rect 8889 19193 8901 19196
rect 8843 19187 8901 19193
rect 9674 19184 9680 19196
rect 9732 19184 9738 19236
rect 12519 19156 12547 19255
rect 13998 19252 14004 19264
rect 14056 19292 14062 19304
rect 14093 19295 14151 19301
rect 14093 19292 14105 19295
rect 14056 19264 14105 19292
rect 14056 19252 14062 19264
rect 14093 19261 14105 19264
rect 14139 19261 14151 19295
rect 14093 19255 14151 19261
rect 15289 19295 15347 19301
rect 15289 19261 15301 19295
rect 15335 19292 15347 19295
rect 15416 19295 15474 19301
rect 15416 19292 15428 19295
rect 15335 19264 15428 19292
rect 15335 19261 15347 19264
rect 15289 19255 15347 19261
rect 15416 19261 15428 19264
rect 15462 19292 15474 19295
rect 15654 19292 15660 19304
rect 15462 19264 15660 19292
rect 15462 19261 15474 19264
rect 15416 19255 15474 19261
rect 15654 19252 15660 19264
rect 15712 19252 15718 19304
rect 17129 19295 17187 19301
rect 17129 19261 17141 19295
rect 17175 19292 17187 19295
rect 17678 19292 17684 19304
rect 17175 19264 17684 19292
rect 17175 19261 17187 19264
rect 17129 19255 17187 19261
rect 17678 19252 17684 19264
rect 17736 19252 17742 19304
rect 12575 19227 12633 19233
rect 12575 19193 12587 19227
rect 12621 19224 12633 19227
rect 13538 19224 13544 19236
rect 12621 19196 13544 19224
rect 12621 19193 12633 19196
rect 12575 19187 12633 19193
rect 13538 19184 13544 19196
rect 13596 19184 13602 19236
rect 15519 19227 15577 19233
rect 15519 19193 15531 19227
rect 15565 19224 15577 19227
rect 16482 19224 16488 19236
rect 15565 19196 16488 19224
rect 15565 19193 15577 19196
rect 15519 19187 15577 19193
rect 16482 19184 16488 19196
rect 16540 19184 16546 19236
rect 16574 19184 16580 19236
rect 16632 19224 16638 19236
rect 17494 19224 17500 19236
rect 16632 19196 16677 19224
rect 17407 19196 17500 19224
rect 16632 19184 16638 19196
rect 17494 19184 17500 19196
rect 17552 19224 17558 19236
rect 20640 19233 20668 19332
rect 21136 19295 21194 19301
rect 21136 19261 21148 19295
rect 21182 19292 21194 19295
rect 21634 19292 21640 19304
rect 21182 19264 21640 19292
rect 21182 19261 21194 19264
rect 21136 19255 21194 19261
rect 21634 19252 21640 19264
rect 21692 19252 21698 19304
rect 19429 19227 19487 19233
rect 19429 19224 19441 19227
rect 17552 19196 19441 19224
rect 17552 19184 17558 19196
rect 19429 19193 19441 19196
rect 19475 19224 19487 19227
rect 19705 19227 19763 19233
rect 19705 19224 19717 19227
rect 19475 19196 19717 19224
rect 19475 19193 19487 19196
rect 19429 19187 19487 19193
rect 19705 19193 19717 19196
rect 19751 19193 19763 19227
rect 19705 19187 19763 19193
rect 20625 19227 20683 19233
rect 20625 19193 20637 19227
rect 20671 19224 20683 19227
rect 21223 19227 21281 19233
rect 21223 19224 21235 19227
rect 20671 19196 21235 19224
rect 20671 19193 20683 19196
rect 20625 19187 20683 19193
rect 21223 19193 21235 19196
rect 21269 19193 21281 19227
rect 21223 19187 21281 19193
rect 12802 19156 12808 19168
rect 12519 19128 12808 19156
rect 12802 19116 12808 19128
rect 12860 19156 12866 19168
rect 12897 19159 12955 19165
rect 12897 19156 12909 19159
rect 12860 19128 12909 19156
rect 12860 19116 12866 19128
rect 12897 19125 12909 19128
rect 12943 19125 12955 19159
rect 12897 19119 12955 19125
rect 15838 19116 15844 19168
rect 15896 19156 15902 19168
rect 16025 19159 16083 19165
rect 16025 19156 16037 19159
rect 15896 19128 16037 19156
rect 15896 19116 15902 19128
rect 16025 19125 16037 19128
rect 16071 19156 16083 19159
rect 18230 19156 18236 19168
rect 16071 19128 18236 19156
rect 16071 19125 16083 19128
rect 16025 19119 16083 19125
rect 18230 19116 18236 19128
rect 18288 19116 18294 19168
rect 18509 19159 18567 19165
rect 18509 19125 18521 19159
rect 18555 19156 18567 19159
rect 18782 19156 18788 19168
rect 18555 19128 18788 19156
rect 18555 19125 18567 19128
rect 18509 19119 18567 19125
rect 18782 19116 18788 19128
rect 18840 19116 18846 19168
rect 18874 19116 18880 19168
rect 18932 19156 18938 19168
rect 18969 19159 19027 19165
rect 18969 19156 18981 19159
rect 18932 19128 18981 19156
rect 18932 19116 18938 19128
rect 18969 19125 18981 19128
rect 19015 19125 19027 19159
rect 18969 19119 19027 19125
rect 1104 19066 22816 19088
rect 1104 19014 8982 19066
rect 9034 19014 9046 19066
rect 9098 19014 9110 19066
rect 9162 19014 9174 19066
rect 9226 19014 16982 19066
rect 17034 19014 17046 19066
rect 17098 19014 17110 19066
rect 17162 19014 17174 19066
rect 17226 19014 22816 19066
rect 1104 18992 22816 19014
rect 10686 18952 10692 18964
rect 10647 18924 10692 18952
rect 10686 18912 10692 18924
rect 10744 18912 10750 18964
rect 13538 18952 13544 18964
rect 13499 18924 13544 18952
rect 13538 18912 13544 18924
rect 13596 18912 13602 18964
rect 14323 18955 14381 18961
rect 14323 18921 14335 18955
rect 14369 18952 14381 18955
rect 16206 18952 16212 18964
rect 14369 18924 16212 18952
rect 14369 18921 14381 18924
rect 14323 18915 14381 18921
rect 16206 18912 16212 18924
rect 16264 18912 16270 18964
rect 16482 18952 16488 18964
rect 16443 18924 16488 18952
rect 16482 18912 16488 18924
rect 16540 18912 16546 18964
rect 9674 18844 9680 18896
rect 9732 18884 9738 18896
rect 10090 18887 10148 18893
rect 10090 18884 10102 18887
rect 9732 18856 10102 18884
rect 9732 18844 9738 18856
rect 10090 18853 10102 18856
rect 10136 18853 10148 18887
rect 10090 18847 10148 18853
rect 11606 18844 11612 18896
rect 11664 18884 11670 18896
rect 11701 18887 11759 18893
rect 11701 18884 11713 18887
rect 11664 18856 11713 18884
rect 11664 18844 11670 18856
rect 11701 18853 11713 18856
rect 11747 18853 11759 18887
rect 12250 18884 12256 18896
rect 12211 18856 12256 18884
rect 11701 18847 11759 18853
rect 12250 18844 12256 18856
rect 12308 18844 12314 18896
rect 15470 18844 15476 18896
rect 15528 18884 15534 18896
rect 15610 18887 15668 18893
rect 15610 18884 15622 18887
rect 15528 18856 15622 18884
rect 15528 18844 15534 18856
rect 15610 18853 15622 18856
rect 15656 18853 15668 18887
rect 15610 18847 15668 18853
rect 16298 18844 16304 18896
rect 16356 18884 16362 18896
rect 17126 18884 17132 18896
rect 16356 18856 17132 18884
rect 16356 18844 16362 18856
rect 17126 18844 17132 18856
rect 17184 18844 17190 18896
rect 17221 18887 17279 18893
rect 17221 18853 17233 18887
rect 17267 18884 17279 18887
rect 17494 18884 17500 18896
rect 17267 18856 17500 18884
rect 17267 18853 17279 18856
rect 17221 18847 17279 18853
rect 17494 18844 17500 18856
rect 17552 18844 17558 18896
rect 18874 18884 18880 18896
rect 18835 18856 18880 18884
rect 18874 18844 18880 18856
rect 18932 18844 18938 18896
rect 1302 18776 1308 18828
rect 1360 18816 1366 18828
rect 1432 18819 1490 18825
rect 1432 18816 1444 18819
rect 1360 18788 1444 18816
rect 1360 18776 1366 18788
rect 1432 18785 1444 18788
rect 1478 18785 1490 18819
rect 1432 18779 1490 18785
rect 12710 18776 12716 18828
rect 12768 18816 12774 18828
rect 13116 18819 13174 18825
rect 13116 18816 13128 18819
rect 12768 18788 13128 18816
rect 12768 18776 12774 18788
rect 13116 18785 13128 18788
rect 13162 18785 13174 18819
rect 13116 18779 13174 18785
rect 14090 18776 14096 18828
rect 14148 18816 14154 18828
rect 14220 18819 14278 18825
rect 14220 18816 14232 18819
rect 14148 18788 14232 18816
rect 14148 18776 14154 18788
rect 14220 18785 14232 18788
rect 14266 18785 14278 18819
rect 14220 18779 14278 18785
rect 9766 18748 9772 18760
rect 9727 18720 9772 18748
rect 9766 18708 9772 18720
rect 9824 18708 9830 18760
rect 11238 18708 11244 18760
rect 11296 18748 11302 18760
rect 11609 18751 11667 18757
rect 11609 18748 11621 18751
rect 11296 18720 11621 18748
rect 11296 18708 11302 18720
rect 11609 18717 11621 18720
rect 11655 18748 11667 18751
rect 13219 18751 13277 18757
rect 13219 18748 13231 18751
rect 11655 18720 13231 18748
rect 11655 18717 11667 18720
rect 11609 18711 11667 18717
rect 13219 18717 13231 18720
rect 13265 18717 13277 18751
rect 13219 18711 13277 18717
rect 15289 18751 15347 18757
rect 15289 18717 15301 18751
rect 15335 18748 15347 18751
rect 15838 18748 15844 18760
rect 15335 18720 15844 18748
rect 15335 18717 15347 18720
rect 15289 18711 15347 18717
rect 15838 18708 15844 18720
rect 15896 18708 15902 18760
rect 18782 18748 18788 18760
rect 18743 18720 18788 18748
rect 18782 18708 18788 18720
rect 18840 18708 18846 18760
rect 19058 18748 19064 18760
rect 19019 18720 19064 18748
rect 19058 18708 19064 18720
rect 19116 18708 19122 18760
rect 16209 18683 16267 18689
rect 16209 18649 16221 18683
rect 16255 18680 16267 18683
rect 17494 18680 17500 18692
rect 16255 18652 17500 18680
rect 16255 18649 16267 18652
rect 16209 18643 16267 18649
rect 17494 18640 17500 18652
rect 17552 18640 17558 18692
rect 17678 18680 17684 18692
rect 17639 18652 17684 18680
rect 17678 18640 17684 18652
rect 17736 18640 17742 18692
rect 1535 18615 1593 18621
rect 1535 18581 1547 18615
rect 1581 18612 1593 18615
rect 7650 18612 7656 18624
rect 1581 18584 7656 18612
rect 1581 18581 1593 18584
rect 1535 18575 1593 18581
rect 7650 18572 7656 18584
rect 7708 18572 7714 18624
rect 8570 18612 8576 18624
rect 8531 18584 8576 18612
rect 8570 18572 8576 18584
rect 8628 18572 8634 18624
rect 19702 18612 19708 18624
rect 19663 18584 19708 18612
rect 19702 18572 19708 18584
rect 19760 18572 19766 18624
rect 1104 18522 22816 18544
rect 1104 18470 4982 18522
rect 5034 18470 5046 18522
rect 5098 18470 5110 18522
rect 5162 18470 5174 18522
rect 5226 18470 12982 18522
rect 13034 18470 13046 18522
rect 13098 18470 13110 18522
rect 13162 18470 13174 18522
rect 13226 18470 20982 18522
rect 21034 18470 21046 18522
rect 21098 18470 21110 18522
rect 21162 18470 21174 18522
rect 21226 18470 22816 18522
rect 1104 18448 22816 18470
rect 1302 18368 1308 18420
rect 1360 18408 1366 18420
rect 1857 18411 1915 18417
rect 1857 18408 1869 18411
rect 1360 18380 1869 18408
rect 1360 18368 1366 18380
rect 1857 18377 1869 18380
rect 1903 18377 1915 18411
rect 7650 18408 7656 18420
rect 7611 18380 7656 18408
rect 1857 18371 1915 18377
rect 7650 18368 7656 18380
rect 7708 18368 7714 18420
rect 9306 18408 9312 18420
rect 9219 18380 9312 18408
rect 9306 18368 9312 18380
rect 9364 18408 9370 18420
rect 9766 18408 9772 18420
rect 9364 18380 9772 18408
rect 9364 18368 9370 18380
rect 9766 18368 9772 18380
rect 9824 18368 9830 18420
rect 11238 18408 11244 18420
rect 11199 18380 11244 18408
rect 11238 18368 11244 18380
rect 11296 18368 11302 18420
rect 11606 18368 11612 18420
rect 11664 18408 11670 18420
rect 12161 18411 12219 18417
rect 12161 18408 12173 18411
rect 11664 18380 12173 18408
rect 11664 18368 11670 18380
rect 12161 18377 12173 18380
rect 12207 18377 12219 18411
rect 12161 18371 12219 18377
rect 15197 18411 15255 18417
rect 15197 18377 15209 18411
rect 15243 18408 15255 18411
rect 16574 18408 16580 18420
rect 15243 18380 16580 18408
rect 15243 18377 15255 18380
rect 15197 18371 15255 18377
rect 16574 18368 16580 18380
rect 16632 18368 16638 18420
rect 17126 18368 17132 18420
rect 17184 18408 17190 18420
rect 17681 18411 17739 18417
rect 17681 18408 17693 18411
rect 17184 18380 17693 18408
rect 17184 18368 17190 18380
rect 17681 18377 17693 18380
rect 17727 18377 17739 18411
rect 17681 18371 17739 18377
rect 18782 18368 18788 18420
rect 18840 18408 18846 18420
rect 19245 18411 19303 18417
rect 19245 18408 19257 18411
rect 18840 18380 19257 18408
rect 18840 18368 18846 18380
rect 19245 18377 19257 18380
rect 19291 18377 19303 18411
rect 19245 18371 19303 18377
rect 21177 18411 21235 18417
rect 21177 18377 21189 18411
rect 21223 18408 21235 18411
rect 21266 18408 21272 18420
rect 21223 18380 21272 18408
rect 21223 18377 21235 18380
rect 21177 18371 21235 18377
rect 21266 18368 21272 18380
rect 21324 18368 21330 18420
rect 2866 18232 2872 18284
rect 2924 18272 2930 18284
rect 7668 18272 7696 18368
rect 8113 18343 8171 18349
rect 8113 18309 8125 18343
rect 8159 18340 8171 18343
rect 8386 18340 8392 18352
rect 8159 18312 8392 18340
rect 8159 18309 8171 18312
rect 8113 18303 8171 18309
rect 8386 18300 8392 18312
rect 8444 18300 8450 18352
rect 10318 18300 10324 18352
rect 10376 18340 10382 18352
rect 11974 18340 11980 18352
rect 10376 18312 11980 18340
rect 10376 18300 10382 18312
rect 11974 18300 11980 18312
rect 12032 18340 12038 18352
rect 13081 18343 13139 18349
rect 13081 18340 13093 18343
rect 12032 18312 13093 18340
rect 12032 18300 12038 18312
rect 13081 18309 13093 18312
rect 13127 18309 13139 18343
rect 16390 18340 16396 18352
rect 13081 18303 13139 18309
rect 13924 18312 16396 18340
rect 8297 18275 8355 18281
rect 8297 18272 8309 18275
rect 2924 18244 4154 18272
rect 7668 18244 8309 18272
rect 2924 18232 2930 18244
rect 1464 18207 1522 18213
rect 1464 18173 1476 18207
rect 1510 18204 1522 18207
rect 2222 18204 2228 18216
rect 1510 18176 2228 18204
rect 1510 18173 1522 18176
rect 1464 18167 1522 18173
rect 2222 18164 2228 18176
rect 2280 18164 2286 18216
rect 4126 18136 4154 18244
rect 8297 18241 8309 18244
rect 8343 18241 8355 18275
rect 8297 18235 8355 18241
rect 8941 18275 8999 18281
rect 8941 18241 8953 18275
rect 8987 18272 8999 18275
rect 10137 18275 10195 18281
rect 10137 18272 10149 18275
rect 8987 18244 10149 18272
rect 8987 18241 8999 18244
rect 8941 18235 8999 18241
rect 10137 18241 10149 18244
rect 10183 18272 10195 18275
rect 11146 18272 11152 18284
rect 10183 18244 11152 18272
rect 10183 18241 10195 18244
rect 10137 18235 10195 18241
rect 11146 18232 11152 18244
rect 11204 18232 11210 18284
rect 13924 18272 13952 18312
rect 16390 18300 16396 18312
rect 16448 18300 16454 18352
rect 11900 18244 13952 18272
rect 14001 18275 14059 18281
rect 11400 18207 11458 18213
rect 11400 18173 11412 18207
rect 11446 18204 11458 18207
rect 11900 18204 11928 18244
rect 14001 18241 14013 18275
rect 14047 18272 14059 18275
rect 16592 18272 16620 18368
rect 17405 18343 17463 18349
rect 17405 18309 17417 18343
rect 17451 18340 17463 18343
rect 17494 18340 17500 18352
rect 17451 18312 17500 18340
rect 17451 18309 17463 18312
rect 17405 18303 17463 18309
rect 17494 18300 17500 18312
rect 17552 18300 17558 18352
rect 18233 18275 18291 18281
rect 18233 18272 18245 18275
rect 14047 18244 14641 18272
rect 16592 18244 18245 18272
rect 14047 18241 14059 18244
rect 14001 18235 14059 18241
rect 11446 18176 11928 18204
rect 11446 18173 11458 18176
rect 11400 18167 11458 18173
rect 4126 18108 8340 18136
rect 1535 18071 1593 18077
rect 1535 18037 1547 18071
rect 1581 18068 1593 18071
rect 1762 18068 1768 18080
rect 1581 18040 1768 18068
rect 1581 18037 1593 18040
rect 1535 18031 1593 18037
rect 1762 18028 1768 18040
rect 1820 18028 1826 18080
rect 8312 18068 8340 18108
rect 8386 18096 8392 18148
rect 8444 18136 8450 18148
rect 8754 18136 8760 18148
rect 8444 18108 8760 18136
rect 8444 18096 8450 18108
rect 8754 18096 8760 18108
rect 8812 18096 8818 18148
rect 9861 18139 9919 18145
rect 9861 18136 9873 18139
rect 9048 18108 9873 18136
rect 9048 18068 9076 18108
rect 9861 18105 9873 18108
rect 9907 18105 9919 18139
rect 9861 18099 9919 18105
rect 9674 18068 9680 18080
rect 8312 18040 9076 18068
rect 9635 18040 9680 18068
rect 9674 18028 9680 18040
rect 9732 18028 9738 18080
rect 9876 18068 9904 18099
rect 9950 18096 9956 18148
rect 10008 18136 10014 18148
rect 10008 18108 10053 18136
rect 10008 18096 10014 18108
rect 10781 18071 10839 18077
rect 10781 18068 10793 18071
rect 9876 18040 10793 18068
rect 10781 18037 10793 18040
rect 10827 18037 10839 18071
rect 10781 18031 10839 18037
rect 11238 18028 11244 18080
rect 11296 18068 11302 18080
rect 11900 18077 11928 18176
rect 12504 18207 12562 18213
rect 12504 18173 12516 18207
rect 12550 18204 12562 18207
rect 12802 18204 12808 18216
rect 12550 18176 12808 18204
rect 12550 18173 12562 18176
rect 12504 18167 12562 18173
rect 12802 18164 12808 18176
rect 12860 18204 12866 18216
rect 13081 18207 13139 18213
rect 12860 18176 13032 18204
rect 12860 18164 12866 18176
rect 13004 18145 13032 18176
rect 13081 18173 13093 18207
rect 13127 18204 13139 18207
rect 13127 18176 13814 18204
rect 13127 18173 13139 18176
rect 13081 18167 13139 18173
rect 12989 18139 13047 18145
rect 12989 18105 13001 18139
rect 13035 18136 13047 18139
rect 13446 18136 13452 18148
rect 13035 18108 13452 18136
rect 13035 18105 13047 18108
rect 12989 18099 13047 18105
rect 13446 18096 13452 18108
rect 13504 18096 13510 18148
rect 13786 18136 13814 18176
rect 14182 18164 14188 18216
rect 14240 18204 14246 18216
rect 14277 18207 14335 18213
rect 14277 18204 14289 18207
rect 14240 18176 14289 18204
rect 14240 18164 14246 18176
rect 14277 18173 14289 18176
rect 14323 18173 14335 18207
rect 14277 18167 14335 18173
rect 14090 18136 14096 18148
rect 13786 18108 14096 18136
rect 14090 18096 14096 18108
rect 14148 18136 14154 18148
rect 14613 18145 14641 18244
rect 18233 18241 18245 18244
rect 18279 18272 18291 18275
rect 18874 18272 18880 18284
rect 18279 18244 18880 18272
rect 18279 18241 18291 18244
rect 18233 18235 18291 18241
rect 18874 18232 18880 18244
rect 18932 18232 18938 18284
rect 19518 18272 19524 18284
rect 19479 18244 19524 18272
rect 19518 18232 19524 18244
rect 19576 18232 19582 18284
rect 19978 18272 19984 18284
rect 19939 18244 19984 18272
rect 19978 18232 19984 18244
rect 20036 18232 20042 18284
rect 15562 18164 15568 18216
rect 15620 18204 15626 18216
rect 16520 18207 16578 18213
rect 16520 18204 16532 18207
rect 15620 18176 16532 18204
rect 15620 18164 15626 18176
rect 16520 18173 16532 18176
rect 16566 18204 16578 18207
rect 16945 18207 17003 18213
rect 16945 18204 16957 18207
rect 16566 18176 16957 18204
rect 16566 18173 16578 18176
rect 16520 18167 16578 18173
rect 16945 18173 16957 18176
rect 16991 18173 17003 18207
rect 16945 18167 17003 18173
rect 18484 18207 18542 18213
rect 18484 18173 18496 18207
rect 18530 18204 18542 18207
rect 20993 18207 21051 18213
rect 18530 18176 19012 18204
rect 18530 18173 18542 18176
rect 18484 18167 18542 18173
rect 14598 18139 14656 18145
rect 14148 18108 14228 18136
rect 14148 18096 14154 18108
rect 11471 18071 11529 18077
rect 11471 18068 11483 18071
rect 11296 18040 11483 18068
rect 11296 18028 11302 18040
rect 11471 18037 11483 18040
rect 11517 18037 11529 18071
rect 11471 18031 11529 18037
rect 11885 18071 11943 18077
rect 11885 18037 11897 18071
rect 11931 18068 11943 18071
rect 11974 18068 11980 18080
rect 11931 18040 11980 18068
rect 11931 18037 11943 18040
rect 11885 18031 11943 18037
rect 11974 18028 11980 18040
rect 12032 18028 12038 18080
rect 12250 18028 12256 18080
rect 12308 18068 12314 18080
rect 12575 18071 12633 18077
rect 12575 18068 12587 18071
rect 12308 18040 12587 18068
rect 12308 18028 12314 18040
rect 12575 18037 12587 18040
rect 12621 18037 12633 18071
rect 12575 18031 12633 18037
rect 12710 18028 12716 18080
rect 12768 18068 12774 18080
rect 13265 18071 13323 18077
rect 13265 18068 13277 18071
rect 12768 18040 13277 18068
rect 12768 18028 12774 18040
rect 13265 18037 13277 18040
rect 13311 18037 13323 18071
rect 13722 18068 13728 18080
rect 13635 18040 13728 18068
rect 13265 18031 13323 18037
rect 13722 18028 13728 18040
rect 13780 18068 13786 18080
rect 14200 18077 14228 18108
rect 14598 18105 14610 18139
rect 14644 18136 14656 18139
rect 14826 18136 14832 18148
rect 14644 18108 14832 18136
rect 14644 18105 14656 18108
rect 14598 18099 14656 18105
rect 14826 18096 14832 18108
rect 14884 18136 14890 18148
rect 15470 18136 15476 18148
rect 14884 18108 15476 18136
rect 14884 18096 14890 18108
rect 15470 18096 15476 18108
rect 15528 18096 15534 18148
rect 14001 18071 14059 18077
rect 14001 18068 14013 18071
rect 13780 18040 14013 18068
rect 13780 18028 13786 18040
rect 14001 18037 14013 18040
rect 14047 18037 14059 18071
rect 14001 18031 14059 18037
rect 14185 18071 14243 18077
rect 14185 18037 14197 18071
rect 14231 18068 14243 18071
rect 15102 18068 15108 18080
rect 14231 18040 15108 18068
rect 14231 18037 14243 18040
rect 14185 18031 14243 18037
rect 15102 18028 15108 18040
rect 15160 18028 15166 18080
rect 15838 18068 15844 18080
rect 15799 18040 15844 18068
rect 15838 18028 15844 18040
rect 15896 18028 15902 18080
rect 16623 18071 16681 18077
rect 16623 18037 16635 18071
rect 16669 18068 16681 18071
rect 16850 18068 16856 18080
rect 16669 18040 16856 18068
rect 16669 18037 16681 18040
rect 16623 18031 16681 18037
rect 16850 18028 16856 18040
rect 16908 18028 16914 18080
rect 18555 18071 18613 18077
rect 18555 18037 18567 18071
rect 18601 18068 18613 18071
rect 18782 18068 18788 18080
rect 18601 18040 18788 18068
rect 18601 18037 18613 18040
rect 18555 18031 18613 18037
rect 18782 18028 18788 18040
rect 18840 18028 18846 18080
rect 18984 18077 19012 18176
rect 20993 18173 21005 18207
rect 21039 18173 21051 18207
rect 20993 18167 21051 18173
rect 19613 18139 19671 18145
rect 19613 18105 19625 18139
rect 19659 18136 19671 18139
rect 19702 18136 19708 18148
rect 19659 18108 19708 18136
rect 19659 18105 19671 18108
rect 19613 18099 19671 18105
rect 19702 18096 19708 18108
rect 19760 18096 19766 18148
rect 18969 18071 19027 18077
rect 18969 18037 18981 18071
rect 19015 18068 19027 18071
rect 19150 18068 19156 18080
rect 19015 18040 19156 18068
rect 19015 18037 19027 18040
rect 18969 18031 19027 18037
rect 19150 18028 19156 18040
rect 19208 18068 19214 18080
rect 21008 18068 21036 18167
rect 21545 18071 21603 18077
rect 21545 18068 21557 18071
rect 19208 18040 21557 18068
rect 19208 18028 19214 18040
rect 21545 18037 21557 18040
rect 21591 18037 21603 18071
rect 21545 18031 21603 18037
rect 1104 17978 22816 18000
rect 1104 17926 8982 17978
rect 9034 17926 9046 17978
rect 9098 17926 9110 17978
rect 9162 17926 9174 17978
rect 9226 17926 16982 17978
rect 17034 17926 17046 17978
rect 17098 17926 17110 17978
rect 17162 17926 17174 17978
rect 17226 17926 22816 17978
rect 1104 17904 22816 17926
rect 1762 17824 1768 17876
rect 1820 17864 1826 17876
rect 2225 17867 2283 17873
rect 2225 17864 2237 17867
rect 1820 17836 2237 17864
rect 1820 17824 1826 17836
rect 2225 17833 2237 17836
rect 2271 17864 2283 17867
rect 2314 17864 2320 17876
rect 2271 17836 2320 17864
rect 2271 17833 2283 17836
rect 2225 17827 2283 17833
rect 2314 17824 2320 17836
rect 2372 17824 2378 17876
rect 9674 17824 9680 17876
rect 9732 17864 9738 17876
rect 10226 17864 10232 17876
rect 9732 17836 10232 17864
rect 9732 17824 9738 17836
rect 10226 17824 10232 17836
rect 10284 17864 10290 17876
rect 13722 17864 13728 17876
rect 10284 17836 13728 17864
rect 10284 17824 10290 17836
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 16960 17836 19104 17864
rect 16960 17808 16988 17836
rect 9950 17796 9956 17808
rect 9863 17768 9956 17796
rect 9950 17756 9956 17768
rect 10008 17796 10014 17808
rect 11698 17796 11704 17808
rect 10008 17768 11704 17796
rect 10008 17756 10014 17768
rect 11698 17756 11704 17768
rect 11756 17756 11762 17808
rect 14369 17799 14427 17805
rect 14369 17765 14381 17799
rect 14415 17796 14427 17799
rect 15838 17796 15844 17808
rect 14415 17768 15844 17796
rect 14415 17765 14427 17768
rect 14369 17759 14427 17765
rect 15838 17756 15844 17768
rect 15896 17756 15902 17808
rect 16850 17796 16856 17808
rect 16811 17768 16856 17796
rect 16850 17756 16856 17768
rect 16908 17756 16914 17808
rect 16942 17756 16948 17808
rect 17000 17796 17006 17808
rect 17000 17768 17093 17796
rect 17000 17756 17006 17768
rect 18782 17756 18788 17808
rect 18840 17796 18846 17808
rect 19076 17805 19104 17836
rect 19518 17824 19524 17876
rect 19576 17864 19582 17876
rect 19889 17867 19947 17873
rect 19889 17864 19901 17867
rect 19576 17836 19901 17864
rect 19576 17824 19582 17836
rect 19889 17833 19901 17836
rect 19935 17833 19947 17867
rect 19889 17827 19947 17833
rect 21085 17867 21143 17873
rect 21085 17833 21097 17867
rect 21131 17864 21143 17867
rect 21726 17864 21732 17876
rect 21131 17836 21732 17864
rect 21131 17833 21143 17836
rect 21085 17827 21143 17833
rect 21726 17824 21732 17836
rect 21784 17824 21790 17876
rect 18969 17799 19027 17805
rect 18969 17796 18981 17799
rect 18840 17768 18981 17796
rect 18840 17756 18846 17768
rect 18969 17765 18981 17768
rect 19015 17765 19027 17799
rect 18969 17759 19027 17765
rect 19061 17799 19119 17805
rect 19061 17765 19073 17799
rect 19107 17796 19119 17799
rect 19242 17796 19248 17808
rect 19107 17768 19248 17796
rect 19107 17765 19119 17768
rect 19061 17759 19119 17765
rect 19242 17756 19248 17768
rect 19300 17796 19306 17808
rect 19702 17796 19708 17808
rect 19300 17768 19708 17796
rect 19300 17756 19306 17768
rect 19702 17756 19708 17768
rect 19760 17756 19766 17808
rect 4798 17688 4804 17740
rect 4856 17728 4862 17740
rect 4893 17731 4951 17737
rect 4893 17728 4905 17731
rect 4856 17700 4905 17728
rect 4856 17688 4862 17700
rect 4893 17697 4905 17700
rect 4939 17697 4951 17731
rect 4893 17691 4951 17697
rect 5353 17731 5411 17737
rect 5353 17697 5365 17731
rect 5399 17728 5411 17731
rect 5534 17728 5540 17740
rect 5399 17700 5540 17728
rect 5399 17697 5411 17700
rect 5353 17691 5411 17697
rect 5534 17688 5540 17700
rect 5592 17688 5598 17740
rect 6457 17731 6515 17737
rect 6457 17697 6469 17731
rect 6503 17728 6515 17731
rect 6638 17728 6644 17740
rect 6503 17700 6644 17728
rect 6503 17697 6515 17700
rect 6457 17691 6515 17697
rect 6638 17688 6644 17700
rect 6696 17688 6702 17740
rect 10318 17728 10324 17740
rect 10279 17700 10324 17728
rect 10318 17688 10324 17700
rect 10376 17688 10382 17740
rect 13354 17688 13360 17740
rect 13412 17728 13418 17740
rect 13633 17731 13691 17737
rect 13633 17728 13645 17731
rect 13412 17700 13645 17728
rect 13412 17688 13418 17700
rect 13633 17697 13645 17700
rect 13679 17697 13691 17731
rect 13633 17691 13691 17697
rect 14093 17731 14151 17737
rect 14093 17697 14105 17731
rect 14139 17697 14151 17731
rect 14093 17691 14151 17697
rect 5442 17660 5448 17672
rect 5403 17632 5448 17660
rect 5442 17620 5448 17632
rect 5500 17620 5506 17672
rect 8573 17663 8631 17669
rect 8573 17629 8585 17663
rect 8619 17660 8631 17663
rect 10778 17660 10784 17672
rect 8619 17632 10784 17660
rect 8619 17629 8631 17632
rect 8573 17623 8631 17629
rect 10778 17620 10784 17632
rect 10836 17660 10842 17672
rect 10873 17663 10931 17669
rect 10873 17660 10885 17663
rect 10836 17632 10885 17660
rect 10836 17620 10842 17632
rect 10873 17629 10885 17632
rect 10919 17629 10931 17663
rect 10873 17623 10931 17629
rect 11609 17663 11667 17669
rect 11609 17629 11621 17663
rect 11655 17629 11667 17663
rect 11882 17660 11888 17672
rect 11843 17632 11888 17660
rect 11609 17623 11667 17629
rect 106 17552 112 17604
rect 164 17592 170 17604
rect 10505 17595 10563 17601
rect 10505 17592 10517 17595
rect 164 17564 10517 17592
rect 164 17552 170 17564
rect 10505 17561 10517 17564
rect 10551 17561 10563 17595
rect 11624 17592 11652 17623
rect 11882 17620 11888 17632
rect 11940 17620 11946 17672
rect 12250 17592 12256 17604
rect 11624 17564 12256 17592
rect 10505 17555 10563 17561
rect 12250 17552 12256 17564
rect 12308 17552 12314 17604
rect 6687 17527 6745 17533
rect 6687 17493 6699 17527
rect 6733 17524 6745 17527
rect 6914 17524 6920 17536
rect 6733 17496 6920 17524
rect 6733 17493 6745 17496
rect 6687 17487 6745 17493
rect 6914 17484 6920 17496
rect 6972 17484 6978 17536
rect 8478 17524 8484 17536
rect 8439 17496 8484 17524
rect 8478 17484 8484 17496
rect 8536 17484 8542 17536
rect 12158 17484 12164 17536
rect 12216 17524 12222 17536
rect 12529 17527 12587 17533
rect 12529 17524 12541 17527
rect 12216 17496 12541 17524
rect 12216 17484 12222 17496
rect 12529 17493 12541 17496
rect 12575 17493 12587 17527
rect 12529 17487 12587 17493
rect 13541 17527 13599 17533
rect 13541 17493 13553 17527
rect 13587 17524 13599 17527
rect 13906 17524 13912 17536
rect 13587 17496 13912 17524
rect 13587 17493 13599 17496
rect 13541 17487 13599 17493
rect 13906 17484 13912 17496
rect 13964 17524 13970 17536
rect 14108 17524 14136 17691
rect 15194 17688 15200 17740
rect 15252 17728 15258 17740
rect 15324 17731 15382 17737
rect 15324 17728 15336 17731
rect 15252 17700 15336 17728
rect 15252 17688 15258 17700
rect 15324 17697 15336 17700
rect 15370 17697 15382 17731
rect 15324 17691 15382 17697
rect 19794 17688 19800 17740
rect 19852 17728 19858 17740
rect 20901 17731 20959 17737
rect 20901 17728 20913 17731
rect 19852 17700 20913 17728
rect 19852 17688 19858 17700
rect 20901 17697 20913 17700
rect 20947 17728 20959 17731
rect 21726 17728 21732 17740
rect 20947 17700 21732 17728
rect 20947 17697 20959 17700
rect 20901 17691 20959 17697
rect 21726 17688 21732 17700
rect 21784 17688 21790 17740
rect 18322 17660 18328 17672
rect 18235 17632 18328 17660
rect 18322 17620 18328 17632
rect 18380 17660 18386 17672
rect 19058 17660 19064 17672
rect 18380 17632 19064 17660
rect 18380 17620 18386 17632
rect 19058 17620 19064 17632
rect 19116 17660 19122 17672
rect 19245 17663 19303 17669
rect 19245 17660 19257 17663
rect 19116 17632 19257 17660
rect 19116 17620 19122 17632
rect 19245 17629 19257 17632
rect 19291 17629 19303 17663
rect 19245 17623 19303 17629
rect 17405 17595 17463 17601
rect 17405 17561 17417 17595
rect 17451 17592 17463 17595
rect 17678 17592 17684 17604
rect 17451 17564 17684 17592
rect 17451 17561 17463 17564
rect 17405 17555 17463 17561
rect 17678 17552 17684 17564
rect 17736 17592 17742 17604
rect 18690 17592 18696 17604
rect 17736 17564 18696 17592
rect 17736 17552 17742 17564
rect 18690 17552 18696 17564
rect 18748 17552 18754 17604
rect 13964 17496 14136 17524
rect 13964 17484 13970 17496
rect 14182 17484 14188 17536
rect 14240 17524 14246 17536
rect 14645 17527 14703 17533
rect 14645 17524 14657 17527
rect 14240 17496 14657 17524
rect 14240 17484 14246 17496
rect 14645 17493 14657 17496
rect 14691 17493 14703 17527
rect 14645 17487 14703 17493
rect 14918 17484 14924 17536
rect 14976 17524 14982 17536
rect 15427 17527 15485 17533
rect 15427 17524 15439 17527
rect 14976 17496 15439 17524
rect 14976 17484 14982 17496
rect 15427 17493 15439 17496
rect 15473 17493 15485 17527
rect 15746 17524 15752 17536
rect 15707 17496 15752 17524
rect 15427 17487 15485 17493
rect 15746 17484 15752 17496
rect 15804 17484 15810 17536
rect 1104 17434 22816 17456
rect 1104 17382 4982 17434
rect 5034 17382 5046 17434
rect 5098 17382 5110 17434
rect 5162 17382 5174 17434
rect 5226 17382 12982 17434
rect 13034 17382 13046 17434
rect 13098 17382 13110 17434
rect 13162 17382 13174 17434
rect 13226 17382 20982 17434
rect 21034 17382 21046 17434
rect 21098 17382 21110 17434
rect 21162 17382 21174 17434
rect 21226 17382 22816 17434
rect 1104 17360 22816 17382
rect 4798 17320 4804 17332
rect 4126 17292 4804 17320
rect 3142 17212 3148 17264
rect 3200 17252 3206 17264
rect 4126 17252 4154 17292
rect 4798 17280 4804 17292
rect 4856 17320 4862 17332
rect 5077 17323 5135 17329
rect 5077 17320 5089 17323
rect 4856 17292 5089 17320
rect 4856 17280 4862 17292
rect 5077 17289 5089 17292
rect 5123 17289 5135 17323
rect 10318 17320 10324 17332
rect 10279 17292 10324 17320
rect 5077 17283 5135 17289
rect 10318 17280 10324 17292
rect 10376 17280 10382 17332
rect 12161 17323 12219 17329
rect 12161 17289 12173 17323
rect 12207 17320 12219 17323
rect 12250 17320 12256 17332
rect 12207 17292 12256 17320
rect 12207 17289 12219 17292
rect 12161 17283 12219 17289
rect 12250 17280 12256 17292
rect 12308 17280 12314 17332
rect 14826 17320 14832 17332
rect 14787 17292 14832 17320
rect 14826 17280 14832 17292
rect 14884 17280 14890 17332
rect 15194 17320 15200 17332
rect 15155 17292 15200 17320
rect 15194 17280 15200 17292
rect 15252 17280 15258 17332
rect 16850 17280 16856 17332
rect 16908 17320 16914 17332
rect 17129 17323 17187 17329
rect 17129 17320 17141 17323
rect 16908 17292 17141 17320
rect 16908 17280 16914 17292
rect 17129 17289 17141 17292
rect 17175 17289 17187 17323
rect 17129 17283 17187 17289
rect 18782 17280 18788 17332
rect 18840 17320 18846 17332
rect 19613 17323 19671 17329
rect 19613 17320 19625 17323
rect 18840 17292 19625 17320
rect 18840 17280 18846 17292
rect 19613 17289 19625 17292
rect 19659 17289 19671 17323
rect 21450 17320 21456 17332
rect 21411 17292 21456 17320
rect 19613 17283 19671 17289
rect 21450 17280 21456 17292
rect 21508 17280 21514 17332
rect 21726 17320 21732 17332
rect 21687 17292 21732 17320
rect 21726 17280 21732 17292
rect 21784 17280 21790 17332
rect 3200 17224 4154 17252
rect 3200 17212 3206 17224
rect 6178 17212 6184 17264
rect 6236 17252 6242 17264
rect 8205 17255 8263 17261
rect 8205 17252 8217 17255
rect 6236 17224 8217 17252
rect 6236 17212 6242 17224
rect 8205 17221 8217 17224
rect 8251 17252 8263 17255
rect 13262 17252 13268 17264
rect 8251 17224 13268 17252
rect 8251 17221 8263 17224
rect 8205 17215 8263 17221
rect 2314 17184 2320 17196
rect 2275 17156 2320 17184
rect 2314 17144 2320 17156
rect 2372 17144 2378 17196
rect 2498 17144 2504 17196
rect 2556 17184 2562 17196
rect 2593 17187 2651 17193
rect 2593 17184 2605 17187
rect 2556 17156 2605 17184
rect 2556 17144 2562 17156
rect 2593 17153 2605 17156
rect 2639 17153 2651 17187
rect 4614 17184 4620 17196
rect 4575 17156 4620 17184
rect 2593 17147 2651 17153
rect 4614 17144 4620 17156
rect 4672 17144 4678 17196
rect 6273 17187 6331 17193
rect 6273 17153 6285 17187
rect 6319 17184 6331 17187
rect 6917 17187 6975 17193
rect 6917 17184 6929 17187
rect 6319 17156 6929 17184
rect 6319 17153 6331 17156
rect 6273 17147 6331 17153
rect 6917 17153 6929 17156
rect 6963 17184 6975 17187
rect 7190 17184 7196 17196
rect 6963 17156 7196 17184
rect 6963 17153 6975 17156
rect 6917 17147 6975 17153
rect 7190 17144 7196 17156
rect 7248 17144 7254 17196
rect 8220 17116 8248 17215
rect 13262 17212 13268 17224
rect 13320 17252 13326 17264
rect 16209 17255 16267 17261
rect 13320 17224 13492 17252
rect 13320 17212 13326 17224
rect 10778 17184 10784 17196
rect 10739 17156 10784 17184
rect 10778 17144 10784 17156
rect 10836 17144 10842 17196
rect 11425 17187 11483 17193
rect 11425 17153 11437 17187
rect 11471 17184 11483 17187
rect 11882 17184 11888 17196
rect 11471 17156 11888 17184
rect 11471 17153 11483 17156
rect 11425 17147 11483 17153
rect 11882 17144 11888 17156
rect 11940 17144 11946 17196
rect 8389 17119 8447 17125
rect 8389 17116 8401 17119
rect 8220 17088 8401 17116
rect 8389 17085 8401 17088
rect 8435 17085 8447 17119
rect 8389 17079 8447 17085
rect 8478 17076 8484 17128
rect 8536 17116 8542 17128
rect 8849 17119 8907 17125
rect 8849 17116 8861 17119
rect 8536 17088 8861 17116
rect 8536 17076 8542 17088
rect 8849 17085 8861 17088
rect 8895 17085 8907 17119
rect 8849 17079 8907 17085
rect 12158 17076 12164 17128
rect 12216 17116 12222 17128
rect 13464 17125 13492 17224
rect 16209 17221 16221 17255
rect 16255 17252 16267 17255
rect 19242 17252 19248 17264
rect 16255 17224 16896 17252
rect 19203 17224 19248 17252
rect 16255 17221 16267 17224
rect 16209 17215 16267 17221
rect 14182 17184 14188 17196
rect 14143 17156 14188 17184
rect 14182 17144 14188 17156
rect 14240 17144 14246 17196
rect 15289 17187 15347 17193
rect 15289 17153 15301 17187
rect 15335 17184 15347 17187
rect 15746 17184 15752 17196
rect 15335 17156 15752 17184
rect 15335 17153 15347 17156
rect 15289 17147 15347 17153
rect 15746 17144 15752 17156
rect 15804 17144 15810 17196
rect 16868 17193 16896 17224
rect 19242 17212 19248 17224
rect 19300 17212 19306 17264
rect 16853 17187 16911 17193
rect 16853 17153 16865 17187
rect 16899 17184 16911 17187
rect 16942 17184 16948 17196
rect 16899 17156 16948 17184
rect 16899 17153 16911 17156
rect 16853 17147 16911 17153
rect 16942 17144 16948 17156
rect 17000 17144 17006 17196
rect 18322 17184 18328 17196
rect 18283 17156 18328 17184
rect 18322 17144 18328 17156
rect 18380 17144 18386 17196
rect 12472 17119 12530 17125
rect 12472 17116 12484 17119
rect 12216 17088 12484 17116
rect 12216 17076 12222 17088
rect 12472 17085 12484 17088
rect 12518 17085 12530 17119
rect 12472 17079 12530 17085
rect 13449 17119 13507 17125
rect 13449 17085 13461 17119
rect 13495 17085 13507 17119
rect 13906 17116 13912 17128
rect 13867 17088 13912 17116
rect 13449 17079 13507 17085
rect 13906 17076 13912 17088
rect 13964 17076 13970 17128
rect 20968 17119 21026 17125
rect 20968 17085 20980 17119
rect 21014 17116 21026 17119
rect 21450 17116 21456 17128
rect 21014 17088 21456 17116
rect 21014 17085 21026 17088
rect 20968 17079 21026 17085
rect 21450 17076 21456 17088
rect 21508 17076 21514 17128
rect 2409 17051 2467 17057
rect 2409 17017 2421 17051
rect 2455 17017 2467 17051
rect 2409 17011 2467 17017
rect 3605 17051 3663 17057
rect 3605 17017 3617 17051
rect 3651 17048 3663 17051
rect 3970 17048 3976 17060
rect 3651 17020 3976 17048
rect 3651 17017 3663 17020
rect 3605 17011 3663 17017
rect 2133 16983 2191 16989
rect 2133 16949 2145 16983
rect 2179 16980 2191 16983
rect 2424 16980 2452 17011
rect 3970 17008 3976 17020
rect 4028 17048 4034 17060
rect 4157 17051 4215 17057
rect 4157 17048 4169 17051
rect 4028 17020 4169 17048
rect 4028 17008 4034 17020
rect 4157 17017 4169 17020
rect 4203 17017 4215 17051
rect 4157 17011 4215 17017
rect 4249 17051 4307 17057
rect 4249 17017 4261 17051
rect 4295 17017 4307 17051
rect 4249 17011 4307 17017
rect 3694 16980 3700 16992
rect 2179 16952 3700 16980
rect 2179 16949 2191 16952
rect 2133 16943 2191 16949
rect 3694 16940 3700 16952
rect 3752 16980 3758 16992
rect 3881 16983 3939 16989
rect 3881 16980 3893 16983
rect 3752 16952 3893 16980
rect 3752 16940 3758 16952
rect 3881 16949 3893 16952
rect 3927 16980 3939 16983
rect 4264 16980 4292 17011
rect 7006 17008 7012 17060
rect 7064 17048 7070 17060
rect 7558 17048 7564 17060
rect 7064 17020 7109 17048
rect 7519 17020 7564 17048
rect 7064 17008 7070 17020
rect 7558 17008 7564 17020
rect 7616 17008 7622 17060
rect 10873 17051 10931 17057
rect 10873 17048 10885 17051
rect 9968 17020 10885 17048
rect 5534 16980 5540 16992
rect 3927 16952 4292 16980
rect 5495 16952 5540 16980
rect 3927 16949 3939 16952
rect 3881 16943 3939 16949
rect 5534 16940 5540 16952
rect 5592 16940 5598 16992
rect 6638 16980 6644 16992
rect 6599 16952 6644 16980
rect 6638 16940 6644 16952
rect 6696 16940 6702 16992
rect 8478 16980 8484 16992
rect 8439 16952 8484 16980
rect 8478 16940 8484 16952
rect 8536 16940 8542 16992
rect 8754 16940 8760 16992
rect 8812 16980 8818 16992
rect 9858 16980 9864 16992
rect 8812 16952 9864 16980
rect 8812 16940 8818 16952
rect 9858 16940 9864 16952
rect 9916 16980 9922 16992
rect 9968 16989 9996 17020
rect 10873 17017 10885 17020
rect 10919 17017 10931 17051
rect 10873 17011 10931 17017
rect 12989 17051 13047 17057
rect 12989 17017 13001 17051
rect 13035 17048 13047 17051
rect 13354 17048 13360 17060
rect 13035 17020 13360 17048
rect 13035 17017 13047 17020
rect 12989 17011 13047 17017
rect 13354 17008 13360 17020
rect 13412 17008 13418 17060
rect 14826 17008 14832 17060
rect 14884 17048 14890 17060
rect 15610 17051 15668 17057
rect 15610 17048 15622 17051
rect 14884 17020 15622 17048
rect 14884 17008 14890 17020
rect 15610 17017 15622 17020
rect 15656 17048 15668 17051
rect 16022 17048 16028 17060
rect 15656 17020 16028 17048
rect 15656 17017 15668 17020
rect 15610 17011 15668 17017
rect 16022 17008 16028 17020
rect 16080 17008 16086 17060
rect 18417 17051 18475 17057
rect 18417 17017 18429 17051
rect 18463 17017 18475 17051
rect 18417 17011 18475 17017
rect 18969 17051 19027 17057
rect 18969 17017 18981 17051
rect 19015 17048 19027 17051
rect 19058 17048 19064 17060
rect 19015 17020 19064 17048
rect 19015 17017 19027 17020
rect 18969 17011 19027 17017
rect 9953 16983 10011 16989
rect 9953 16980 9965 16983
rect 9916 16952 9965 16980
rect 9916 16940 9922 16952
rect 9953 16949 9965 16952
rect 9999 16949 10011 16983
rect 11698 16980 11704 16992
rect 11659 16952 11704 16980
rect 9953 16943 10011 16949
rect 11698 16940 11704 16952
rect 11756 16940 11762 16992
rect 12575 16983 12633 16989
rect 12575 16949 12587 16983
rect 12621 16980 12633 16983
rect 12802 16980 12808 16992
rect 12621 16952 12808 16980
rect 12621 16949 12633 16952
rect 12575 16943 12633 16949
rect 12802 16940 12808 16952
rect 12860 16940 12866 16992
rect 17862 16980 17868 16992
rect 17823 16952 17868 16980
rect 17862 16940 17868 16952
rect 17920 16980 17926 16992
rect 18432 16980 18460 17011
rect 19058 17008 19064 17020
rect 19116 17008 19122 17060
rect 17920 16952 18460 16980
rect 17920 16940 17926 16952
rect 19334 16940 19340 16992
rect 19392 16980 19398 16992
rect 21039 16983 21097 16989
rect 21039 16980 21051 16983
rect 19392 16952 21051 16980
rect 19392 16940 19398 16952
rect 21039 16949 21051 16952
rect 21085 16949 21097 16983
rect 21039 16943 21097 16949
rect 1104 16890 22816 16912
rect 1104 16838 8982 16890
rect 9034 16838 9046 16890
rect 9098 16838 9110 16890
rect 9162 16838 9174 16890
rect 9226 16838 16982 16890
rect 17034 16838 17046 16890
rect 17098 16838 17110 16890
rect 17162 16838 17174 16890
rect 17226 16838 22816 16890
rect 1104 16816 22816 16838
rect 8754 16776 8760 16788
rect 8715 16748 8760 16776
rect 8754 16736 8760 16748
rect 8812 16736 8818 16788
rect 10226 16736 10232 16788
rect 10284 16776 10290 16788
rect 10321 16779 10379 16785
rect 10321 16776 10333 16779
rect 10284 16748 10333 16776
rect 10284 16736 10290 16748
rect 10321 16745 10333 16748
rect 10367 16745 10379 16779
rect 10321 16739 10379 16745
rect 10873 16779 10931 16785
rect 10873 16745 10885 16779
rect 10919 16776 10931 16779
rect 15565 16779 15623 16785
rect 10919 16748 11928 16776
rect 10919 16745 10931 16748
rect 10873 16739 10931 16745
rect 3970 16668 3976 16720
rect 4028 16708 4034 16720
rect 4203 16711 4261 16717
rect 4203 16708 4215 16711
rect 4028 16680 4215 16708
rect 4028 16668 4034 16680
rect 4203 16677 4215 16680
rect 4249 16677 4261 16711
rect 4203 16671 4261 16677
rect 5626 16668 5632 16720
rect 5684 16708 5690 16720
rect 5807 16711 5865 16717
rect 5807 16708 5819 16711
rect 5684 16680 5819 16708
rect 5684 16668 5690 16680
rect 5807 16677 5819 16680
rect 5853 16708 5865 16711
rect 7926 16708 7932 16720
rect 5853 16680 7932 16708
rect 5853 16677 5865 16680
rect 5807 16671 5865 16677
rect 7926 16668 7932 16680
rect 7984 16708 7990 16720
rect 8199 16711 8257 16717
rect 8199 16708 8211 16711
rect 7984 16680 8211 16708
rect 7984 16668 7990 16680
rect 8199 16677 8211 16680
rect 8245 16708 8257 16711
rect 10244 16708 10272 16736
rect 11900 16720 11928 16748
rect 15565 16745 15577 16779
rect 15611 16776 15623 16779
rect 15746 16776 15752 16788
rect 15611 16748 15752 16776
rect 15611 16745 15623 16748
rect 15565 16739 15623 16745
rect 15746 16736 15752 16748
rect 15804 16736 15810 16788
rect 17313 16779 17371 16785
rect 17313 16745 17325 16779
rect 17359 16776 17371 16779
rect 17402 16776 17408 16788
rect 17359 16748 17408 16776
rect 17359 16745 17371 16748
rect 17313 16739 17371 16745
rect 17402 16736 17408 16748
rect 17460 16736 17466 16788
rect 17862 16776 17868 16788
rect 17823 16748 17868 16776
rect 17862 16736 17868 16748
rect 17920 16736 17926 16788
rect 21085 16779 21143 16785
rect 21085 16745 21097 16779
rect 21131 16776 21143 16779
rect 21726 16776 21732 16788
rect 21131 16748 21732 16776
rect 21131 16745 21143 16748
rect 21085 16739 21143 16745
rect 21726 16736 21732 16748
rect 21784 16736 21790 16788
rect 11882 16708 11888 16720
rect 8245 16680 10272 16708
rect 11795 16680 11888 16708
rect 8245 16677 8257 16680
rect 8199 16671 8257 16677
rect 11882 16668 11888 16680
rect 11940 16668 11946 16720
rect 17420 16708 17448 16736
rect 18325 16711 18383 16717
rect 18325 16708 18337 16711
rect 17420 16680 18337 16708
rect 18325 16677 18337 16680
rect 18371 16677 18383 16711
rect 18874 16708 18880 16720
rect 18835 16680 18880 16708
rect 18325 16671 18383 16677
rect 18874 16668 18880 16680
rect 18932 16668 18938 16720
rect 4111 16643 4169 16649
rect 4111 16609 4123 16643
rect 4157 16609 4169 16643
rect 5442 16640 5448 16652
rect 5403 16612 5448 16640
rect 4111 16603 4169 16609
rect 4126 16504 4154 16603
rect 5442 16600 5448 16612
rect 5500 16600 5506 16652
rect 10870 16640 10876 16652
rect 9646 16612 10876 16640
rect 7837 16575 7895 16581
rect 7837 16541 7849 16575
rect 7883 16572 7895 16575
rect 8478 16572 8484 16584
rect 7883 16544 8484 16572
rect 7883 16541 7895 16544
rect 7837 16535 7895 16541
rect 8478 16532 8484 16544
rect 8536 16532 8542 16584
rect 4430 16504 4436 16516
rect 4126 16476 4436 16504
rect 4430 16464 4436 16476
rect 4488 16504 4494 16516
rect 9646 16504 9674 16612
rect 10870 16600 10876 16612
rect 10928 16600 10934 16652
rect 13538 16600 13544 16652
rect 13596 16640 13602 16652
rect 13633 16643 13691 16649
rect 13633 16640 13645 16643
rect 13596 16612 13645 16640
rect 13596 16600 13602 16612
rect 13633 16609 13645 16612
rect 13679 16609 13691 16643
rect 13633 16603 13691 16609
rect 13906 16600 13912 16652
rect 13964 16640 13970 16652
rect 14093 16643 14151 16649
rect 14093 16640 14105 16643
rect 13964 16612 14105 16640
rect 13964 16600 13970 16612
rect 14093 16609 14105 16612
rect 14139 16609 14151 16643
rect 15286 16640 15292 16652
rect 15247 16612 15292 16640
rect 14093 16603 14151 16609
rect 15286 16600 15292 16612
rect 15344 16600 15350 16652
rect 15746 16640 15752 16652
rect 15707 16612 15752 16640
rect 15746 16600 15752 16612
rect 15804 16600 15810 16652
rect 20898 16640 20904 16652
rect 20859 16612 20904 16640
rect 20898 16600 20904 16612
rect 20956 16640 20962 16652
rect 21266 16640 21272 16652
rect 20956 16612 21272 16640
rect 20956 16600 20962 16612
rect 21266 16600 21272 16612
rect 21324 16600 21330 16652
rect 9766 16532 9772 16584
rect 9824 16572 9830 16584
rect 9953 16575 10011 16581
rect 9953 16572 9965 16575
rect 9824 16544 9965 16572
rect 9824 16532 9830 16544
rect 9953 16541 9965 16544
rect 9999 16541 10011 16575
rect 11790 16572 11796 16584
rect 11751 16544 11796 16572
rect 9953 16535 10011 16541
rect 11790 16532 11796 16544
rect 11848 16532 11854 16584
rect 12158 16572 12164 16584
rect 12119 16544 12164 16572
rect 12158 16532 12164 16544
rect 12216 16532 12222 16584
rect 14366 16572 14372 16584
rect 14327 16544 14372 16572
rect 14366 16532 14372 16544
rect 14424 16532 14430 16584
rect 16942 16572 16948 16584
rect 16855 16544 16948 16572
rect 16942 16532 16948 16544
rect 17000 16572 17006 16584
rect 17770 16572 17776 16584
rect 17000 16544 17776 16572
rect 17000 16532 17006 16544
rect 17770 16532 17776 16544
rect 17828 16532 17834 16584
rect 18782 16572 18788 16584
rect 18743 16544 18788 16572
rect 18782 16532 18788 16544
rect 18840 16532 18846 16584
rect 19058 16572 19064 16584
rect 19019 16544 19064 16572
rect 19058 16532 19064 16544
rect 19116 16532 19122 16584
rect 4488 16476 9674 16504
rect 4488 16464 4494 16476
rect 2593 16439 2651 16445
rect 2593 16405 2605 16439
rect 2639 16436 2651 16439
rect 3142 16436 3148 16448
rect 2639 16408 3148 16436
rect 2639 16405 2651 16408
rect 2593 16399 2651 16405
rect 3142 16396 3148 16408
rect 3200 16396 3206 16448
rect 6362 16436 6368 16448
rect 6323 16408 6368 16436
rect 6362 16396 6368 16408
rect 6420 16436 6426 16448
rect 6825 16439 6883 16445
rect 6825 16436 6837 16439
rect 6420 16408 6837 16436
rect 6420 16396 6426 16408
rect 6825 16405 6837 16408
rect 6871 16436 6883 16439
rect 7006 16436 7012 16448
rect 6871 16408 7012 16436
rect 6871 16405 6883 16408
rect 6825 16399 6883 16405
rect 7006 16396 7012 16408
rect 7064 16396 7070 16448
rect 13446 16436 13452 16448
rect 13407 16408 13452 16436
rect 13446 16396 13452 16408
rect 13504 16436 13510 16448
rect 13906 16436 13912 16448
rect 13504 16408 13912 16436
rect 13504 16396 13510 16408
rect 13906 16396 13912 16408
rect 13964 16396 13970 16448
rect 1104 16346 22816 16368
rect 1104 16294 4982 16346
rect 5034 16294 5046 16346
rect 5098 16294 5110 16346
rect 5162 16294 5174 16346
rect 5226 16294 12982 16346
rect 13034 16294 13046 16346
rect 13098 16294 13110 16346
rect 13162 16294 13174 16346
rect 13226 16294 20982 16346
rect 21034 16294 21046 16346
rect 21098 16294 21110 16346
rect 21162 16294 21174 16346
rect 21226 16294 22816 16346
rect 1104 16272 22816 16294
rect 5442 16192 5448 16244
rect 5500 16232 5506 16244
rect 5813 16235 5871 16241
rect 5813 16232 5825 16235
rect 5500 16204 5825 16232
rect 5500 16192 5506 16204
rect 5813 16201 5825 16204
rect 5859 16201 5871 16235
rect 7926 16232 7932 16244
rect 7887 16204 7932 16232
rect 5813 16195 5871 16201
rect 7926 16192 7932 16204
rect 7984 16192 7990 16244
rect 8297 16235 8355 16241
rect 8297 16201 8309 16235
rect 8343 16232 8355 16235
rect 8478 16232 8484 16244
rect 8343 16204 8484 16232
rect 8343 16201 8355 16204
rect 8297 16195 8355 16201
rect 8478 16192 8484 16204
rect 8536 16192 8542 16244
rect 10137 16235 10195 16241
rect 10137 16201 10149 16235
rect 10183 16232 10195 16235
rect 10226 16232 10232 16244
rect 10183 16204 10232 16232
rect 10183 16201 10195 16204
rect 10137 16195 10195 16201
rect 10226 16192 10232 16204
rect 10284 16192 10290 16244
rect 11882 16232 11888 16244
rect 11843 16204 11888 16232
rect 11882 16192 11888 16204
rect 11940 16192 11946 16244
rect 13357 16235 13415 16241
rect 13357 16201 13369 16235
rect 13403 16232 13415 16235
rect 13446 16232 13452 16244
rect 13403 16204 13452 16232
rect 13403 16201 13415 16204
rect 13357 16195 13415 16201
rect 13446 16192 13452 16204
rect 13504 16192 13510 16244
rect 15286 16232 15292 16244
rect 15247 16204 15292 16232
rect 15286 16192 15292 16204
rect 15344 16192 15350 16244
rect 16022 16232 16028 16244
rect 15983 16204 16028 16232
rect 16022 16192 16028 16204
rect 16080 16192 16086 16244
rect 17129 16235 17187 16241
rect 17129 16201 17141 16235
rect 17175 16232 17187 16235
rect 18874 16232 18880 16244
rect 17175 16204 18880 16232
rect 17175 16201 17187 16204
rect 17129 16195 17187 16201
rect 18874 16192 18880 16204
rect 18932 16232 18938 16244
rect 19521 16235 19579 16241
rect 19521 16232 19533 16235
rect 18932 16204 19533 16232
rect 18932 16192 18938 16204
rect 19521 16201 19533 16204
rect 19567 16201 19579 16235
rect 19521 16195 19579 16201
rect 21177 16235 21235 16241
rect 21177 16201 21189 16235
rect 21223 16232 21235 16235
rect 21266 16232 21272 16244
rect 21223 16204 21272 16232
rect 21223 16201 21235 16204
rect 21177 16195 21235 16201
rect 21266 16192 21272 16204
rect 21324 16192 21330 16244
rect 106 16124 112 16176
rect 164 16164 170 16176
rect 1581 16167 1639 16173
rect 1581 16164 1593 16167
rect 164 16136 1593 16164
rect 164 16124 170 16136
rect 1581 16133 1593 16136
rect 1627 16133 1639 16167
rect 4338 16164 4344 16176
rect 1581 16127 1639 16133
rect 2976 16136 4344 16164
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 1578 16028 1584 16040
rect 1443 16000 1584 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 1578 15988 1584 16000
rect 1636 16028 1642 16040
rect 1949 16031 2007 16037
rect 1949 16028 1961 16031
rect 1636 16000 1961 16028
rect 1636 15988 1642 16000
rect 1949 15997 1961 16000
rect 1995 15997 2007 16031
rect 1949 15991 2007 15997
rect 2409 16031 2467 16037
rect 2409 15997 2421 16031
rect 2455 16028 2467 16031
rect 2777 16031 2835 16037
rect 2777 16028 2789 16031
rect 2455 16000 2789 16028
rect 2455 15997 2467 16000
rect 2409 15991 2467 15997
rect 2777 15997 2789 16000
rect 2823 16028 2835 16031
rect 2976 16028 3004 16136
rect 4338 16124 4344 16136
rect 4396 16164 4402 16176
rect 11425 16167 11483 16173
rect 4396 16136 8984 16164
rect 4396 16124 4402 16136
rect 3973 16099 4031 16105
rect 3973 16065 3985 16099
rect 4019 16096 4031 16099
rect 4430 16096 4436 16108
rect 4019 16068 4436 16096
rect 4019 16065 4031 16068
rect 3973 16059 4031 16065
rect 4430 16056 4436 16068
rect 4488 16056 4494 16108
rect 5537 16099 5595 16105
rect 5537 16065 5549 16099
rect 5583 16096 5595 16099
rect 5626 16096 5632 16108
rect 5583 16068 5632 16096
rect 5583 16065 5595 16068
rect 5537 16059 5595 16065
rect 2823 16000 3004 16028
rect 3053 16031 3111 16037
rect 2823 15997 2835 16000
rect 2777 15991 2835 15997
rect 3053 15997 3065 16031
rect 3099 16028 3111 16031
rect 3142 16028 3148 16040
rect 3099 16000 3148 16028
rect 3099 15997 3111 16000
rect 3053 15991 3111 15997
rect 3142 15988 3148 16000
rect 3200 15988 3206 16040
rect 3237 16031 3295 16037
rect 3237 15997 3249 16031
rect 3283 16028 3295 16031
rect 4065 16031 4123 16037
rect 4065 16028 4077 16031
rect 3283 16000 4077 16028
rect 3283 15997 3295 16000
rect 3237 15991 3295 15997
rect 4065 15997 4077 16000
rect 4111 16028 4123 16031
rect 4246 16028 4252 16040
rect 4111 16000 4252 16028
rect 4111 15997 4123 16000
rect 4065 15991 4123 15997
rect 4246 15988 4252 16000
rect 4304 15988 4310 16040
rect 3605 15963 3663 15969
rect 3605 15929 3617 15963
rect 3651 15960 3663 15963
rect 4154 15960 4160 15972
rect 3651 15932 4160 15960
rect 3651 15929 3663 15932
rect 3605 15923 3663 15929
rect 4154 15920 4160 15932
rect 4212 15960 4218 15972
rect 4427 15963 4485 15969
rect 4427 15960 4439 15963
rect 4212 15932 4439 15960
rect 4212 15920 4218 15932
rect 4427 15929 4439 15932
rect 4473 15960 4485 15963
rect 5552 15960 5580 16059
rect 5626 16056 5632 16068
rect 5684 16056 5690 16108
rect 6273 16099 6331 16105
rect 6273 16065 6285 16099
rect 6319 16096 6331 16099
rect 6914 16096 6920 16108
rect 6319 16068 6920 16096
rect 6319 16065 6331 16068
rect 6273 16059 6331 16065
rect 6914 16056 6920 16068
rect 6972 16056 6978 16108
rect 7190 16096 7196 16108
rect 7151 16068 7196 16096
rect 7190 16056 7196 16068
rect 7248 16056 7254 16108
rect 8956 16037 8984 16136
rect 9646 16136 11376 16164
rect 9646 16096 9674 16136
rect 9324 16068 9674 16096
rect 10873 16099 10931 16105
rect 9324 16037 9352 16068
rect 10873 16065 10885 16099
rect 10919 16096 10931 16099
rect 11238 16096 11244 16108
rect 10919 16068 11244 16096
rect 10919 16065 10931 16068
rect 10873 16059 10931 16065
rect 11238 16056 11244 16068
rect 11296 16056 11302 16108
rect 11348 16096 11376 16136
rect 11425 16133 11437 16167
rect 11471 16164 11483 16167
rect 11790 16164 11796 16176
rect 11471 16136 11796 16164
rect 11471 16133 11483 16136
rect 11425 16127 11483 16133
rect 11790 16124 11796 16136
rect 11848 16164 11854 16176
rect 12161 16167 12219 16173
rect 12161 16164 12173 16167
rect 11848 16136 12173 16164
rect 11848 16124 11854 16136
rect 12161 16133 12173 16136
rect 12207 16133 12219 16167
rect 12161 16127 12219 16133
rect 14366 16124 14372 16176
rect 14424 16164 14430 16176
rect 17773 16167 17831 16173
rect 17773 16164 17785 16167
rect 14424 16136 17785 16164
rect 14424 16124 14430 16136
rect 17773 16133 17785 16136
rect 17819 16133 17831 16167
rect 17773 16127 17831 16133
rect 14921 16099 14979 16105
rect 11348 16068 12848 16096
rect 12820 16040 12848 16068
rect 13786 16068 14688 16096
rect 8941 16031 8999 16037
rect 8941 15997 8953 16031
rect 8987 16028 8999 16031
rect 9309 16031 9367 16037
rect 9309 16028 9321 16031
rect 8987 16000 9321 16028
rect 8987 15997 8999 16000
rect 8941 15991 8999 15997
rect 9309 15997 9321 16000
rect 9355 15997 9367 16031
rect 9490 16028 9496 16040
rect 9451 16000 9496 16028
rect 9309 15991 9367 15997
rect 9490 15988 9496 16000
rect 9548 15988 9554 16040
rect 12802 15988 12808 16040
rect 12860 15988 12866 16040
rect 4473 15932 5580 15960
rect 7009 15963 7067 15969
rect 4473 15929 4485 15932
rect 4427 15923 4485 15929
rect 7009 15929 7021 15963
rect 7055 15929 7067 15963
rect 9766 15960 9772 15972
rect 9727 15932 9772 15960
rect 7009 15923 7067 15929
rect 4982 15892 4988 15904
rect 4943 15864 4988 15892
rect 4982 15852 4988 15864
rect 5040 15852 5046 15904
rect 6362 15852 6368 15904
rect 6420 15892 6426 15904
rect 6549 15895 6607 15901
rect 6549 15892 6561 15895
rect 6420 15864 6561 15892
rect 6420 15852 6426 15864
rect 6549 15861 6561 15864
rect 6595 15892 6607 15895
rect 7024 15892 7052 15923
rect 9766 15920 9772 15932
rect 9824 15920 9830 15972
rect 10594 15920 10600 15972
rect 10652 15960 10658 15972
rect 10689 15963 10747 15969
rect 10689 15960 10701 15963
rect 10652 15932 10701 15960
rect 10652 15920 10658 15932
rect 10689 15929 10701 15932
rect 10735 15960 10747 15963
rect 10965 15963 11023 15969
rect 10965 15960 10977 15963
rect 10735 15932 10977 15960
rect 10735 15929 10747 15932
rect 10689 15923 10747 15929
rect 10965 15929 10977 15932
rect 11011 15929 11023 15963
rect 10965 15923 11023 15929
rect 13446 15920 13452 15972
rect 13504 15960 13510 15972
rect 13786 15960 13814 16068
rect 14660 16040 14688 16068
rect 14921 16065 14933 16099
rect 14967 16096 14979 16099
rect 16942 16096 16948 16108
rect 14967 16068 16948 16096
rect 14967 16065 14979 16068
rect 14921 16059 14979 16065
rect 16942 16056 16948 16068
rect 17000 16056 17006 16108
rect 17788 16096 17816 16127
rect 19058 16124 19064 16176
rect 19116 16164 19122 16176
rect 19116 16136 20484 16164
rect 19116 16124 19122 16136
rect 18325 16099 18383 16105
rect 18325 16096 18337 16099
rect 17788 16068 18337 16096
rect 18325 16065 18337 16068
rect 18371 16065 18383 16099
rect 18325 16059 18383 16065
rect 19978 16056 19984 16108
rect 20036 16096 20042 16108
rect 20456 16105 20484 16136
rect 20165 16099 20223 16105
rect 20165 16096 20177 16099
rect 20036 16068 20177 16096
rect 20036 16056 20042 16068
rect 20165 16065 20177 16068
rect 20211 16065 20223 16099
rect 20165 16059 20223 16065
rect 20441 16099 20499 16105
rect 20441 16065 20453 16099
rect 20487 16065 20499 16099
rect 20441 16059 20499 16065
rect 14185 16031 14243 16037
rect 14185 16028 14197 16031
rect 13504 15932 13814 15960
rect 14016 16000 14197 16028
rect 13504 15920 13510 15932
rect 14016 15904 14044 16000
rect 14185 15997 14197 16000
rect 14231 15997 14243 16031
rect 14642 16028 14648 16040
rect 14603 16000 14648 16028
rect 14185 15991 14243 15997
rect 14642 15988 14648 16000
rect 14700 16028 14706 16040
rect 15657 16031 15715 16037
rect 15657 16028 15669 16031
rect 14700 16000 15669 16028
rect 14700 15988 14706 16000
rect 15657 15997 15669 16000
rect 15703 16028 15715 16031
rect 15746 16028 15752 16040
rect 15703 16000 15752 16028
rect 15703 15997 15715 16000
rect 15657 15991 15715 15997
rect 15746 15988 15752 16000
rect 15804 15988 15810 16040
rect 16206 16028 16212 16040
rect 16167 16000 16212 16028
rect 16206 15988 16212 16000
rect 16264 15988 16270 16040
rect 19245 16031 19303 16037
rect 19245 15997 19257 16031
rect 19291 16028 19303 16031
rect 19889 16031 19947 16037
rect 19889 16028 19901 16031
rect 19291 16000 19901 16028
rect 19291 15997 19303 16000
rect 19245 15991 19303 15997
rect 19889 15997 19901 16000
rect 19935 15997 19947 16031
rect 19889 15991 19947 15997
rect 16022 15920 16028 15972
rect 16080 15960 16086 15972
rect 16530 15963 16588 15969
rect 16530 15960 16542 15963
rect 16080 15932 16542 15960
rect 16080 15920 16086 15932
rect 16530 15929 16542 15932
rect 16576 15960 16588 15963
rect 17402 15960 17408 15972
rect 16576 15932 17408 15960
rect 16576 15929 16588 15932
rect 16530 15923 16588 15929
rect 17402 15920 17408 15932
rect 17460 15960 17466 15972
rect 18646 15963 18704 15969
rect 18646 15960 18658 15963
rect 17460 15932 18658 15960
rect 17460 15920 17466 15932
rect 18646 15929 18658 15932
rect 18692 15929 18704 15963
rect 18646 15923 18704 15929
rect 6595 15864 7052 15892
rect 6595 15861 6607 15864
rect 6549 15855 6607 15861
rect 13538 15852 13544 15904
rect 13596 15892 13602 15904
rect 13633 15895 13691 15901
rect 13633 15892 13645 15895
rect 13596 15864 13645 15892
rect 13596 15852 13602 15864
rect 13633 15861 13645 15864
rect 13679 15861 13691 15895
rect 13998 15892 14004 15904
rect 13959 15864 14004 15892
rect 13633 15855 13691 15861
rect 13998 15852 14004 15864
rect 14056 15852 14062 15904
rect 19904 15892 19932 15991
rect 20257 15963 20315 15969
rect 20257 15929 20269 15963
rect 20303 15929 20315 15963
rect 20257 15923 20315 15929
rect 20272 15892 20300 15923
rect 19904 15864 20300 15892
rect 1104 15802 22816 15824
rect 1104 15750 8982 15802
rect 9034 15750 9046 15802
rect 9098 15750 9110 15802
rect 9162 15750 9174 15802
rect 9226 15750 16982 15802
rect 17034 15750 17046 15802
rect 17098 15750 17110 15802
rect 17162 15750 17174 15802
rect 17226 15750 22816 15802
rect 1104 15728 22816 15750
rect 4246 15688 4252 15700
rect 4207 15660 4252 15688
rect 4246 15648 4252 15660
rect 4304 15648 4310 15700
rect 8386 15688 8392 15700
rect 8347 15660 8392 15688
rect 8386 15648 8392 15660
rect 8444 15688 8450 15700
rect 8846 15688 8852 15700
rect 8444 15660 8852 15688
rect 8444 15648 8450 15660
rect 8846 15648 8852 15660
rect 8904 15688 8910 15700
rect 9033 15691 9091 15697
rect 9033 15688 9045 15691
rect 8904 15660 9045 15688
rect 8904 15648 8910 15660
rect 9033 15657 9045 15660
rect 9079 15688 9091 15691
rect 9490 15688 9496 15700
rect 9079 15660 9496 15688
rect 9079 15657 9091 15660
rect 9033 15651 9091 15657
rect 9490 15648 9496 15660
rect 9548 15648 9554 15700
rect 9766 15648 9772 15700
rect 9824 15688 9830 15700
rect 10689 15691 10747 15697
rect 10689 15688 10701 15691
rect 9824 15660 10701 15688
rect 9824 15648 9830 15660
rect 10689 15657 10701 15660
rect 10735 15657 10747 15691
rect 10689 15651 10747 15657
rect 11149 15691 11207 15697
rect 11149 15657 11161 15691
rect 11195 15688 11207 15691
rect 11238 15688 11244 15700
rect 11195 15660 11244 15688
rect 11195 15657 11207 15660
rect 11149 15651 11207 15657
rect 11238 15648 11244 15660
rect 11296 15648 11302 15700
rect 16574 15688 16580 15700
rect 16535 15660 16580 15688
rect 16574 15648 16580 15660
rect 16632 15648 16638 15700
rect 17770 15688 17776 15700
rect 17731 15660 17776 15688
rect 17770 15648 17776 15660
rect 17828 15648 17834 15700
rect 18782 15688 18788 15700
rect 18743 15660 18788 15688
rect 18782 15648 18788 15660
rect 18840 15648 18846 15700
rect 19978 15648 19984 15700
rect 20036 15688 20042 15700
rect 20073 15691 20131 15697
rect 20073 15688 20085 15691
rect 20036 15660 20085 15688
rect 20036 15648 20042 15660
rect 20073 15657 20085 15660
rect 20119 15657 20131 15691
rect 20073 15651 20131 15657
rect 2590 15620 2596 15632
rect 2551 15592 2596 15620
rect 2590 15580 2596 15592
rect 2648 15580 2654 15632
rect 4062 15580 4068 15632
rect 4120 15620 4126 15632
rect 4709 15623 4767 15629
rect 4709 15620 4721 15623
rect 4120 15592 4721 15620
rect 4120 15580 4126 15592
rect 4709 15589 4721 15592
rect 4755 15620 4767 15623
rect 4982 15620 4988 15632
rect 4755 15592 4988 15620
rect 4755 15589 4767 15592
rect 4709 15583 4767 15589
rect 4982 15580 4988 15592
rect 5040 15580 5046 15632
rect 6546 15620 6552 15632
rect 6507 15592 6552 15620
rect 6546 15580 6552 15592
rect 6604 15580 6610 15632
rect 9508 15620 9536 15648
rect 11606 15620 11612 15632
rect 9508 15592 10180 15620
rect 11567 15592 11612 15620
rect 1464 15555 1522 15561
rect 1464 15521 1476 15555
rect 1510 15552 1522 15555
rect 9674 15552 9680 15564
rect 1510 15524 2360 15552
rect 9635 15524 9680 15552
rect 1510 15521 1522 15524
rect 1464 15515 1522 15521
rect 1578 15484 1584 15496
rect 1550 15444 1584 15484
rect 1636 15444 1642 15496
rect 1550 15357 1578 15444
rect 2332 15425 2360 15524
rect 9674 15512 9680 15524
rect 9732 15512 9738 15564
rect 10152 15561 10180 15592
rect 11606 15580 11612 15592
rect 11664 15580 11670 15632
rect 14369 15623 14427 15629
rect 14369 15589 14381 15623
rect 14415 15620 14427 15623
rect 16206 15620 16212 15632
rect 14415 15592 16212 15620
rect 14415 15589 14427 15592
rect 14369 15583 14427 15589
rect 16206 15580 16212 15592
rect 16264 15580 16270 15632
rect 16850 15580 16856 15632
rect 16908 15620 16914 15632
rect 16945 15623 17003 15629
rect 16945 15620 16957 15623
rect 16908 15592 16957 15620
rect 16908 15580 16914 15592
rect 16945 15589 16957 15592
rect 16991 15589 17003 15623
rect 16945 15583 17003 15589
rect 10137 15555 10195 15561
rect 10137 15521 10149 15555
rect 10183 15521 10195 15555
rect 13630 15552 13636 15564
rect 13591 15524 13636 15552
rect 10137 15515 10195 15521
rect 13630 15512 13636 15524
rect 13688 15512 13694 15564
rect 14182 15552 14188 15564
rect 14143 15524 14188 15552
rect 14182 15512 14188 15524
rect 14240 15552 14246 15564
rect 14642 15552 14648 15564
rect 14240 15524 14648 15552
rect 14240 15512 14246 15524
rect 14642 15512 14648 15524
rect 14700 15512 14706 15564
rect 15657 15555 15715 15561
rect 15657 15521 15669 15555
rect 15703 15552 15715 15555
rect 15746 15552 15752 15564
rect 15703 15524 15752 15552
rect 15703 15521 15715 15524
rect 15657 15515 15715 15521
rect 15746 15512 15752 15524
rect 15804 15512 15810 15564
rect 18322 15552 18328 15564
rect 18283 15524 18328 15552
rect 18322 15512 18328 15524
rect 18380 15512 18386 15564
rect 19058 15512 19064 15564
rect 19116 15552 19122 15564
rect 19372 15555 19430 15561
rect 19372 15552 19384 15555
rect 19116 15524 19384 15552
rect 19116 15512 19122 15524
rect 19372 15521 19384 15524
rect 19418 15521 19430 15555
rect 19372 15515 19430 15521
rect 2498 15484 2504 15496
rect 2459 15456 2504 15484
rect 2498 15444 2504 15456
rect 2556 15444 2562 15496
rect 4614 15484 4620 15496
rect 4575 15456 4620 15484
rect 4614 15444 4620 15456
rect 4672 15444 4678 15496
rect 4893 15487 4951 15493
rect 4893 15453 4905 15487
rect 4939 15453 4951 15487
rect 6454 15484 6460 15496
rect 6367 15456 6460 15484
rect 4893 15447 4951 15453
rect 2317 15419 2375 15425
rect 2317 15385 2329 15419
rect 2363 15416 2375 15419
rect 3053 15419 3111 15425
rect 3053 15416 3065 15419
rect 2363 15388 3065 15416
rect 2363 15385 2375 15388
rect 2317 15379 2375 15385
rect 3053 15385 3065 15388
rect 3099 15416 3111 15419
rect 4798 15416 4804 15428
rect 3099 15388 4804 15416
rect 3099 15385 3111 15388
rect 3053 15379 3111 15385
rect 4798 15376 4804 15388
rect 4856 15416 4862 15428
rect 4908 15416 4936 15447
rect 6454 15444 6460 15456
rect 6512 15484 6518 15496
rect 7929 15487 7987 15493
rect 7929 15484 7941 15487
rect 6512 15456 7941 15484
rect 6512 15444 6518 15456
rect 7929 15453 7941 15456
rect 7975 15453 7987 15487
rect 10410 15484 10416 15496
rect 10371 15456 10416 15484
rect 7929 15447 7987 15453
rect 10410 15444 10416 15456
rect 10468 15444 10474 15496
rect 11146 15444 11152 15496
rect 11204 15484 11210 15496
rect 11517 15487 11575 15493
rect 11517 15484 11529 15487
rect 11204 15456 11529 15484
rect 11204 15444 11210 15456
rect 11517 15453 11529 15456
rect 11563 15484 11575 15487
rect 11790 15484 11796 15496
rect 11563 15456 11796 15484
rect 11563 15453 11575 15456
rect 11517 15447 11575 15453
rect 11790 15444 11796 15456
rect 11848 15444 11854 15496
rect 12158 15484 12164 15496
rect 12119 15456 12164 15484
rect 12158 15444 12164 15456
rect 12216 15444 12222 15496
rect 16842 15487 16900 15493
rect 16842 15484 16854 15487
rect 16776 15456 16854 15484
rect 4856 15388 4936 15416
rect 7009 15419 7067 15425
rect 4856 15376 4862 15388
rect 7009 15385 7021 15419
rect 7055 15416 7067 15419
rect 7190 15416 7196 15428
rect 7055 15388 7196 15416
rect 7055 15385 7067 15388
rect 7009 15379 7067 15385
rect 1535 15351 1593 15357
rect 1535 15317 1547 15351
rect 1581 15317 1593 15351
rect 1854 15348 1860 15360
rect 1815 15320 1860 15348
rect 1535 15311 1593 15317
rect 1854 15308 1860 15320
rect 1912 15308 1918 15360
rect 4614 15308 4620 15360
rect 4672 15348 4678 15360
rect 7024 15348 7052 15379
rect 7190 15376 7196 15388
rect 7248 15376 7254 15428
rect 12526 15348 12532 15360
rect 4672 15320 7052 15348
rect 12487 15320 12532 15348
rect 4672 15308 4678 15320
rect 12526 15308 12532 15320
rect 12584 15308 12590 15360
rect 15887 15351 15945 15357
rect 15887 15317 15899 15351
rect 15933 15348 15945 15351
rect 16482 15348 16488 15360
rect 15933 15320 16488 15348
rect 15933 15317 15945 15320
rect 15887 15311 15945 15317
rect 16482 15308 16488 15320
rect 16540 15308 16546 15360
rect 16776 15348 16804 15456
rect 16842 15453 16854 15456
rect 16888 15453 16900 15487
rect 17310 15484 17316 15496
rect 17271 15456 17316 15484
rect 16842 15447 16900 15453
rect 17310 15444 17316 15456
rect 17368 15444 17374 15496
rect 16850 15348 16856 15360
rect 16763 15320 16856 15348
rect 16850 15308 16856 15320
rect 16908 15348 16914 15360
rect 18463 15351 18521 15357
rect 18463 15348 18475 15351
rect 16908 15320 18475 15348
rect 16908 15308 16914 15320
rect 18463 15317 18475 15320
rect 18509 15317 18521 15351
rect 18463 15311 18521 15317
rect 19475 15351 19533 15357
rect 19475 15317 19487 15351
rect 19521 15348 19533 15351
rect 19794 15348 19800 15360
rect 19521 15320 19800 15348
rect 19521 15317 19533 15320
rect 19475 15311 19533 15317
rect 19794 15308 19800 15320
rect 19852 15308 19858 15360
rect 1104 15258 22816 15280
rect 1104 15206 4982 15258
rect 5034 15206 5046 15258
rect 5098 15206 5110 15258
rect 5162 15206 5174 15258
rect 5226 15206 12982 15258
rect 13034 15206 13046 15258
rect 13098 15206 13110 15258
rect 13162 15206 13174 15258
rect 13226 15206 20982 15258
rect 21034 15206 21046 15258
rect 21098 15206 21110 15258
rect 21162 15206 21174 15258
rect 21226 15206 22816 15258
rect 1104 15184 22816 15206
rect 2590 15104 2596 15156
rect 2648 15144 2654 15156
rect 2685 15147 2743 15153
rect 2685 15144 2697 15147
rect 2648 15116 2697 15144
rect 2648 15104 2654 15116
rect 2685 15113 2697 15116
rect 2731 15144 2743 15147
rect 2961 15147 3019 15153
rect 2961 15144 2973 15147
rect 2731 15116 2973 15144
rect 2731 15113 2743 15116
rect 2685 15107 2743 15113
rect 2961 15113 2973 15116
rect 3007 15113 3019 15147
rect 4062 15144 4068 15156
rect 4023 15116 4068 15144
rect 2961 15107 3019 15113
rect 4062 15104 4068 15116
rect 4120 15104 4126 15156
rect 6454 15144 6460 15156
rect 4540 15116 6316 15144
rect 6415 15116 6460 15144
rect 2498 15036 2504 15088
rect 2556 15076 2562 15088
rect 3329 15079 3387 15085
rect 3329 15076 3341 15079
rect 2556 15048 3341 15076
rect 2556 15036 2562 15048
rect 3329 15045 3341 15048
rect 3375 15076 3387 15079
rect 4540 15076 4568 15116
rect 5350 15076 5356 15088
rect 3375 15048 4568 15076
rect 4632 15048 5356 15076
rect 3375 15045 3387 15048
rect 3329 15039 3387 15045
rect 1765 15011 1823 15017
rect 1765 14977 1777 15011
rect 1811 15008 1823 15011
rect 1854 15008 1860 15020
rect 1811 14980 1860 15008
rect 1811 14977 1823 14980
rect 1765 14971 1823 14977
rect 1854 14968 1860 14980
rect 1912 14968 1918 15020
rect 4632 15017 4660 15048
rect 5350 15036 5356 15048
rect 5408 15036 5414 15088
rect 6288 15076 6316 15116
rect 6454 15104 6460 15116
rect 6512 15104 6518 15156
rect 9861 15147 9919 15153
rect 9861 15113 9873 15147
rect 9907 15144 9919 15147
rect 10226 15144 10232 15156
rect 9907 15116 10232 15144
rect 9907 15113 9919 15116
rect 9861 15107 9919 15113
rect 10226 15104 10232 15116
rect 10284 15104 10290 15156
rect 10873 15147 10931 15153
rect 10873 15113 10885 15147
rect 10919 15144 10931 15147
rect 11517 15147 11575 15153
rect 11517 15144 11529 15147
rect 10919 15116 11529 15144
rect 10919 15113 10931 15116
rect 10873 15107 10931 15113
rect 11517 15113 11529 15116
rect 11563 15144 11575 15147
rect 11606 15144 11612 15156
rect 11563 15116 11612 15144
rect 11563 15113 11575 15116
rect 11517 15107 11575 15113
rect 11606 15104 11612 15116
rect 11664 15104 11670 15156
rect 11790 15144 11796 15156
rect 11751 15116 11796 15144
rect 11790 15104 11796 15116
rect 11848 15104 11854 15156
rect 14182 15104 14188 15156
rect 14240 15144 14246 15156
rect 15013 15147 15071 15153
rect 15013 15144 15025 15147
rect 14240 15116 15025 15144
rect 14240 15104 14246 15116
rect 15013 15113 15025 15116
rect 15059 15113 15071 15147
rect 15746 15144 15752 15156
rect 15707 15116 15752 15144
rect 15013 15107 15071 15113
rect 15746 15104 15752 15116
rect 15804 15104 15810 15156
rect 18322 15144 18328 15156
rect 18283 15116 18328 15144
rect 18322 15104 18328 15116
rect 18380 15104 18386 15156
rect 19058 15104 19064 15156
rect 19116 15144 19122 15156
rect 19521 15147 19579 15153
rect 19521 15144 19533 15147
rect 19116 15116 19533 15144
rect 19116 15104 19122 15116
rect 19521 15113 19533 15116
rect 19567 15113 19579 15147
rect 21450 15144 21456 15156
rect 21411 15116 21456 15144
rect 19521 15107 19579 15113
rect 21450 15104 21456 15116
rect 21508 15104 21514 15156
rect 7469 15079 7527 15085
rect 7469 15076 7481 15079
rect 6288 15048 7481 15076
rect 7469 15045 7481 15048
rect 7515 15076 7527 15079
rect 7558 15076 7564 15088
rect 7515 15048 7564 15076
rect 7515 15045 7527 15048
rect 7469 15039 7527 15045
rect 7558 15036 7564 15048
rect 7616 15036 7622 15088
rect 16574 15076 16580 15088
rect 16224 15048 16580 15076
rect 4617 15011 4675 15017
rect 4617 14977 4629 15011
rect 4663 14977 4675 15011
rect 4617 14971 4675 14977
rect 4798 14968 4804 15020
rect 4856 15008 4862 15020
rect 4893 15011 4951 15017
rect 4893 15008 4905 15011
rect 4856 14980 4905 15008
rect 4856 14968 4862 14980
rect 4893 14977 4905 14980
rect 4939 14977 4951 15011
rect 4893 14971 4951 14977
rect 6917 15011 6975 15017
rect 6917 14977 6929 15011
rect 6963 15008 6975 15011
rect 7190 15008 7196 15020
rect 6963 14980 7196 15008
rect 6963 14977 6975 14980
rect 6917 14971 6975 14977
rect 7190 14968 7196 14980
rect 7248 15008 7254 15020
rect 7837 15011 7895 15017
rect 7837 15008 7849 15011
rect 7248 14980 7849 15008
rect 7248 14968 7254 14980
rect 7837 14977 7849 14980
rect 7883 14977 7895 15011
rect 7837 14971 7895 14977
rect 12158 14968 12164 15020
rect 12216 15008 12222 15020
rect 12805 15011 12863 15017
rect 12805 15008 12817 15011
rect 12216 14980 12817 15008
rect 12216 14968 12222 14980
rect 12805 14977 12817 14980
rect 12851 14977 12863 15011
rect 14366 15008 14372 15020
rect 14279 14980 14372 15008
rect 12805 14971 12863 14977
rect 8389 14943 8447 14949
rect 8389 14909 8401 14943
rect 8435 14909 8447 14943
rect 8846 14940 8852 14952
rect 8807 14912 8852 14940
rect 8389 14903 8447 14909
rect 1673 14875 1731 14881
rect 1673 14841 1685 14875
rect 1719 14872 1731 14875
rect 1762 14872 1768 14884
rect 1719 14844 1768 14872
rect 1719 14841 1731 14844
rect 1673 14835 1731 14841
rect 1762 14832 1768 14844
rect 1820 14872 1826 14884
rect 2086 14875 2144 14881
rect 2086 14872 2098 14875
rect 1820 14844 2098 14872
rect 1820 14832 1826 14844
rect 2086 14841 2098 14844
rect 2132 14841 2144 14875
rect 2086 14835 2144 14841
rect 4709 14875 4767 14881
rect 4709 14841 4721 14875
rect 4755 14841 4767 14875
rect 4709 14835 4767 14841
rect 6089 14875 6147 14881
rect 6089 14841 6101 14875
rect 6135 14872 6147 14875
rect 6546 14872 6552 14884
rect 6135 14844 6552 14872
rect 6135 14841 6147 14844
rect 6089 14835 6147 14841
rect 4433 14807 4491 14813
rect 4433 14773 4445 14807
rect 4479 14804 4491 14807
rect 4724 14804 4752 14835
rect 6546 14832 6552 14844
rect 6604 14872 6610 14884
rect 7006 14872 7012 14884
rect 6604 14844 7012 14872
rect 6604 14832 6610 14844
rect 7006 14832 7012 14844
rect 7064 14832 7070 14884
rect 8202 14872 8208 14884
rect 8163 14844 8208 14872
rect 8202 14832 8208 14844
rect 8260 14872 8266 14884
rect 8404 14872 8432 14903
rect 8846 14900 8852 14912
rect 8904 14900 8910 14952
rect 9125 14943 9183 14949
rect 9125 14909 9137 14943
rect 9171 14940 9183 14943
rect 9950 14940 9956 14952
rect 9171 14912 9956 14940
rect 9171 14909 9183 14912
rect 9125 14903 9183 14909
rect 9950 14900 9956 14912
rect 10008 14900 10014 14952
rect 14292 14949 14320 14980
rect 14366 14968 14372 14980
rect 14424 15008 14430 15020
rect 15286 15008 15292 15020
rect 14424 14980 15292 15008
rect 14424 14968 14430 14980
rect 15286 14968 15292 14980
rect 15344 14968 15350 15020
rect 14277 14943 14335 14949
rect 14277 14909 14289 14943
rect 14323 14909 14335 14943
rect 14458 14940 14464 14952
rect 14419 14912 14464 14940
rect 14277 14903 14335 14909
rect 14458 14900 14464 14912
rect 14516 14900 14522 14952
rect 12526 14872 12532 14884
rect 8260 14844 8432 14872
rect 12487 14844 12532 14872
rect 8260 14832 8266 14844
rect 12526 14832 12532 14844
rect 12584 14832 12590 14884
rect 12621 14875 12679 14881
rect 12621 14841 12633 14875
rect 12667 14841 12679 14875
rect 14734 14872 14740 14884
rect 14695 14844 14740 14872
rect 12621 14835 12679 14841
rect 4982 14804 4988 14816
rect 4479 14776 4988 14804
rect 4479 14773 4491 14776
rect 4433 14767 4491 14773
rect 4982 14764 4988 14776
rect 5040 14764 5046 14816
rect 5350 14764 5356 14816
rect 5408 14804 5414 14816
rect 5629 14807 5687 14813
rect 5629 14804 5641 14807
rect 5408 14776 5641 14804
rect 5408 14764 5414 14776
rect 5629 14773 5641 14776
rect 5675 14804 5687 14807
rect 6822 14804 6828 14816
rect 5675 14776 6828 14804
rect 5675 14773 5687 14776
rect 5629 14767 5687 14773
rect 6822 14764 6828 14776
rect 6880 14764 6886 14816
rect 7742 14764 7748 14816
rect 7800 14804 7806 14816
rect 9401 14807 9459 14813
rect 9401 14804 9413 14807
rect 7800 14776 9413 14804
rect 7800 14764 7806 14776
rect 9401 14773 9413 14776
rect 9447 14804 9459 14807
rect 9674 14804 9680 14816
rect 9447 14776 9680 14804
rect 9447 14773 9459 14776
rect 9401 14767 9459 14773
rect 9674 14764 9680 14776
rect 9732 14764 9738 14816
rect 10226 14764 10232 14816
rect 10284 14804 10290 14816
rect 10321 14807 10379 14813
rect 10321 14804 10333 14807
rect 10284 14776 10333 14804
rect 10284 14764 10290 14776
rect 10321 14773 10333 14776
rect 10367 14773 10379 14807
rect 12158 14804 12164 14816
rect 12119 14776 12164 14804
rect 10321 14767 10379 14773
rect 12158 14764 12164 14776
rect 12216 14804 12222 14816
rect 12636 14804 12664 14835
rect 14734 14832 14740 14844
rect 14792 14832 14798 14884
rect 16224 14872 16252 15048
rect 16574 15036 16580 15048
rect 16632 15036 16638 15088
rect 16390 14968 16396 15020
rect 16448 15008 16454 15020
rect 16669 15011 16727 15017
rect 16669 15008 16681 15011
rect 16448 14980 16681 15008
rect 16448 14968 16454 14980
rect 16669 14977 16681 14980
rect 16715 14977 16727 15011
rect 16669 14971 16727 14977
rect 20968 14943 21026 14949
rect 20968 14909 20980 14943
rect 21014 14940 21026 14943
rect 21450 14940 21456 14952
rect 21014 14912 21456 14940
rect 21014 14909 21026 14912
rect 20968 14903 21026 14909
rect 21450 14900 21456 14912
rect 21508 14900 21514 14952
rect 16393 14875 16451 14881
rect 16393 14872 16405 14875
rect 16224 14844 16405 14872
rect 16393 14841 16405 14844
rect 16439 14841 16451 14875
rect 16393 14835 16451 14841
rect 16485 14875 16543 14881
rect 16485 14841 16497 14875
rect 16531 14841 16543 14875
rect 16485 14835 16543 14841
rect 13630 14804 13636 14816
rect 12216 14776 12664 14804
rect 13591 14776 13636 14804
rect 12216 14764 12222 14776
rect 13630 14764 13636 14776
rect 13688 14764 13694 14816
rect 16206 14804 16212 14816
rect 16167 14776 16212 14804
rect 16206 14764 16212 14776
rect 16264 14804 16270 14816
rect 16500 14804 16528 14835
rect 16264 14776 16528 14804
rect 16264 14764 16270 14776
rect 16758 14764 16764 14816
rect 16816 14804 16822 14816
rect 17313 14807 17371 14813
rect 17313 14804 17325 14807
rect 16816 14776 17325 14804
rect 16816 14764 16822 14776
rect 17313 14773 17325 14776
rect 17359 14804 17371 14807
rect 18230 14804 18236 14816
rect 17359 14776 18236 14804
rect 17359 14773 17371 14776
rect 17313 14767 17371 14773
rect 18230 14764 18236 14776
rect 18288 14764 18294 14816
rect 19058 14804 19064 14816
rect 19019 14776 19064 14804
rect 19058 14764 19064 14776
rect 19116 14764 19122 14816
rect 20714 14764 20720 14816
rect 20772 14804 20778 14816
rect 21039 14807 21097 14813
rect 21039 14804 21051 14807
rect 20772 14776 21051 14804
rect 20772 14764 20778 14776
rect 21039 14773 21051 14776
rect 21085 14773 21097 14807
rect 21039 14767 21097 14773
rect 1104 14714 22816 14736
rect 1104 14662 8982 14714
rect 9034 14662 9046 14714
rect 9098 14662 9110 14714
rect 9162 14662 9174 14714
rect 9226 14662 16982 14714
rect 17034 14662 17046 14714
rect 17098 14662 17110 14714
rect 17162 14662 17174 14714
rect 17226 14662 22816 14714
rect 1104 14640 22816 14662
rect 1854 14560 1860 14612
rect 1912 14600 1918 14612
rect 1949 14603 2007 14609
rect 1949 14600 1961 14603
rect 1912 14572 1961 14600
rect 1912 14560 1918 14572
rect 1949 14569 1961 14572
rect 1995 14569 2007 14603
rect 4982 14600 4988 14612
rect 4943 14572 4988 14600
rect 1949 14563 2007 14569
rect 4982 14560 4988 14572
rect 5040 14560 5046 14612
rect 8018 14600 8024 14612
rect 7979 14572 8024 14600
rect 8018 14560 8024 14572
rect 8076 14560 8082 14612
rect 8846 14560 8852 14612
rect 8904 14600 8910 14612
rect 9861 14603 9919 14609
rect 9861 14600 9873 14603
rect 8904 14572 9873 14600
rect 8904 14560 8910 14572
rect 9861 14569 9873 14572
rect 9907 14569 9919 14603
rect 9861 14563 9919 14569
rect 9950 14560 9956 14612
rect 10008 14600 10014 14612
rect 10229 14603 10287 14609
rect 10229 14600 10241 14603
rect 10008 14572 10241 14600
rect 10008 14560 10014 14572
rect 10229 14569 10241 14572
rect 10275 14569 10287 14603
rect 10229 14563 10287 14569
rect 11425 14603 11483 14609
rect 11425 14569 11437 14603
rect 11471 14600 11483 14603
rect 12158 14600 12164 14612
rect 11471 14572 12164 14600
rect 11471 14569 11483 14572
rect 11425 14563 11483 14569
rect 12158 14560 12164 14572
rect 12216 14560 12222 14612
rect 14366 14600 14372 14612
rect 14327 14572 14372 14600
rect 14366 14560 14372 14572
rect 14424 14560 14430 14612
rect 15010 14560 15016 14612
rect 15068 14600 15074 14612
rect 15657 14603 15715 14609
rect 15657 14600 15669 14603
rect 15068 14572 15669 14600
rect 15068 14560 15074 14572
rect 15657 14569 15669 14572
rect 15703 14569 15715 14603
rect 16206 14600 16212 14612
rect 16167 14572 16212 14600
rect 15657 14563 15715 14569
rect 16206 14560 16212 14572
rect 16264 14560 16270 14612
rect 16850 14600 16856 14612
rect 16811 14572 16856 14600
rect 16850 14560 16856 14572
rect 16908 14560 16914 14612
rect 18230 14560 18236 14612
rect 18288 14600 18294 14612
rect 18288 14572 19380 14600
rect 18288 14560 18294 14572
rect 3786 14492 3792 14544
rect 3844 14532 3850 14544
rect 4154 14532 4160 14544
rect 3844 14504 4160 14532
rect 3844 14492 3850 14504
rect 4154 14492 4160 14504
rect 4212 14532 4218 14544
rect 4386 14535 4444 14541
rect 4386 14532 4398 14535
rect 4212 14504 4398 14532
rect 4212 14492 4218 14504
rect 4386 14501 4398 14504
rect 4432 14501 4444 14535
rect 4386 14495 4444 14501
rect 4614 14492 4620 14544
rect 4672 14532 4678 14544
rect 5261 14535 5319 14541
rect 5261 14532 5273 14535
rect 4672 14504 5273 14532
rect 4672 14492 4678 14504
rect 5261 14501 5273 14504
rect 5307 14501 5319 14535
rect 5261 14495 5319 14501
rect 6273 14535 6331 14541
rect 6273 14501 6285 14535
rect 6319 14532 6331 14535
rect 6362 14532 6368 14544
rect 6319 14504 6368 14532
rect 6319 14501 6331 14504
rect 6273 14495 6331 14501
rect 6362 14492 6368 14504
rect 6420 14492 6426 14544
rect 1946 14464 1952 14476
rect 1907 14436 1952 14464
rect 1946 14424 1952 14436
rect 2004 14424 2010 14476
rect 2225 14467 2283 14473
rect 2225 14433 2237 14467
rect 2271 14464 2283 14467
rect 3510 14464 3516 14476
rect 2271 14436 3516 14464
rect 2271 14433 2283 14436
rect 2225 14427 2283 14433
rect 3510 14424 3516 14436
rect 3568 14424 3574 14476
rect 7834 14424 7840 14476
rect 7892 14464 7898 14476
rect 8021 14467 8079 14473
rect 8021 14464 8033 14467
rect 7892 14436 8033 14464
rect 7892 14424 7898 14436
rect 8021 14433 8033 14436
rect 8067 14464 8079 14467
rect 8110 14464 8116 14476
rect 8067 14436 8116 14464
rect 8067 14433 8079 14436
rect 8021 14427 8079 14433
rect 8110 14424 8116 14436
rect 8168 14424 8174 14476
rect 8294 14464 8300 14476
rect 8207 14436 8300 14464
rect 8294 14424 8300 14436
rect 8352 14464 8358 14476
rect 8864 14464 8892 14560
rect 10318 14492 10324 14544
rect 10376 14532 10382 14544
rect 10826 14535 10884 14541
rect 10826 14532 10838 14535
rect 10376 14504 10838 14532
rect 10376 14492 10382 14504
rect 10826 14501 10838 14504
rect 10872 14501 10884 14535
rect 16224 14532 16252 14560
rect 17221 14535 17279 14541
rect 17221 14532 17233 14535
rect 16224 14504 17233 14532
rect 10826 14495 10884 14501
rect 17221 14501 17233 14504
rect 17267 14501 17279 14535
rect 17221 14495 17279 14501
rect 19058 14492 19064 14544
rect 19116 14532 19122 14544
rect 19352 14541 19380 14572
rect 19245 14535 19303 14541
rect 19245 14532 19257 14535
rect 19116 14504 19257 14532
rect 19116 14492 19122 14504
rect 19245 14501 19257 14504
rect 19291 14501 19303 14535
rect 19245 14495 19303 14501
rect 19337 14535 19395 14541
rect 19337 14501 19349 14535
rect 19383 14532 19395 14535
rect 19610 14532 19616 14544
rect 19383 14504 19616 14532
rect 19383 14501 19395 14504
rect 19337 14495 19395 14501
rect 19610 14492 19616 14504
rect 19668 14492 19674 14544
rect 8352 14436 8892 14464
rect 8352 14424 8358 14436
rect 10410 14424 10416 14476
rect 10468 14464 10474 14476
rect 10505 14467 10563 14473
rect 10505 14464 10517 14467
rect 10468 14436 10517 14464
rect 10468 14424 10474 14436
rect 10505 14433 10517 14436
rect 10551 14464 10563 14467
rect 10551 14436 10916 14464
rect 10551 14433 10563 14436
rect 10505 14427 10563 14433
rect 10888 14408 10916 14436
rect 13262 14424 13268 14476
rect 13320 14464 13326 14476
rect 13357 14467 13415 14473
rect 13357 14464 13369 14467
rect 13320 14436 13369 14464
rect 13320 14424 13326 14436
rect 13357 14433 13369 14436
rect 13403 14433 13415 14467
rect 13357 14427 13415 14433
rect 13909 14467 13967 14473
rect 13909 14433 13921 14467
rect 13955 14433 13967 14467
rect 13909 14427 13967 14433
rect 4062 14396 4068 14408
rect 4023 14368 4068 14396
rect 4062 14356 4068 14368
rect 4120 14356 4126 14408
rect 6181 14399 6239 14405
rect 6181 14396 6193 14399
rect 5920 14368 6193 14396
rect 5920 14272 5948 14368
rect 6181 14365 6193 14368
rect 6227 14365 6239 14399
rect 6822 14396 6828 14408
rect 6783 14368 6828 14396
rect 6181 14359 6239 14365
rect 6822 14356 6828 14368
rect 6880 14356 6886 14408
rect 10870 14356 10876 14408
rect 10928 14356 10934 14408
rect 9674 14288 9680 14340
rect 9732 14328 9738 14340
rect 13630 14328 13636 14340
rect 9732 14300 13636 14328
rect 9732 14288 9738 14300
rect 13630 14288 13636 14300
rect 13688 14288 13694 14340
rect 13924 14328 13952 14427
rect 14734 14424 14740 14476
rect 14792 14464 14798 14476
rect 15289 14467 15347 14473
rect 15289 14464 15301 14467
rect 14792 14436 15301 14464
rect 14792 14424 14798 14436
rect 15289 14433 15301 14436
rect 15335 14464 15347 14467
rect 15654 14464 15660 14476
rect 15335 14436 15660 14464
rect 15335 14433 15347 14436
rect 15289 14427 15347 14433
rect 15654 14424 15660 14436
rect 15712 14424 15718 14476
rect 14090 14396 14096 14408
rect 14051 14368 14096 14396
rect 14090 14356 14096 14368
rect 14148 14356 14154 14408
rect 16482 14356 16488 14408
rect 16540 14396 16546 14408
rect 17129 14399 17187 14405
rect 17129 14396 17141 14399
rect 16540 14368 17141 14396
rect 16540 14356 16546 14368
rect 17129 14365 17141 14368
rect 17175 14396 17187 14399
rect 17586 14396 17592 14408
rect 17175 14368 17592 14396
rect 17175 14365 17187 14368
rect 17129 14359 17187 14365
rect 17586 14356 17592 14368
rect 17644 14356 17650 14408
rect 17773 14399 17831 14405
rect 17773 14365 17785 14399
rect 17819 14396 17831 14399
rect 18874 14396 18880 14408
rect 17819 14368 18880 14396
rect 17819 14365 17831 14368
rect 17773 14359 17831 14365
rect 18874 14356 18880 14368
rect 18932 14356 18938 14408
rect 19521 14399 19579 14405
rect 19521 14396 19533 14399
rect 19306 14368 19533 14396
rect 19306 14340 19334 14368
rect 19521 14365 19533 14368
rect 19567 14365 19579 14399
rect 19521 14359 19579 14365
rect 14458 14328 14464 14340
rect 13924 14300 14464 14328
rect 14458 14288 14464 14300
rect 14516 14328 14522 14340
rect 14516 14300 14780 14328
rect 14516 14288 14522 14300
rect 14752 14272 14780 14300
rect 16298 14288 16304 14340
rect 16356 14328 16362 14340
rect 19242 14328 19248 14340
rect 16356 14300 19248 14328
rect 16356 14288 16362 14300
rect 19242 14288 19248 14300
rect 19300 14300 19334 14340
rect 19300 14288 19306 14300
rect 2682 14260 2688 14272
rect 2643 14232 2688 14260
rect 2682 14220 2688 14232
rect 2740 14220 2746 14272
rect 3878 14260 3884 14272
rect 3839 14232 3884 14260
rect 3878 14220 3884 14232
rect 3936 14220 3942 14272
rect 5902 14260 5908 14272
rect 5863 14232 5908 14260
rect 5902 14220 5908 14232
rect 5960 14220 5966 14272
rect 7006 14220 7012 14272
rect 7064 14260 7070 14272
rect 7101 14263 7159 14269
rect 7101 14260 7113 14263
rect 7064 14232 7113 14260
rect 7064 14220 7070 14232
rect 7101 14229 7113 14232
rect 7147 14229 7159 14263
rect 12526 14260 12532 14272
rect 12487 14232 12532 14260
rect 7101 14223 7159 14229
rect 12526 14220 12532 14232
rect 12584 14220 12590 14272
rect 14734 14260 14740 14272
rect 14695 14232 14740 14260
rect 14734 14220 14740 14232
rect 14792 14220 14798 14272
rect 1104 14170 22816 14192
rect 1104 14118 4982 14170
rect 5034 14118 5046 14170
rect 5098 14118 5110 14170
rect 5162 14118 5174 14170
rect 5226 14118 12982 14170
rect 13034 14118 13046 14170
rect 13098 14118 13110 14170
rect 13162 14118 13174 14170
rect 13226 14118 20982 14170
rect 21034 14118 21046 14170
rect 21098 14118 21110 14170
rect 21162 14118 21174 14170
rect 21226 14118 22816 14170
rect 1104 14096 22816 14118
rect 1762 14056 1768 14068
rect 1723 14028 1768 14056
rect 1762 14016 1768 14028
rect 1820 14056 1826 14068
rect 2130 14056 2136 14068
rect 1820 14028 2136 14056
rect 1820 14016 1826 14028
rect 2130 14016 2136 14028
rect 2188 14056 2194 14068
rect 3786 14056 3792 14068
rect 2188 14028 3792 14056
rect 2188 14016 2194 14028
rect 3786 14016 3792 14028
rect 3844 14016 3850 14068
rect 4062 14016 4068 14068
rect 4120 14056 4126 14068
rect 5353 14059 5411 14065
rect 5353 14056 5365 14059
rect 4120 14028 5365 14056
rect 4120 14016 4126 14028
rect 5353 14025 5365 14028
rect 5399 14025 5411 14059
rect 6362 14056 6368 14068
rect 6323 14028 6368 14056
rect 5353 14019 5411 14025
rect 6362 14016 6368 14028
rect 6420 14016 6426 14068
rect 10226 14056 10232 14068
rect 10187 14028 10232 14056
rect 10226 14016 10232 14028
rect 10284 14016 10290 14068
rect 10594 14016 10600 14068
rect 10652 14056 10658 14068
rect 12161 14059 12219 14065
rect 12161 14056 12173 14059
rect 10652 14028 12173 14056
rect 10652 14016 10658 14028
rect 12161 14025 12173 14028
rect 12207 14056 12219 14059
rect 12618 14056 12624 14068
rect 12207 14028 12624 14056
rect 12207 14025 12219 14028
rect 12161 14019 12219 14025
rect 12618 14016 12624 14028
rect 12676 14016 12682 14068
rect 15654 14056 15660 14068
rect 15615 14028 15660 14056
rect 15654 14016 15660 14028
rect 15712 14016 15718 14068
rect 16206 14056 16212 14068
rect 16167 14028 16212 14056
rect 16206 14016 16212 14028
rect 16264 14056 16270 14068
rect 16574 14056 16580 14068
rect 16264 14028 16580 14056
rect 16264 14016 16270 14028
rect 16574 14016 16580 14028
rect 16632 14056 16638 14068
rect 17405 14059 17463 14065
rect 17405 14056 17417 14059
rect 16632 14028 17417 14056
rect 16632 14016 16638 14028
rect 17405 14025 17417 14028
rect 17451 14025 17463 14059
rect 17405 14019 17463 14025
rect 17586 14016 17592 14068
rect 17644 14056 17650 14068
rect 17773 14059 17831 14065
rect 17773 14056 17785 14059
rect 17644 14028 17785 14056
rect 17644 14016 17650 14028
rect 17773 14025 17785 14028
rect 17819 14025 17831 14059
rect 17773 14019 17831 14025
rect 19058 14016 19064 14068
rect 19116 14056 19122 14068
rect 19153 14059 19211 14065
rect 19153 14056 19165 14059
rect 19116 14028 19165 14056
rect 19116 14016 19122 14028
rect 19153 14025 19165 14028
rect 19199 14025 19211 14059
rect 19153 14019 19211 14025
rect 5675 13991 5733 13997
rect 5675 13988 5687 13991
rect 4080 13960 5687 13988
rect 1857 13923 1915 13929
rect 1857 13889 1869 13923
rect 1903 13920 1915 13923
rect 2222 13920 2228 13932
rect 1903 13892 2228 13920
rect 1903 13889 1915 13892
rect 1857 13883 1915 13889
rect 2222 13880 2228 13892
rect 2280 13920 2286 13932
rect 2682 13920 2688 13932
rect 2280 13892 2688 13920
rect 2280 13880 2286 13892
rect 2682 13880 2688 13892
rect 2740 13880 2746 13932
rect 3878 13880 3884 13932
rect 3936 13920 3942 13932
rect 4080 13929 4108 13960
rect 5675 13957 5687 13960
rect 5721 13957 5733 13991
rect 5675 13951 5733 13957
rect 8941 13991 8999 13997
rect 8941 13957 8953 13991
rect 8987 13988 8999 13991
rect 9858 13988 9864 14000
rect 8987 13960 9352 13988
rect 9819 13960 9864 13988
rect 8987 13957 8999 13960
rect 8941 13951 8999 13957
rect 4054 13923 4112 13929
rect 4054 13920 4066 13923
rect 3936 13892 4066 13920
rect 3936 13880 3942 13892
rect 4054 13889 4066 13892
rect 4100 13889 4112 13923
rect 4054 13883 4112 13889
rect 4709 13923 4767 13929
rect 4709 13889 4721 13923
rect 4755 13920 4767 13923
rect 5350 13920 5356 13932
rect 4755 13892 5356 13920
rect 4755 13889 4767 13892
rect 4709 13883 4767 13889
rect 5350 13880 5356 13892
rect 5408 13880 5414 13932
rect 8018 13920 8024 13932
rect 5603 13892 6040 13920
rect 7979 13892 8024 13920
rect 5603 13861 5631 13892
rect 2777 13855 2835 13861
rect 2777 13821 2789 13855
rect 2823 13852 2835 13855
rect 5588 13855 5646 13861
rect 2823 13824 2857 13852
rect 2823 13821 2835 13824
rect 2777 13815 2835 13821
rect 5588 13821 5600 13855
rect 5634 13821 5646 13855
rect 5588 13815 5646 13821
rect 2130 13784 2136 13796
rect 2091 13756 2136 13784
rect 2130 13744 2136 13756
rect 2188 13744 2194 13796
rect 2792 13784 2820 13815
rect 3694 13784 3700 13796
rect 2792 13756 3700 13784
rect 3694 13744 3700 13756
rect 3752 13784 3758 13796
rect 4157 13787 4215 13793
rect 4157 13784 4169 13787
rect 3752 13756 4169 13784
rect 3752 13744 3758 13756
rect 4157 13753 4169 13756
rect 4203 13784 4215 13787
rect 4985 13787 5043 13793
rect 4985 13784 4997 13787
rect 4203 13756 4997 13784
rect 4203 13753 4215 13756
rect 4157 13747 4215 13753
rect 4985 13753 4997 13756
rect 5031 13753 5043 13787
rect 4985 13747 5043 13753
rect 1946 13676 1952 13728
rect 2004 13716 2010 13728
rect 3142 13716 3148 13728
rect 2004 13688 3148 13716
rect 2004 13676 2010 13688
rect 3142 13676 3148 13688
rect 3200 13676 3206 13728
rect 3510 13716 3516 13728
rect 3423 13688 3516 13716
rect 3510 13676 3516 13688
rect 3568 13716 3574 13728
rect 3878 13716 3884 13728
rect 3568 13688 3884 13716
rect 3568 13676 3574 13688
rect 3878 13676 3884 13688
rect 3936 13676 3942 13728
rect 6012 13725 6040 13892
rect 8018 13880 8024 13892
rect 8076 13920 8082 13932
rect 9217 13923 9275 13929
rect 9217 13920 9229 13923
rect 8076 13892 9229 13920
rect 8076 13880 8082 13892
rect 9217 13889 9229 13892
rect 9263 13889 9275 13923
rect 9217 13883 9275 13889
rect 6454 13812 6460 13864
rect 6512 13852 6518 13864
rect 6876 13855 6934 13861
rect 6876 13852 6888 13855
rect 6512 13824 6888 13852
rect 6512 13812 6518 13824
rect 6876 13821 6888 13824
rect 6922 13852 6934 13855
rect 7285 13855 7343 13861
rect 7285 13852 7297 13855
rect 6922 13824 7297 13852
rect 6922 13821 6934 13824
rect 6876 13815 6934 13821
rect 7285 13821 7297 13824
rect 7331 13821 7343 13855
rect 7285 13815 7343 13821
rect 9324 13784 9352 13960
rect 9858 13948 9864 13960
rect 9916 13948 9922 14000
rect 11057 13991 11115 13997
rect 11057 13957 11069 13991
rect 11103 13988 11115 13991
rect 11514 13988 11520 14000
rect 11103 13960 11520 13988
rect 11103 13957 11115 13960
rect 11057 13951 11115 13957
rect 11514 13948 11520 13960
rect 11572 13988 11578 14000
rect 12434 13988 12440 14000
rect 11572 13960 12440 13988
rect 11572 13948 11578 13960
rect 12434 13948 12440 13960
rect 12492 13948 12498 14000
rect 13262 13948 13268 14000
rect 13320 13988 13326 14000
rect 13449 13991 13507 13997
rect 13449 13988 13461 13991
rect 13320 13960 13461 13988
rect 13320 13948 13326 13960
rect 13449 13957 13461 13960
rect 13495 13957 13507 13991
rect 13449 13951 13507 13957
rect 15013 13991 15071 13997
rect 15013 13957 15025 13991
rect 15059 13988 15071 13991
rect 16758 13988 16764 14000
rect 15059 13960 16764 13988
rect 15059 13957 15071 13960
rect 15013 13951 15071 13957
rect 16758 13948 16764 13960
rect 16816 13948 16822 14000
rect 9876 13852 9904 13948
rect 10502 13920 10508 13932
rect 10415 13892 10508 13920
rect 10502 13880 10508 13892
rect 10560 13920 10566 13932
rect 11425 13923 11483 13929
rect 11425 13920 11437 13923
rect 10560 13892 11437 13920
rect 10560 13880 10566 13892
rect 11425 13889 11437 13892
rect 11471 13889 11483 13923
rect 11425 13883 11483 13889
rect 11790 13880 11796 13932
rect 11848 13920 11854 13932
rect 12805 13923 12863 13929
rect 12805 13920 12817 13923
rect 11848 13892 12817 13920
rect 11848 13880 11854 13892
rect 12805 13889 12817 13892
rect 12851 13889 12863 13923
rect 14090 13920 14096 13932
rect 14051 13892 14096 13920
rect 12805 13883 12863 13889
rect 14090 13880 14096 13892
rect 14148 13880 14154 13932
rect 17129 13923 17187 13929
rect 17129 13889 17141 13923
rect 17175 13920 17187 13923
rect 17310 13920 17316 13932
rect 17175 13892 17316 13920
rect 17175 13889 17187 13892
rect 17129 13883 17187 13889
rect 17310 13880 17316 13892
rect 17368 13880 17374 13932
rect 18360 13855 18418 13861
rect 18360 13852 18372 13855
rect 9692 13824 9904 13852
rect 17972 13824 18372 13852
rect 9398 13784 9404 13796
rect 9324 13756 9404 13784
rect 9398 13744 9404 13756
rect 9456 13744 9462 13796
rect 9692 13784 9720 13824
rect 10597 13787 10655 13793
rect 10597 13784 10609 13787
rect 9692 13756 10609 13784
rect 10597 13753 10609 13756
rect 10643 13753 10655 13787
rect 12526 13784 12532 13796
rect 12487 13756 12532 13784
rect 10597 13747 10655 13753
rect 12526 13744 12532 13756
rect 12584 13744 12590 13796
rect 12618 13744 12624 13796
rect 12676 13784 12682 13796
rect 14001 13787 14059 13793
rect 14001 13784 14013 13787
rect 12676 13756 12721 13784
rect 13786 13756 14013 13784
rect 12676 13744 12682 13756
rect 5997 13719 6055 13725
rect 5997 13716 6009 13719
rect 5907 13688 6009 13716
rect 5997 13685 6009 13688
rect 6043 13716 6055 13719
rect 6086 13716 6092 13728
rect 6043 13688 6092 13716
rect 6043 13685 6055 13688
rect 5997 13679 6055 13685
rect 6086 13676 6092 13688
rect 6144 13676 6150 13728
rect 6730 13676 6736 13728
rect 6788 13716 6794 13728
rect 6963 13719 7021 13725
rect 6963 13716 6975 13719
rect 6788 13688 6975 13716
rect 6788 13676 6794 13688
rect 6963 13685 6975 13688
rect 7009 13685 7021 13719
rect 6963 13679 7021 13685
rect 7929 13719 7987 13725
rect 7929 13685 7941 13719
rect 7975 13716 7987 13719
rect 8386 13716 8392 13728
rect 7975 13688 8392 13716
rect 7975 13685 7987 13688
rect 7929 13679 7987 13685
rect 8386 13676 8392 13688
rect 8444 13676 8450 13728
rect 10226 13676 10232 13728
rect 10284 13716 10290 13728
rect 13786 13716 13814 13756
rect 14001 13753 14013 13756
rect 14047 13784 14059 13787
rect 14455 13787 14513 13793
rect 14455 13784 14467 13787
rect 14047 13756 14467 13784
rect 14047 13753 14059 13756
rect 14001 13747 14059 13753
rect 14455 13753 14467 13756
rect 14501 13784 14513 13787
rect 16482 13784 16488 13796
rect 14501 13756 15056 13784
rect 16443 13756 16488 13784
rect 14501 13753 14513 13756
rect 14455 13747 14513 13753
rect 15028 13728 15056 13756
rect 16482 13744 16488 13756
rect 16540 13744 16546 13796
rect 16574 13744 16580 13796
rect 16632 13784 16638 13796
rect 16632 13756 16677 13784
rect 16632 13744 16638 13756
rect 10284 13688 13814 13716
rect 10284 13676 10290 13688
rect 15010 13676 15016 13728
rect 15068 13716 15074 13728
rect 15286 13716 15292 13728
rect 15068 13688 15292 13716
rect 15068 13676 15074 13688
rect 15286 13676 15292 13688
rect 15344 13676 15350 13728
rect 15378 13676 15384 13728
rect 15436 13716 15442 13728
rect 17972 13716 18000 13824
rect 18340 13821 18372 13824
rect 18406 13821 18418 13855
rect 18340 13815 18418 13821
rect 18463 13855 18521 13861
rect 18463 13821 18475 13855
rect 18509 13852 18521 13855
rect 18782 13852 18788 13864
rect 18509 13824 18788 13852
rect 18509 13821 18521 13824
rect 18463 13815 18521 13821
rect 18340 13784 18368 13815
rect 18782 13812 18788 13824
rect 18840 13812 18846 13864
rect 20968 13855 21026 13861
rect 20968 13821 20980 13855
rect 21014 13852 21026 13855
rect 21014 13824 21496 13852
rect 21014 13821 21026 13824
rect 20968 13815 21026 13821
rect 18877 13787 18935 13793
rect 18877 13784 18889 13787
rect 18340 13756 18889 13784
rect 18877 13753 18889 13756
rect 18923 13753 18935 13787
rect 19426 13784 19432 13796
rect 19387 13756 19432 13784
rect 18877 13747 18935 13753
rect 15436 13688 18000 13716
rect 18892 13716 18920 13747
rect 19426 13744 19432 13756
rect 19484 13744 19490 13796
rect 19521 13787 19579 13793
rect 19521 13753 19533 13787
rect 19567 13753 19579 13787
rect 20070 13784 20076 13796
rect 20031 13756 20076 13784
rect 19521 13747 19579 13753
rect 19334 13716 19340 13728
rect 18892 13688 19340 13716
rect 15436 13676 15442 13688
rect 19334 13676 19340 13688
rect 19392 13676 19398 13728
rect 19536 13716 19564 13747
rect 20070 13744 20076 13756
rect 20128 13744 20134 13796
rect 20530 13744 20536 13796
rect 20588 13784 20594 13796
rect 20806 13784 20812 13796
rect 20588 13756 20812 13784
rect 20588 13744 20594 13756
rect 20806 13744 20812 13756
rect 20864 13744 20870 13796
rect 21468 13793 21496 13824
rect 21453 13787 21511 13793
rect 21453 13784 21465 13787
rect 21363 13756 21465 13784
rect 21453 13753 21465 13756
rect 21499 13784 21511 13787
rect 21726 13784 21732 13796
rect 21499 13756 21732 13784
rect 21499 13753 21511 13756
rect 21453 13747 21511 13753
rect 21726 13744 21732 13756
rect 21784 13744 21790 13796
rect 19610 13716 19616 13728
rect 19523 13688 19616 13716
rect 19610 13676 19616 13688
rect 19668 13716 19674 13728
rect 20349 13719 20407 13725
rect 20349 13716 20361 13719
rect 19668 13688 20361 13716
rect 19668 13676 19674 13688
rect 20349 13685 20361 13688
rect 20395 13685 20407 13719
rect 20349 13679 20407 13685
rect 20438 13676 20444 13728
rect 20496 13716 20502 13728
rect 21039 13719 21097 13725
rect 21039 13716 21051 13719
rect 20496 13688 21051 13716
rect 20496 13676 20502 13688
rect 21039 13685 21051 13688
rect 21085 13685 21097 13719
rect 21039 13679 21097 13685
rect 1104 13626 22816 13648
rect 1104 13574 8982 13626
rect 9034 13574 9046 13626
rect 9098 13574 9110 13626
rect 9162 13574 9174 13626
rect 9226 13574 16982 13626
rect 17034 13574 17046 13626
rect 17098 13574 17110 13626
rect 17162 13574 17174 13626
rect 17226 13574 22816 13626
rect 1104 13552 22816 13574
rect 4062 13472 4068 13524
rect 4120 13512 4126 13524
rect 4157 13515 4215 13521
rect 4157 13512 4169 13515
rect 4120 13484 4169 13512
rect 4120 13472 4126 13484
rect 4157 13481 4169 13484
rect 4203 13481 4215 13515
rect 4157 13475 4215 13481
rect 6825 13515 6883 13521
rect 6825 13481 6837 13515
rect 6871 13512 6883 13515
rect 7006 13512 7012 13524
rect 6871 13484 7012 13512
rect 6871 13481 6883 13484
rect 6825 13475 6883 13481
rect 7006 13472 7012 13484
rect 7064 13512 7070 13524
rect 7101 13515 7159 13521
rect 7101 13512 7113 13515
rect 7064 13484 7113 13512
rect 7064 13472 7070 13484
rect 7101 13481 7113 13484
rect 7147 13481 7159 13515
rect 7834 13512 7840 13524
rect 7795 13484 7840 13512
rect 7101 13475 7159 13481
rect 7834 13472 7840 13484
rect 7892 13472 7898 13524
rect 8202 13472 8208 13524
rect 8260 13512 8266 13524
rect 10594 13512 10600 13524
rect 8260 13484 10247 13512
rect 10555 13484 10600 13512
rect 8260 13472 8266 13484
rect 2222 13444 2228 13456
rect 2183 13416 2228 13444
rect 2222 13404 2228 13416
rect 2280 13404 2286 13456
rect 6267 13447 6325 13453
rect 6267 13413 6279 13447
rect 6313 13444 6325 13447
rect 6546 13444 6552 13456
rect 6313 13416 6552 13444
rect 6313 13413 6325 13416
rect 6267 13407 6325 13413
rect 6546 13404 6552 13416
rect 6604 13444 6610 13456
rect 8386 13444 8392 13456
rect 6604 13416 8392 13444
rect 6604 13404 6610 13416
rect 8386 13404 8392 13416
rect 8444 13444 8450 13456
rect 9926 13447 9984 13453
rect 9926 13444 9938 13447
rect 8444 13416 9938 13444
rect 8444 13404 8450 13416
rect 9926 13413 9938 13416
rect 9972 13444 9984 13447
rect 10042 13444 10048 13456
rect 9972 13416 10048 13444
rect 9972 13413 9984 13416
rect 9926 13407 9984 13413
rect 10042 13404 10048 13416
rect 10100 13404 10106 13456
rect 10219 13444 10247 13484
rect 10594 13472 10600 13484
rect 10652 13472 10658 13524
rect 10870 13512 10876 13524
rect 10831 13484 10876 13512
rect 10870 13472 10876 13484
rect 10928 13472 10934 13524
rect 11882 13512 11888 13524
rect 11624 13484 11888 13512
rect 11624 13444 11652 13484
rect 11882 13472 11888 13484
rect 11940 13512 11946 13524
rect 13538 13512 13544 13524
rect 11940 13484 13544 13512
rect 11940 13472 11946 13484
rect 13538 13472 13544 13484
rect 13596 13472 13602 13524
rect 14090 13512 14096 13524
rect 14051 13484 14096 13512
rect 14090 13472 14096 13484
rect 14148 13472 14154 13524
rect 17402 13472 17408 13524
rect 17460 13512 17466 13524
rect 18049 13515 18107 13521
rect 18049 13512 18061 13515
rect 17460 13484 18061 13512
rect 17460 13472 17466 13484
rect 18049 13481 18061 13484
rect 18095 13512 18107 13515
rect 18138 13512 18144 13524
rect 18095 13484 18144 13512
rect 18095 13481 18107 13484
rect 18049 13475 18107 13481
rect 18138 13472 18144 13484
rect 18196 13512 18202 13524
rect 19610 13512 19616 13524
rect 18196 13484 19288 13512
rect 19571 13484 19616 13512
rect 18196 13472 18202 13484
rect 10219 13416 11652 13444
rect 11701 13447 11759 13453
rect 11701 13413 11713 13447
rect 11747 13444 11759 13447
rect 11790 13444 11796 13456
rect 11747 13416 11796 13444
rect 11747 13413 11759 13416
rect 11701 13407 11759 13413
rect 11790 13404 11796 13416
rect 11848 13404 11854 13456
rect 12253 13447 12311 13453
rect 12253 13413 12265 13447
rect 12299 13444 12311 13447
rect 12434 13444 12440 13456
rect 12299 13416 12440 13444
rect 12299 13413 12311 13416
rect 12253 13407 12311 13413
rect 12434 13404 12440 13416
rect 12492 13404 12498 13456
rect 16850 13444 16856 13456
rect 16811 13416 16856 13444
rect 16850 13404 16856 13416
rect 16908 13404 16914 13456
rect 18693 13447 18751 13453
rect 18693 13413 18705 13447
rect 18739 13444 18751 13447
rect 19058 13444 19064 13456
rect 18739 13416 19064 13444
rect 18739 13413 18751 13416
rect 18693 13407 18751 13413
rect 19058 13404 19064 13416
rect 19116 13404 19122 13456
rect 19260 13453 19288 13484
rect 19610 13472 19616 13484
rect 19668 13472 19674 13524
rect 20070 13472 20076 13524
rect 20128 13512 20134 13524
rect 20128 13484 21220 13512
rect 20128 13472 20134 13484
rect 19245 13447 19303 13453
rect 19245 13413 19257 13447
rect 19291 13413 19303 13447
rect 19245 13407 19303 13413
rect 20806 13404 20812 13456
rect 20864 13444 20870 13456
rect 21085 13447 21143 13453
rect 21085 13444 21097 13447
rect 20864 13416 21097 13444
rect 20864 13404 20870 13416
rect 21085 13413 21097 13416
rect 21131 13413 21143 13447
rect 21192 13444 21220 13484
rect 21637 13447 21695 13453
rect 21637 13444 21649 13447
rect 21192 13416 21649 13444
rect 21085 13407 21143 13413
rect 21637 13413 21649 13416
rect 21683 13413 21695 13447
rect 21637 13407 21695 13413
rect 1765 13379 1823 13385
rect 1765 13345 1777 13379
rect 1811 13376 1823 13379
rect 1854 13376 1860 13388
rect 1811 13348 1860 13376
rect 1811 13345 1823 13348
rect 1765 13339 1823 13345
rect 1854 13336 1860 13348
rect 1912 13336 1918 13388
rect 2041 13379 2099 13385
rect 2041 13345 2053 13379
rect 2087 13376 2099 13379
rect 2498 13376 2504 13388
rect 2087 13348 2504 13376
rect 2087 13345 2099 13348
rect 2041 13339 2099 13345
rect 2498 13336 2504 13348
rect 2556 13336 2562 13388
rect 4154 13336 4160 13388
rect 4212 13376 4218 13388
rect 4614 13376 4620 13388
rect 4212 13348 4257 13376
rect 4575 13348 4620 13376
rect 4212 13336 4218 13348
rect 4614 13336 4620 13348
rect 4672 13336 4678 13388
rect 8478 13336 8484 13388
rect 8536 13376 8542 13388
rect 8608 13379 8666 13385
rect 8608 13376 8620 13379
rect 8536 13348 8620 13376
rect 8536 13336 8542 13348
rect 8608 13345 8620 13348
rect 8654 13345 8666 13379
rect 8608 13339 8666 13345
rect 8711 13379 8769 13385
rect 8711 13345 8723 13379
rect 8757 13376 8769 13379
rect 10502 13376 10508 13388
rect 8757 13348 10508 13376
rect 8757 13345 8769 13348
rect 8711 13339 8769 13345
rect 10502 13336 10508 13348
rect 10560 13336 10566 13388
rect 15562 13336 15568 13388
rect 15620 13376 15626 13388
rect 15692 13379 15750 13385
rect 15692 13376 15704 13379
rect 15620 13348 15704 13376
rect 15620 13336 15626 13348
rect 15692 13345 15704 13348
rect 15738 13345 15750 13379
rect 15692 13339 15750 13345
rect 5905 13311 5963 13317
rect 5905 13277 5917 13311
rect 5951 13277 5963 13311
rect 9674 13308 9680 13320
rect 9635 13280 9680 13308
rect 5905 13271 5963 13277
rect 2314 13200 2320 13252
rect 2372 13240 2378 13252
rect 2869 13243 2927 13249
rect 2869 13240 2881 13243
rect 2372 13212 2881 13240
rect 2372 13200 2378 13212
rect 2869 13209 2881 13212
rect 2915 13209 2927 13243
rect 2869 13203 2927 13209
rect 1854 13132 1860 13184
rect 1912 13172 1918 13184
rect 2501 13175 2559 13181
rect 2501 13172 2513 13175
rect 1912 13144 2513 13172
rect 1912 13132 1918 13144
rect 2501 13141 2513 13144
rect 2547 13141 2559 13175
rect 3786 13172 3792 13184
rect 3747 13144 3792 13172
rect 2501 13135 2559 13141
rect 3786 13132 3792 13144
rect 3844 13132 3850 13184
rect 5718 13172 5724 13184
rect 5679 13144 5724 13172
rect 5718 13132 5724 13144
rect 5776 13172 5782 13184
rect 5920 13172 5948 13271
rect 9674 13268 9680 13280
rect 9732 13268 9738 13320
rect 11606 13308 11612 13320
rect 11567 13280 11612 13308
rect 11606 13268 11612 13280
rect 11664 13268 11670 13320
rect 16761 13311 16819 13317
rect 16761 13277 16773 13311
rect 16807 13308 16819 13311
rect 16942 13308 16948 13320
rect 16807 13280 16948 13308
rect 16807 13277 16819 13280
rect 16761 13271 16819 13277
rect 16942 13268 16948 13280
rect 17000 13268 17006 13320
rect 17402 13308 17408 13320
rect 17315 13280 17408 13308
rect 17402 13268 17408 13280
rect 17460 13308 17466 13320
rect 18414 13308 18420 13320
rect 17460 13280 18420 13308
rect 17460 13268 17466 13280
rect 18414 13268 18420 13280
rect 18472 13268 18478 13320
rect 18601 13311 18659 13317
rect 18601 13277 18613 13311
rect 18647 13308 18659 13311
rect 18782 13308 18788 13320
rect 18647 13280 18788 13308
rect 18647 13277 18659 13280
rect 18601 13271 18659 13277
rect 18782 13268 18788 13280
rect 18840 13268 18846 13320
rect 20993 13311 21051 13317
rect 20993 13277 21005 13311
rect 21039 13277 21051 13311
rect 20993 13271 21051 13277
rect 15795 13243 15853 13249
rect 15795 13209 15807 13243
rect 15841 13240 15853 13243
rect 21008 13240 21036 13271
rect 21450 13240 21456 13252
rect 15841 13212 21456 13240
rect 15841 13209 15853 13212
rect 15795 13203 15853 13209
rect 21450 13200 21456 13212
rect 21508 13200 21514 13252
rect 5776 13144 5948 13172
rect 8205 13175 8263 13181
rect 5776 13132 5782 13144
rect 8205 13141 8217 13175
rect 8251 13172 8263 13175
rect 8294 13172 8300 13184
rect 8251 13144 8300 13172
rect 8251 13141 8263 13144
rect 8205 13135 8263 13141
rect 8294 13132 8300 13144
rect 8352 13172 8358 13184
rect 9125 13175 9183 13181
rect 9125 13172 9137 13175
rect 8352 13144 9137 13172
rect 8352 13132 8358 13144
rect 9125 13141 9137 13144
rect 9171 13172 9183 13175
rect 9398 13172 9404 13184
rect 9171 13144 9404 13172
rect 9171 13141 9183 13144
rect 9125 13135 9183 13141
rect 9398 13132 9404 13144
rect 9456 13132 9462 13184
rect 13449 13175 13507 13181
rect 13449 13141 13461 13175
rect 13495 13172 13507 13175
rect 13817 13175 13875 13181
rect 13817 13172 13829 13175
rect 13495 13144 13829 13172
rect 13495 13141 13507 13144
rect 13449 13135 13507 13141
rect 13817 13141 13829 13144
rect 13863 13172 13875 13175
rect 14090 13172 14096 13184
rect 13863 13144 14096 13172
rect 13863 13141 13875 13144
rect 13817 13135 13875 13141
rect 14090 13132 14096 13144
rect 14148 13172 14154 13184
rect 14734 13172 14740 13184
rect 14148 13144 14740 13172
rect 14148 13132 14154 13144
rect 14734 13132 14740 13144
rect 14792 13132 14798 13184
rect 16482 13172 16488 13184
rect 16395 13144 16488 13172
rect 16482 13132 16488 13144
rect 16540 13172 16546 13184
rect 17586 13172 17592 13184
rect 16540 13144 17592 13172
rect 16540 13132 16546 13144
rect 17586 13132 17592 13144
rect 17644 13132 17650 13184
rect 19426 13132 19432 13184
rect 19484 13172 19490 13184
rect 19981 13175 20039 13181
rect 19981 13172 19993 13175
rect 19484 13144 19993 13172
rect 19484 13132 19490 13144
rect 19981 13141 19993 13144
rect 20027 13172 20039 13175
rect 20070 13172 20076 13184
rect 20027 13144 20076 13172
rect 20027 13141 20039 13144
rect 19981 13135 20039 13141
rect 20070 13132 20076 13144
rect 20128 13132 20134 13184
rect 1104 13082 22816 13104
rect 1104 13030 4982 13082
rect 5034 13030 5046 13082
rect 5098 13030 5110 13082
rect 5162 13030 5174 13082
rect 5226 13030 12982 13082
rect 13034 13030 13046 13082
rect 13098 13030 13110 13082
rect 13162 13030 13174 13082
rect 13226 13030 20982 13082
rect 21034 13030 21046 13082
rect 21098 13030 21110 13082
rect 21162 13030 21174 13082
rect 21226 13030 22816 13082
rect 1104 13008 22816 13030
rect 3142 12968 3148 12980
rect 3055 12940 3148 12968
rect 3142 12928 3148 12940
rect 3200 12968 3206 12980
rect 4154 12968 4160 12980
rect 3200 12940 4160 12968
rect 3200 12928 3206 12940
rect 4126 12928 4160 12940
rect 4212 12928 4218 12980
rect 5767 12971 5825 12977
rect 5767 12937 5779 12971
rect 5813 12968 5825 12971
rect 5902 12968 5908 12980
rect 5813 12940 5908 12968
rect 5813 12937 5825 12940
rect 5767 12931 5825 12937
rect 5902 12928 5908 12940
rect 5960 12928 5966 12980
rect 8205 12971 8263 12977
rect 8205 12968 8217 12971
rect 6282 12940 8217 12968
rect 14 12860 20 12912
rect 72 12900 78 12912
rect 1765 12903 1823 12909
rect 1765 12900 1777 12903
rect 72 12872 1777 12900
rect 72 12860 78 12872
rect 1765 12869 1777 12872
rect 1811 12900 1823 12903
rect 1854 12900 1860 12912
rect 1811 12872 1860 12900
rect 1811 12869 1823 12872
rect 1765 12863 1823 12869
rect 1854 12860 1860 12872
rect 1912 12860 1918 12912
rect 4126 12900 4154 12928
rect 4890 12900 4896 12912
rect 4126 12872 4896 12900
rect 4890 12860 4896 12872
rect 4948 12860 4954 12912
rect 5626 12860 5632 12912
rect 5684 12900 5690 12912
rect 6282 12900 6310 12940
rect 8205 12937 8217 12940
rect 8251 12937 8263 12971
rect 8205 12931 8263 12937
rect 6546 12900 6552 12912
rect 5684 12872 6310 12900
rect 6507 12872 6552 12900
rect 5684 12860 5690 12872
rect 6546 12860 6552 12872
rect 6604 12860 6610 12912
rect 6822 12860 6828 12912
rect 6880 12900 6886 12912
rect 7469 12903 7527 12909
rect 7469 12900 7481 12903
rect 6880 12872 7481 12900
rect 6880 12860 6886 12872
rect 7469 12869 7481 12872
rect 7515 12869 7527 12903
rect 7469 12863 7527 12869
rect 4522 12832 4528 12844
rect 4435 12804 4528 12832
rect 4522 12792 4528 12804
rect 4580 12832 4586 12844
rect 5350 12832 5356 12844
rect 4580 12804 5356 12832
rect 4580 12792 4586 12804
rect 5350 12792 5356 12804
rect 5408 12792 5414 12844
rect 6730 12792 6736 12844
rect 6788 12832 6794 12844
rect 6917 12835 6975 12841
rect 6917 12832 6929 12835
rect 6788 12804 6929 12832
rect 6788 12792 6794 12804
rect 6917 12801 6929 12804
rect 6963 12832 6975 12835
rect 7837 12835 7895 12841
rect 7837 12832 7849 12835
rect 6963 12804 7849 12832
rect 6963 12801 6975 12804
rect 6917 12795 6975 12801
rect 7837 12801 7849 12804
rect 7883 12801 7895 12835
rect 7837 12795 7895 12801
rect 1670 12764 1676 12776
rect 1631 12736 1676 12764
rect 1670 12724 1676 12736
rect 1728 12724 1734 12776
rect 1949 12767 2007 12773
rect 1949 12733 1961 12767
rect 1995 12764 2007 12767
rect 2314 12764 2320 12776
rect 1995 12736 2320 12764
rect 1995 12733 2007 12736
rect 1949 12727 2007 12733
rect 2314 12724 2320 12736
rect 2372 12724 2378 12776
rect 3786 12764 3792 12776
rect 3747 12736 3792 12764
rect 3786 12724 3792 12736
rect 3844 12724 3850 12776
rect 3881 12767 3939 12773
rect 3881 12733 3893 12767
rect 3927 12764 3939 12767
rect 3970 12764 3976 12776
rect 3927 12736 3976 12764
rect 3927 12733 3939 12736
rect 3881 12727 3939 12733
rect 3970 12724 3976 12736
rect 4028 12724 4034 12776
rect 4065 12767 4123 12773
rect 4065 12733 4077 12767
rect 4111 12733 4123 12767
rect 4065 12727 4123 12733
rect 5696 12767 5754 12773
rect 5696 12733 5708 12767
rect 5742 12764 5754 12767
rect 8220 12764 8248 12931
rect 8478 12928 8484 12980
rect 8536 12968 8542 12980
rect 8573 12971 8631 12977
rect 8573 12968 8585 12971
rect 8536 12940 8585 12968
rect 8536 12928 8542 12940
rect 8573 12937 8585 12940
rect 8619 12968 8631 12971
rect 8754 12968 8760 12980
rect 8619 12940 8760 12968
rect 8619 12937 8631 12940
rect 8573 12931 8631 12937
rect 8754 12928 8760 12940
rect 8812 12928 8818 12980
rect 10594 12968 10600 12980
rect 10555 12940 10600 12968
rect 10594 12928 10600 12940
rect 10652 12928 10658 12980
rect 11606 12928 11612 12980
rect 11664 12968 11670 12980
rect 12161 12971 12219 12977
rect 12161 12968 12173 12971
rect 11664 12940 12173 12968
rect 11664 12928 11670 12940
rect 12161 12937 12173 12940
rect 12207 12968 12219 12971
rect 12575 12971 12633 12977
rect 12575 12968 12587 12971
rect 12207 12940 12587 12968
rect 12207 12937 12219 12940
rect 12161 12931 12219 12937
rect 12575 12937 12587 12940
rect 12621 12937 12633 12971
rect 12575 12931 12633 12937
rect 13449 12971 13507 12977
rect 13449 12937 13461 12971
rect 13495 12968 13507 12971
rect 13538 12968 13544 12980
rect 13495 12940 13544 12968
rect 13495 12937 13507 12940
rect 13449 12931 13507 12937
rect 13538 12928 13544 12940
rect 13596 12928 13602 12980
rect 16761 12971 16819 12977
rect 16761 12937 16773 12971
rect 16807 12968 16819 12971
rect 16850 12968 16856 12980
rect 16807 12940 16856 12968
rect 16807 12937 16819 12940
rect 16761 12931 16819 12937
rect 16850 12928 16856 12940
rect 16908 12928 16914 12980
rect 16942 12928 16948 12980
rect 17000 12968 17006 12980
rect 17405 12971 17463 12977
rect 17405 12968 17417 12971
rect 17000 12940 17417 12968
rect 17000 12928 17006 12940
rect 17405 12937 17417 12940
rect 17451 12968 17463 12971
rect 18874 12968 18880 12980
rect 17451 12940 18880 12968
rect 17451 12937 17463 12940
rect 17405 12931 17463 12937
rect 18874 12928 18880 12940
rect 18932 12928 18938 12980
rect 19521 12971 19579 12977
rect 19521 12937 19533 12971
rect 19567 12968 19579 12971
rect 20806 12968 20812 12980
rect 19567 12940 20812 12968
rect 19567 12937 19579 12940
rect 19521 12931 19579 12937
rect 11790 12900 11796 12912
rect 11751 12872 11796 12900
rect 11790 12860 11796 12872
rect 11848 12860 11854 12912
rect 16025 12903 16083 12909
rect 16025 12869 16037 12903
rect 16071 12900 16083 12903
rect 17773 12903 17831 12909
rect 17773 12900 17785 12903
rect 16071 12872 17785 12900
rect 16071 12869 16083 12872
rect 16025 12863 16083 12869
rect 17773 12869 17785 12872
rect 17819 12900 17831 12903
rect 18230 12900 18236 12912
rect 17819 12872 18236 12900
rect 17819 12869 17831 12872
rect 17773 12863 17831 12869
rect 18230 12860 18236 12872
rect 18288 12860 18294 12912
rect 9585 12835 9643 12841
rect 9585 12801 9597 12835
rect 9631 12832 9643 12835
rect 9674 12832 9680 12844
rect 9631 12804 9680 12832
rect 9631 12801 9643 12804
rect 9585 12795 9643 12801
rect 9674 12792 9680 12804
rect 9732 12832 9738 12844
rect 10229 12835 10287 12841
rect 10229 12832 10241 12835
rect 9732 12804 10241 12832
rect 9732 12792 9738 12804
rect 10229 12801 10241 12804
rect 10275 12801 10287 12835
rect 11514 12832 11520 12844
rect 11475 12804 11520 12832
rect 10229 12795 10287 12801
rect 11514 12792 11520 12804
rect 11572 12792 11578 12844
rect 18138 12832 18144 12844
rect 18099 12804 18144 12832
rect 18138 12792 18144 12804
rect 18196 12792 18202 12844
rect 18414 12832 18420 12844
rect 18375 12804 18420 12832
rect 18414 12792 18420 12804
rect 18472 12792 18478 12844
rect 8849 12767 8907 12773
rect 8849 12764 8861 12767
rect 5742 12736 6040 12764
rect 8220 12736 8861 12764
rect 5742 12733 5754 12736
rect 5696 12727 5754 12733
rect 2409 12699 2467 12705
rect 2409 12665 2421 12699
rect 2455 12696 2467 12699
rect 3510 12696 3516 12708
rect 2455 12668 3516 12696
rect 2455 12665 2467 12668
rect 2409 12659 2467 12665
rect 3510 12656 3516 12668
rect 3568 12656 3574 12708
rect 4080 12640 4108 12727
rect 4614 12656 4620 12708
rect 4672 12696 4678 12708
rect 4672 12668 5304 12696
rect 4672 12656 4678 12668
rect 2682 12628 2688 12640
rect 2643 12600 2688 12628
rect 2682 12588 2688 12600
rect 2740 12588 2746 12640
rect 3694 12628 3700 12640
rect 3607 12600 3700 12628
rect 3694 12588 3700 12600
rect 3752 12628 3758 12640
rect 4062 12628 4068 12640
rect 3752 12600 4068 12628
rect 3752 12588 3758 12600
rect 4062 12588 4068 12600
rect 4120 12588 4126 12640
rect 4890 12628 4896 12640
rect 4851 12600 4896 12628
rect 4890 12588 4896 12600
rect 4948 12588 4954 12640
rect 5276 12637 5304 12668
rect 6012 12640 6040 12736
rect 8849 12733 8861 12736
rect 8895 12733 8907 12767
rect 9398 12764 9404 12776
rect 9359 12736 9404 12764
rect 8849 12727 8907 12733
rect 7006 12656 7012 12708
rect 7064 12696 7070 12708
rect 8864 12696 8892 12727
rect 9398 12724 9404 12736
rect 9456 12724 9462 12776
rect 12504 12767 12562 12773
rect 12504 12733 12516 12767
rect 12550 12764 12562 12767
rect 12989 12767 13047 12773
rect 12989 12764 13001 12767
rect 12550 12736 13001 12764
rect 12550 12733 12562 12736
rect 12504 12727 12562 12733
rect 12989 12733 13001 12736
rect 13035 12764 13047 12767
rect 13354 12764 13360 12776
rect 13035 12736 13360 12764
rect 13035 12733 13047 12736
rect 12989 12727 13047 12733
rect 13354 12724 13360 12736
rect 13412 12724 13418 12776
rect 13538 12764 13544 12776
rect 13499 12736 13544 12764
rect 13538 12724 13544 12736
rect 13596 12724 13602 12776
rect 14090 12764 14096 12776
rect 14051 12736 14096 12764
rect 14090 12724 14096 12736
rect 14148 12724 14154 12776
rect 14277 12767 14335 12773
rect 14277 12733 14289 12767
rect 14323 12764 14335 12767
rect 14645 12767 14703 12773
rect 14645 12764 14657 12767
rect 14323 12736 14657 12764
rect 14323 12733 14335 12736
rect 14277 12727 14335 12733
rect 14645 12733 14657 12736
rect 14691 12764 14703 12767
rect 15105 12767 15163 12773
rect 15105 12764 15117 12767
rect 14691 12736 15117 12764
rect 14691 12733 14703 12736
rect 14645 12727 14703 12733
rect 15105 12733 15117 12736
rect 15151 12733 15163 12767
rect 15105 12727 15163 12733
rect 16920 12767 16978 12773
rect 16920 12733 16932 12767
rect 16966 12764 16978 12767
rect 17402 12764 17408 12776
rect 16966 12736 17408 12764
rect 16966 12733 16978 12736
rect 16920 12727 16978 12733
rect 17402 12724 17408 12736
rect 17460 12724 17466 12776
rect 19058 12724 19064 12776
rect 19116 12764 19122 12776
rect 19153 12767 19211 12773
rect 19153 12764 19165 12767
rect 19116 12736 19165 12764
rect 19116 12724 19122 12736
rect 19153 12733 19165 12736
rect 19199 12764 19211 12767
rect 19536 12764 19564 12931
rect 20806 12928 20812 12940
rect 20864 12968 20870 12980
rect 20901 12971 20959 12977
rect 20901 12968 20913 12971
rect 20864 12940 20913 12968
rect 20864 12928 20870 12940
rect 20901 12937 20913 12940
rect 20947 12937 20959 12971
rect 20901 12931 20959 12937
rect 21450 12928 21456 12980
rect 21508 12968 21514 12980
rect 22097 12971 22155 12977
rect 22097 12968 22109 12971
rect 21508 12940 22109 12968
rect 21508 12928 21514 12940
rect 22097 12937 22109 12940
rect 22143 12937 22155 12971
rect 22097 12931 22155 12937
rect 20254 12900 20260 12912
rect 20215 12872 20260 12900
rect 20254 12860 20260 12872
rect 20312 12860 20318 12912
rect 21358 12900 21364 12912
rect 21319 12872 21364 12900
rect 21358 12860 21364 12872
rect 21416 12860 21422 12912
rect 19705 12835 19763 12841
rect 19705 12801 19717 12835
rect 19751 12832 19763 12835
rect 20438 12832 20444 12844
rect 19751 12804 20444 12832
rect 19751 12801 19763 12804
rect 19705 12795 19763 12801
rect 20438 12792 20444 12804
rect 20496 12792 20502 12844
rect 19199 12736 19564 12764
rect 19199 12733 19211 12736
rect 19153 12727 19211 12733
rect 10502 12696 10508 12708
rect 7064 12668 7109 12696
rect 8864 12668 10508 12696
rect 7064 12656 7070 12668
rect 10502 12656 10508 12668
rect 10560 12656 10566 12708
rect 10870 12696 10876 12708
rect 10831 12668 10876 12696
rect 10870 12656 10876 12668
rect 10928 12656 10934 12708
rect 10965 12699 11023 12705
rect 10965 12665 10977 12699
rect 11011 12665 11023 12699
rect 10965 12659 11023 12665
rect 15013 12699 15071 12705
rect 15013 12665 15025 12699
rect 15059 12696 15071 12699
rect 15286 12696 15292 12708
rect 15059 12668 15292 12696
rect 15059 12665 15071 12668
rect 15013 12659 15071 12665
rect 5261 12631 5319 12637
rect 5261 12597 5273 12631
rect 5307 12628 5319 12631
rect 5810 12628 5816 12640
rect 5307 12600 5816 12628
rect 5307 12597 5319 12600
rect 5261 12591 5319 12597
rect 5810 12588 5816 12600
rect 5868 12588 5874 12640
rect 5994 12588 6000 12640
rect 6052 12628 6058 12640
rect 6089 12631 6147 12637
rect 6089 12628 6101 12631
rect 6052 12600 6101 12628
rect 6052 12588 6058 12600
rect 6089 12597 6101 12600
rect 6135 12597 6147 12631
rect 6089 12591 6147 12597
rect 9953 12631 10011 12637
rect 9953 12597 9965 12631
rect 9999 12628 10011 12631
rect 10226 12628 10232 12640
rect 9999 12600 10232 12628
rect 9999 12597 10011 12600
rect 9953 12591 10011 12597
rect 10226 12588 10232 12600
rect 10284 12628 10290 12640
rect 10410 12628 10416 12640
rect 10284 12600 10416 12628
rect 10284 12588 10290 12600
rect 10410 12588 10416 12600
rect 10468 12588 10474 12640
rect 10594 12588 10600 12640
rect 10652 12628 10658 12640
rect 10980 12628 11008 12659
rect 15286 12656 15292 12668
rect 15344 12696 15350 12708
rect 15467 12699 15525 12705
rect 15467 12696 15479 12699
rect 15344 12668 15479 12696
rect 15344 12656 15350 12668
rect 15467 12665 15479 12668
rect 15513 12696 15525 12699
rect 16022 12696 16028 12708
rect 15513 12668 16028 12696
rect 15513 12665 15525 12668
rect 15467 12659 15525 12665
rect 16022 12656 16028 12668
rect 16080 12656 16086 12708
rect 18230 12656 18236 12708
rect 18288 12696 18294 12708
rect 19536 12696 19564 12736
rect 20806 12724 20812 12776
rect 20864 12764 20870 12776
rect 21177 12767 21235 12773
rect 21177 12764 21189 12767
rect 20864 12736 21189 12764
rect 20864 12724 20870 12736
rect 21177 12733 21189 12736
rect 21223 12764 21235 12767
rect 21729 12767 21787 12773
rect 21729 12764 21741 12767
rect 21223 12736 21741 12764
rect 21223 12733 21235 12736
rect 21177 12727 21235 12733
rect 21729 12733 21741 12736
rect 21775 12733 21787 12767
rect 21729 12727 21787 12733
rect 19797 12699 19855 12705
rect 19797 12696 19809 12699
rect 18288 12668 18333 12696
rect 19536 12668 19809 12696
rect 18288 12656 18294 12668
rect 19797 12665 19809 12668
rect 19843 12665 19855 12699
rect 19797 12659 19855 12665
rect 10652 12600 11008 12628
rect 10652 12588 10658 12600
rect 15562 12588 15568 12640
rect 15620 12628 15626 12640
rect 16301 12631 16359 12637
rect 16301 12628 16313 12631
rect 15620 12600 16313 12628
rect 15620 12588 15626 12600
rect 16301 12597 16313 12600
rect 16347 12597 16359 12631
rect 16301 12591 16359 12597
rect 16758 12588 16764 12640
rect 16816 12628 16822 12640
rect 16991 12631 17049 12637
rect 16991 12628 17003 12631
rect 16816 12600 17003 12628
rect 16816 12588 16822 12600
rect 16991 12597 17003 12600
rect 17037 12597 17049 12631
rect 16991 12591 17049 12597
rect 1104 12538 22816 12560
rect 1104 12486 8982 12538
rect 9034 12486 9046 12538
rect 9098 12486 9110 12538
rect 9162 12486 9174 12538
rect 9226 12486 16982 12538
rect 17034 12486 17046 12538
rect 17098 12486 17110 12538
rect 17162 12486 17174 12538
rect 17226 12486 22816 12538
rect 1104 12464 22816 12486
rect 1854 12384 1860 12436
rect 1912 12424 1918 12436
rect 3789 12427 3847 12433
rect 3789 12424 3801 12427
rect 1912 12396 3801 12424
rect 1912 12384 1918 12396
rect 3789 12393 3801 12396
rect 3835 12424 3847 12427
rect 3970 12424 3976 12436
rect 3835 12396 3976 12424
rect 3835 12393 3847 12396
rect 3789 12387 3847 12393
rect 3970 12384 3976 12396
rect 4028 12424 4034 12436
rect 4154 12424 4160 12436
rect 4028 12396 4160 12424
rect 4028 12384 4034 12396
rect 4154 12384 4160 12396
rect 4212 12384 4218 12436
rect 5718 12424 5724 12436
rect 5679 12396 5724 12424
rect 5718 12384 5724 12396
rect 5776 12384 5782 12436
rect 8113 12427 8171 12433
rect 8113 12424 8125 12427
rect 5920 12396 8125 12424
rect 1670 12316 1676 12368
rect 1728 12356 1734 12368
rect 2682 12356 2688 12368
rect 1728 12328 2688 12356
rect 1728 12316 1734 12328
rect 1780 12297 1808 12328
rect 2682 12316 2688 12328
rect 2740 12316 2746 12368
rect 2869 12359 2927 12365
rect 2869 12325 2881 12359
rect 2915 12356 2927 12359
rect 5626 12356 5632 12368
rect 2915 12328 5632 12356
rect 2915 12325 2927 12328
rect 2869 12319 2927 12325
rect 1765 12291 1823 12297
rect 1765 12257 1777 12291
rect 1811 12257 1823 12291
rect 1765 12251 1823 12257
rect 1854 12248 1860 12300
rect 1912 12288 1918 12300
rect 2038 12288 2044 12300
rect 1912 12260 1957 12288
rect 1999 12260 2044 12288
rect 1912 12248 1918 12260
rect 2038 12248 2044 12260
rect 2096 12248 2102 12300
rect 2498 12288 2504 12300
rect 2411 12260 2504 12288
rect 2498 12248 2504 12260
rect 2556 12288 2562 12300
rect 2884 12288 2912 12319
rect 5626 12316 5632 12328
rect 5684 12316 5690 12368
rect 4154 12288 4160 12300
rect 2556 12260 2912 12288
rect 4115 12260 4160 12288
rect 2556 12248 2562 12260
rect 4154 12248 4160 12260
rect 4212 12248 4218 12300
rect 4890 12248 4896 12300
rect 4948 12288 4954 12300
rect 5718 12288 5724 12300
rect 4948 12260 5724 12288
rect 4948 12248 4954 12260
rect 5718 12248 5724 12260
rect 5776 12288 5782 12300
rect 5920 12297 5948 12396
rect 8113 12393 8125 12396
rect 8159 12393 8171 12427
rect 8113 12387 8171 12393
rect 10275 12427 10333 12433
rect 10275 12393 10287 12427
rect 10321 12424 10333 12427
rect 10870 12424 10876 12436
rect 10321 12396 10876 12424
rect 10321 12393 10333 12396
rect 10275 12387 10333 12393
rect 10870 12384 10876 12396
rect 10928 12384 10934 12436
rect 16301 12427 16359 12433
rect 16301 12393 16313 12427
rect 16347 12424 16359 12427
rect 16850 12424 16856 12436
rect 16347 12396 16856 12424
rect 16347 12393 16359 12396
rect 16301 12387 16359 12393
rect 16850 12384 16856 12396
rect 16908 12384 16914 12436
rect 17037 12427 17095 12433
rect 17037 12393 17049 12427
rect 17083 12424 17095 12427
rect 17402 12424 17408 12436
rect 17083 12396 17408 12424
rect 17083 12393 17095 12396
rect 17037 12387 17095 12393
rect 17402 12384 17408 12396
rect 17460 12384 17466 12436
rect 18782 12424 18788 12436
rect 18743 12396 18788 12424
rect 18782 12384 18788 12396
rect 18840 12384 18846 12436
rect 20349 12427 20407 12433
rect 20349 12393 20361 12427
rect 20395 12424 20407 12427
rect 20438 12424 20444 12436
rect 20395 12396 20444 12424
rect 20395 12393 20407 12396
rect 20349 12387 20407 12393
rect 20438 12384 20444 12396
rect 20496 12384 20502 12436
rect 12434 12316 12440 12368
rect 12492 12356 12498 12368
rect 12802 12356 12808 12368
rect 12492 12328 12808 12356
rect 12492 12316 12498 12328
rect 12802 12316 12808 12328
rect 12860 12316 12866 12368
rect 15743 12359 15801 12365
rect 15743 12325 15755 12359
rect 15789 12356 15801 12359
rect 16022 12356 16028 12368
rect 15789 12328 16028 12356
rect 15789 12325 15801 12328
rect 15743 12319 15801 12325
rect 16022 12316 16028 12328
rect 16080 12316 16086 12368
rect 17951 12359 18009 12365
rect 17951 12325 17963 12359
rect 17997 12356 18009 12359
rect 18138 12356 18144 12368
rect 17997 12328 18144 12356
rect 17997 12325 18009 12328
rect 17951 12319 18009 12325
rect 18138 12316 18144 12328
rect 18196 12316 18202 12368
rect 20714 12316 20720 12368
rect 20772 12356 20778 12368
rect 20993 12359 21051 12365
rect 20993 12356 21005 12359
rect 20772 12328 21005 12356
rect 20772 12316 20778 12328
rect 20993 12325 21005 12328
rect 21039 12325 21051 12359
rect 20993 12319 21051 12325
rect 21085 12359 21143 12365
rect 21085 12325 21097 12359
rect 21131 12356 21143 12359
rect 21266 12356 21272 12368
rect 21131 12328 21272 12356
rect 21131 12325 21143 12328
rect 21085 12319 21143 12325
rect 21266 12316 21272 12328
rect 21324 12316 21330 12368
rect 5905 12291 5963 12297
rect 5905 12288 5917 12291
rect 5776 12260 5917 12288
rect 5776 12248 5782 12260
rect 5905 12257 5917 12260
rect 5951 12257 5963 12291
rect 6178 12288 6184 12300
rect 6139 12260 6184 12288
rect 5905 12251 5963 12257
rect 6178 12248 6184 12260
rect 6236 12248 6242 12300
rect 6917 12291 6975 12297
rect 6917 12257 6929 12291
rect 6963 12288 6975 12291
rect 7282 12288 7288 12300
rect 6963 12260 7288 12288
rect 6963 12257 6975 12260
rect 6917 12251 6975 12257
rect 7282 12248 7288 12260
rect 7340 12248 7346 12300
rect 7653 12291 7711 12297
rect 7653 12257 7665 12291
rect 7699 12288 7711 12291
rect 7834 12288 7840 12300
rect 7699 12260 7840 12288
rect 7699 12257 7711 12260
rect 7653 12251 7711 12257
rect 7834 12248 7840 12260
rect 7892 12248 7898 12300
rect 7929 12291 7987 12297
rect 7929 12257 7941 12291
rect 7975 12288 7987 12291
rect 8018 12288 8024 12300
rect 7975 12260 8024 12288
rect 7975 12257 7987 12260
rect 7929 12251 7987 12257
rect 8018 12248 8024 12260
rect 8076 12248 8082 12300
rect 10204 12291 10262 12297
rect 10204 12257 10216 12291
rect 10250 12288 10262 12291
rect 10594 12288 10600 12300
rect 10250 12260 10600 12288
rect 10250 12257 10262 12260
rect 10204 12251 10262 12257
rect 10594 12248 10600 12260
rect 10652 12248 10658 12300
rect 11882 12288 11888 12300
rect 11843 12260 11888 12288
rect 11882 12248 11888 12260
rect 11940 12248 11946 12300
rect 12066 12288 12072 12300
rect 12027 12260 12072 12288
rect 12066 12248 12072 12260
rect 12124 12248 12130 12300
rect 13630 12288 13636 12300
rect 13591 12260 13636 12288
rect 13630 12248 13636 12260
rect 13688 12248 13694 12300
rect 14090 12248 14096 12300
rect 14148 12288 14154 12300
rect 14185 12291 14243 12297
rect 14185 12288 14197 12291
rect 14148 12260 14197 12288
rect 14148 12248 14154 12260
rect 14185 12257 14197 12260
rect 14231 12288 14243 12291
rect 14458 12288 14464 12300
rect 14231 12260 14464 12288
rect 14231 12257 14243 12260
rect 14185 12251 14243 12257
rect 14458 12248 14464 12260
rect 14516 12248 14522 12300
rect 18509 12291 18567 12297
rect 18509 12257 18521 12291
rect 18555 12288 18567 12291
rect 19058 12288 19064 12300
rect 18555 12260 19064 12288
rect 18555 12257 18567 12260
rect 18509 12251 18567 12257
rect 19058 12248 19064 12260
rect 19116 12248 19122 12300
rect 19334 12248 19340 12300
rect 19392 12288 19398 12300
rect 19702 12288 19708 12300
rect 19392 12260 19708 12288
rect 19392 12248 19398 12260
rect 19702 12248 19708 12260
rect 19760 12248 19766 12300
rect 1673 12223 1731 12229
rect 1673 12189 1685 12223
rect 1719 12220 1731 12223
rect 2056 12220 2084 12248
rect 1719 12192 2084 12220
rect 1719 12189 1731 12192
rect 1673 12183 1731 12189
rect 3970 12180 3976 12232
rect 4028 12220 4034 12232
rect 4801 12223 4859 12229
rect 4801 12220 4813 12223
rect 4028 12192 4813 12220
rect 4028 12180 4034 12192
rect 4801 12189 4813 12192
rect 4847 12220 4859 12223
rect 12158 12220 12164 12232
rect 4847 12192 6960 12220
rect 12119 12192 12164 12220
rect 4847 12189 4859 12192
rect 4801 12183 4859 12189
rect 6932 12096 6960 12192
rect 12158 12180 12164 12192
rect 12216 12180 12222 12232
rect 12713 12223 12771 12229
rect 12713 12189 12725 12223
rect 12759 12220 12771 12223
rect 12802 12220 12808 12232
rect 12759 12192 12808 12220
rect 12759 12189 12771 12192
rect 12713 12183 12771 12189
rect 12802 12180 12808 12192
rect 12860 12180 12866 12232
rect 14369 12223 14427 12229
rect 14369 12189 14381 12223
rect 14415 12220 14427 12223
rect 15381 12223 15439 12229
rect 15381 12220 15393 12223
rect 14415 12192 15393 12220
rect 14415 12189 14427 12192
rect 14369 12183 14427 12189
rect 15381 12189 15393 12192
rect 15427 12220 15439 12223
rect 15746 12220 15752 12232
rect 15427 12192 15752 12220
rect 15427 12189 15439 12192
rect 15381 12183 15439 12189
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 16942 12180 16948 12232
rect 17000 12220 17006 12232
rect 17589 12223 17647 12229
rect 17589 12220 17601 12223
rect 17000 12192 17601 12220
rect 17000 12180 17006 12192
rect 17589 12189 17601 12192
rect 17635 12189 17647 12223
rect 21634 12220 21640 12232
rect 21595 12192 21640 12220
rect 17589 12183 17647 12189
rect 21634 12180 21640 12192
rect 21692 12180 21698 12232
rect 7745 12155 7803 12161
rect 7745 12121 7757 12155
rect 7791 12152 7803 12155
rect 8202 12152 8208 12164
rect 7791 12124 8208 12152
rect 7791 12121 7803 12124
rect 7745 12115 7803 12121
rect 8202 12112 8208 12124
rect 8260 12152 8266 12164
rect 8757 12155 8815 12161
rect 8757 12152 8769 12155
rect 8260 12124 8769 12152
rect 8260 12112 8266 12124
rect 8757 12121 8769 12124
rect 8803 12121 8815 12155
rect 19886 12152 19892 12164
rect 19847 12124 19892 12152
rect 8757 12115 8815 12121
rect 19886 12112 19892 12124
rect 19944 12112 19950 12164
rect 6914 12044 6920 12096
rect 6972 12084 6978 12096
rect 7193 12087 7251 12093
rect 7193 12084 7205 12087
rect 6972 12056 7205 12084
rect 6972 12044 6978 12056
rect 7193 12053 7205 12056
rect 7239 12053 7251 12087
rect 9122 12084 9128 12096
rect 9083 12056 9128 12084
rect 7193 12047 7251 12053
rect 9122 12044 9128 12056
rect 9180 12044 9186 12096
rect 12710 12044 12716 12096
rect 12768 12084 12774 12096
rect 12989 12087 13047 12093
rect 12989 12084 13001 12087
rect 12768 12056 13001 12084
rect 12768 12044 12774 12056
rect 12989 12053 13001 12056
rect 13035 12053 13047 12087
rect 12989 12047 13047 12053
rect 16482 12044 16488 12096
rect 16540 12084 16546 12096
rect 16577 12087 16635 12093
rect 16577 12084 16589 12087
rect 16540 12056 16589 12084
rect 16540 12044 16546 12056
rect 16577 12053 16589 12056
rect 16623 12053 16635 12087
rect 16577 12047 16635 12053
rect 19978 12044 19984 12096
rect 20036 12084 20042 12096
rect 23566 12084 23572 12096
rect 20036 12056 23572 12084
rect 20036 12044 20042 12056
rect 23566 12044 23572 12056
rect 23624 12044 23630 12096
rect 1104 11994 22816 12016
rect 1104 11942 4982 11994
rect 5034 11942 5046 11994
rect 5098 11942 5110 11994
rect 5162 11942 5174 11994
rect 5226 11942 12982 11994
rect 13034 11942 13046 11994
rect 13098 11942 13110 11994
rect 13162 11942 13174 11994
rect 13226 11942 20982 11994
rect 21034 11942 21046 11994
rect 21098 11942 21110 11994
rect 21162 11942 21174 11994
rect 21226 11942 22816 11994
rect 1104 11920 22816 11942
rect 3053 11883 3111 11889
rect 3053 11849 3065 11883
rect 3099 11880 3111 11883
rect 3694 11880 3700 11892
rect 3099 11852 3700 11880
rect 3099 11849 3111 11852
rect 3053 11843 3111 11849
rect 3068 11812 3096 11843
rect 3694 11840 3700 11852
rect 3752 11840 3758 11892
rect 4246 11840 4252 11892
rect 4304 11880 4310 11892
rect 4893 11883 4951 11889
rect 4893 11880 4905 11883
rect 4304 11852 4905 11880
rect 4304 11840 4310 11852
rect 4893 11849 4905 11852
rect 4939 11849 4951 11883
rect 5718 11880 5724 11892
rect 5679 11852 5724 11880
rect 4893 11843 4951 11849
rect 5718 11840 5724 11852
rect 5776 11840 5782 11892
rect 5810 11840 5816 11892
rect 5868 11880 5874 11892
rect 5868 11852 7604 11880
rect 5868 11840 5874 11852
rect 2516 11784 3096 11812
rect 3421 11815 3479 11821
rect 2038 11636 2044 11688
rect 2096 11676 2102 11688
rect 2225 11679 2283 11685
rect 2225 11676 2237 11679
rect 2096 11648 2237 11676
rect 2096 11636 2102 11648
rect 2225 11645 2237 11648
rect 2271 11676 2283 11679
rect 2516 11676 2544 11784
rect 3421 11781 3433 11815
rect 3467 11812 3479 11815
rect 3970 11812 3976 11824
rect 3467 11784 3976 11812
rect 3467 11781 3479 11784
rect 3421 11775 3479 11781
rect 3970 11772 3976 11784
rect 4028 11772 4034 11824
rect 4154 11772 4160 11824
rect 4212 11812 4218 11824
rect 6178 11812 6184 11824
rect 4212 11784 6184 11812
rect 4212 11772 4218 11784
rect 6178 11772 6184 11784
rect 6236 11772 6242 11824
rect 6914 11812 6920 11824
rect 6875 11784 6920 11812
rect 6914 11772 6920 11784
rect 6972 11772 6978 11824
rect 2682 11744 2688 11756
rect 2595 11716 2688 11744
rect 2682 11704 2688 11716
rect 2740 11744 2746 11756
rect 2740 11716 4016 11744
rect 2740 11704 2746 11716
rect 2271 11648 2544 11676
rect 2271 11645 2283 11648
rect 2225 11639 2283 11645
rect 3694 11636 3700 11688
rect 3752 11676 3758 11688
rect 3881 11679 3939 11685
rect 3881 11676 3893 11679
rect 3752 11648 3893 11676
rect 3752 11636 3758 11648
rect 3881 11645 3893 11648
rect 3927 11645 3939 11679
rect 3881 11639 3939 11645
rect 2314 11608 2320 11620
rect 2275 11580 2320 11608
rect 2314 11568 2320 11580
rect 2372 11568 2378 11620
rect 3988 11608 4016 11716
rect 4062 11704 4068 11756
rect 4120 11744 4126 11756
rect 4120 11716 7144 11744
rect 4120 11704 4126 11716
rect 4172 11685 4200 11716
rect 4157 11679 4215 11685
rect 4157 11645 4169 11679
rect 4203 11645 4215 11679
rect 6549 11679 6607 11685
rect 6549 11676 6561 11679
rect 4157 11639 4215 11645
rect 4448 11648 6561 11676
rect 4448 11608 4476 11648
rect 6549 11645 6561 11648
rect 6595 11676 6607 11679
rect 6822 11676 6828 11688
rect 6595 11648 6828 11676
rect 6595 11645 6607 11648
rect 6549 11639 6607 11645
rect 6822 11636 6828 11648
rect 6880 11636 6886 11688
rect 7116 11685 7144 11716
rect 7101 11679 7159 11685
rect 7101 11645 7113 11679
rect 7147 11676 7159 11679
rect 7282 11676 7288 11688
rect 7147 11648 7288 11676
rect 7147 11645 7159 11648
rect 7101 11639 7159 11645
rect 7282 11636 7288 11648
rect 7340 11636 7346 11688
rect 7576 11685 7604 11852
rect 11882 11840 11888 11892
rect 11940 11880 11946 11892
rect 12161 11883 12219 11889
rect 12161 11880 12173 11883
rect 11940 11852 12173 11880
rect 11940 11840 11946 11852
rect 12161 11849 12173 11852
rect 12207 11849 12219 11883
rect 13630 11880 13636 11892
rect 13591 11852 13636 11880
rect 12161 11843 12219 11849
rect 13630 11840 13636 11852
rect 13688 11840 13694 11892
rect 15746 11880 15752 11892
rect 15707 11852 15752 11880
rect 15746 11840 15752 11852
rect 15804 11840 15810 11892
rect 19702 11880 19708 11892
rect 19663 11852 19708 11880
rect 19702 11840 19708 11852
rect 19760 11840 19766 11892
rect 20714 11840 20720 11892
rect 20772 11880 20778 11892
rect 21361 11883 21419 11889
rect 21361 11880 21373 11883
rect 20772 11852 21373 11880
rect 20772 11840 20778 11852
rect 21361 11849 21373 11852
rect 21407 11849 21419 11883
rect 21361 11843 21419 11849
rect 11054 11772 11060 11824
rect 11112 11812 11118 11824
rect 11241 11815 11299 11821
rect 11241 11812 11253 11815
rect 11112 11784 11253 11812
rect 11112 11772 11118 11784
rect 11241 11781 11253 11784
rect 11287 11812 11299 11815
rect 12066 11812 12072 11824
rect 11287 11784 12072 11812
rect 11287 11781 11299 11784
rect 11241 11775 11299 11781
rect 12066 11772 12072 11784
rect 12124 11772 12130 11824
rect 12618 11772 12624 11824
rect 12676 11812 12682 11824
rect 15473 11815 15531 11821
rect 12676 11784 12848 11812
rect 12676 11772 12682 11784
rect 7745 11747 7803 11753
rect 7745 11713 7757 11747
rect 7791 11744 7803 11747
rect 8573 11747 8631 11753
rect 8573 11744 8585 11747
rect 7791 11716 8585 11744
rect 7791 11713 7803 11716
rect 7745 11707 7803 11713
rect 8573 11713 8585 11716
rect 8619 11744 8631 11747
rect 11471 11747 11529 11753
rect 8619 11716 9996 11744
rect 8619 11713 8631 11716
rect 8573 11707 8631 11713
rect 9968 11688 9996 11716
rect 11471 11713 11483 11747
rect 11517 11744 11529 11747
rect 12529 11747 12587 11753
rect 12529 11744 12541 11747
rect 11517 11716 12541 11744
rect 11517 11713 11529 11716
rect 11471 11707 11529 11713
rect 12529 11713 12541 11716
rect 12575 11744 12587 11747
rect 12710 11744 12716 11756
rect 12575 11716 12716 11744
rect 12575 11713 12587 11716
rect 12529 11707 12587 11713
rect 12710 11704 12716 11716
rect 12768 11704 12774 11756
rect 12820 11753 12848 11784
rect 15473 11781 15485 11815
rect 15519 11812 15531 11815
rect 16022 11812 16028 11824
rect 15519 11784 16028 11812
rect 15519 11781 15531 11784
rect 15473 11775 15531 11781
rect 16022 11772 16028 11784
rect 16080 11772 16086 11824
rect 18233 11815 18291 11821
rect 18233 11812 18245 11815
rect 16960 11784 18245 11812
rect 16960 11756 16988 11784
rect 18233 11781 18245 11784
rect 18279 11781 18291 11815
rect 18233 11775 18291 11781
rect 12805 11747 12863 11753
rect 12805 11713 12817 11747
rect 12851 11713 12863 11747
rect 12805 11707 12863 11713
rect 14737 11747 14795 11753
rect 14737 11713 14749 11747
rect 14783 11744 14795 11747
rect 16942 11744 16948 11756
rect 14783 11716 16948 11744
rect 14783 11713 14795 11716
rect 14737 11707 14795 11713
rect 16942 11704 16948 11716
rect 17000 11704 17006 11756
rect 17129 11747 17187 11753
rect 17129 11713 17141 11747
rect 17175 11744 17187 11747
rect 17402 11744 17408 11756
rect 17175 11716 17408 11744
rect 17175 11713 17187 11716
rect 17129 11707 17187 11713
rect 17402 11704 17408 11716
rect 17460 11704 17466 11756
rect 19720 11744 19748 11840
rect 19978 11772 19984 11824
rect 20036 11812 20042 11824
rect 21085 11815 21143 11821
rect 21085 11812 21097 11815
rect 20036 11784 21097 11812
rect 20036 11772 20042 11784
rect 21085 11781 21097 11784
rect 21131 11812 21143 11815
rect 21266 11812 21272 11824
rect 21131 11784 21272 11812
rect 21131 11781 21143 11784
rect 21085 11775 21143 11781
rect 21266 11772 21272 11784
rect 21324 11772 21330 11824
rect 19720 11716 21312 11744
rect 7561 11679 7619 11685
rect 7561 11645 7573 11679
rect 7607 11676 7619 11679
rect 7834 11676 7840 11688
rect 7607 11648 7840 11676
rect 7607 11645 7619 11648
rect 7561 11639 7619 11645
rect 7834 11636 7840 11648
rect 7892 11636 7898 11688
rect 8110 11636 8116 11688
rect 8168 11676 8174 11688
rect 8757 11679 8815 11685
rect 8757 11676 8769 11679
rect 8168 11648 8769 11676
rect 8168 11636 8174 11648
rect 8757 11645 8769 11648
rect 8803 11676 8815 11679
rect 9122 11676 9128 11688
rect 8803 11648 9128 11676
rect 8803 11645 8815 11648
rect 8757 11639 8815 11645
rect 9122 11636 9128 11648
rect 9180 11636 9186 11688
rect 9217 11679 9275 11685
rect 9217 11645 9229 11679
rect 9263 11645 9275 11679
rect 9582 11676 9588 11688
rect 9543 11648 9588 11676
rect 9217 11639 9275 11645
rect 3988 11580 4476 11608
rect 6089 11611 6147 11617
rect 6089 11577 6101 11611
rect 6135 11608 6147 11611
rect 6178 11608 6184 11620
rect 6135 11580 6184 11608
rect 6135 11577 6147 11580
rect 6089 11571 6147 11577
rect 6178 11568 6184 11580
rect 6236 11608 6242 11620
rect 7650 11608 7656 11620
rect 6236 11580 7656 11608
rect 6236 11568 6242 11580
rect 7650 11568 7656 11580
rect 7708 11568 7714 11620
rect 9232 11608 9260 11639
rect 9582 11636 9588 11648
rect 9640 11636 9646 11688
rect 9950 11676 9956 11688
rect 9863 11648 9956 11676
rect 9950 11636 9956 11648
rect 10008 11636 10014 11688
rect 11330 11676 11336 11688
rect 11294 11648 11336 11676
rect 11330 11636 11336 11648
rect 11388 11685 11394 11688
rect 11388 11679 11442 11685
rect 11388 11645 11396 11679
rect 11430 11676 11442 11679
rect 11882 11676 11888 11688
rect 11430 11648 11888 11676
rect 11430 11645 11442 11648
rect 11388 11639 11442 11645
rect 11388 11636 11394 11639
rect 11882 11636 11888 11648
rect 11940 11636 11946 11688
rect 14001 11679 14059 11685
rect 14001 11645 14013 11679
rect 14047 11645 14059 11679
rect 14458 11676 14464 11688
rect 14419 11648 14464 11676
rect 14001 11639 14059 11645
rect 8220 11580 9260 11608
rect 8220 11552 8248 11580
rect 10502 11568 10508 11620
rect 10560 11608 10566 11620
rect 12621 11611 12679 11617
rect 10560 11580 12157 11608
rect 10560 11568 10566 11580
rect 1762 11500 1768 11552
rect 1820 11540 1826 11552
rect 2682 11540 2688 11552
rect 1820 11512 2688 11540
rect 1820 11500 1826 11512
rect 2682 11500 2688 11512
rect 2740 11500 2746 11552
rect 4338 11540 4344 11552
rect 4299 11512 4344 11540
rect 4338 11500 4344 11512
rect 4396 11500 4402 11552
rect 6822 11500 6828 11552
rect 6880 11540 6886 11552
rect 7745 11543 7803 11549
rect 7745 11540 7757 11543
rect 6880 11512 7757 11540
rect 6880 11500 6886 11512
rect 7745 11509 7757 11512
rect 7791 11509 7803 11543
rect 7745 11503 7803 11509
rect 7929 11543 7987 11549
rect 7929 11509 7941 11543
rect 7975 11540 7987 11543
rect 8018 11540 8024 11552
rect 7975 11512 8024 11540
rect 7975 11509 7987 11512
rect 7929 11503 7987 11509
rect 8018 11500 8024 11512
rect 8076 11500 8082 11552
rect 8202 11540 8208 11552
rect 8163 11512 8208 11540
rect 8202 11500 8208 11512
rect 8260 11500 8266 11552
rect 9033 11543 9091 11549
rect 9033 11509 9045 11543
rect 9079 11540 9091 11543
rect 9306 11540 9312 11552
rect 9079 11512 9312 11540
rect 9079 11509 9091 11512
rect 9033 11503 9091 11509
rect 9306 11500 9312 11512
rect 9364 11500 9370 11552
rect 10594 11540 10600 11552
rect 10507 11512 10600 11540
rect 10594 11500 10600 11512
rect 10652 11540 10658 11552
rect 11238 11540 11244 11552
rect 10652 11512 11244 11540
rect 10652 11500 10658 11512
rect 11238 11500 11244 11512
rect 11296 11500 11302 11552
rect 11882 11540 11888 11552
rect 11843 11512 11888 11540
rect 11882 11500 11888 11512
rect 11940 11500 11946 11552
rect 12129 11540 12157 11580
rect 12621 11577 12633 11611
rect 12667 11608 12679 11611
rect 12802 11608 12808 11620
rect 12667 11580 12808 11608
rect 12667 11577 12679 11580
rect 12621 11571 12679 11577
rect 12802 11568 12808 11580
rect 12860 11568 12866 11620
rect 14016 11552 14044 11639
rect 14458 11636 14464 11648
rect 14516 11636 14522 11688
rect 21284 11676 21312 11716
rect 21580 11679 21638 11685
rect 21580 11676 21592 11679
rect 21284 11648 21592 11676
rect 21580 11645 21592 11648
rect 21626 11676 21638 11679
rect 22005 11679 22063 11685
rect 22005 11676 22017 11679
rect 21626 11648 22017 11676
rect 21626 11645 21638 11648
rect 21580 11639 21638 11645
rect 22005 11645 22017 11648
rect 22051 11645 22063 11679
rect 22005 11639 22063 11645
rect 16482 11608 16488 11620
rect 16443 11580 16488 11608
rect 16482 11568 16488 11580
rect 16540 11568 16546 11620
rect 16574 11568 16580 11620
rect 16632 11608 16638 11620
rect 20073 11611 20131 11617
rect 16632 11580 16677 11608
rect 16632 11568 16638 11580
rect 20073 11577 20085 11611
rect 20119 11577 20131 11611
rect 20073 11571 20131 11577
rect 13446 11540 13452 11552
rect 12129 11512 13452 11540
rect 13446 11500 13452 11512
rect 13504 11540 13510 11552
rect 13998 11540 14004 11552
rect 13504 11512 14004 11540
rect 13504 11500 13510 11512
rect 13998 11500 14004 11512
rect 14056 11500 14062 11552
rect 16298 11540 16304 11552
rect 16259 11512 16304 11540
rect 16298 11500 16304 11512
rect 16356 11500 16362 11552
rect 17681 11543 17739 11549
rect 17681 11509 17693 11543
rect 17727 11540 17739 11543
rect 18138 11540 18144 11552
rect 17727 11512 18144 11540
rect 17727 11509 17739 11512
rect 17681 11503 17739 11509
rect 18138 11500 18144 11512
rect 18196 11500 18202 11552
rect 18966 11540 18972 11552
rect 18927 11512 18972 11540
rect 18966 11500 18972 11512
rect 19024 11500 19030 11552
rect 20088 11540 20116 11571
rect 20162 11568 20168 11620
rect 20220 11608 20226 11620
rect 20714 11608 20720 11620
rect 20220 11580 20265 11608
rect 20675 11580 20720 11608
rect 20220 11568 20226 11580
rect 20714 11568 20720 11580
rect 20772 11568 20778 11620
rect 20622 11540 20628 11552
rect 20088 11512 20628 11540
rect 20622 11500 20628 11512
rect 20680 11500 20686 11552
rect 21542 11500 21548 11552
rect 21600 11540 21606 11552
rect 21683 11543 21741 11549
rect 21683 11540 21695 11543
rect 21600 11512 21695 11540
rect 21600 11500 21606 11512
rect 21683 11509 21695 11512
rect 21729 11509 21741 11543
rect 21683 11503 21741 11509
rect 1104 11450 22816 11472
rect 1104 11398 8982 11450
rect 9034 11398 9046 11450
rect 9098 11398 9110 11450
rect 9162 11398 9174 11450
rect 9226 11398 16982 11450
rect 17034 11398 17046 11450
rect 17098 11398 17110 11450
rect 17162 11398 17174 11450
rect 17226 11398 22816 11450
rect 1104 11376 22816 11398
rect 1762 11336 1768 11348
rect 1723 11308 1768 11336
rect 1762 11296 1768 11308
rect 1820 11296 1826 11348
rect 2406 11296 2412 11348
rect 2464 11336 2470 11348
rect 2869 11339 2927 11345
rect 2869 11336 2881 11339
rect 2464 11308 2881 11336
rect 2464 11296 2470 11308
rect 2869 11305 2881 11308
rect 2915 11305 2927 11339
rect 2869 11299 2927 11305
rect 6546 11296 6552 11348
rect 6604 11336 6610 11348
rect 6641 11339 6699 11345
rect 6641 11336 6653 11339
rect 6604 11308 6653 11336
rect 6604 11296 6610 11308
rect 6641 11305 6653 11308
rect 6687 11305 6699 11339
rect 8846 11336 8852 11348
rect 6641 11299 6699 11305
rect 8036 11308 8852 11336
rect 2498 11268 2504 11280
rect 1780 11240 2504 11268
rect 1780 11209 1808 11240
rect 2498 11228 2504 11240
rect 2556 11228 2562 11280
rect 3786 11228 3792 11280
rect 3844 11268 3850 11280
rect 3844 11240 5028 11268
rect 3844 11228 3850 11240
rect 1765 11203 1823 11209
rect 1765 11169 1777 11203
rect 1811 11169 1823 11203
rect 2038 11200 2044 11212
rect 1999 11172 2044 11200
rect 1765 11163 1823 11169
rect 2038 11160 2044 11172
rect 2096 11160 2102 11212
rect 4706 11200 4712 11212
rect 4667 11172 4712 11200
rect 4706 11160 4712 11172
rect 4764 11160 4770 11212
rect 5000 11200 5028 11240
rect 8036 11209 8064 11308
rect 8846 11296 8852 11308
rect 8904 11336 8910 11348
rect 9125 11339 9183 11345
rect 9125 11336 9137 11339
rect 8904 11308 9137 11336
rect 8904 11296 8910 11308
rect 9125 11305 9137 11308
rect 9171 11336 9183 11339
rect 9582 11336 9588 11348
rect 9171 11308 9588 11336
rect 9171 11305 9183 11308
rect 9125 11299 9183 11305
rect 9582 11296 9588 11308
rect 9640 11296 9646 11348
rect 11333 11339 11391 11345
rect 11333 11305 11345 11339
rect 11379 11336 11391 11339
rect 12342 11336 12348 11348
rect 11379 11308 12348 11336
rect 11379 11305 11391 11308
rect 11333 11299 11391 11305
rect 12342 11296 12348 11308
rect 12400 11336 12406 11348
rect 12802 11336 12808 11348
rect 12400 11308 12808 11336
rect 12400 11296 12406 11308
rect 12802 11296 12808 11308
rect 12860 11296 12866 11348
rect 13998 11336 14004 11348
rect 13959 11308 14004 11336
rect 13998 11296 14004 11308
rect 14056 11296 14062 11348
rect 16022 11336 16028 11348
rect 15983 11308 16028 11336
rect 16022 11296 16028 11308
rect 16080 11296 16086 11348
rect 16298 11296 16304 11348
rect 16356 11336 16362 11348
rect 16574 11336 16580 11348
rect 16356 11308 16580 11336
rect 16356 11296 16362 11308
rect 16574 11296 16580 11308
rect 16632 11296 16638 11348
rect 8757 11271 8815 11277
rect 8757 11237 8769 11271
rect 8803 11268 8815 11271
rect 9398 11268 9404 11280
rect 8803 11240 9404 11268
rect 8803 11237 8815 11240
rect 8757 11231 8815 11237
rect 9398 11228 9404 11240
rect 9456 11228 9462 11280
rect 10410 11228 10416 11280
rect 10468 11268 10474 11280
rect 10775 11271 10833 11277
rect 10775 11268 10787 11271
rect 10468 11240 10787 11268
rect 10468 11228 10474 11240
rect 10775 11237 10787 11240
rect 10821 11268 10833 11271
rect 12250 11268 12256 11280
rect 10821 11240 12256 11268
rect 10821 11237 10833 11240
rect 10775 11231 10833 11237
rect 12250 11228 12256 11240
rect 12308 11268 12314 11280
rect 12482 11271 12540 11277
rect 12482 11268 12494 11271
rect 12308 11240 12494 11268
rect 12308 11228 12314 11240
rect 12482 11237 12494 11240
rect 12528 11237 12540 11271
rect 20162 11268 20168 11280
rect 12482 11231 12540 11237
rect 19904 11240 20168 11268
rect 5169 11203 5227 11209
rect 5169 11200 5181 11203
rect 5000 11172 5181 11200
rect 5169 11169 5181 11172
rect 5215 11169 5227 11203
rect 5169 11163 5227 11169
rect 8021 11203 8079 11209
rect 8021 11169 8033 11203
rect 8067 11169 8079 11203
rect 8021 11163 8079 11169
rect 8297 11203 8355 11209
rect 8297 11169 8309 11203
rect 8343 11169 8355 11203
rect 12158 11200 12164 11212
rect 12119 11172 12164 11200
rect 8297 11163 8355 11169
rect 1854 11092 1860 11144
rect 1912 11132 1918 11144
rect 2501 11135 2559 11141
rect 2501 11132 2513 11135
rect 1912 11104 2513 11132
rect 1912 11092 1918 11104
rect 2501 11101 2513 11104
rect 2547 11101 2559 11135
rect 2501 11095 2559 11101
rect 5445 11135 5503 11141
rect 5445 11101 5457 11135
rect 5491 11132 5503 11135
rect 5902 11132 5908 11144
rect 5491 11104 5908 11132
rect 5491 11101 5503 11104
rect 5445 11095 5503 11101
rect 5902 11092 5908 11104
rect 5960 11132 5966 11144
rect 6273 11135 6331 11141
rect 6273 11132 6285 11135
rect 5960 11104 6285 11132
rect 5960 11092 5966 11104
rect 6273 11101 6285 11104
rect 6319 11101 6331 11135
rect 8312 11132 8340 11163
rect 12158 11160 12164 11172
rect 12216 11160 12222 11212
rect 17862 11160 17868 11212
rect 17920 11200 17926 11212
rect 19904 11209 19932 11240
rect 20162 11228 20168 11240
rect 20220 11268 20226 11280
rect 20349 11271 20407 11277
rect 20349 11268 20361 11271
rect 20220 11240 20361 11268
rect 20220 11228 20226 11240
rect 20349 11237 20361 11240
rect 20395 11268 20407 11271
rect 21085 11271 21143 11277
rect 21085 11268 21097 11271
rect 20395 11240 21097 11268
rect 20395 11237 20407 11240
rect 20349 11231 20407 11237
rect 21085 11237 21097 11240
rect 21131 11268 21143 11271
rect 21266 11268 21272 11280
rect 21131 11240 21272 11268
rect 21131 11237 21143 11240
rect 21085 11231 21143 11237
rect 21266 11228 21272 11240
rect 21324 11228 21330 11280
rect 21634 11268 21640 11280
rect 21595 11240 21640 11268
rect 21634 11228 21640 11240
rect 21692 11228 21698 11280
rect 18268 11203 18326 11209
rect 18268 11200 18280 11203
rect 17920 11172 18280 11200
rect 17920 11160 17926 11172
rect 18268 11169 18280 11172
rect 18314 11169 18326 11203
rect 18268 11163 18326 11169
rect 19889 11203 19947 11209
rect 19889 11169 19901 11203
rect 19935 11169 19947 11203
rect 19889 11163 19947 11169
rect 19978 11160 19984 11212
rect 20036 11200 20042 11212
rect 20036 11172 20081 11200
rect 20036 11160 20042 11172
rect 6273 11095 6331 11101
rect 8036 11104 8340 11132
rect 10413 11135 10471 11141
rect 8036 11076 8064 11104
rect 10413 11101 10425 11135
rect 10459 11132 10471 11135
rect 10870 11132 10876 11144
rect 10459 11104 10876 11132
rect 10459 11101 10471 11104
rect 10413 11095 10471 11101
rect 10870 11092 10876 11104
rect 10928 11092 10934 11144
rect 15654 11132 15660 11144
rect 15615 11104 15660 11132
rect 15654 11092 15660 11104
rect 15712 11092 15718 11144
rect 20993 11135 21051 11141
rect 20993 11101 21005 11135
rect 21039 11132 21051 11135
rect 21450 11132 21456 11144
rect 21039 11104 21456 11132
rect 21039 11101 21051 11104
rect 20993 11095 21051 11101
rect 21450 11092 21456 11104
rect 21508 11092 21514 11144
rect 8018 11024 8024 11076
rect 8076 11024 8082 11076
rect 8113 11067 8171 11073
rect 8113 11033 8125 11067
rect 8159 11064 8171 11067
rect 8202 11064 8208 11076
rect 8159 11036 8208 11064
rect 8159 11033 8171 11036
rect 8113 11027 8171 11033
rect 8202 11024 8208 11036
rect 8260 11024 8266 11076
rect 13725 11067 13783 11073
rect 13725 11033 13737 11067
rect 13771 11064 13783 11067
rect 14458 11064 14464 11076
rect 13771 11036 14464 11064
rect 13771 11033 13783 11036
rect 13725 11027 13783 11033
rect 14458 11024 14464 11036
rect 14516 11064 14522 11076
rect 15838 11064 15844 11076
rect 14516 11036 15844 11064
rect 14516 11024 14522 11036
rect 15838 11024 15844 11036
rect 15896 11024 15902 11076
rect 3234 10956 3240 11008
rect 3292 10996 3298 11008
rect 3694 10996 3700 11008
rect 3292 10968 3700 10996
rect 3292 10956 3298 10968
rect 3694 10956 3700 10968
rect 3752 10996 3758 11008
rect 4341 10999 4399 11005
rect 4341 10996 4353 10999
rect 3752 10968 4353 10996
rect 3752 10956 3758 10968
rect 4341 10965 4353 10968
rect 4387 10996 4399 10999
rect 5718 10996 5724 11008
rect 4387 10968 5724 10996
rect 4387 10965 4399 10968
rect 4341 10959 4399 10965
rect 5718 10956 5724 10968
rect 5776 10956 5782 11008
rect 7193 10999 7251 11005
rect 7193 10965 7205 10999
rect 7239 10996 7251 10999
rect 7374 10996 7380 11008
rect 7239 10968 7380 10996
rect 7239 10965 7251 10968
rect 7193 10959 7251 10965
rect 7374 10956 7380 10968
rect 7432 10956 7438 11008
rect 7745 10999 7803 11005
rect 7745 10965 7757 10999
rect 7791 10996 7803 10999
rect 7926 10996 7932 11008
rect 7791 10968 7932 10996
rect 7791 10965 7803 10968
rect 7745 10959 7803 10965
rect 7926 10956 7932 10968
rect 7984 10956 7990 11008
rect 12802 10956 12808 11008
rect 12860 10996 12866 11008
rect 13081 10999 13139 11005
rect 13081 10996 13093 10999
rect 12860 10968 13093 10996
rect 12860 10956 12866 10968
rect 13081 10965 13093 10968
rect 13127 10965 13139 10999
rect 13081 10959 13139 10965
rect 15565 10999 15623 11005
rect 15565 10965 15577 10999
rect 15611 10996 15623 10999
rect 15930 10996 15936 11008
rect 15611 10968 15936 10996
rect 15611 10965 15623 10968
rect 15565 10959 15623 10965
rect 15930 10956 15936 10968
rect 15988 10956 15994 11008
rect 18138 10996 18144 11008
rect 18099 10968 18144 10996
rect 18138 10956 18144 10968
rect 18196 10956 18202 11008
rect 18371 10999 18429 11005
rect 18371 10965 18383 10999
rect 18417 10996 18429 10999
rect 18506 10996 18512 11008
rect 18417 10968 18512 10996
rect 18417 10965 18429 10968
rect 18371 10959 18429 10965
rect 18506 10956 18512 10968
rect 18564 10956 18570 11008
rect 20622 10996 20628 11008
rect 20583 10968 20628 10996
rect 20622 10956 20628 10968
rect 20680 10956 20686 11008
rect 1104 10906 22816 10928
rect 1104 10854 4982 10906
rect 5034 10854 5046 10906
rect 5098 10854 5110 10906
rect 5162 10854 5174 10906
rect 5226 10854 12982 10906
rect 13034 10854 13046 10906
rect 13098 10854 13110 10906
rect 13162 10854 13174 10906
rect 13226 10854 20982 10906
rect 21034 10854 21046 10906
rect 21098 10854 21110 10906
rect 21162 10854 21174 10906
rect 21226 10854 22816 10906
rect 1104 10832 22816 10854
rect 1578 10792 1584 10804
rect 1539 10764 1584 10792
rect 1578 10752 1584 10764
rect 1636 10752 1642 10804
rect 2409 10795 2467 10801
rect 2409 10761 2421 10795
rect 2455 10792 2467 10795
rect 2498 10792 2504 10804
rect 2455 10764 2504 10792
rect 2455 10761 2467 10764
rect 2409 10755 2467 10761
rect 2498 10752 2504 10764
rect 2556 10752 2562 10804
rect 4338 10752 4344 10804
rect 4396 10792 4402 10804
rect 4433 10795 4491 10801
rect 4433 10792 4445 10795
rect 4396 10764 4445 10792
rect 4396 10752 4402 10764
rect 4433 10761 4445 10764
rect 4479 10761 4491 10795
rect 5902 10792 5908 10804
rect 5863 10764 5908 10792
rect 4433 10755 4491 10761
rect 2041 10727 2099 10733
rect 2041 10693 2053 10727
rect 2087 10724 2099 10727
rect 4062 10724 4068 10736
rect 2087 10696 4068 10724
rect 2087 10693 2099 10696
rect 2041 10687 2099 10693
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10588 1455 10591
rect 2056 10588 2084 10687
rect 4062 10684 4068 10696
rect 4120 10684 4126 10736
rect 2406 10616 2412 10668
rect 2464 10656 2470 10668
rect 2685 10659 2743 10665
rect 2685 10656 2697 10659
rect 2464 10628 2697 10656
rect 2464 10616 2470 10628
rect 2685 10625 2697 10628
rect 2731 10625 2743 10659
rect 2958 10656 2964 10668
rect 2919 10628 2964 10656
rect 2685 10619 2743 10625
rect 2958 10616 2964 10628
rect 3016 10616 3022 10668
rect 1443 10560 2084 10588
rect 4448 10588 4476 10755
rect 5902 10752 5908 10764
rect 5960 10752 5966 10804
rect 6365 10795 6423 10801
rect 6365 10761 6377 10795
rect 6411 10792 6423 10795
rect 6546 10792 6552 10804
rect 6411 10764 6552 10792
rect 6411 10761 6423 10764
rect 6365 10755 6423 10761
rect 6546 10752 6552 10764
rect 6604 10752 6610 10804
rect 10410 10792 10416 10804
rect 10371 10764 10416 10792
rect 10410 10752 10416 10764
rect 10468 10752 10474 10804
rect 11885 10795 11943 10801
rect 11885 10761 11897 10795
rect 11931 10792 11943 10795
rect 12158 10792 12164 10804
rect 11931 10764 12164 10792
rect 11931 10761 11943 10764
rect 11885 10755 11943 10761
rect 12158 10752 12164 10764
rect 12216 10752 12222 10804
rect 18969 10795 19027 10801
rect 18969 10761 18981 10795
rect 19015 10792 19027 10795
rect 19337 10795 19395 10801
rect 19337 10792 19349 10795
rect 19015 10764 19349 10792
rect 19015 10761 19027 10764
rect 18969 10755 19027 10761
rect 19337 10761 19349 10764
rect 19383 10792 19395 10795
rect 20162 10792 20168 10804
rect 19383 10764 20168 10792
rect 19383 10761 19395 10764
rect 19337 10755 19395 10761
rect 20162 10752 20168 10764
rect 20220 10752 20226 10804
rect 21266 10792 21272 10804
rect 21227 10764 21272 10792
rect 21266 10752 21272 10764
rect 21324 10752 21330 10804
rect 21542 10792 21548 10804
rect 21503 10764 21548 10792
rect 21542 10752 21548 10764
rect 21600 10752 21606 10804
rect 9950 10684 9956 10736
rect 10008 10724 10014 10736
rect 10594 10724 10600 10736
rect 10008 10696 10600 10724
rect 10008 10684 10014 10696
rect 10594 10684 10600 10696
rect 10652 10724 10658 10736
rect 14921 10727 14979 10733
rect 14921 10724 14933 10727
rect 10652 10696 14933 10724
rect 10652 10684 10658 10696
rect 14921 10693 14933 10696
rect 14967 10693 14979 10727
rect 19978 10724 19984 10736
rect 19939 10696 19984 10724
rect 14921 10687 14979 10693
rect 7239 10659 7297 10665
rect 7239 10625 7251 10659
rect 7285 10656 7297 10659
rect 10318 10656 10324 10668
rect 7285 10628 10324 10656
rect 7285 10625 7297 10628
rect 7239 10619 7297 10625
rect 10318 10616 10324 10628
rect 10376 10616 10382 10668
rect 14936 10656 14964 10687
rect 19978 10684 19984 10696
rect 20036 10684 20042 10736
rect 14936 10628 16344 10656
rect 16316 10600 16344 10628
rect 18966 10616 18972 10668
rect 19024 10656 19030 10668
rect 20254 10656 20260 10668
rect 19024 10628 20260 10656
rect 19024 10616 19030 10628
rect 20254 10616 20260 10628
rect 20312 10616 20318 10668
rect 20714 10656 20720 10668
rect 20675 10628 20720 10656
rect 20714 10616 20720 10628
rect 20772 10616 20778 10668
rect 4617 10591 4675 10597
rect 4617 10588 4629 10591
rect 4448 10560 4629 10588
rect 1443 10557 1455 10560
rect 1397 10551 1455 10557
rect 4617 10557 4629 10560
rect 4663 10557 4675 10591
rect 5077 10591 5135 10597
rect 5077 10588 5089 10591
rect 4617 10551 4675 10557
rect 5000 10560 5089 10588
rect 2774 10520 2780 10532
rect 2735 10492 2780 10520
rect 2774 10480 2780 10492
rect 2832 10480 2838 10532
rect 5000 10520 5028 10560
rect 5077 10557 5089 10560
rect 5123 10557 5135 10591
rect 5077 10551 5135 10557
rect 7152 10591 7210 10597
rect 7152 10557 7164 10591
rect 7198 10588 7210 10591
rect 7558 10588 7564 10600
rect 7198 10560 7564 10588
rect 7198 10557 7210 10560
rect 7152 10551 7210 10557
rect 7558 10548 7564 10560
rect 7616 10548 7622 10600
rect 8110 10588 8116 10600
rect 8071 10560 8116 10588
rect 8110 10548 8116 10560
rect 8168 10548 8174 10600
rect 8202 10548 8208 10600
rect 8260 10588 8266 10600
rect 8573 10591 8631 10597
rect 8573 10588 8585 10591
rect 8260 10560 8585 10588
rect 8260 10548 8266 10560
rect 8573 10557 8585 10560
rect 8619 10557 8631 10591
rect 8573 10551 8631 10557
rect 8846 10548 8852 10600
rect 8904 10588 8910 10600
rect 8941 10591 8999 10597
rect 8941 10588 8953 10591
rect 8904 10560 8953 10588
rect 8904 10548 8910 10560
rect 8941 10557 8953 10560
rect 8987 10557 8999 10591
rect 9306 10588 9312 10600
rect 9267 10560 9312 10588
rect 8941 10551 8999 10557
rect 9306 10548 9312 10560
rect 9364 10548 9370 10600
rect 10502 10588 10508 10600
rect 10463 10560 10508 10588
rect 10502 10548 10508 10560
rect 10560 10548 10566 10600
rect 11054 10588 11060 10600
rect 11015 10560 11060 10588
rect 11054 10548 11060 10560
rect 11112 10548 11118 10600
rect 14277 10591 14335 10597
rect 14277 10557 14289 10591
rect 14323 10588 14335 10591
rect 15010 10588 15016 10600
rect 14323 10560 15016 10588
rect 14323 10557 14335 10560
rect 14277 10551 14335 10557
rect 15010 10548 15016 10560
rect 15068 10588 15074 10600
rect 15105 10591 15163 10597
rect 15105 10588 15117 10591
rect 15068 10560 15117 10588
rect 15068 10548 15074 10560
rect 15105 10557 15117 10560
rect 15151 10557 15163 10591
rect 15105 10551 15163 10557
rect 15565 10591 15623 10597
rect 15565 10557 15577 10591
rect 15611 10557 15623 10591
rect 15930 10588 15936 10600
rect 15891 10560 15936 10588
rect 15565 10551 15623 10557
rect 4356 10492 5028 10520
rect 5353 10523 5411 10529
rect 3786 10452 3792 10464
rect 3747 10424 3792 10452
rect 3786 10412 3792 10424
rect 3844 10452 3850 10464
rect 4065 10455 4123 10461
rect 4065 10452 4077 10455
rect 3844 10424 4077 10452
rect 3844 10412 3850 10424
rect 4065 10421 4077 10424
rect 4111 10452 4123 10455
rect 4356 10452 4384 10492
rect 5353 10489 5365 10523
rect 5399 10520 5411 10523
rect 5442 10520 5448 10532
rect 5399 10492 5448 10520
rect 5399 10489 5411 10492
rect 5353 10483 5411 10489
rect 5442 10480 5448 10492
rect 5500 10480 5506 10532
rect 7653 10523 7711 10529
rect 7653 10489 7665 10523
rect 7699 10520 7711 10523
rect 8220 10520 8248 10548
rect 7699 10492 8248 10520
rect 7699 10489 7711 10492
rect 7653 10483 7711 10489
rect 9490 10480 9496 10532
rect 9548 10520 9554 10532
rect 10045 10523 10103 10529
rect 10045 10520 10057 10523
rect 9548 10492 10057 10520
rect 9548 10480 9554 10492
rect 10045 10489 10057 10492
rect 10091 10520 10103 10523
rect 11072 10520 11100 10548
rect 10091 10492 11100 10520
rect 10091 10489 10103 10492
rect 10045 10483 10103 10489
rect 12618 10480 12624 10532
rect 12676 10520 12682 10532
rect 12805 10523 12863 10529
rect 12805 10520 12817 10523
rect 12676 10492 12817 10520
rect 12676 10480 12682 10492
rect 12805 10489 12817 10492
rect 12851 10489 12863 10523
rect 12805 10483 12863 10489
rect 12894 10480 12900 10532
rect 12952 10520 12958 10532
rect 13446 10520 13452 10532
rect 12952 10492 12997 10520
rect 13407 10492 13452 10520
rect 12952 10480 12958 10492
rect 13446 10480 13452 10492
rect 13504 10520 13510 10532
rect 13906 10520 13912 10532
rect 13504 10492 13912 10520
rect 13504 10480 13510 10492
rect 13906 10480 13912 10492
rect 13964 10480 13970 10532
rect 13998 10480 14004 10532
rect 14056 10520 14062 10532
rect 14553 10523 14611 10529
rect 14553 10520 14565 10523
rect 14056 10492 14565 10520
rect 14056 10480 14062 10492
rect 14553 10489 14565 10492
rect 14599 10520 14611 10523
rect 15580 10520 15608 10551
rect 15930 10548 15936 10560
rect 15988 10548 15994 10600
rect 16298 10588 16304 10600
rect 16211 10560 16304 10588
rect 16298 10548 16304 10560
rect 16356 10548 16362 10600
rect 16577 10591 16635 10597
rect 16577 10557 16589 10591
rect 16623 10588 16635 10591
rect 17405 10591 17463 10597
rect 17405 10588 17417 10591
rect 16623 10560 17417 10588
rect 16623 10557 16635 10560
rect 16577 10551 16635 10557
rect 17405 10557 17417 10560
rect 17451 10588 17463 10591
rect 18049 10591 18107 10597
rect 18049 10588 18061 10591
rect 17451 10560 18061 10588
rect 17451 10557 17463 10560
rect 17405 10551 17463 10557
rect 18049 10557 18061 10560
rect 18095 10557 18107 10591
rect 18049 10551 18107 10557
rect 14599 10492 15608 10520
rect 14599 10489 14611 10492
rect 14553 10483 14611 10489
rect 15654 10480 15660 10532
rect 15712 10520 15718 10532
rect 16853 10523 16911 10529
rect 16853 10520 16865 10523
rect 15712 10492 16865 10520
rect 15712 10480 15718 10492
rect 16853 10489 16865 10492
rect 16899 10489 16911 10523
rect 17862 10520 17868 10532
rect 17823 10492 17868 10520
rect 16853 10483 16911 10489
rect 17862 10480 17868 10492
rect 17920 10480 17926 10532
rect 19978 10480 19984 10532
rect 20036 10520 20042 10532
rect 20349 10523 20407 10529
rect 20349 10520 20361 10523
rect 20036 10492 20361 10520
rect 20036 10480 20042 10492
rect 20349 10489 20361 10492
rect 20395 10489 20407 10523
rect 20349 10483 20407 10489
rect 8018 10452 8024 10464
rect 4111 10424 4384 10452
rect 7979 10424 8024 10452
rect 4111 10421 4123 10424
rect 4065 10415 4123 10421
rect 8018 10412 8024 10424
rect 8076 10412 8082 10464
rect 8389 10455 8447 10461
rect 8389 10421 8401 10455
rect 8435 10452 8447 10455
rect 8570 10452 8576 10464
rect 8435 10424 8576 10452
rect 8435 10421 8447 10424
rect 8389 10415 8447 10421
rect 8570 10412 8576 10424
rect 8628 10412 8634 10464
rect 10781 10455 10839 10461
rect 10781 10421 10793 10455
rect 10827 10452 10839 10455
rect 10870 10452 10876 10464
rect 10827 10424 10876 10452
rect 10827 10421 10839 10424
rect 10781 10415 10839 10421
rect 10870 10412 10876 10424
rect 10928 10412 10934 10464
rect 12250 10452 12256 10464
rect 12211 10424 12256 10452
rect 12250 10412 12256 10424
rect 12308 10412 12314 10464
rect 18138 10412 18144 10464
rect 18196 10452 18202 10464
rect 18417 10455 18475 10461
rect 18417 10452 18429 10455
rect 18196 10424 18429 10452
rect 18196 10412 18202 10424
rect 18417 10421 18429 10424
rect 18463 10421 18475 10455
rect 18417 10415 18475 10421
rect 1104 10362 22816 10384
rect 1104 10310 8982 10362
rect 9034 10310 9046 10362
rect 9098 10310 9110 10362
rect 9162 10310 9174 10362
rect 9226 10310 16982 10362
rect 17034 10310 17046 10362
rect 17098 10310 17110 10362
rect 17162 10310 17174 10362
rect 17226 10310 22816 10362
rect 1104 10288 22816 10310
rect 2593 10251 2651 10257
rect 2593 10217 2605 10251
rect 2639 10217 2651 10251
rect 4706 10248 4712 10260
rect 4667 10220 4712 10248
rect 2593 10211 2651 10217
rect 2035 10183 2093 10189
rect 2035 10149 2047 10183
rect 2081 10180 2093 10183
rect 2130 10180 2136 10192
rect 2081 10152 2136 10180
rect 2081 10149 2093 10152
rect 2035 10143 2093 10149
rect 2130 10140 2136 10152
rect 2188 10140 2194 10192
rect 2608 10180 2636 10211
rect 4706 10208 4712 10220
rect 4764 10208 4770 10260
rect 8665 10251 8723 10257
rect 8665 10217 8677 10251
rect 8711 10248 8723 10251
rect 8846 10248 8852 10260
rect 8711 10220 8852 10248
rect 8711 10217 8723 10220
rect 8665 10211 8723 10217
rect 8846 10208 8852 10220
rect 8904 10208 8910 10260
rect 10502 10248 10508 10260
rect 10463 10220 10508 10248
rect 10502 10208 10508 10220
rect 10560 10208 10566 10260
rect 10870 10248 10876 10260
rect 10831 10220 10876 10248
rect 10870 10208 10876 10220
rect 10928 10208 10934 10260
rect 12802 10248 12808 10260
rect 12763 10220 12808 10248
rect 12802 10208 12808 10220
rect 12860 10208 12866 10260
rect 15565 10251 15623 10257
rect 15565 10217 15577 10251
rect 15611 10248 15623 10251
rect 15654 10248 15660 10260
rect 15611 10220 15660 10248
rect 15611 10217 15623 10220
rect 15565 10211 15623 10217
rect 15654 10208 15660 10220
rect 15712 10208 15718 10260
rect 16022 10208 16028 10260
rect 16080 10248 16086 10260
rect 16393 10251 16451 10257
rect 16393 10248 16405 10251
rect 16080 10220 16405 10248
rect 16080 10208 16086 10220
rect 16393 10217 16405 10220
rect 16439 10248 16451 10251
rect 18138 10248 18144 10260
rect 16439 10220 18144 10248
rect 16439 10217 16451 10220
rect 16393 10211 16451 10217
rect 18138 10208 18144 10220
rect 18196 10208 18202 10260
rect 19843 10251 19901 10257
rect 19843 10217 19855 10251
rect 19889 10248 19901 10251
rect 20622 10248 20628 10260
rect 19889 10220 20628 10248
rect 19889 10217 19901 10220
rect 19843 10211 19901 10217
rect 20622 10208 20628 10220
rect 20680 10208 20686 10260
rect 21085 10251 21143 10257
rect 21085 10217 21097 10251
rect 21131 10248 21143 10251
rect 21358 10248 21364 10260
rect 21131 10220 21364 10248
rect 21131 10217 21143 10220
rect 21085 10211 21143 10217
rect 21358 10208 21364 10220
rect 21416 10208 21422 10260
rect 2774 10180 2780 10192
rect 2608 10152 2780 10180
rect 2774 10140 2780 10152
rect 2832 10180 2838 10192
rect 2961 10183 3019 10189
rect 2961 10180 2973 10183
rect 2832 10152 2973 10180
rect 2832 10140 2838 10152
rect 2961 10149 2973 10152
rect 3007 10180 3019 10183
rect 3970 10180 3976 10192
rect 3007 10152 3976 10180
rect 3007 10149 3019 10152
rect 2961 10143 3019 10149
rect 3970 10140 3976 10152
rect 4028 10180 4034 10192
rect 5810 10189 5816 10192
rect 5077 10183 5135 10189
rect 5077 10180 5089 10183
rect 4028 10152 5089 10180
rect 4028 10140 4034 10152
rect 5077 10149 5089 10152
rect 5123 10149 5135 10183
rect 5807 10180 5816 10189
rect 5723 10152 5816 10180
rect 5077 10143 5135 10149
rect 5807 10143 5816 10152
rect 5868 10180 5874 10192
rect 6546 10180 6552 10192
rect 5868 10152 6552 10180
rect 5810 10140 5816 10143
rect 5868 10140 5874 10152
rect 6546 10140 6552 10152
rect 6604 10140 6610 10192
rect 7374 10180 7380 10192
rect 7335 10152 7380 10180
rect 7374 10140 7380 10152
rect 7432 10140 7438 10192
rect 11422 10180 11428 10192
rect 11383 10152 11428 10180
rect 11422 10140 11428 10152
rect 11480 10140 11486 10192
rect 14001 10183 14059 10189
rect 14001 10149 14013 10183
rect 14047 10180 14059 10183
rect 14182 10180 14188 10192
rect 14047 10152 14188 10180
rect 14047 10149 14059 10152
rect 14001 10143 14059 10149
rect 14182 10140 14188 10152
rect 14240 10140 14246 10192
rect 17494 10140 17500 10192
rect 17552 10180 17558 10192
rect 18049 10183 18107 10189
rect 18049 10180 18061 10183
rect 17552 10152 18061 10180
rect 17552 10140 17558 10152
rect 18049 10149 18061 10152
rect 18095 10149 18107 10183
rect 20254 10180 20260 10192
rect 20215 10152 20260 10180
rect 18049 10143 18107 10149
rect 20254 10140 20260 10152
rect 20312 10140 20318 10192
rect 1673 10115 1731 10121
rect 1673 10081 1685 10115
rect 1719 10112 1731 10115
rect 1762 10112 1768 10124
rect 1719 10084 1768 10112
rect 1719 10081 1731 10084
rect 1673 10075 1731 10081
rect 1762 10072 1768 10084
rect 1820 10112 1826 10124
rect 3237 10115 3295 10121
rect 3237 10112 3249 10115
rect 1820 10084 3249 10112
rect 1820 10072 1826 10084
rect 3237 10081 3249 10084
rect 3283 10081 3295 10115
rect 3237 10075 3295 10081
rect 3881 10115 3939 10121
rect 3881 10081 3893 10115
rect 3927 10112 3939 10115
rect 4062 10112 4068 10124
rect 3927 10084 4068 10112
rect 3927 10081 3939 10084
rect 3881 10075 3939 10081
rect 4062 10072 4068 10084
rect 4120 10072 4126 10124
rect 6365 10115 6423 10121
rect 6365 10081 6377 10115
rect 6411 10112 6423 10115
rect 7006 10112 7012 10124
rect 6411 10084 7012 10112
rect 6411 10081 6423 10084
rect 6365 10075 6423 10081
rect 7006 10072 7012 10084
rect 7064 10072 7070 10124
rect 13262 10112 13268 10124
rect 13223 10084 13268 10112
rect 13262 10072 13268 10084
rect 13320 10072 13326 10124
rect 13538 10112 13544 10124
rect 13499 10084 13544 10112
rect 13538 10072 13544 10084
rect 13596 10072 13602 10124
rect 15470 10112 15476 10124
rect 15431 10084 15476 10112
rect 15470 10072 15476 10084
rect 15528 10072 15534 10124
rect 15838 10112 15844 10124
rect 15799 10084 15844 10112
rect 15838 10072 15844 10084
rect 15896 10072 15902 10124
rect 16850 10112 16856 10124
rect 16811 10084 16856 10112
rect 16850 10072 16856 10084
rect 16908 10072 16914 10124
rect 19150 10072 19156 10124
rect 19208 10112 19214 10124
rect 19518 10112 19524 10124
rect 19208 10084 19524 10112
rect 19208 10072 19214 10084
rect 19518 10072 19524 10084
rect 19576 10112 19582 10124
rect 19740 10115 19798 10121
rect 19740 10112 19752 10115
rect 19576 10084 19752 10112
rect 19576 10072 19582 10084
rect 19740 10081 19752 10084
rect 19786 10081 19798 10115
rect 20898 10112 20904 10124
rect 20859 10084 20904 10112
rect 19740 10075 19798 10081
rect 20898 10072 20904 10084
rect 20956 10112 20962 10124
rect 21542 10112 21548 10124
rect 20956 10084 21548 10112
rect 20956 10072 20962 10084
rect 21542 10072 21548 10084
rect 21600 10072 21606 10124
rect 5442 10044 5448 10056
rect 5403 10016 5448 10044
rect 5442 10004 5448 10016
rect 5500 10004 5506 10056
rect 7098 10004 7104 10056
rect 7156 10044 7162 10056
rect 7285 10047 7343 10053
rect 7285 10044 7297 10047
rect 7156 10016 7297 10044
rect 7156 10004 7162 10016
rect 7285 10013 7297 10016
rect 7331 10013 7343 10047
rect 7558 10044 7564 10056
rect 7519 10016 7564 10044
rect 7285 10007 7343 10013
rect 7558 10004 7564 10016
rect 7616 10004 7622 10056
rect 11330 10044 11336 10056
rect 11291 10016 11336 10044
rect 11330 10004 11336 10016
rect 11388 10004 11394 10056
rect 11606 10044 11612 10056
rect 11567 10016 11612 10044
rect 11606 10004 11612 10016
rect 11664 10044 11670 10056
rect 12618 10044 12624 10056
rect 11664 10016 12624 10044
rect 11664 10004 11670 10016
rect 12618 10004 12624 10016
rect 12676 10044 12682 10056
rect 13081 10047 13139 10053
rect 13081 10044 13093 10047
rect 12676 10016 13093 10044
rect 12676 10004 12682 10016
rect 13081 10013 13093 10016
rect 13127 10013 13139 10047
rect 17954 10044 17960 10056
rect 17915 10016 17960 10044
rect 13081 10007 13139 10013
rect 17954 10004 17960 10016
rect 18012 10004 18018 10056
rect 18601 10047 18659 10053
rect 18601 10013 18613 10047
rect 18647 10044 18659 10047
rect 18782 10044 18788 10056
rect 18647 10016 18788 10044
rect 18647 10013 18659 10016
rect 18601 10007 18659 10013
rect 18782 10004 18788 10016
rect 18840 10004 18846 10056
rect 3694 9936 3700 9988
rect 3752 9976 3758 9988
rect 4203 9979 4261 9985
rect 4203 9976 4215 9979
rect 3752 9948 4215 9976
rect 3752 9936 3758 9948
rect 4203 9945 4215 9948
rect 4249 9945 4261 9979
rect 4203 9939 4261 9945
rect 6733 9979 6791 9985
rect 6733 9945 6745 9979
rect 6779 9976 6791 9979
rect 7576 9976 7604 10004
rect 6779 9948 7604 9976
rect 13357 9979 13415 9985
rect 6779 9945 6791 9948
rect 6733 9939 6791 9945
rect 13357 9945 13369 9979
rect 13403 9976 13415 9979
rect 13906 9976 13912 9988
rect 13403 9948 13912 9976
rect 13403 9945 13415 9948
rect 13357 9939 13415 9945
rect 13906 9936 13912 9948
rect 13964 9936 13970 9988
rect 3602 9908 3608 9920
rect 3563 9880 3608 9908
rect 3602 9868 3608 9880
rect 3660 9868 3666 9920
rect 3878 9868 3884 9920
rect 3936 9908 3942 9920
rect 4706 9908 4712 9920
rect 3936 9880 4712 9908
rect 3936 9868 3942 9880
rect 4706 9868 4712 9880
rect 4764 9868 4770 9920
rect 7098 9908 7104 9920
rect 7059 9880 7104 9908
rect 7098 9868 7104 9880
rect 7156 9868 7162 9920
rect 8202 9908 8208 9920
rect 8163 9880 8208 9908
rect 8202 9868 8208 9880
rect 8260 9868 8266 9920
rect 9033 9911 9091 9917
rect 9033 9877 9045 9911
rect 9079 9908 9091 9911
rect 9306 9908 9312 9920
rect 9079 9880 9312 9908
rect 9079 9877 9091 9880
rect 9033 9871 9091 9877
rect 9306 9868 9312 9880
rect 9364 9868 9370 9920
rect 14826 9868 14832 9920
rect 14884 9908 14890 9920
rect 15013 9911 15071 9917
rect 15013 9908 15025 9911
rect 14884 9880 15025 9908
rect 14884 9868 14890 9880
rect 15013 9877 15025 9880
rect 15059 9877 15071 9911
rect 15013 9871 15071 9877
rect 16991 9911 17049 9917
rect 16991 9877 17003 9911
rect 17037 9908 17049 9911
rect 18138 9908 18144 9920
rect 17037 9880 18144 9908
rect 17037 9877 17049 9880
rect 16991 9871 17049 9877
rect 18138 9868 18144 9880
rect 18196 9908 18202 9920
rect 18877 9911 18935 9917
rect 18877 9908 18889 9911
rect 18196 9880 18889 9908
rect 18196 9868 18202 9880
rect 18877 9877 18889 9880
rect 18923 9877 18935 9911
rect 18877 9871 18935 9877
rect 1104 9818 22816 9840
rect 1104 9766 4982 9818
rect 5034 9766 5046 9818
rect 5098 9766 5110 9818
rect 5162 9766 5174 9818
rect 5226 9766 12982 9818
rect 13034 9766 13046 9818
rect 13098 9766 13110 9818
rect 13162 9766 13174 9818
rect 13226 9766 20982 9818
rect 21034 9766 21046 9818
rect 21098 9766 21110 9818
rect 21162 9766 21174 9818
rect 21226 9766 22816 9818
rect 1104 9744 22816 9766
rect 2041 9707 2099 9713
rect 2041 9673 2053 9707
rect 2087 9704 2099 9707
rect 2130 9704 2136 9716
rect 2087 9676 2136 9704
rect 2087 9673 2099 9676
rect 2041 9667 2099 9673
rect 2130 9664 2136 9676
rect 2188 9664 2194 9716
rect 3602 9704 3608 9716
rect 2240 9676 3608 9704
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 2240 9500 2268 9676
rect 3602 9664 3608 9676
rect 3660 9664 3666 9716
rect 5442 9664 5448 9716
rect 5500 9704 5506 9716
rect 5813 9707 5871 9713
rect 5813 9704 5825 9707
rect 5500 9676 5825 9704
rect 5500 9664 5506 9676
rect 5813 9673 5825 9676
rect 5859 9673 5871 9707
rect 5813 9667 5871 9673
rect 6641 9707 6699 9713
rect 6641 9673 6653 9707
rect 6687 9704 6699 9707
rect 7374 9704 7380 9716
rect 6687 9676 7380 9704
rect 6687 9673 6699 9676
rect 6641 9667 6699 9673
rect 7374 9664 7380 9676
rect 7432 9664 7438 9716
rect 7742 9664 7748 9716
rect 7800 9704 7806 9716
rect 8113 9707 8171 9713
rect 8113 9704 8125 9707
rect 7800 9676 8125 9704
rect 7800 9664 7806 9676
rect 8113 9673 8125 9676
rect 8159 9704 8171 9707
rect 8846 9704 8852 9716
rect 8159 9676 8852 9704
rect 8159 9673 8171 9676
rect 8113 9667 8171 9673
rect 8846 9664 8852 9676
rect 8904 9664 8910 9716
rect 11422 9664 11428 9716
rect 11480 9704 11486 9716
rect 11609 9707 11667 9713
rect 11609 9704 11621 9707
rect 11480 9676 11621 9704
rect 11480 9664 11486 9676
rect 11609 9673 11621 9676
rect 11655 9673 11667 9707
rect 16850 9704 16856 9716
rect 16811 9676 16856 9704
rect 11609 9667 11667 9673
rect 16850 9664 16856 9676
rect 16908 9664 16914 9716
rect 21542 9704 21548 9716
rect 21503 9676 21548 9704
rect 21542 9664 21548 9676
rect 21600 9664 21606 9716
rect 2958 9596 2964 9648
rect 3016 9636 3022 9648
rect 6089 9639 6147 9645
rect 6089 9636 6101 9639
rect 3016 9608 6101 9636
rect 3016 9596 3022 9608
rect 6089 9605 6101 9608
rect 6135 9605 6147 9639
rect 6089 9599 6147 9605
rect 8018 9596 8024 9648
rect 8076 9636 8082 9648
rect 13449 9639 13507 9645
rect 13449 9636 13461 9639
rect 8076 9608 13461 9636
rect 8076 9596 8082 9608
rect 13449 9605 13461 9608
rect 13495 9636 13507 9639
rect 13538 9636 13544 9648
rect 13495 9608 13544 9636
rect 13495 9605 13507 9608
rect 13449 9599 13507 9605
rect 13538 9596 13544 9608
rect 13596 9596 13602 9648
rect 14550 9636 14556 9648
rect 14511 9608 14556 9636
rect 14550 9596 14556 9608
rect 14608 9596 14614 9648
rect 14826 9596 14832 9648
rect 14884 9636 14890 9648
rect 14884 9608 16068 9636
rect 14884 9596 14890 9608
rect 2869 9571 2927 9577
rect 2869 9537 2881 9571
rect 2915 9568 2927 9571
rect 3694 9568 3700 9580
rect 2915 9540 3700 9568
rect 2915 9537 2927 9540
rect 2869 9531 2927 9537
rect 3694 9528 3700 9540
rect 3752 9528 3758 9580
rect 4430 9528 4436 9580
rect 4488 9568 4494 9580
rect 5534 9568 5540 9580
rect 4488 9540 5540 9568
rect 4488 9528 4494 9540
rect 5534 9528 5540 9540
rect 5592 9528 5598 9580
rect 11333 9571 11391 9577
rect 11333 9537 11345 9571
rect 11379 9568 11391 9571
rect 11606 9568 11612 9580
rect 11379 9540 11612 9568
rect 11379 9537 11391 9540
rect 11333 9531 11391 9537
rect 11606 9528 11612 9540
rect 11664 9528 11670 9580
rect 15378 9568 15384 9580
rect 12452 9540 15384 9568
rect 12452 9512 12480 9540
rect 15378 9528 15384 9540
rect 15436 9528 15442 9580
rect 4062 9500 4068 9512
rect 1443 9472 2268 9500
rect 4023 9472 4068 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 4062 9460 4068 9472
rect 4120 9460 4126 9512
rect 7650 9460 7656 9512
rect 7708 9500 7714 9512
rect 8849 9503 8907 9509
rect 8849 9500 8861 9503
rect 7708 9472 8861 9500
rect 7708 9460 7714 9472
rect 8849 9469 8861 9472
rect 8895 9500 8907 9503
rect 8941 9503 8999 9509
rect 8941 9500 8953 9503
rect 8895 9472 8953 9500
rect 8895 9469 8907 9472
rect 8849 9463 8907 9469
rect 8941 9469 8953 9472
rect 8987 9469 8999 9503
rect 9490 9500 9496 9512
rect 9451 9472 9496 9500
rect 8941 9463 8999 9469
rect 9490 9460 9496 9472
rect 9548 9460 9554 9512
rect 12253 9503 12311 9509
rect 12253 9469 12265 9503
rect 12299 9500 12311 9503
rect 12434 9500 12440 9512
rect 12299 9472 12440 9500
rect 12299 9469 12311 9472
rect 12253 9463 12311 9469
rect 12434 9460 12440 9472
rect 12492 9460 12498 9512
rect 12894 9500 12900 9512
rect 12855 9472 12900 9500
rect 12894 9460 12900 9472
rect 12952 9460 12958 9512
rect 14052 9503 14110 9509
rect 14052 9469 14064 9503
rect 14098 9500 14110 9503
rect 14550 9500 14556 9512
rect 14098 9472 14556 9500
rect 14098 9469 14110 9472
rect 14052 9463 14110 9469
rect 14550 9460 14556 9472
rect 14608 9460 14614 9512
rect 15010 9500 15016 9512
rect 14971 9472 15016 9500
rect 15010 9460 15016 9472
rect 15068 9460 15074 9512
rect 15473 9503 15531 9509
rect 15473 9469 15485 9503
rect 15519 9469 15531 9503
rect 15841 9503 15899 9509
rect 15841 9500 15853 9503
rect 15473 9463 15531 9469
rect 15580 9472 15853 9500
rect 2961 9435 3019 9441
rect 2961 9401 2973 9435
rect 3007 9401 3019 9435
rect 3510 9432 3516 9444
rect 3471 9404 3516 9432
rect 2961 9395 3019 9401
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 2038 9324 2044 9376
rect 2096 9364 2102 9376
rect 2317 9367 2375 9373
rect 2317 9364 2329 9367
rect 2096 9336 2329 9364
rect 2096 9324 2102 9336
rect 2317 9333 2329 9336
rect 2363 9333 2375 9367
rect 2976 9364 3004 9395
rect 3510 9392 3516 9404
rect 3568 9392 3574 9444
rect 3970 9392 3976 9444
rect 4028 9432 4034 9444
rect 4430 9432 4436 9444
rect 4028 9404 4154 9432
rect 4391 9404 4436 9432
rect 4028 9392 4034 9404
rect 3142 9364 3148 9376
rect 2976 9336 3148 9364
rect 2317 9327 2375 9333
rect 3142 9324 3148 9336
rect 3200 9364 3206 9376
rect 3988 9364 4016 9392
rect 3200 9336 4016 9364
rect 4126 9364 4154 9404
rect 4430 9392 4436 9404
rect 4488 9392 4494 9444
rect 4525 9435 4583 9441
rect 4525 9401 4537 9435
rect 4571 9401 4583 9435
rect 4525 9395 4583 9401
rect 5077 9435 5135 9441
rect 5077 9401 5089 9435
rect 5123 9432 5135 9435
rect 6730 9432 6736 9444
rect 5123 9404 6736 9432
rect 5123 9401 5135 9404
rect 5077 9395 5135 9401
rect 4540 9364 4568 9395
rect 6730 9392 6736 9404
rect 6788 9392 6794 9444
rect 6914 9432 6920 9444
rect 6875 9404 6920 9432
rect 6914 9392 6920 9404
rect 6972 9392 6978 9444
rect 7006 9392 7012 9444
rect 7064 9432 7070 9444
rect 7558 9432 7564 9444
rect 7064 9404 7109 9432
rect 7519 9404 7564 9432
rect 7064 9392 7070 9404
rect 7558 9392 7564 9404
rect 7616 9392 7622 9444
rect 9674 9432 9680 9444
rect 9635 9404 9680 9432
rect 9674 9392 9680 9404
rect 9732 9392 9738 9444
rect 10137 9435 10195 9441
rect 10137 9401 10149 9435
rect 10183 9432 10195 9435
rect 10686 9432 10692 9444
rect 10183 9404 10692 9432
rect 10183 9401 10195 9404
rect 10137 9395 10195 9401
rect 10686 9392 10692 9404
rect 10744 9392 10750 9444
rect 10781 9435 10839 9441
rect 10781 9401 10793 9435
rect 10827 9401 10839 9435
rect 10781 9395 10839 9401
rect 4126 9336 4568 9364
rect 5537 9367 5595 9373
rect 3200 9324 3206 9336
rect 5537 9333 5549 9367
rect 5583 9364 5595 9367
rect 5810 9364 5816 9376
rect 5583 9336 5816 9364
rect 5583 9333 5595 9336
rect 5537 9327 5595 9333
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 6089 9367 6147 9373
rect 6089 9333 6101 9367
rect 6135 9364 6147 9367
rect 6273 9367 6331 9373
rect 6273 9364 6285 9367
rect 6135 9336 6285 9364
rect 6135 9333 6147 9336
rect 6089 9327 6147 9333
rect 6273 9333 6285 9336
rect 6319 9364 6331 9367
rect 6932 9364 6960 9392
rect 6319 9336 6960 9364
rect 6319 9333 6331 9336
rect 6273 9327 6331 9333
rect 8110 9324 8116 9376
rect 8168 9364 8174 9376
rect 8478 9364 8484 9376
rect 8168 9336 8484 9364
rect 8168 9324 8174 9336
rect 8478 9324 8484 9336
rect 8536 9324 8542 9376
rect 10226 9324 10232 9376
rect 10284 9364 10290 9376
rect 10413 9367 10471 9373
rect 10413 9364 10425 9367
rect 10284 9336 10425 9364
rect 10284 9324 10290 9336
rect 10413 9333 10425 9336
rect 10459 9364 10471 9367
rect 10796 9364 10824 9395
rect 11330 9392 11336 9444
rect 11388 9432 11394 9444
rect 14139 9435 14197 9441
rect 14139 9432 14151 9435
rect 11388 9404 14151 9432
rect 11388 9392 11394 9404
rect 14139 9401 14151 9404
rect 14185 9401 14197 9435
rect 14829 9435 14887 9441
rect 14829 9432 14841 9435
rect 14139 9395 14197 9401
rect 14384 9404 14841 9432
rect 12710 9364 12716 9376
rect 10459 9336 10824 9364
rect 12671 9336 12716 9364
rect 10459 9333 10471 9336
rect 10413 9327 10471 9333
rect 12710 9324 12716 9336
rect 12768 9324 12774 9376
rect 13814 9324 13820 9376
rect 13872 9364 13878 9376
rect 14384 9364 14412 9404
rect 14829 9401 14841 9404
rect 14875 9432 14887 9435
rect 15488 9432 15516 9463
rect 14875 9404 15516 9432
rect 14875 9401 14887 9404
rect 14829 9395 14887 9401
rect 13872 9336 14412 9364
rect 13872 9324 13878 9336
rect 15102 9324 15108 9376
rect 15160 9364 15166 9376
rect 15580 9364 15608 9472
rect 15841 9469 15853 9472
rect 15887 9500 15899 9503
rect 15930 9500 15936 9512
rect 15887 9472 15936 9500
rect 15887 9469 15899 9472
rect 15841 9463 15899 9469
rect 15930 9460 15936 9472
rect 15988 9460 15994 9512
rect 16040 9500 16068 9608
rect 17954 9596 17960 9648
rect 18012 9636 18018 9648
rect 19061 9639 19119 9645
rect 19061 9636 19073 9639
rect 18012 9608 19073 9636
rect 18012 9596 18018 9608
rect 19061 9605 19073 9608
rect 19107 9605 19119 9639
rect 19061 9599 19119 9605
rect 18138 9568 18144 9580
rect 18099 9540 18144 9568
rect 18138 9528 18144 9540
rect 18196 9528 18202 9580
rect 20625 9571 20683 9577
rect 20625 9537 20637 9571
rect 20671 9568 20683 9571
rect 20714 9568 20720 9580
rect 20671 9540 20720 9568
rect 20671 9537 20683 9540
rect 20625 9531 20683 9537
rect 20714 9528 20720 9540
rect 20772 9528 20778 9580
rect 16209 9503 16267 9509
rect 16209 9500 16221 9503
rect 16040 9472 16221 9500
rect 16209 9469 16221 9472
rect 16255 9500 16267 9503
rect 16482 9500 16488 9512
rect 16255 9472 16488 9500
rect 16255 9469 16267 9472
rect 16209 9463 16267 9469
rect 16482 9460 16488 9472
rect 16540 9460 16546 9512
rect 18233 9435 18291 9441
rect 18233 9401 18245 9435
rect 18279 9401 18291 9435
rect 18782 9432 18788 9444
rect 18743 9404 18788 9432
rect 18233 9395 18291 9401
rect 15160 9336 15608 9364
rect 15160 9324 15166 9336
rect 16022 9324 16028 9376
rect 16080 9364 16086 9376
rect 16209 9367 16267 9373
rect 16209 9364 16221 9367
rect 16080 9336 16221 9364
rect 16080 9324 16086 9336
rect 16209 9333 16221 9336
rect 16255 9333 16267 9367
rect 17494 9364 17500 9376
rect 17455 9336 17500 9364
rect 16209 9327 16267 9333
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 17862 9364 17868 9376
rect 17823 9336 17868 9364
rect 17862 9324 17868 9336
rect 17920 9364 17926 9376
rect 18248 9364 18276 9395
rect 18782 9392 18788 9404
rect 18840 9392 18846 9444
rect 20441 9435 20499 9441
rect 20441 9401 20453 9435
rect 20487 9432 20499 9435
rect 20717 9435 20775 9441
rect 20717 9432 20729 9435
rect 20487 9404 20729 9432
rect 20487 9401 20499 9404
rect 20441 9395 20499 9401
rect 20717 9401 20729 9404
rect 20763 9432 20775 9435
rect 20806 9432 20812 9444
rect 20763 9404 20812 9432
rect 20763 9401 20775 9404
rect 20717 9395 20775 9401
rect 20806 9392 20812 9404
rect 20864 9392 20870 9444
rect 21266 9432 21272 9444
rect 21227 9404 21272 9432
rect 21266 9392 21272 9404
rect 21324 9392 21330 9444
rect 17920 9336 18276 9364
rect 17920 9324 17926 9336
rect 19518 9324 19524 9376
rect 19576 9364 19582 9376
rect 19705 9367 19763 9373
rect 19705 9364 19717 9367
rect 19576 9336 19717 9364
rect 19576 9324 19582 9336
rect 19705 9333 19717 9336
rect 19751 9333 19763 9367
rect 19705 9327 19763 9333
rect 1104 9274 22816 9296
rect 1104 9222 8982 9274
rect 9034 9222 9046 9274
rect 9098 9222 9110 9274
rect 9162 9222 9174 9274
rect 9226 9222 16982 9274
rect 17034 9222 17046 9274
rect 17098 9222 17110 9274
rect 17162 9222 17174 9274
rect 17226 9222 22816 9274
rect 1104 9200 22816 9222
rect 3142 9160 3148 9172
rect 3103 9132 3148 9160
rect 3142 9120 3148 9132
rect 3200 9120 3206 9172
rect 3513 9163 3571 9169
rect 3513 9129 3525 9163
rect 3559 9160 3571 9163
rect 3694 9160 3700 9172
rect 3559 9132 3700 9160
rect 3559 9129 3571 9132
rect 3513 9123 3571 9129
rect 3694 9120 3700 9132
rect 3752 9120 3758 9172
rect 3881 9163 3939 9169
rect 3881 9129 3893 9163
rect 3927 9160 3939 9163
rect 4203 9163 4261 9169
rect 4203 9160 4215 9163
rect 3927 9132 4215 9160
rect 3927 9129 3939 9132
rect 3881 9123 3939 9129
rect 4203 9129 4215 9132
rect 4249 9160 4261 9163
rect 4430 9160 4436 9172
rect 4249 9132 4436 9160
rect 4249 9129 4261 9132
rect 4203 9123 4261 9129
rect 4430 9120 4436 9132
rect 4488 9120 4494 9172
rect 6917 9163 6975 9169
rect 6917 9129 6929 9163
rect 6963 9160 6975 9163
rect 7006 9160 7012 9172
rect 6963 9132 7012 9160
rect 6963 9129 6975 9132
rect 6917 9123 6975 9129
rect 7006 9120 7012 9132
rect 7064 9120 7070 9172
rect 8570 9120 8576 9172
rect 8628 9160 8634 9172
rect 9033 9163 9091 9169
rect 9033 9160 9045 9163
rect 8628 9132 9045 9160
rect 8628 9120 8634 9132
rect 9033 9129 9045 9132
rect 9079 9160 9091 9163
rect 9490 9160 9496 9172
rect 9079 9132 9496 9160
rect 9079 9129 9091 9132
rect 9033 9123 9091 9129
rect 9490 9120 9496 9132
rect 9548 9120 9554 9172
rect 10045 9163 10103 9169
rect 10045 9129 10057 9163
rect 10091 9160 10103 9163
rect 10410 9160 10416 9172
rect 10091 9132 10416 9160
rect 10091 9129 10103 9132
rect 10045 9123 10103 9129
rect 10410 9120 10416 9132
rect 10468 9120 10474 9172
rect 10686 9120 10692 9172
rect 10744 9160 10750 9172
rect 11563 9163 11621 9169
rect 11563 9160 11575 9163
rect 10744 9132 11575 9160
rect 10744 9120 10750 9132
rect 11563 9129 11575 9132
rect 11609 9129 11621 9163
rect 14734 9160 14740 9172
rect 14647 9132 14740 9160
rect 11563 9123 11621 9129
rect 14734 9120 14740 9132
rect 14792 9160 14798 9172
rect 15010 9160 15016 9172
rect 14792 9132 15016 9160
rect 14792 9120 14798 9132
rect 15010 9120 15016 9132
rect 15068 9120 15074 9172
rect 15470 9160 15476 9172
rect 15431 9132 15476 9160
rect 15470 9120 15476 9132
rect 15528 9120 15534 9172
rect 17494 9120 17500 9172
rect 17552 9160 17558 9172
rect 20625 9163 20683 9169
rect 17552 9132 18644 9160
rect 17552 9120 17558 9132
rect 5715 9095 5773 9101
rect 5715 9061 5727 9095
rect 5761 9092 5773 9095
rect 5810 9092 5816 9104
rect 5761 9064 5816 9092
rect 5761 9061 5773 9064
rect 5715 9055 5773 9061
rect 5810 9052 5816 9064
rect 5868 9052 5874 9104
rect 6638 9092 6644 9104
rect 6288 9064 6644 9092
rect 2038 9024 2044 9036
rect 1999 8996 2044 9024
rect 2038 8984 2044 8996
rect 2096 8984 2102 9036
rect 2314 9024 2320 9036
rect 2275 8996 2320 9024
rect 2314 8984 2320 8996
rect 2372 8984 2378 9036
rect 2777 9027 2835 9033
rect 2777 8993 2789 9027
rect 2823 9024 2835 9027
rect 3878 9024 3884 9036
rect 2823 8996 3884 9024
rect 2823 8993 2835 8996
rect 2777 8987 2835 8993
rect 3878 8984 3884 8996
rect 3936 8984 3942 9036
rect 4132 9027 4190 9033
rect 4132 8993 4144 9027
rect 4178 9024 4190 9027
rect 4430 9024 4436 9036
rect 4178 8996 4436 9024
rect 4178 8993 4190 8996
rect 4132 8987 4190 8993
rect 4430 8984 4436 8996
rect 4488 9024 4494 9036
rect 5994 9024 6000 9036
rect 4488 8996 6000 9024
rect 4488 8984 4494 8996
rect 5994 8984 6000 8996
rect 6052 8984 6058 9036
rect 6288 9033 6316 9064
rect 6638 9052 6644 9064
rect 6696 9092 6702 9104
rect 7285 9095 7343 9101
rect 7285 9092 7297 9095
rect 6696 9064 7297 9092
rect 6696 9052 6702 9064
rect 7285 9061 7297 9064
rect 7331 9061 7343 9095
rect 11330 9092 11336 9104
rect 11291 9064 11336 9092
rect 7285 9055 7343 9061
rect 11330 9052 11336 9064
rect 11388 9052 11394 9104
rect 12250 9052 12256 9104
rect 12308 9092 12314 9104
rect 13034 9095 13092 9101
rect 13034 9092 13046 9095
rect 12308 9064 13046 9092
rect 12308 9052 12314 9064
rect 13034 9061 13046 9064
rect 13080 9061 13092 9095
rect 13034 9055 13092 9061
rect 16206 9052 16212 9104
rect 16264 9092 16270 9104
rect 16346 9095 16404 9101
rect 16346 9092 16358 9095
rect 16264 9064 16358 9092
rect 16264 9052 16270 9064
rect 16346 9061 16358 9064
rect 16392 9061 16404 9095
rect 18506 9092 18512 9104
rect 18467 9064 18512 9092
rect 16346 9055 16404 9061
rect 18506 9052 18512 9064
rect 18564 9052 18570 9104
rect 18616 9101 18644 9132
rect 20625 9129 20637 9163
rect 20671 9160 20683 9163
rect 20714 9160 20720 9172
rect 20671 9132 20720 9160
rect 20671 9129 20683 9132
rect 20625 9123 20683 9129
rect 20714 9120 20720 9132
rect 20772 9120 20778 9172
rect 21634 9160 21640 9172
rect 21008 9132 21640 9160
rect 18601 9095 18659 9101
rect 18601 9061 18613 9095
rect 18647 9092 18659 9095
rect 19242 9092 19248 9104
rect 18647 9064 19248 9092
rect 18647 9061 18659 9064
rect 18601 9055 18659 9061
rect 19242 9052 19248 9064
rect 19300 9052 19306 9104
rect 21008 9101 21036 9132
rect 21634 9120 21640 9132
rect 21692 9120 21698 9172
rect 20993 9095 21051 9101
rect 20993 9061 21005 9095
rect 21039 9061 21051 9095
rect 20993 9055 21051 9061
rect 21082 9052 21088 9104
rect 21140 9092 21146 9104
rect 21140 9064 21185 9092
rect 21140 9052 21146 9064
rect 6273 9027 6331 9033
rect 6273 8993 6285 9027
rect 6319 8993 6331 9027
rect 9674 9024 9680 9036
rect 9635 8996 9680 9024
rect 6273 8987 6331 8993
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 11238 8984 11244 9036
rect 11296 9024 11302 9036
rect 11460 9027 11518 9033
rect 11460 9024 11472 9027
rect 11296 8996 11472 9024
rect 11296 8984 11302 8996
rect 11460 8993 11472 8996
rect 11506 8993 11518 9027
rect 12710 9024 12716 9036
rect 12671 8996 12716 9024
rect 11460 8987 11518 8993
rect 12710 8984 12716 8996
rect 12768 8984 12774 9036
rect 1854 8916 1860 8968
rect 1912 8956 1918 8968
rect 2133 8959 2191 8965
rect 2133 8956 2145 8959
rect 1912 8928 2145 8956
rect 1912 8916 1918 8928
rect 2133 8925 2145 8928
rect 2179 8925 2191 8959
rect 3786 8956 3792 8968
rect 2133 8919 2191 8925
rect 3114 8928 3792 8956
rect 1673 8823 1731 8829
rect 1673 8789 1685 8823
rect 1719 8820 1731 8823
rect 1946 8820 1952 8832
rect 1719 8792 1952 8820
rect 1719 8789 1731 8792
rect 1673 8783 1731 8789
rect 1946 8780 1952 8792
rect 2004 8820 2010 8832
rect 3114 8820 3142 8928
rect 3786 8916 3792 8928
rect 3844 8956 3850 8968
rect 5350 8956 5356 8968
rect 3844 8928 4844 8956
rect 5311 8928 5356 8956
rect 3844 8916 3850 8928
rect 4816 8832 4844 8928
rect 5350 8916 5356 8928
rect 5408 8916 5414 8968
rect 6730 8916 6736 8968
rect 6788 8956 6794 8968
rect 7193 8959 7251 8965
rect 7193 8956 7205 8959
rect 6788 8928 7205 8956
rect 6788 8916 6794 8928
rect 7193 8925 7205 8928
rect 7239 8956 7251 8959
rect 7374 8956 7380 8968
rect 7239 8928 7380 8956
rect 7239 8925 7251 8928
rect 7193 8919 7251 8925
rect 7374 8916 7380 8928
rect 7432 8916 7438 8968
rect 7558 8956 7564 8968
rect 7519 8928 7564 8956
rect 7558 8916 7564 8928
rect 7616 8916 7622 8968
rect 11054 8916 11060 8968
rect 11112 8956 11118 8968
rect 12437 8959 12495 8965
rect 12437 8956 12449 8959
rect 11112 8928 12449 8956
rect 11112 8916 11118 8928
rect 12437 8925 12449 8928
rect 12483 8956 12495 8959
rect 12894 8956 12900 8968
rect 12483 8928 12900 8956
rect 12483 8925 12495 8928
rect 12437 8919 12495 8925
rect 12894 8916 12900 8928
rect 12952 8916 12958 8968
rect 13262 8916 13268 8968
rect 13320 8956 13326 8968
rect 13909 8959 13967 8965
rect 13909 8956 13921 8959
rect 13320 8928 13921 8956
rect 13320 8916 13326 8928
rect 13909 8925 13921 8928
rect 13955 8925 13967 8959
rect 15010 8956 15016 8968
rect 14971 8928 15016 8956
rect 13909 8919 13967 8925
rect 15010 8916 15016 8928
rect 15068 8916 15074 8968
rect 16022 8956 16028 8968
rect 15983 8928 16028 8956
rect 16022 8916 16028 8928
rect 16080 8916 16086 8968
rect 18966 8956 18972 8968
rect 18927 8928 18972 8956
rect 18966 8916 18972 8928
rect 19024 8916 19030 8968
rect 21266 8956 21272 8968
rect 21227 8928 21272 8956
rect 21266 8916 21272 8928
rect 21324 8916 21330 8968
rect 10686 8848 10692 8900
rect 10744 8888 10750 8900
rect 13280 8888 13308 8916
rect 10744 8860 13308 8888
rect 16945 8891 17003 8897
rect 10744 8848 10750 8860
rect 16945 8857 16957 8891
rect 16991 8888 17003 8891
rect 20714 8888 20720 8900
rect 16991 8860 20720 8888
rect 16991 8857 17003 8860
rect 16945 8851 17003 8857
rect 20714 8848 20720 8860
rect 20772 8888 20778 8900
rect 21082 8888 21088 8900
rect 20772 8860 21088 8888
rect 20772 8848 20778 8860
rect 21082 8848 21088 8860
rect 21140 8848 21146 8900
rect 4706 8820 4712 8832
rect 2004 8792 3142 8820
rect 4667 8792 4712 8820
rect 2004 8780 2010 8792
rect 4706 8780 4712 8792
rect 4764 8780 4770 8832
rect 4798 8780 4804 8832
rect 4856 8820 4862 8832
rect 4985 8823 5043 8829
rect 4985 8820 4997 8823
rect 4856 8792 4997 8820
rect 4856 8780 4862 8792
rect 4985 8789 4997 8792
rect 5031 8789 5043 8823
rect 4985 8783 5043 8789
rect 10226 8780 10232 8832
rect 10284 8820 10290 8832
rect 10597 8823 10655 8829
rect 10597 8820 10609 8823
rect 10284 8792 10609 8820
rect 10284 8780 10290 8792
rect 10597 8789 10609 8792
rect 10643 8789 10655 8823
rect 13630 8820 13636 8832
rect 13591 8792 13636 8820
rect 10597 8783 10655 8789
rect 13630 8780 13636 8792
rect 13688 8780 13694 8832
rect 15838 8820 15844 8832
rect 15799 8792 15844 8820
rect 15838 8780 15844 8792
rect 15896 8780 15902 8832
rect 18230 8820 18236 8832
rect 18191 8792 18236 8820
rect 18230 8780 18236 8792
rect 18288 8780 18294 8832
rect 1104 8730 22816 8752
rect 1104 8678 4982 8730
rect 5034 8678 5046 8730
rect 5098 8678 5110 8730
rect 5162 8678 5174 8730
rect 5226 8678 12982 8730
rect 13034 8678 13046 8730
rect 13098 8678 13110 8730
rect 13162 8678 13174 8730
rect 13226 8678 20982 8730
rect 21034 8678 21046 8730
rect 21098 8678 21110 8730
rect 21162 8678 21174 8730
rect 21226 8678 22816 8730
rect 1104 8656 22816 8678
rect 2314 8576 2320 8628
rect 2372 8616 2378 8628
rect 2869 8619 2927 8625
rect 2869 8616 2881 8619
rect 2372 8588 2881 8616
rect 2372 8576 2378 8588
rect 2869 8585 2881 8588
rect 2915 8585 2927 8619
rect 2869 8579 2927 8585
rect 4065 8619 4123 8625
rect 4065 8585 4077 8619
rect 4111 8616 4123 8619
rect 6086 8616 6092 8628
rect 4111 8588 6092 8616
rect 4111 8585 4123 8588
rect 4065 8579 4123 8585
rect 2038 8508 2044 8560
rect 2096 8548 2102 8560
rect 3234 8548 3240 8560
rect 2096 8520 3240 8548
rect 2096 8508 2102 8520
rect 3234 8508 3240 8520
rect 3292 8508 3298 8560
rect 1854 8440 1860 8492
rect 1912 8480 1918 8492
rect 2501 8483 2559 8489
rect 2501 8480 2513 8483
rect 1912 8452 2513 8480
rect 1912 8440 1918 8452
rect 2501 8449 2513 8452
rect 2547 8449 2559 8483
rect 2501 8443 2559 8449
rect 1670 8412 1676 8424
rect 1631 8384 1676 8412
rect 1670 8372 1676 8384
rect 1728 8372 1734 8424
rect 1946 8412 1952 8424
rect 1907 8384 1952 8412
rect 1946 8372 1952 8384
rect 2004 8372 2010 8424
rect 3580 8415 3638 8421
rect 3580 8381 3592 8415
rect 3626 8412 3638 8415
rect 4080 8412 4108 8579
rect 6086 8576 6092 8588
rect 6144 8576 6150 8628
rect 6638 8616 6644 8628
rect 6599 8588 6644 8616
rect 6638 8576 6644 8588
rect 6696 8576 6702 8628
rect 10318 8576 10324 8628
rect 10376 8616 10382 8628
rect 10505 8619 10563 8625
rect 10505 8616 10517 8619
rect 10376 8588 10517 8616
rect 10376 8576 10382 8588
rect 10505 8585 10517 8588
rect 10551 8616 10563 8619
rect 11422 8616 11428 8628
rect 10551 8588 11428 8616
rect 10551 8585 10563 8588
rect 10505 8579 10563 8585
rect 11422 8576 11428 8588
rect 11480 8576 11486 8628
rect 11885 8619 11943 8625
rect 11885 8585 11897 8619
rect 11931 8616 11943 8619
rect 12710 8616 12716 8628
rect 11931 8588 12716 8616
rect 11931 8585 11943 8588
rect 11885 8579 11943 8585
rect 12710 8576 12716 8588
rect 12768 8576 12774 8628
rect 15473 8619 15531 8625
rect 15473 8616 15485 8619
rect 13096 8588 15485 8616
rect 4522 8508 4528 8560
rect 4580 8548 4586 8560
rect 7837 8551 7895 8557
rect 7837 8548 7849 8551
rect 4580 8520 7849 8548
rect 4580 8508 4586 8520
rect 7837 8517 7849 8520
rect 7883 8517 7895 8551
rect 7837 8511 7895 8517
rect 5350 8480 5356 8492
rect 5263 8452 5356 8480
rect 5350 8440 5356 8452
rect 5408 8480 5414 8492
rect 5997 8483 6055 8489
rect 5997 8480 6009 8483
rect 5408 8452 6009 8480
rect 5408 8440 5414 8452
rect 5997 8449 6009 8452
rect 6043 8449 6055 8483
rect 5997 8443 6055 8449
rect 4706 8412 4712 8424
rect 3626 8384 4108 8412
rect 4667 8384 4712 8412
rect 3626 8381 3638 8384
rect 3580 8375 3638 8381
rect 4706 8372 4712 8384
rect 4764 8372 4770 8424
rect 4798 8372 4804 8424
rect 4856 8412 4862 8424
rect 5077 8415 5135 8421
rect 5077 8412 5089 8415
rect 4856 8384 5089 8412
rect 4856 8372 4862 8384
rect 5077 8381 5089 8384
rect 5123 8381 5135 8415
rect 5077 8375 5135 8381
rect 5721 8415 5779 8421
rect 5721 8381 5733 8415
rect 5767 8412 5779 8415
rect 5810 8412 5816 8424
rect 5767 8384 5816 8412
rect 5767 8381 5779 8384
rect 5721 8375 5779 8381
rect 5810 8372 5816 8384
rect 5868 8372 5874 8424
rect 6892 8415 6950 8421
rect 6892 8381 6904 8415
rect 6938 8412 6950 8415
rect 7852 8412 7880 8511
rect 11238 8440 11244 8492
rect 11296 8480 11302 8492
rect 11425 8483 11483 8489
rect 11425 8480 11437 8483
rect 11296 8452 11437 8480
rect 11296 8440 11302 8452
rect 11425 8449 11437 8452
rect 11471 8449 11483 8483
rect 11425 8443 11483 8449
rect 12250 8440 12256 8492
rect 12308 8480 12314 8492
rect 12713 8483 12771 8489
rect 12713 8480 12725 8483
rect 12308 8452 12725 8480
rect 12308 8440 12314 8452
rect 12713 8449 12725 8452
rect 12759 8480 12771 8483
rect 13096 8480 13124 8588
rect 15473 8585 15485 8588
rect 15519 8616 15531 8619
rect 15841 8619 15899 8625
rect 15841 8616 15853 8619
rect 15519 8588 15853 8616
rect 15519 8585 15531 8588
rect 15473 8579 15531 8585
rect 15841 8585 15853 8588
rect 15887 8585 15899 8619
rect 15841 8579 15899 8585
rect 13538 8548 13544 8560
rect 13188 8520 13544 8548
rect 13188 8489 13216 8520
rect 13538 8508 13544 8520
rect 13596 8508 13602 8560
rect 12759 8452 13124 8480
rect 13173 8483 13231 8489
rect 12759 8449 12771 8452
rect 12713 8443 12771 8449
rect 13173 8449 13185 8483
rect 13219 8449 13231 8483
rect 13446 8480 13452 8492
rect 13407 8452 13452 8480
rect 13173 8443 13231 8449
rect 13446 8440 13452 8452
rect 13504 8440 13510 8492
rect 15856 8480 15884 8579
rect 16022 8576 16028 8628
rect 16080 8616 16086 8628
rect 17221 8619 17279 8625
rect 17221 8616 17233 8619
rect 16080 8588 17233 8616
rect 16080 8576 16086 8588
rect 17221 8585 17233 8588
rect 17267 8585 17279 8619
rect 17221 8579 17279 8585
rect 20714 8576 20720 8628
rect 20772 8616 20778 8628
rect 20901 8619 20959 8625
rect 20901 8616 20913 8619
rect 20772 8588 20913 8616
rect 20772 8576 20778 8588
rect 20901 8585 20913 8588
rect 20947 8585 20959 8619
rect 20901 8579 20959 8585
rect 21634 8576 21640 8628
rect 21692 8616 21698 8628
rect 21729 8619 21787 8625
rect 21729 8616 21741 8619
rect 21692 8588 21741 8616
rect 21692 8576 21698 8588
rect 21729 8585 21741 8588
rect 21775 8585 21787 8619
rect 21729 8579 21787 8585
rect 16945 8551 17003 8557
rect 16945 8517 16957 8551
rect 16991 8548 17003 8551
rect 17494 8548 17500 8560
rect 16991 8520 17500 8548
rect 16991 8517 17003 8520
rect 16945 8511 17003 8517
rect 17494 8508 17500 8520
rect 17552 8508 17558 8560
rect 16206 8480 16212 8492
rect 15856 8452 16212 8480
rect 16206 8440 16212 8452
rect 16264 8480 16270 8492
rect 18230 8480 18236 8492
rect 16264 8452 16389 8480
rect 18143 8452 18236 8480
rect 16264 8440 16270 8452
rect 8021 8415 8079 8421
rect 8021 8412 8033 8415
rect 6938 8384 7420 8412
rect 7852 8384 8033 8412
rect 6938 8381 6950 8384
rect 6892 8375 6950 8381
rect 1762 8276 1768 8288
rect 1723 8248 1768 8276
rect 1762 8236 1768 8248
rect 1820 8236 1826 8288
rect 3651 8279 3709 8285
rect 3651 8245 3663 8279
rect 3697 8276 3709 8279
rect 3878 8276 3884 8288
rect 3697 8248 3884 8276
rect 3697 8245 3709 8248
rect 3651 8239 3709 8245
rect 3878 8236 3884 8248
rect 3936 8236 3942 8288
rect 4430 8276 4436 8288
rect 4391 8248 4436 8276
rect 4430 8236 4436 8248
rect 4488 8236 4494 8288
rect 6730 8236 6736 8288
rect 6788 8276 6794 8288
rect 7392 8285 7420 8384
rect 8021 8381 8033 8384
rect 8067 8381 8079 8415
rect 8570 8412 8576 8424
rect 8531 8384 8576 8412
rect 8021 8375 8079 8381
rect 8570 8372 8576 8384
rect 8628 8372 8634 8424
rect 8757 8415 8815 8421
rect 8757 8381 8769 8415
rect 8803 8412 8815 8415
rect 9585 8415 9643 8421
rect 9585 8412 9597 8415
rect 8803 8384 9597 8412
rect 8803 8381 8815 8384
rect 8757 8375 8815 8381
rect 9585 8381 9597 8384
rect 9631 8412 9643 8415
rect 10781 8415 10839 8421
rect 10781 8412 10793 8415
rect 9631 8384 10793 8412
rect 9631 8381 9643 8384
rect 9585 8375 9643 8381
rect 10781 8381 10793 8384
rect 10827 8381 10839 8415
rect 16025 8415 16083 8421
rect 16025 8412 16037 8415
rect 10781 8375 10839 8381
rect 15396 8384 16037 8412
rect 9947 8347 10005 8353
rect 9947 8344 9959 8347
rect 9646 8316 9959 8344
rect 6963 8279 7021 8285
rect 6963 8276 6975 8279
rect 6788 8248 6975 8276
rect 6788 8236 6794 8248
rect 6963 8245 6975 8248
rect 7009 8245 7021 8279
rect 6963 8239 7021 8245
rect 7377 8279 7435 8285
rect 7377 8245 7389 8279
rect 7423 8276 7435 8279
rect 7558 8276 7564 8288
rect 7423 8248 7564 8276
rect 7423 8245 7435 8248
rect 7377 8239 7435 8245
rect 7558 8236 7564 8248
rect 7616 8236 7622 8288
rect 9125 8279 9183 8285
rect 9125 8245 9137 8279
rect 9171 8276 9183 8279
rect 9493 8279 9551 8285
rect 9493 8276 9505 8279
rect 9171 8248 9505 8276
rect 9171 8245 9183 8248
rect 9125 8239 9183 8245
rect 9493 8245 9505 8248
rect 9539 8276 9551 8279
rect 9646 8276 9674 8316
rect 9947 8313 9959 8316
rect 9993 8344 10005 8347
rect 10410 8344 10416 8356
rect 9993 8316 10416 8344
rect 9993 8313 10005 8316
rect 9947 8307 10005 8313
rect 10410 8304 10416 8316
rect 10468 8304 10474 8356
rect 12253 8347 12311 8353
rect 12253 8313 12265 8347
rect 12299 8344 12311 8347
rect 13265 8347 13323 8353
rect 12299 8316 13077 8344
rect 12299 8313 12311 8316
rect 12253 8307 12311 8313
rect 9539 8248 9674 8276
rect 13049 8276 13077 8316
rect 13265 8313 13277 8347
rect 13311 8344 13323 8347
rect 13630 8344 13636 8356
rect 13311 8316 13636 8344
rect 13311 8313 13323 8316
rect 13265 8307 13323 8313
rect 13280 8276 13308 8307
rect 13630 8304 13636 8316
rect 13688 8304 13694 8356
rect 15396 8288 15424 8384
rect 16025 8381 16037 8384
rect 16071 8381 16083 8415
rect 16025 8375 16083 8381
rect 16361 8353 16389 8452
rect 18230 8440 18236 8452
rect 18288 8480 18294 8492
rect 19610 8480 19616 8492
rect 18288 8452 19616 8480
rect 18288 8440 18294 8452
rect 19610 8440 19616 8452
rect 19668 8440 19674 8492
rect 19242 8412 19248 8424
rect 19155 8384 19248 8412
rect 19242 8372 19248 8384
rect 19300 8412 19306 8424
rect 19521 8415 19579 8421
rect 19521 8412 19533 8415
rect 19300 8384 19533 8412
rect 19300 8372 19306 8384
rect 19521 8381 19533 8384
rect 19567 8412 19579 8415
rect 19797 8415 19855 8421
rect 19797 8412 19809 8415
rect 19567 8384 19809 8412
rect 19567 8381 19579 8384
rect 19521 8375 19579 8381
rect 19797 8381 19809 8384
rect 19843 8381 19855 8415
rect 19797 8375 19855 8381
rect 21177 8415 21235 8421
rect 21177 8381 21189 8415
rect 21223 8412 21235 8415
rect 21266 8412 21272 8424
rect 21223 8384 21272 8412
rect 21223 8381 21235 8384
rect 21177 8375 21235 8381
rect 21266 8372 21272 8384
rect 21324 8412 21330 8424
rect 22097 8415 22155 8421
rect 22097 8412 22109 8415
rect 21324 8384 22109 8412
rect 21324 8372 21330 8384
rect 22097 8381 22109 8384
rect 22143 8381 22155 8415
rect 22097 8375 22155 8381
rect 16346 8347 16404 8353
rect 16346 8313 16358 8347
rect 16392 8344 16404 8347
rect 17678 8344 17684 8356
rect 16392 8316 17684 8344
rect 16392 8313 16404 8316
rect 16346 8307 16404 8313
rect 17678 8304 17684 8316
rect 17736 8304 17742 8356
rect 17862 8344 17868 8356
rect 17775 8316 17868 8344
rect 17862 8304 17868 8316
rect 17920 8344 17926 8356
rect 18325 8347 18383 8353
rect 18325 8344 18337 8347
rect 17920 8316 18337 8344
rect 17920 8304 17926 8316
rect 18325 8313 18337 8316
rect 18371 8313 18383 8347
rect 18325 8307 18383 8313
rect 18877 8347 18935 8353
rect 18877 8313 18889 8347
rect 18923 8344 18935 8347
rect 18966 8344 18972 8356
rect 18923 8316 18972 8344
rect 18923 8313 18935 8316
rect 18877 8307 18935 8313
rect 13049 8248 13308 8276
rect 15197 8279 15255 8285
rect 9539 8245 9551 8248
rect 9493 8239 9551 8245
rect 15197 8245 15209 8279
rect 15243 8276 15255 8279
rect 15378 8276 15384 8288
rect 15243 8248 15384 8276
rect 15243 8245 15255 8248
rect 15197 8239 15255 8245
rect 15378 8236 15384 8248
rect 15436 8236 15442 8288
rect 18340 8276 18368 8307
rect 18966 8304 18972 8316
rect 19024 8304 19030 8356
rect 19705 8347 19763 8353
rect 19705 8344 19717 8347
rect 19076 8316 19717 8344
rect 19076 8276 19104 8316
rect 19705 8313 19717 8316
rect 19751 8313 19763 8347
rect 19705 8307 19763 8313
rect 18340 8248 19104 8276
rect 19150 8236 19156 8288
rect 19208 8276 19214 8288
rect 21407 8279 21465 8285
rect 21407 8276 21419 8279
rect 19208 8248 21419 8276
rect 19208 8236 19214 8248
rect 21407 8245 21419 8248
rect 21453 8245 21465 8279
rect 21407 8239 21465 8245
rect 1104 8186 22816 8208
rect 1104 8134 8982 8186
rect 9034 8134 9046 8186
rect 9098 8134 9110 8186
rect 9162 8134 9174 8186
rect 9226 8134 16982 8186
rect 17034 8134 17046 8186
rect 17098 8134 17110 8186
rect 17162 8134 17174 8186
rect 17226 8134 22816 8186
rect 1104 8112 22816 8134
rect 1670 8072 1676 8084
rect 1631 8044 1676 8072
rect 1670 8032 1676 8044
rect 1728 8032 1734 8084
rect 2130 8072 2136 8084
rect 2091 8044 2136 8072
rect 2130 8032 2136 8044
rect 2188 8032 2194 8084
rect 2685 8075 2743 8081
rect 2685 8041 2697 8075
rect 2731 8072 2743 8075
rect 2731 8044 4292 8072
rect 2731 8041 2743 8044
rect 2685 8035 2743 8041
rect 4264 8016 4292 8044
rect 4706 8032 4712 8084
rect 4764 8072 4770 8084
rect 4764 8044 7006 8072
rect 4764 8032 4770 8044
rect 3878 7964 3884 8016
rect 3936 8004 3942 8016
rect 4157 8007 4215 8013
rect 4157 8004 4169 8007
rect 3936 7976 4169 8004
rect 3936 7964 3942 7976
rect 4157 7973 4169 7976
rect 4203 7973 4215 8007
rect 4157 7967 4215 7973
rect 4246 7964 4252 8016
rect 4304 8004 4310 8016
rect 6549 8007 6607 8013
rect 4304 7976 4349 8004
rect 4304 7964 4310 7976
rect 6549 7973 6561 8007
rect 6595 8004 6607 8007
rect 6730 8004 6736 8016
rect 6595 7976 6736 8004
rect 6595 7973 6607 7976
rect 6549 7967 6607 7973
rect 6730 7964 6736 7976
rect 6788 7964 6794 8016
rect 6822 7964 6828 8016
rect 6880 8004 6886 8016
rect 6978 8004 7006 8044
rect 7374 8032 7380 8084
rect 7432 8072 7438 8084
rect 7653 8075 7711 8081
rect 7653 8072 7665 8075
rect 7432 8044 7665 8072
rect 7432 8032 7438 8044
rect 7653 8041 7665 8044
rect 7699 8041 7711 8075
rect 7653 8035 7711 8041
rect 8113 8075 8171 8081
rect 8113 8041 8125 8075
rect 8159 8072 8171 8075
rect 8570 8072 8576 8084
rect 8159 8044 8576 8072
rect 8159 8041 8171 8044
rect 8113 8035 8171 8041
rect 8570 8032 8576 8044
rect 8628 8032 8634 8084
rect 9493 8075 9551 8081
rect 9493 8041 9505 8075
rect 9539 8072 9551 8075
rect 9674 8072 9680 8084
rect 9539 8044 9680 8072
rect 9539 8041 9551 8044
rect 9493 8035 9551 8041
rect 9674 8032 9680 8044
rect 9732 8032 9738 8084
rect 15378 8072 15384 8084
rect 15339 8044 15384 8072
rect 15378 8032 15384 8044
rect 15436 8032 15442 8084
rect 18506 8032 18512 8084
rect 18564 8072 18570 8084
rect 19061 8075 19119 8081
rect 19061 8072 19073 8075
rect 18564 8044 19073 8072
rect 18564 8032 18570 8044
rect 19061 8041 19073 8044
rect 19107 8041 19119 8075
rect 19610 8072 19616 8084
rect 19571 8044 19616 8072
rect 19061 8035 19119 8041
rect 19610 8032 19616 8044
rect 19668 8032 19674 8084
rect 7834 8004 7840 8016
rect 6880 7976 6925 8004
rect 6978 7976 7840 8004
rect 6880 7964 6886 7976
rect 7834 7964 7840 7976
rect 7892 8004 7898 8016
rect 7892 7976 11008 8004
rect 7892 7964 7898 7976
rect 5696 7939 5754 7945
rect 5696 7905 5708 7939
rect 5742 7936 5754 7939
rect 6454 7936 6460 7948
rect 5742 7908 6460 7936
rect 5742 7905 5754 7908
rect 5696 7899 5754 7905
rect 6454 7896 6460 7908
rect 6512 7896 6518 7948
rect 10980 7945 11008 7976
rect 12250 7964 12256 8016
rect 12308 8004 12314 8016
rect 12618 8004 12624 8016
rect 12308 7976 12624 8004
rect 12308 7964 12314 7976
rect 12618 7964 12624 7976
rect 12676 8013 12682 8016
rect 12676 8007 12724 8013
rect 12676 7973 12678 8007
rect 12712 7973 12724 8007
rect 18230 8004 18236 8016
rect 18191 7976 18236 8004
rect 12676 7967 12724 7973
rect 12676 7964 12682 7967
rect 18230 7964 18236 7976
rect 18288 7964 18294 8016
rect 20806 7964 20812 8016
rect 20864 8004 20870 8016
rect 20901 8007 20959 8013
rect 20901 8004 20913 8007
rect 20864 7976 20913 8004
rect 20864 7964 20870 7976
rect 20901 7973 20913 7976
rect 20947 7973 20959 8007
rect 20901 7967 20959 7973
rect 10965 7939 11023 7945
rect 10965 7905 10977 7939
rect 11011 7905 11023 7939
rect 10965 7899 11023 7905
rect 1762 7868 1768 7880
rect 1723 7840 1768 7868
rect 1762 7828 1768 7840
rect 1820 7828 1826 7880
rect 3510 7828 3516 7880
rect 3568 7868 3574 7880
rect 4433 7871 4491 7877
rect 4433 7868 4445 7871
rect 3568 7840 4445 7868
rect 3568 7828 3574 7840
rect 4433 7837 4445 7840
rect 4479 7868 4491 7871
rect 7009 7871 7067 7877
rect 7009 7868 7021 7871
rect 4479 7840 7021 7868
rect 4479 7837 4491 7840
rect 4433 7831 4491 7837
rect 7009 7837 7021 7840
rect 7055 7868 7067 7871
rect 7098 7868 7104 7880
rect 7055 7840 7104 7868
rect 7055 7837 7067 7840
rect 7009 7831 7067 7837
rect 7098 7828 7104 7840
rect 7156 7828 7162 7880
rect 9769 7871 9827 7877
rect 9769 7837 9781 7871
rect 9815 7868 9827 7871
rect 10413 7871 10471 7877
rect 10413 7868 10425 7871
rect 9815 7840 10425 7868
rect 9815 7837 9827 7840
rect 9769 7831 9827 7837
rect 10413 7837 10425 7840
rect 10459 7868 10471 7871
rect 10502 7868 10508 7880
rect 10459 7840 10508 7868
rect 10459 7837 10471 7840
rect 10413 7831 10471 7837
rect 10502 7828 10508 7840
rect 10560 7828 10566 7880
rect 10980 7868 11008 7899
rect 11054 7896 11060 7948
rect 11112 7936 11118 7948
rect 11241 7939 11299 7945
rect 11241 7936 11253 7939
rect 11112 7908 11253 7936
rect 11112 7896 11118 7908
rect 11241 7905 11253 7908
rect 11287 7905 11299 7939
rect 15286 7936 15292 7948
rect 15247 7908 15292 7936
rect 11241 7899 11299 7905
rect 15286 7896 15292 7908
rect 15344 7896 15350 7948
rect 15746 7936 15752 7948
rect 15707 7908 15752 7936
rect 15746 7896 15752 7908
rect 15804 7896 15810 7948
rect 15930 7896 15936 7948
rect 15988 7936 15994 7948
rect 16117 7939 16175 7945
rect 16117 7936 16129 7939
rect 15988 7908 16129 7936
rect 15988 7896 15994 7908
rect 16117 7905 16129 7908
rect 16163 7905 16175 7939
rect 16117 7899 16175 7905
rect 16298 7896 16304 7948
rect 16356 7936 16362 7948
rect 16485 7939 16543 7945
rect 16485 7936 16497 7939
rect 16356 7908 16497 7936
rect 16356 7896 16362 7908
rect 16485 7905 16497 7908
rect 16531 7905 16543 7939
rect 16485 7899 16543 7905
rect 20714 7896 20720 7948
rect 20772 7936 20778 7948
rect 20993 7939 21051 7945
rect 20993 7936 21005 7939
rect 20772 7908 21005 7936
rect 20772 7896 20778 7908
rect 20993 7905 21005 7908
rect 21039 7905 21051 7939
rect 20993 7899 21051 7905
rect 11422 7868 11428 7880
rect 10980 7840 11428 7868
rect 11422 7828 11428 7840
rect 11480 7828 11486 7880
rect 11517 7871 11575 7877
rect 11517 7837 11529 7871
rect 11563 7868 11575 7871
rect 11790 7868 11796 7880
rect 11563 7840 11796 7868
rect 11563 7837 11575 7840
rect 11517 7831 11575 7837
rect 11790 7828 11796 7840
rect 11848 7868 11854 7880
rect 12345 7871 12403 7877
rect 12345 7868 12357 7871
rect 11848 7840 12357 7868
rect 11848 7828 11854 7840
rect 12345 7837 12357 7840
rect 12391 7837 12403 7871
rect 12345 7831 12403 7837
rect 18141 7871 18199 7877
rect 18141 7837 18153 7871
rect 18187 7868 18199 7871
rect 18782 7868 18788 7880
rect 18187 7840 18788 7868
rect 18187 7837 18199 7840
rect 18141 7831 18199 7837
rect 18782 7828 18788 7840
rect 18840 7828 18846 7880
rect 13262 7800 13268 7812
rect 13223 7772 13268 7800
rect 13262 7760 13268 7772
rect 13320 7760 13326 7812
rect 18690 7800 18696 7812
rect 18651 7772 18696 7800
rect 18690 7760 18696 7772
rect 18748 7760 18754 7812
rect 5767 7735 5825 7741
rect 5767 7701 5779 7735
rect 5813 7732 5825 7735
rect 6914 7732 6920 7744
rect 5813 7704 6920 7732
rect 5813 7701 5825 7704
rect 5767 7695 5825 7701
rect 6914 7692 6920 7704
rect 6972 7692 6978 7744
rect 8478 7692 8484 7744
rect 8536 7732 8542 7744
rect 8849 7735 8907 7741
rect 8849 7732 8861 7735
rect 8536 7704 8861 7732
rect 8536 7692 8542 7704
rect 8849 7701 8861 7704
rect 8895 7732 8907 7735
rect 9398 7732 9404 7744
rect 8895 7704 9404 7732
rect 8895 7701 8907 7704
rect 8849 7695 8907 7701
rect 9398 7692 9404 7704
rect 9456 7692 9462 7744
rect 13538 7732 13544 7744
rect 13499 7704 13544 7732
rect 13538 7692 13544 7704
rect 13596 7692 13602 7744
rect 1104 7642 22816 7664
rect 1104 7590 4982 7642
rect 5034 7590 5046 7642
rect 5098 7590 5110 7642
rect 5162 7590 5174 7642
rect 5226 7590 12982 7642
rect 13034 7590 13046 7642
rect 13098 7590 13110 7642
rect 13162 7590 13174 7642
rect 13226 7590 20982 7642
rect 21034 7590 21046 7642
rect 21098 7590 21110 7642
rect 21162 7590 21174 7642
rect 21226 7590 22816 7642
rect 1104 7568 22816 7590
rect 1762 7488 1768 7540
rect 1820 7528 1826 7540
rect 2869 7531 2927 7537
rect 2869 7528 2881 7531
rect 1820 7500 2881 7528
rect 1820 7488 1826 7500
rect 2869 7497 2881 7500
rect 2915 7497 2927 7531
rect 2869 7491 2927 7497
rect 6273 7531 6331 7537
rect 6273 7497 6285 7531
rect 6319 7528 6331 7531
rect 6454 7528 6460 7540
rect 6319 7500 6460 7528
rect 6319 7497 6331 7500
rect 6273 7491 6331 7497
rect 6454 7488 6460 7500
rect 6512 7528 6518 7540
rect 7650 7528 7656 7540
rect 6512 7500 7656 7528
rect 6512 7488 6518 7500
rect 7650 7488 7656 7500
rect 7708 7488 7714 7540
rect 8665 7531 8723 7537
rect 8665 7497 8677 7531
rect 8711 7528 8723 7531
rect 8846 7528 8852 7540
rect 8711 7500 8852 7528
rect 8711 7497 8723 7500
rect 8665 7491 8723 7497
rect 1854 7420 1860 7472
rect 1912 7420 1918 7472
rect 6380 7432 7420 7460
rect 1765 7395 1823 7401
rect 1765 7361 1777 7395
rect 1811 7392 1823 7395
rect 1872 7392 1900 7420
rect 2130 7392 2136 7404
rect 1811 7364 2136 7392
rect 1811 7361 1823 7364
rect 1765 7355 1823 7361
rect 2130 7352 2136 7364
rect 2188 7352 2194 7404
rect 2593 7395 2651 7401
rect 2593 7361 2605 7395
rect 2639 7392 2651 7395
rect 2958 7392 2964 7404
rect 2639 7364 2964 7392
rect 2639 7361 2651 7364
rect 2593 7355 2651 7361
rect 2958 7352 2964 7364
rect 3016 7352 3022 7404
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7392 4215 7395
rect 6380 7392 6408 7432
rect 7392 7404 7420 7432
rect 6914 7392 6920 7404
rect 4203 7364 6408 7392
rect 6875 7364 6920 7392
rect 4203 7361 4215 7364
rect 4157 7355 4215 7361
rect 6914 7352 6920 7364
rect 6972 7352 6978 7404
rect 7374 7392 7380 7404
rect 7335 7364 7380 7392
rect 7374 7352 7380 7364
rect 7432 7352 7438 7404
rect 4525 7327 4583 7333
rect 4525 7293 4537 7327
rect 4571 7324 4583 7327
rect 4706 7324 4712 7336
rect 4571 7296 4712 7324
rect 4571 7293 4583 7296
rect 4525 7287 4583 7293
rect 4706 7284 4712 7296
rect 4764 7324 4770 7336
rect 4985 7327 5043 7333
rect 4985 7324 4997 7327
rect 4764 7296 4997 7324
rect 4764 7284 4770 7296
rect 4985 7293 4997 7296
rect 5031 7293 5043 7327
rect 4985 7287 5043 7293
rect 5905 7327 5963 7333
rect 5905 7293 5917 7327
rect 5951 7324 5963 7327
rect 5951 7296 6684 7324
rect 5951 7293 5963 7296
rect 5905 7287 5963 7293
rect 1946 7256 1952 7268
rect 1907 7228 1952 7256
rect 1946 7216 1952 7228
rect 2004 7216 2010 7268
rect 2038 7216 2044 7268
rect 2096 7256 2102 7268
rect 3510 7256 3516 7268
rect 2096 7228 2141 7256
rect 3471 7228 3516 7256
rect 2096 7216 2102 7228
rect 3510 7216 3516 7228
rect 3568 7216 3574 7268
rect 3605 7259 3663 7265
rect 3605 7225 3617 7259
rect 3651 7225 3663 7259
rect 3605 7219 3663 7225
rect 4893 7259 4951 7265
rect 4893 7225 4905 7259
rect 4939 7256 4951 7259
rect 5347 7259 5405 7265
rect 5347 7256 5359 7259
rect 4939 7228 5359 7256
rect 4939 7225 4951 7228
rect 4893 7219 4951 7225
rect 5347 7225 5359 7228
rect 5393 7256 5405 7259
rect 5810 7256 5816 7268
rect 5393 7228 5816 7256
rect 5393 7225 5405 7228
rect 5347 7219 5405 7225
rect 3326 7188 3332 7200
rect 3239 7160 3332 7188
rect 3326 7148 3332 7160
rect 3384 7188 3390 7200
rect 3620 7188 3648 7219
rect 5810 7216 5816 7228
rect 5868 7216 5874 7268
rect 4246 7188 4252 7200
rect 3384 7160 4252 7188
rect 3384 7148 3390 7160
rect 4246 7148 4252 7160
rect 4304 7148 4310 7200
rect 6656 7197 6684 7296
rect 7558 7284 7564 7336
rect 7616 7324 7622 7336
rect 8772 7333 8800 7500
rect 8846 7488 8852 7500
rect 8904 7488 8910 7540
rect 10321 7531 10379 7537
rect 10321 7497 10333 7531
rect 10367 7528 10379 7531
rect 11054 7528 11060 7540
rect 10367 7500 11060 7528
rect 10367 7497 10379 7500
rect 10321 7491 10379 7497
rect 9493 7395 9551 7401
rect 9493 7361 9505 7395
rect 9539 7392 9551 7395
rect 10336 7392 10364 7491
rect 11054 7488 11060 7500
rect 11112 7488 11118 7540
rect 11422 7528 11428 7540
rect 11383 7500 11428 7528
rect 11422 7488 11428 7500
rect 11480 7488 11486 7540
rect 11790 7528 11796 7540
rect 11751 7500 11796 7528
rect 11790 7488 11796 7500
rect 11848 7488 11854 7540
rect 12618 7528 12624 7540
rect 12579 7500 12624 7528
rect 12618 7488 12624 7500
rect 12676 7488 12682 7540
rect 15930 7488 15936 7540
rect 15988 7528 15994 7540
rect 16025 7531 16083 7537
rect 16025 7528 16037 7531
rect 15988 7500 16037 7528
rect 15988 7488 15994 7500
rect 16025 7497 16037 7500
rect 16071 7497 16083 7531
rect 16025 7491 16083 7497
rect 17083 7531 17141 7537
rect 17083 7497 17095 7531
rect 17129 7528 17141 7531
rect 17954 7528 17960 7540
rect 17129 7500 17960 7528
rect 17129 7497 17141 7500
rect 17083 7491 17141 7497
rect 17954 7488 17960 7500
rect 18012 7488 18018 7540
rect 21085 7531 21143 7537
rect 21085 7497 21097 7531
rect 21131 7528 21143 7531
rect 21266 7528 21272 7540
rect 21131 7500 21272 7528
rect 21131 7497 21143 7500
rect 21085 7491 21143 7497
rect 21266 7488 21272 7500
rect 21324 7488 21330 7540
rect 13446 7460 13452 7472
rect 13407 7432 13452 7460
rect 13446 7420 13452 7432
rect 13504 7420 13510 7472
rect 15381 7463 15439 7469
rect 15381 7429 15393 7463
rect 15427 7460 15439 7463
rect 16298 7460 16304 7472
rect 15427 7432 16304 7460
rect 15427 7429 15439 7432
rect 15381 7423 15439 7429
rect 16298 7420 16304 7432
rect 16356 7420 16362 7472
rect 18230 7420 18236 7472
rect 18288 7460 18294 7472
rect 19058 7460 19064 7472
rect 18288 7432 19064 7460
rect 18288 7420 18294 7432
rect 19058 7420 19064 7432
rect 19116 7460 19122 7472
rect 19245 7463 19303 7469
rect 19245 7460 19257 7463
rect 19116 7432 19257 7460
rect 19116 7420 19122 7432
rect 19245 7429 19257 7432
rect 19291 7429 19303 7463
rect 19245 7423 19303 7429
rect 20714 7420 20720 7472
rect 20772 7460 20778 7472
rect 21453 7463 21511 7469
rect 21453 7460 21465 7463
rect 20772 7432 21465 7460
rect 20772 7420 20778 7432
rect 21453 7429 21465 7432
rect 21499 7429 21511 7463
rect 21453 7423 21511 7429
rect 10502 7392 10508 7404
rect 9539 7364 10364 7392
rect 10463 7364 10508 7392
rect 9539 7361 9551 7364
rect 9493 7355 9551 7361
rect 10502 7352 10508 7364
rect 10560 7352 10566 7404
rect 10962 7392 10968 7404
rect 10923 7364 10968 7392
rect 10962 7352 10968 7364
rect 11020 7352 11026 7404
rect 12253 7395 12311 7401
rect 12253 7361 12265 7395
rect 12299 7392 12311 7395
rect 13262 7392 13268 7404
rect 12299 7364 13268 7392
rect 12299 7361 12311 7364
rect 12253 7355 12311 7361
rect 13262 7352 13268 7364
rect 13320 7352 13326 7404
rect 14550 7352 14556 7404
rect 14608 7392 14614 7404
rect 18325 7395 18383 7401
rect 14608 7364 16389 7392
rect 14608 7352 14614 7364
rect 8757 7327 8815 7333
rect 8757 7324 8769 7327
rect 7616 7296 8769 7324
rect 7616 7284 7622 7296
rect 8757 7293 8769 7296
rect 8803 7293 8815 7327
rect 8757 7287 8815 7293
rect 8846 7284 8852 7336
rect 8904 7324 8910 7336
rect 9033 7327 9091 7333
rect 8904 7296 8949 7324
rect 8904 7284 8910 7296
rect 9033 7293 9045 7327
rect 9079 7324 9091 7327
rect 9398 7324 9404 7336
rect 9079 7296 9404 7324
rect 9079 7293 9091 7296
rect 9033 7287 9091 7293
rect 9398 7284 9404 7296
rect 9456 7284 9462 7336
rect 9953 7327 10011 7333
rect 9953 7293 9965 7327
rect 9999 7324 10011 7327
rect 10226 7324 10232 7336
rect 9999 7296 10232 7324
rect 9999 7293 10011 7296
rect 9953 7287 10011 7293
rect 10226 7284 10232 7296
rect 10284 7284 10290 7336
rect 14826 7284 14832 7336
rect 14884 7324 14890 7336
rect 14921 7327 14979 7333
rect 14921 7324 14933 7327
rect 14884 7296 14933 7324
rect 14884 7284 14890 7296
rect 14921 7293 14933 7296
rect 14967 7293 14979 7327
rect 14921 7287 14979 7293
rect 15286 7284 15292 7336
rect 15344 7324 15350 7336
rect 15657 7327 15715 7333
rect 15657 7324 15669 7327
rect 15344 7296 15669 7324
rect 15344 7284 15350 7296
rect 15657 7293 15669 7296
rect 15703 7293 15715 7327
rect 16361 7324 16389 7364
rect 18325 7361 18337 7395
rect 18371 7392 18383 7395
rect 18966 7392 18972 7404
rect 18371 7364 18972 7392
rect 18371 7361 18383 7364
rect 18325 7355 18383 7361
rect 18966 7352 18972 7364
rect 19024 7392 19030 7404
rect 19613 7395 19671 7401
rect 19613 7392 19625 7395
rect 19024 7364 19625 7392
rect 19024 7352 19030 7364
rect 19613 7361 19625 7364
rect 19659 7361 19671 7395
rect 19613 7355 19671 7361
rect 16980 7327 17038 7333
rect 16980 7324 16992 7327
rect 16361 7296 16992 7324
rect 15657 7287 15715 7293
rect 16980 7293 16992 7296
rect 17026 7324 17038 7327
rect 17405 7327 17463 7333
rect 17405 7324 17417 7327
rect 17026 7296 17417 7324
rect 17026 7293 17038 7296
rect 16980 7287 17038 7293
rect 17405 7293 17417 7296
rect 17451 7293 17463 7327
rect 17405 7287 17463 7293
rect 19935 7327 19993 7333
rect 19935 7293 19947 7327
rect 19981 7293 19993 7327
rect 19935 7287 19993 7293
rect 20901 7327 20959 7333
rect 20901 7293 20913 7327
rect 20947 7293 20959 7327
rect 20901 7287 20959 7293
rect 7009 7259 7067 7265
rect 7009 7225 7021 7259
rect 7055 7225 7067 7259
rect 7009 7219 7067 7225
rect 8297 7259 8355 7265
rect 8297 7225 8309 7259
rect 8343 7256 8355 7259
rect 8662 7256 8668 7268
rect 8343 7228 8668 7256
rect 8343 7225 8355 7228
rect 8297 7219 8355 7225
rect 6641 7191 6699 7197
rect 6641 7157 6653 7191
rect 6687 7188 6699 7191
rect 6730 7188 6736 7200
rect 6687 7160 6736 7188
rect 6687 7157 6699 7160
rect 6641 7151 6699 7157
rect 6730 7148 6736 7160
rect 6788 7188 6794 7200
rect 7024 7188 7052 7219
rect 8662 7216 8668 7228
rect 8720 7256 8726 7268
rect 8864 7256 8892 7284
rect 8720 7228 8892 7256
rect 10244 7256 10272 7284
rect 10597 7259 10655 7265
rect 10597 7256 10609 7259
rect 10244 7228 10609 7256
rect 8720 7216 8726 7228
rect 10597 7225 10609 7228
rect 10643 7225 10655 7259
rect 12894 7256 12900 7268
rect 12855 7228 12900 7256
rect 10597 7219 10655 7225
rect 12894 7216 12900 7228
rect 12952 7216 12958 7268
rect 12989 7259 13047 7265
rect 12989 7225 13001 7259
rect 13035 7256 13047 7259
rect 13262 7256 13268 7268
rect 13035 7228 13268 7256
rect 13035 7225 13047 7228
rect 12989 7219 13047 7225
rect 13262 7216 13268 7228
rect 13320 7216 13326 7268
rect 18414 7216 18420 7268
rect 18472 7256 18478 7268
rect 18472 7228 18517 7256
rect 18472 7216 18478 7228
rect 18690 7216 18696 7268
rect 18748 7256 18754 7268
rect 18969 7259 19027 7265
rect 18969 7256 18981 7259
rect 18748 7228 18981 7256
rect 18748 7216 18754 7228
rect 18969 7225 18981 7228
rect 19015 7225 19027 7259
rect 18969 7219 19027 7225
rect 7837 7191 7895 7197
rect 7837 7188 7849 7191
rect 6788 7160 7849 7188
rect 6788 7148 6794 7160
rect 7837 7157 7849 7160
rect 7883 7157 7895 7191
rect 7837 7151 7895 7157
rect 17865 7191 17923 7197
rect 17865 7157 17877 7191
rect 17911 7188 17923 7191
rect 18432 7188 18460 7216
rect 17911 7160 18460 7188
rect 19950 7188 19978 7287
rect 20027 7259 20085 7265
rect 20027 7225 20039 7259
rect 20073 7256 20085 7259
rect 20717 7259 20775 7265
rect 20717 7256 20729 7259
rect 20073 7228 20729 7256
rect 20073 7225 20085 7228
rect 20027 7219 20085 7225
rect 20717 7225 20729 7228
rect 20763 7256 20775 7259
rect 20916 7256 20944 7287
rect 20763 7228 20944 7256
rect 20763 7225 20775 7228
rect 20717 7219 20775 7225
rect 20441 7191 20499 7197
rect 20441 7188 20453 7191
rect 19950 7160 20453 7188
rect 17911 7157 17923 7160
rect 17865 7151 17923 7157
rect 20441 7157 20453 7160
rect 20487 7188 20499 7191
rect 20806 7188 20812 7200
rect 20487 7160 20812 7188
rect 20487 7157 20499 7160
rect 20441 7151 20499 7157
rect 20806 7148 20812 7160
rect 20864 7148 20870 7200
rect 1104 7098 22816 7120
rect 1104 7046 8982 7098
rect 9034 7046 9046 7098
rect 9098 7046 9110 7098
rect 9162 7046 9174 7098
rect 9226 7046 16982 7098
rect 17034 7046 17046 7098
rect 17098 7046 17110 7098
rect 17162 7046 17174 7098
rect 17226 7046 22816 7098
rect 1104 7024 22816 7046
rect 1578 6984 1584 6996
rect 1539 6956 1584 6984
rect 1578 6944 1584 6956
rect 1636 6944 1642 6996
rect 1946 6984 1952 6996
rect 1907 6956 1952 6984
rect 1946 6944 1952 6956
rect 2004 6984 2010 6996
rect 2501 6987 2559 6993
rect 2501 6984 2513 6987
rect 2004 6956 2513 6984
rect 2004 6944 2010 6956
rect 2501 6953 2513 6956
rect 2547 6953 2559 6987
rect 3878 6984 3884 6996
rect 3839 6956 3884 6984
rect 2501 6947 2559 6953
rect 3878 6944 3884 6956
rect 3936 6944 3942 6996
rect 4246 6984 4252 6996
rect 4207 6956 4252 6984
rect 4246 6944 4252 6956
rect 4304 6944 4310 6996
rect 4706 6984 4712 6996
rect 4667 6956 4712 6984
rect 4706 6944 4712 6956
rect 4764 6944 4770 6996
rect 6914 6944 6920 6996
rect 6972 6984 6978 6996
rect 7561 6987 7619 6993
rect 7561 6984 7573 6987
rect 6972 6956 7573 6984
rect 6972 6944 6978 6956
rect 7561 6953 7573 6956
rect 7607 6953 7619 6987
rect 7561 6947 7619 6953
rect 14645 6987 14703 6993
rect 14645 6953 14657 6987
rect 14691 6984 14703 6987
rect 14826 6984 14832 6996
rect 14691 6956 14832 6984
rect 14691 6953 14703 6956
rect 14645 6947 14703 6953
rect 14826 6944 14832 6956
rect 14884 6984 14890 6996
rect 15746 6984 15752 6996
rect 14884 6956 15752 6984
rect 14884 6944 14890 6956
rect 15746 6944 15752 6956
rect 15804 6984 15810 6996
rect 15804 6956 15884 6984
rect 15804 6944 15810 6956
rect 2038 6876 2044 6928
rect 2096 6916 2102 6928
rect 2409 6919 2467 6925
rect 2409 6916 2421 6919
rect 2096 6888 2421 6916
rect 2096 6876 2102 6888
rect 2409 6885 2421 6888
rect 2455 6916 2467 6919
rect 3326 6916 3332 6928
rect 2455 6888 3332 6916
rect 2455 6885 2467 6888
rect 2409 6879 2467 6885
rect 3326 6876 3332 6888
rect 3384 6876 3390 6928
rect 6457 6919 6515 6925
rect 6457 6885 6469 6919
rect 6503 6916 6515 6919
rect 6730 6916 6736 6928
rect 6503 6888 6736 6916
rect 6503 6885 6515 6888
rect 6457 6879 6515 6885
rect 6730 6876 6736 6888
rect 6788 6876 6794 6928
rect 8754 6916 8760 6928
rect 8623 6888 8760 6916
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 2866 6848 2872 6860
rect 1443 6820 2872 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 2866 6808 2872 6820
rect 2924 6808 2930 6860
rect 4522 6848 4528 6860
rect 4483 6820 4528 6848
rect 4522 6808 4528 6820
rect 4580 6808 4586 6860
rect 4798 6808 4804 6860
rect 4856 6848 4862 6860
rect 4985 6851 5043 6857
rect 4985 6848 4997 6851
rect 4856 6820 4997 6848
rect 4856 6808 4862 6820
rect 4985 6817 4997 6820
rect 5031 6848 5043 6851
rect 5626 6848 5632 6860
rect 5031 6820 5632 6848
rect 5031 6817 5043 6820
rect 4985 6811 5043 6817
rect 5626 6808 5632 6820
rect 5684 6808 5690 6860
rect 8623 6857 8651 6888
rect 8754 6876 8760 6888
rect 8812 6876 8818 6928
rect 10318 6916 10324 6928
rect 10279 6888 10324 6916
rect 10318 6876 10324 6888
rect 10376 6876 10382 6928
rect 12342 6916 12348 6928
rect 12303 6888 12348 6916
rect 12342 6876 12348 6888
rect 12400 6876 12406 6928
rect 8608 6851 8666 6857
rect 8608 6817 8620 6851
rect 8654 6817 8666 6851
rect 8608 6811 8666 6817
rect 13776 6851 13834 6857
rect 13776 6817 13788 6851
rect 13822 6848 13834 6851
rect 13998 6848 14004 6860
rect 13822 6820 14004 6848
rect 13822 6817 13834 6820
rect 13776 6811 13834 6817
rect 13998 6808 14004 6820
rect 14056 6808 14062 6860
rect 15286 6848 15292 6860
rect 15247 6820 15292 6848
rect 15286 6808 15292 6820
rect 15344 6808 15350 6860
rect 15856 6857 15884 6956
rect 18230 6944 18236 6996
rect 18288 6984 18294 6996
rect 18509 6987 18567 6993
rect 18509 6984 18521 6987
rect 18288 6956 18521 6984
rect 18288 6944 18294 6956
rect 18509 6953 18521 6956
rect 18555 6953 18567 6987
rect 18782 6984 18788 6996
rect 18743 6956 18788 6984
rect 18509 6947 18567 6953
rect 18782 6944 18788 6956
rect 18840 6944 18846 6996
rect 17678 6876 17684 6928
rect 17736 6916 17742 6928
rect 17910 6919 17968 6925
rect 17910 6916 17922 6919
rect 17736 6888 17922 6916
rect 17736 6876 17742 6888
rect 17910 6885 17922 6888
rect 17956 6885 17968 6919
rect 17910 6879 17968 6885
rect 20530 6876 20536 6928
rect 20588 6916 20594 6928
rect 20993 6919 21051 6925
rect 20993 6916 21005 6919
rect 20588 6888 21005 6916
rect 20588 6876 20594 6888
rect 20993 6885 21005 6888
rect 21039 6885 21051 6919
rect 20993 6879 21051 6885
rect 21085 6919 21143 6925
rect 21085 6885 21097 6919
rect 21131 6916 21143 6919
rect 21450 6916 21456 6928
rect 21131 6888 21456 6916
rect 21131 6885 21143 6888
rect 21085 6879 21143 6885
rect 21450 6876 21456 6888
rect 21508 6876 21514 6928
rect 15841 6851 15899 6857
rect 15841 6817 15853 6851
rect 15887 6817 15899 6851
rect 15841 6811 15899 6817
rect 15930 6808 15936 6860
rect 15988 6848 15994 6860
rect 16117 6851 16175 6857
rect 16117 6848 16129 6851
rect 15988 6820 16129 6848
rect 15988 6808 15994 6820
rect 16117 6817 16129 6820
rect 16163 6817 16175 6851
rect 16482 6848 16488 6860
rect 16443 6820 16488 6848
rect 16117 6811 16175 6817
rect 16482 6808 16488 6820
rect 16540 6808 16546 6860
rect 19702 6848 19708 6860
rect 19663 6820 19708 6848
rect 19702 6808 19708 6820
rect 19760 6808 19766 6860
rect 6089 6783 6147 6789
rect 6089 6749 6101 6783
rect 6135 6780 6147 6783
rect 6638 6780 6644 6792
rect 6135 6752 6644 6780
rect 6135 6749 6147 6752
rect 6089 6743 6147 6749
rect 6638 6740 6644 6752
rect 6696 6740 6702 6792
rect 7006 6780 7012 6792
rect 6967 6752 7012 6780
rect 7006 6740 7012 6752
rect 7064 6740 7070 6792
rect 8711 6783 8769 6789
rect 8711 6749 8723 6783
rect 8757 6780 8769 6783
rect 10229 6783 10287 6789
rect 10229 6780 10241 6783
rect 8757 6752 10241 6780
rect 8757 6749 8769 6752
rect 8711 6743 8769 6749
rect 10229 6749 10241 6752
rect 10275 6780 10287 6783
rect 11054 6780 11060 6792
rect 10275 6752 11060 6780
rect 10275 6749 10287 6752
rect 10229 6743 10287 6749
rect 11054 6740 11060 6752
rect 11112 6740 11118 6792
rect 12250 6780 12256 6792
rect 12163 6752 12256 6780
rect 12250 6740 12256 6752
rect 12308 6780 12314 6792
rect 13863 6783 13921 6789
rect 13863 6780 13875 6783
rect 12308 6752 13875 6780
rect 12308 6740 12314 6752
rect 13863 6749 13875 6752
rect 13909 6749 13921 6783
rect 16758 6780 16764 6792
rect 16719 6752 16764 6780
rect 13863 6743 13921 6749
rect 16758 6740 16764 6752
rect 16816 6780 16822 6792
rect 17589 6783 17647 6789
rect 17589 6780 17601 6783
rect 16816 6752 17601 6780
rect 16816 6740 16822 6752
rect 17589 6749 17601 6752
rect 17635 6749 17647 6783
rect 21266 6780 21272 6792
rect 21227 6752 21272 6780
rect 17589 6743 17647 6749
rect 21266 6740 21272 6752
rect 21324 6740 21330 6792
rect 10778 6712 10784 6724
rect 10739 6684 10784 6712
rect 10778 6672 10784 6684
rect 10836 6712 10842 6724
rect 12805 6715 12863 6721
rect 12805 6712 12817 6715
rect 10836 6684 12817 6712
rect 10836 6672 10842 6684
rect 12805 6681 12817 6684
rect 12851 6712 12863 6715
rect 12894 6712 12900 6724
rect 12851 6684 12900 6712
rect 12851 6681 12863 6684
rect 12805 6675 12863 6681
rect 12894 6672 12900 6684
rect 12952 6712 12958 6724
rect 13173 6715 13231 6721
rect 13173 6712 13185 6715
rect 12952 6684 13185 6712
rect 12952 6672 12958 6684
rect 13173 6681 13185 6684
rect 13219 6681 13231 6715
rect 13173 6675 13231 6681
rect 14550 6672 14556 6724
rect 14608 6712 14614 6724
rect 19518 6712 19524 6724
rect 14608 6684 19524 6712
rect 14608 6672 14614 6684
rect 19518 6672 19524 6684
rect 19576 6672 19582 6724
rect 3510 6644 3516 6656
rect 3471 6616 3516 6644
rect 3510 6604 3516 6616
rect 3568 6604 3574 6656
rect 5350 6604 5356 6656
rect 5408 6644 5414 6656
rect 5445 6647 5503 6653
rect 5445 6644 5457 6647
rect 5408 6616 5457 6644
rect 5408 6604 5414 6616
rect 5445 6613 5457 6616
rect 5491 6613 5503 6647
rect 14182 6644 14188 6656
rect 14143 6616 14188 6644
rect 5445 6607 5503 6613
rect 14182 6604 14188 6616
rect 14240 6604 14246 6656
rect 16390 6604 16396 6656
rect 16448 6644 16454 6656
rect 19935 6647 19993 6653
rect 19935 6644 19947 6647
rect 16448 6616 19947 6644
rect 16448 6604 16454 6616
rect 19935 6613 19947 6616
rect 19981 6613 19993 6647
rect 19935 6607 19993 6613
rect 1104 6554 22816 6576
rect 1104 6502 4982 6554
rect 5034 6502 5046 6554
rect 5098 6502 5110 6554
rect 5162 6502 5174 6554
rect 5226 6502 12982 6554
rect 13034 6502 13046 6554
rect 13098 6502 13110 6554
rect 13162 6502 13174 6554
rect 13226 6502 20982 6554
rect 21034 6502 21046 6554
rect 21098 6502 21110 6554
rect 21162 6502 21174 6554
rect 21226 6502 22816 6554
rect 1104 6480 22816 6502
rect 3099 6443 3157 6449
rect 3099 6409 3111 6443
rect 3145 6440 3157 6443
rect 3602 6440 3608 6452
rect 3145 6412 3608 6440
rect 3145 6409 3157 6412
rect 3099 6403 3157 6409
rect 3602 6400 3608 6412
rect 3660 6400 3666 6452
rect 4341 6443 4399 6449
rect 4341 6409 4353 6443
rect 4387 6440 4399 6443
rect 4522 6440 4528 6452
rect 4387 6412 4528 6440
rect 4387 6409 4399 6412
rect 4341 6403 4399 6409
rect 4522 6400 4528 6412
rect 4580 6400 4586 6452
rect 4706 6400 4712 6452
rect 4764 6440 4770 6452
rect 7929 6443 7987 6449
rect 7929 6440 7941 6443
rect 4764 6412 7941 6440
rect 4764 6400 4770 6412
rect 3973 6375 4031 6381
rect 3973 6341 3985 6375
rect 4019 6372 4031 6375
rect 4798 6372 4804 6384
rect 4019 6344 4804 6372
rect 4019 6341 4031 6344
rect 3973 6335 4031 6341
rect 4798 6332 4804 6344
rect 4856 6332 4862 6384
rect 5077 6375 5135 6381
rect 5077 6341 5089 6375
rect 5123 6372 5135 6375
rect 5261 6375 5319 6381
rect 5261 6372 5273 6375
rect 5123 6344 5273 6372
rect 5123 6341 5135 6344
rect 5077 6335 5135 6341
rect 5261 6341 5273 6344
rect 5307 6372 5319 6375
rect 6546 6372 6552 6384
rect 5307 6344 6552 6372
rect 5307 6341 5319 6344
rect 5261 6335 5319 6341
rect 2866 6304 2872 6316
rect 2827 6276 2872 6304
rect 2866 6264 2872 6276
rect 2924 6264 2930 6316
rect 2041 6239 2099 6245
rect 2041 6205 2053 6239
rect 2087 6205 2099 6239
rect 2041 6199 2099 6205
rect 2056 6168 2084 6199
rect 2130 6196 2136 6248
rect 2188 6236 2194 6248
rect 3028 6239 3086 6245
rect 3028 6236 3040 6239
rect 2188 6208 3040 6236
rect 2188 6196 2194 6208
rect 3028 6205 3040 6208
rect 3074 6236 3086 6239
rect 3421 6239 3479 6245
rect 3421 6236 3433 6239
rect 3074 6208 3433 6236
rect 3074 6205 3086 6208
rect 3028 6199 3086 6205
rect 3421 6205 3433 6208
rect 3467 6205 3479 6239
rect 3421 6199 3479 6205
rect 2056 6140 2452 6168
rect 2424 6112 2452 6140
rect 2682 6128 2688 6180
rect 2740 6168 2746 6180
rect 5092 6168 5120 6335
rect 6546 6332 6552 6344
rect 6604 6332 6610 6384
rect 6932 6381 6960 6412
rect 7929 6409 7941 6412
rect 7975 6440 7987 6443
rect 8662 6440 8668 6452
rect 7975 6412 8668 6440
rect 7975 6409 7987 6412
rect 7929 6403 7987 6409
rect 8662 6400 8668 6412
rect 8720 6400 8726 6452
rect 8754 6400 8760 6452
rect 8812 6440 8818 6452
rect 9401 6443 9459 6449
rect 9401 6440 9413 6443
rect 8812 6412 9413 6440
rect 8812 6400 8818 6412
rect 9401 6409 9413 6412
rect 9447 6409 9459 6443
rect 9401 6403 9459 6409
rect 9953 6443 10011 6449
rect 9953 6409 9965 6443
rect 9999 6440 10011 6443
rect 10318 6440 10324 6452
rect 9999 6412 10324 6440
rect 9999 6409 10011 6412
rect 9953 6403 10011 6409
rect 10318 6400 10324 6412
rect 10376 6400 10382 6452
rect 11054 6440 11060 6452
rect 11015 6412 11060 6440
rect 11054 6400 11060 6412
rect 11112 6400 11118 6452
rect 11885 6443 11943 6449
rect 11885 6409 11897 6443
rect 11931 6440 11943 6443
rect 12253 6443 12311 6449
rect 12253 6440 12265 6443
rect 11931 6412 12265 6440
rect 11931 6409 11943 6412
rect 11885 6403 11943 6409
rect 12253 6409 12265 6412
rect 12299 6440 12311 6443
rect 12342 6440 12348 6452
rect 12299 6412 12348 6440
rect 12299 6409 12311 6412
rect 12253 6403 12311 6409
rect 12342 6400 12348 6412
rect 12400 6400 12406 6452
rect 13633 6443 13691 6449
rect 13633 6409 13645 6443
rect 13679 6440 13691 6443
rect 13998 6440 14004 6452
rect 13679 6412 14004 6440
rect 13679 6409 13691 6412
rect 13633 6403 13691 6409
rect 13998 6400 14004 6412
rect 14056 6400 14062 6452
rect 15746 6400 15752 6452
rect 15804 6440 15810 6452
rect 16393 6443 16451 6449
rect 16393 6440 16405 6443
rect 15804 6412 16405 6440
rect 15804 6400 15810 6412
rect 16393 6409 16405 6412
rect 16439 6409 16451 6443
rect 16758 6440 16764 6452
rect 16719 6412 16764 6440
rect 16393 6403 16451 6409
rect 16758 6400 16764 6412
rect 16816 6400 16822 6452
rect 17678 6400 17684 6452
rect 17736 6440 17742 6452
rect 17773 6443 17831 6449
rect 17773 6440 17785 6443
rect 17736 6412 17785 6440
rect 17736 6400 17742 6412
rect 17773 6409 17785 6412
rect 17819 6409 17831 6443
rect 17773 6403 17831 6409
rect 18325 6443 18383 6449
rect 18325 6409 18337 6443
rect 18371 6440 18383 6443
rect 18414 6440 18420 6452
rect 18371 6412 18420 6440
rect 18371 6409 18383 6412
rect 18325 6403 18383 6409
rect 18414 6400 18420 6412
rect 18472 6400 18478 6452
rect 19058 6440 19064 6452
rect 19019 6412 19064 6440
rect 19058 6400 19064 6412
rect 19116 6400 19122 6452
rect 20530 6400 20536 6452
rect 20588 6440 20594 6452
rect 21821 6443 21879 6449
rect 21821 6440 21833 6443
rect 20588 6412 21833 6440
rect 20588 6400 20594 6412
rect 21821 6409 21833 6412
rect 21867 6409 21879 6443
rect 21821 6403 21879 6409
rect 6917 6375 6975 6381
rect 6917 6341 6929 6375
rect 6963 6341 6975 6375
rect 6917 6335 6975 6341
rect 14185 6375 14243 6381
rect 14185 6341 14197 6375
rect 14231 6372 14243 6375
rect 14826 6372 14832 6384
rect 14231 6344 14832 6372
rect 14231 6341 14243 6344
rect 14185 6335 14243 6341
rect 14826 6332 14832 6344
rect 14884 6332 14890 6384
rect 16117 6375 16175 6381
rect 16117 6341 16129 6375
rect 16163 6372 16175 6375
rect 16482 6372 16488 6384
rect 16163 6344 16488 6372
rect 16163 6341 16175 6344
rect 16117 6335 16175 6341
rect 16482 6332 16488 6344
rect 16540 6332 16546 6384
rect 19702 6332 19708 6384
rect 19760 6372 19766 6384
rect 19889 6375 19947 6381
rect 19889 6372 19901 6375
rect 19760 6344 19901 6372
rect 19760 6332 19766 6344
rect 19889 6341 19901 6344
rect 19935 6372 19947 6375
rect 21358 6372 21364 6384
rect 19935 6344 21364 6372
rect 19935 6341 19947 6344
rect 19889 6335 19947 6341
rect 21358 6332 21364 6344
rect 21416 6332 21422 6384
rect 21450 6332 21456 6384
rect 21508 6372 21514 6384
rect 21508 6344 21553 6372
rect 21508 6332 21514 6344
rect 5350 6304 5356 6316
rect 5184 6276 5356 6304
rect 5184 6245 5212 6276
rect 5350 6264 5356 6276
rect 5408 6264 5414 6316
rect 5626 6264 5632 6316
rect 5684 6304 5690 6316
rect 7285 6307 7343 6313
rect 7285 6304 7297 6307
rect 5684 6276 7297 6304
rect 5684 6264 5690 6276
rect 7285 6273 7297 6276
rect 7331 6273 7343 6307
rect 10778 6304 10784 6316
rect 10739 6276 10784 6304
rect 7285 6267 7343 6273
rect 10778 6264 10784 6276
rect 10836 6264 10842 6316
rect 10962 6264 10968 6316
rect 11020 6304 11026 6316
rect 12897 6307 12955 6313
rect 12897 6304 12909 6307
rect 11020 6276 12909 6304
rect 11020 6264 11026 6276
rect 12897 6273 12909 6276
rect 12943 6304 12955 6307
rect 13538 6304 13544 6316
rect 12943 6276 13544 6304
rect 12943 6273 12955 6276
rect 12897 6267 12955 6273
rect 13538 6264 13544 6276
rect 13596 6264 13602 6316
rect 13630 6264 13636 6316
rect 13688 6304 13694 6316
rect 15749 6307 15807 6313
rect 13688 6276 14412 6304
rect 13688 6264 13694 6276
rect 5169 6239 5227 6245
rect 5169 6205 5181 6239
rect 5215 6205 5227 6239
rect 5169 6199 5227 6205
rect 5445 6239 5503 6245
rect 5445 6205 5457 6239
rect 5491 6205 5503 6239
rect 5445 6199 5503 6205
rect 6273 6239 6331 6245
rect 6273 6205 6285 6239
rect 6319 6236 6331 6239
rect 6825 6239 6883 6245
rect 6825 6236 6837 6239
rect 6319 6208 6837 6236
rect 6319 6205 6331 6208
rect 6273 6199 6331 6205
rect 6825 6205 6837 6208
rect 6871 6236 6883 6239
rect 6914 6236 6920 6248
rect 6871 6208 6920 6236
rect 6871 6205 6883 6208
rect 6825 6199 6883 6205
rect 2740 6140 5120 6168
rect 2740 6128 2746 6140
rect 5460 6112 5488 6199
rect 6914 6196 6920 6208
rect 6972 6196 6978 6248
rect 7098 6236 7104 6248
rect 7059 6208 7104 6236
rect 7098 6196 7104 6208
rect 7156 6236 7162 6248
rect 8018 6236 8024 6248
rect 7156 6208 8024 6236
rect 7156 6196 7162 6208
rect 8018 6196 8024 6208
rect 8076 6196 8082 6248
rect 8481 6239 8539 6245
rect 8481 6236 8493 6239
rect 8220 6208 8493 6236
rect 5905 6171 5963 6177
rect 5905 6137 5917 6171
rect 5951 6168 5963 6171
rect 7558 6168 7564 6180
rect 5951 6140 7564 6168
rect 5951 6137 5963 6140
rect 5905 6131 5963 6137
rect 7558 6128 7564 6140
rect 7616 6128 7622 6180
rect 8220 6112 8248 6208
rect 8481 6205 8493 6208
rect 8527 6205 8539 6239
rect 8481 6199 8539 6205
rect 14093 6239 14151 6245
rect 14093 6205 14105 6239
rect 14139 6236 14151 6239
rect 14182 6236 14188 6248
rect 14139 6208 14188 6236
rect 14139 6205 14151 6208
rect 14093 6199 14151 6205
rect 14182 6196 14188 6208
rect 14240 6196 14246 6248
rect 14384 6245 14412 6276
rect 15749 6273 15761 6307
rect 15795 6304 15807 6307
rect 15930 6304 15936 6316
rect 15795 6276 15936 6304
rect 15795 6273 15807 6276
rect 15749 6267 15807 6273
rect 15930 6264 15936 6276
rect 15988 6264 15994 6316
rect 16500 6304 16528 6332
rect 16758 6304 16764 6316
rect 16500 6276 16764 6304
rect 16758 6264 16764 6276
rect 16816 6264 16822 6316
rect 20530 6304 20536 6316
rect 20443 6276 20536 6304
rect 20530 6264 20536 6276
rect 20588 6304 20594 6316
rect 21266 6304 21272 6316
rect 20588 6276 21272 6304
rect 20588 6264 20594 6276
rect 21266 6264 21272 6276
rect 21324 6264 21330 6316
rect 14369 6239 14427 6245
rect 14369 6205 14381 6239
rect 14415 6205 14427 6239
rect 14369 6199 14427 6205
rect 14829 6239 14887 6245
rect 14829 6205 14841 6239
rect 14875 6236 14887 6239
rect 15838 6236 15844 6248
rect 14875 6208 15844 6236
rect 14875 6205 14887 6208
rect 14829 6199 14887 6205
rect 10134 6168 10140 6180
rect 10095 6140 10140 6168
rect 10134 6128 10140 6140
rect 10192 6128 10198 6180
rect 10226 6128 10232 6180
rect 10284 6168 10290 6180
rect 12618 6168 12624 6180
rect 10284 6140 10329 6168
rect 12579 6140 12624 6168
rect 10284 6128 10290 6140
rect 12618 6128 12624 6140
rect 12676 6128 12682 6180
rect 12713 6171 12771 6177
rect 12713 6137 12725 6171
rect 12759 6137 12771 6171
rect 12713 6131 12771 6137
rect 1670 6100 1676 6112
rect 1631 6072 1676 6100
rect 1670 6060 1676 6072
rect 1728 6060 1734 6112
rect 2406 6100 2412 6112
rect 2367 6072 2412 6100
rect 2406 6060 2412 6072
rect 2464 6060 2470 6112
rect 4709 6103 4767 6109
rect 4709 6069 4721 6103
rect 4755 6100 4767 6103
rect 5442 6100 5448 6112
rect 4755 6072 5448 6100
rect 4755 6069 4767 6072
rect 4709 6063 4767 6069
rect 5442 6060 5448 6072
rect 5500 6060 5506 6112
rect 6362 6060 6368 6112
rect 6420 6100 6426 6112
rect 6549 6103 6607 6109
rect 6549 6100 6561 6103
rect 6420 6072 6561 6100
rect 6420 6060 6426 6072
rect 6549 6069 6561 6072
rect 6595 6100 6607 6103
rect 7098 6100 7104 6112
rect 6595 6072 7104 6100
rect 6595 6069 6607 6072
rect 6549 6063 6607 6069
rect 7098 6060 7104 6072
rect 7156 6060 7162 6112
rect 8202 6100 8208 6112
rect 8163 6072 8208 6100
rect 8202 6060 8208 6072
rect 8260 6060 8266 6112
rect 10152 6100 10180 6128
rect 11425 6103 11483 6109
rect 11425 6100 11437 6103
rect 10152 6072 11437 6100
rect 11425 6069 11437 6072
rect 11471 6069 11483 6103
rect 11425 6063 11483 6069
rect 12342 6060 12348 6112
rect 12400 6100 12406 6112
rect 12728 6100 12756 6131
rect 13998 6100 14004 6112
rect 12400 6072 12756 6100
rect 13959 6072 14004 6100
rect 12400 6060 12406 6072
rect 13998 6060 14004 6072
rect 14056 6100 14062 6112
rect 14384 6100 14412 6199
rect 15838 6196 15844 6208
rect 15896 6196 15902 6248
rect 16574 6196 16580 6248
rect 16632 6236 16638 6248
rect 17012 6239 17070 6245
rect 17012 6236 17024 6239
rect 16632 6208 17024 6236
rect 16632 6196 16638 6208
rect 17012 6205 17024 6208
rect 17058 6236 17070 6239
rect 18693 6239 18751 6245
rect 17058 6208 17540 6236
rect 17058 6205 17070 6208
rect 17012 6199 17070 6205
rect 17512 6177 17540 6208
rect 18693 6205 18705 6239
rect 18739 6236 18751 6239
rect 19058 6236 19064 6248
rect 18739 6208 19064 6236
rect 18739 6205 18751 6208
rect 18693 6199 18751 6205
rect 19058 6196 19064 6208
rect 19116 6196 19122 6248
rect 17497 6171 17555 6177
rect 17497 6137 17509 6171
rect 17543 6168 17555 6171
rect 20349 6171 20407 6177
rect 17543 6140 18414 6168
rect 17543 6137 17555 6140
rect 17497 6131 17555 6137
rect 15286 6100 15292 6112
rect 14056 6072 15292 6100
rect 14056 6060 14062 6072
rect 15286 6060 15292 6072
rect 15344 6060 15350 6112
rect 17083 6103 17141 6109
rect 17083 6069 17095 6103
rect 17129 6100 17141 6103
rect 17310 6100 17316 6112
rect 17129 6072 17316 6100
rect 17129 6069 17141 6072
rect 17083 6063 17141 6069
rect 17310 6060 17316 6072
rect 17368 6060 17374 6112
rect 18386 6100 18414 6140
rect 20349 6137 20361 6171
rect 20395 6168 20407 6171
rect 20622 6168 20628 6180
rect 20395 6140 20628 6168
rect 20395 6137 20407 6140
rect 20349 6131 20407 6137
rect 20622 6128 20628 6140
rect 20680 6128 20686 6180
rect 20806 6128 20812 6180
rect 20864 6168 20870 6180
rect 21177 6171 21235 6177
rect 21177 6168 21189 6171
rect 20864 6140 21189 6168
rect 20864 6128 20870 6140
rect 21177 6137 21189 6140
rect 21223 6168 21235 6171
rect 21266 6168 21272 6180
rect 21223 6140 21272 6168
rect 21223 6137 21235 6140
rect 21177 6131 21235 6137
rect 21266 6128 21272 6140
rect 21324 6128 21330 6180
rect 23474 6100 23480 6112
rect 18386 6072 23480 6100
rect 23474 6060 23480 6072
rect 23532 6060 23538 6112
rect 1104 6010 22816 6032
rect 1104 5958 8982 6010
rect 9034 5958 9046 6010
rect 9098 5958 9110 6010
rect 9162 5958 9174 6010
rect 9226 5958 16982 6010
rect 17034 5958 17046 6010
rect 17098 5958 17110 6010
rect 17162 5958 17174 6010
rect 17226 5958 22816 6010
rect 1104 5936 22816 5958
rect 2777 5899 2835 5905
rect 2777 5896 2789 5899
rect 1504 5868 2789 5896
rect 1504 5769 1532 5868
rect 2777 5865 2789 5868
rect 2823 5896 2835 5899
rect 4157 5899 4215 5905
rect 4157 5896 4169 5899
rect 2823 5868 4169 5896
rect 2823 5865 2835 5868
rect 2777 5859 2835 5865
rect 4157 5865 4169 5868
rect 4203 5865 4215 5899
rect 4157 5859 4215 5865
rect 5350 5856 5356 5908
rect 5408 5896 5414 5908
rect 6273 5899 6331 5905
rect 6273 5896 6285 5899
rect 5408 5868 6285 5896
rect 5408 5856 5414 5868
rect 6273 5865 6285 5868
rect 6319 5865 6331 5899
rect 6273 5859 6331 5865
rect 10137 5899 10195 5905
rect 10137 5865 10149 5899
rect 10183 5896 10195 5899
rect 10226 5896 10232 5908
rect 10183 5868 10232 5896
rect 10183 5865 10195 5868
rect 10137 5859 10195 5865
rect 1854 5837 1860 5840
rect 1851 5828 1860 5837
rect 1815 5800 1860 5828
rect 1851 5791 1860 5800
rect 1854 5788 1860 5791
rect 1912 5788 1918 5840
rect 2866 5788 2872 5840
rect 2924 5828 2930 5840
rect 3421 5831 3479 5837
rect 3421 5828 3433 5831
rect 2924 5800 3433 5828
rect 2924 5788 2930 5800
rect 3421 5797 3433 5800
rect 3467 5828 3479 5831
rect 3467 5800 4752 5828
rect 3467 5797 3479 5800
rect 3421 5791 3479 5797
rect 4724 5772 4752 5800
rect 1489 5763 1547 5769
rect 1489 5729 1501 5763
rect 1535 5729 1547 5763
rect 2406 5760 2412 5772
rect 2367 5732 2412 5760
rect 1489 5723 1547 5729
rect 2406 5720 2412 5732
rect 2464 5720 2470 5772
rect 3602 5720 3608 5772
rect 3660 5760 3666 5772
rect 4065 5763 4123 5769
rect 4065 5760 4077 5763
rect 3660 5732 4077 5760
rect 3660 5720 3666 5732
rect 4065 5729 4077 5732
rect 4111 5760 4123 5763
rect 4522 5760 4528 5772
rect 4111 5732 4528 5760
rect 4111 5729 4123 5732
rect 4065 5723 4123 5729
rect 4522 5720 4528 5732
rect 4580 5720 4586 5772
rect 4706 5760 4712 5772
rect 4667 5732 4712 5760
rect 4706 5720 4712 5732
rect 4764 5720 4770 5772
rect 5077 5763 5135 5769
rect 5077 5729 5089 5763
rect 5123 5729 5135 5763
rect 5077 5723 5135 5729
rect 5445 5763 5503 5769
rect 5445 5729 5457 5763
rect 5491 5760 5503 5763
rect 5718 5760 5724 5772
rect 5491 5732 5724 5760
rect 5491 5729 5503 5732
rect 5445 5723 5503 5729
rect 3789 5695 3847 5701
rect 3789 5661 3801 5695
rect 3835 5692 3847 5695
rect 5092 5692 5120 5723
rect 5718 5720 5724 5732
rect 5776 5720 5782 5772
rect 6178 5720 6184 5772
rect 6236 5760 6242 5772
rect 6288 5760 6316 5859
rect 10226 5856 10232 5868
rect 10284 5856 10290 5908
rect 12250 5896 12256 5908
rect 12211 5868 12256 5896
rect 12250 5856 12256 5868
rect 12308 5856 12314 5908
rect 17310 5856 17316 5908
rect 17368 5896 17374 5908
rect 19061 5899 19119 5905
rect 19061 5896 19073 5899
rect 17368 5868 19073 5896
rect 17368 5856 17374 5868
rect 19061 5865 19073 5868
rect 19107 5896 19119 5899
rect 20530 5896 20536 5908
rect 19107 5868 19380 5896
rect 20491 5868 20536 5896
rect 19107 5865 19119 5868
rect 19061 5859 19119 5865
rect 10318 5788 10324 5840
rect 10376 5828 10382 5840
rect 10413 5831 10471 5837
rect 10413 5828 10425 5831
rect 10376 5800 10425 5828
rect 10376 5788 10382 5800
rect 10413 5797 10425 5800
rect 10459 5797 10471 5831
rect 10962 5828 10968 5840
rect 10923 5800 10968 5828
rect 10413 5791 10471 5797
rect 10962 5788 10968 5800
rect 11020 5788 11026 5840
rect 17678 5828 17684 5840
rect 17639 5800 17684 5828
rect 17678 5788 17684 5800
rect 17736 5788 17742 5840
rect 19352 5837 19380 5868
rect 20530 5856 20536 5868
rect 20588 5856 20594 5908
rect 21450 5896 21456 5908
rect 20640 5868 21456 5896
rect 19337 5831 19395 5837
rect 19337 5797 19349 5831
rect 19383 5797 19395 5831
rect 19337 5791 19395 5797
rect 19426 5788 19432 5840
rect 19484 5828 19490 5840
rect 20640 5828 20668 5868
rect 21450 5856 21456 5868
rect 21508 5856 21514 5908
rect 19484 5800 20668 5828
rect 19484 5788 19490 5800
rect 20806 5788 20812 5840
rect 20864 5828 20870 5840
rect 21085 5831 21143 5837
rect 21085 5828 21097 5831
rect 20864 5800 21097 5828
rect 20864 5788 20870 5800
rect 21085 5797 21097 5800
rect 21131 5797 21143 5831
rect 21085 5791 21143 5797
rect 6457 5763 6515 5769
rect 6457 5760 6469 5763
rect 6236 5732 6469 5760
rect 6236 5720 6242 5732
rect 6457 5729 6469 5732
rect 6503 5729 6515 5763
rect 6457 5723 6515 5729
rect 6733 5763 6791 5769
rect 6733 5729 6745 5763
rect 6779 5760 6791 5763
rect 6822 5760 6828 5772
rect 6779 5732 6828 5760
rect 6779 5729 6791 5732
rect 6733 5723 6791 5729
rect 6822 5720 6828 5732
rect 6880 5760 6886 5772
rect 8021 5763 8079 5769
rect 8021 5760 8033 5763
rect 6880 5732 8033 5760
rect 6880 5720 6886 5732
rect 8021 5729 8033 5732
rect 8067 5729 8079 5763
rect 8021 5723 8079 5729
rect 8110 5720 8116 5772
rect 8168 5760 8174 5772
rect 14252 5763 14310 5769
rect 8168 5732 8213 5760
rect 8168 5720 8174 5732
rect 14252 5729 14264 5763
rect 14298 5760 14310 5763
rect 15102 5760 15108 5772
rect 14298 5732 15108 5760
rect 14298 5729 14310 5732
rect 14252 5723 14310 5729
rect 15102 5720 15108 5732
rect 15160 5720 15166 5772
rect 16393 5763 16451 5769
rect 16393 5729 16405 5763
rect 16439 5760 16451 5763
rect 16482 5760 16488 5772
rect 16439 5732 16488 5760
rect 16439 5729 16451 5732
rect 16393 5723 16451 5729
rect 16482 5720 16488 5732
rect 16540 5720 16546 5772
rect 5626 5692 5632 5704
rect 3835 5664 5632 5692
rect 3835 5661 3847 5664
rect 3789 5655 3847 5661
rect 5626 5652 5632 5664
rect 5684 5652 5690 5704
rect 6914 5652 6920 5704
rect 6972 5692 6978 5704
rect 7193 5695 7251 5701
rect 7193 5692 7205 5695
rect 6972 5664 7205 5692
rect 6972 5652 6978 5664
rect 7193 5661 7205 5664
rect 7239 5692 7251 5695
rect 8754 5692 8760 5704
rect 7239 5664 8760 5692
rect 7239 5661 7251 5664
rect 7193 5655 7251 5661
rect 8754 5652 8760 5664
rect 8812 5652 8818 5704
rect 10318 5692 10324 5704
rect 10279 5664 10324 5692
rect 10318 5652 10324 5664
rect 10376 5652 10382 5704
rect 17405 5695 17463 5701
rect 17405 5661 17417 5695
rect 17451 5661 17463 5695
rect 17405 5655 17463 5661
rect 20993 5695 21051 5701
rect 20993 5661 21005 5695
rect 21039 5661 21051 5695
rect 21266 5692 21272 5704
rect 21227 5664 21272 5692
rect 20993 5655 21051 5661
rect 4522 5584 4528 5636
rect 4580 5624 4586 5636
rect 6362 5624 6368 5636
rect 4580 5596 6368 5624
rect 4580 5584 4586 5596
rect 6362 5584 6368 5596
rect 6420 5584 6426 5636
rect 6546 5624 6552 5636
rect 6507 5596 6552 5624
rect 6546 5584 6552 5596
rect 6604 5584 6610 5636
rect 14182 5584 14188 5636
rect 14240 5624 14246 5636
rect 15933 5627 15991 5633
rect 15933 5624 15945 5627
rect 14240 5596 15945 5624
rect 14240 5584 14246 5596
rect 15933 5593 15945 5596
rect 15979 5624 15991 5627
rect 16114 5624 16120 5636
rect 15979 5596 16120 5624
rect 15979 5593 15991 5596
rect 15933 5587 15991 5593
rect 16114 5584 16120 5596
rect 16172 5584 16178 5636
rect 4430 5516 4436 5568
rect 4488 5556 4494 5568
rect 7006 5556 7012 5568
rect 4488 5528 7012 5556
rect 4488 5516 4494 5528
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 7558 5556 7564 5568
rect 7519 5528 7564 5556
rect 7558 5516 7564 5528
rect 7616 5516 7622 5568
rect 12618 5556 12624 5568
rect 12579 5528 12624 5556
rect 12618 5516 12624 5528
rect 12676 5516 12682 5568
rect 14323 5559 14381 5565
rect 14323 5525 14335 5559
rect 14369 5556 14381 5559
rect 15010 5556 15016 5568
rect 14369 5528 15016 5556
rect 14369 5525 14381 5528
rect 14323 5519 14381 5525
rect 15010 5516 15016 5528
rect 15068 5516 15074 5568
rect 15654 5556 15660 5568
rect 15615 5528 15660 5556
rect 15654 5516 15660 5528
rect 15712 5516 15718 5568
rect 16531 5559 16589 5565
rect 16531 5525 16543 5559
rect 16577 5556 16589 5559
rect 16666 5556 16672 5568
rect 16577 5528 16672 5556
rect 16577 5525 16589 5528
rect 16531 5519 16589 5525
rect 16666 5516 16672 5528
rect 16724 5516 16730 5568
rect 17310 5556 17316 5568
rect 17271 5528 17316 5556
rect 17310 5516 17316 5528
rect 17368 5556 17374 5568
rect 17420 5556 17448 5655
rect 18325 5627 18383 5633
rect 18325 5593 18337 5627
rect 18371 5624 18383 5627
rect 18874 5624 18880 5636
rect 18371 5596 18880 5624
rect 18371 5593 18383 5596
rect 18325 5587 18383 5593
rect 18874 5584 18880 5596
rect 18932 5624 18938 5636
rect 19426 5624 19432 5636
rect 18932 5596 19432 5624
rect 18932 5584 18938 5596
rect 19426 5584 19432 5596
rect 19484 5584 19490 5636
rect 19886 5624 19892 5636
rect 19847 5596 19892 5624
rect 19886 5584 19892 5596
rect 19944 5624 19950 5636
rect 21008 5624 21036 5655
rect 21266 5652 21272 5664
rect 21324 5652 21330 5704
rect 21450 5624 21456 5636
rect 19944 5596 21456 5624
rect 19944 5584 19950 5596
rect 21450 5584 21456 5596
rect 21508 5584 21514 5636
rect 17368 5528 17448 5556
rect 17368 5516 17374 5528
rect 1104 5466 22816 5488
rect 1104 5414 4982 5466
rect 5034 5414 5046 5466
rect 5098 5414 5110 5466
rect 5162 5414 5174 5466
rect 5226 5414 12982 5466
rect 13034 5414 13046 5466
rect 13098 5414 13110 5466
rect 13162 5414 13174 5466
rect 13226 5414 20982 5466
rect 21034 5414 21046 5466
rect 21098 5414 21110 5466
rect 21162 5414 21174 5466
rect 21226 5414 22816 5466
rect 1104 5392 22816 5414
rect 2866 5352 2872 5364
rect 2827 5324 2872 5352
rect 2866 5312 2872 5324
rect 2924 5312 2930 5364
rect 5442 5312 5448 5364
rect 5500 5352 5506 5364
rect 6089 5355 6147 5361
rect 6089 5352 6101 5355
rect 5500 5324 6101 5352
rect 5500 5312 5506 5324
rect 6089 5321 6101 5324
rect 6135 5352 6147 5355
rect 6365 5355 6423 5361
rect 6365 5352 6377 5355
rect 6135 5324 6377 5352
rect 6135 5321 6147 5324
rect 6089 5315 6147 5321
rect 6365 5321 6377 5324
rect 6411 5321 6423 5355
rect 6546 5352 6552 5364
rect 6459 5324 6552 5352
rect 6365 5315 6423 5321
rect 6546 5312 6552 5324
rect 6604 5352 6610 5364
rect 7653 5355 7711 5361
rect 7653 5352 7665 5355
rect 6604 5324 7665 5352
rect 6604 5312 6610 5324
rect 7653 5321 7665 5324
rect 7699 5321 7711 5355
rect 7653 5315 7711 5321
rect 7742 5312 7748 5364
rect 7800 5352 7806 5364
rect 10226 5352 10232 5364
rect 7800 5324 7845 5352
rect 10187 5324 10232 5352
rect 7800 5312 7806 5324
rect 10226 5312 10232 5324
rect 10284 5312 10290 5364
rect 10594 5352 10600 5364
rect 10555 5324 10600 5352
rect 10594 5312 10600 5324
rect 10652 5312 10658 5364
rect 17678 5312 17684 5364
rect 17736 5352 17742 5364
rect 17773 5355 17831 5361
rect 17773 5352 17785 5355
rect 17736 5324 17785 5352
rect 17736 5312 17742 5324
rect 17773 5321 17785 5324
rect 17819 5321 17831 5355
rect 17773 5315 17831 5321
rect 20901 5355 20959 5361
rect 20901 5321 20913 5355
rect 20947 5352 20959 5355
rect 21358 5352 21364 5364
rect 20947 5324 21364 5352
rect 20947 5321 20959 5324
rect 20901 5315 20959 5321
rect 21358 5312 21364 5324
rect 21416 5312 21422 5364
rect 21450 5312 21456 5364
rect 21508 5352 21514 5364
rect 22189 5355 22247 5361
rect 22189 5352 22201 5355
rect 21508 5324 22201 5352
rect 21508 5312 21514 5324
rect 22189 5321 22201 5324
rect 22235 5321 22247 5355
rect 22189 5315 22247 5321
rect 1762 5244 1768 5296
rect 1820 5284 1826 5296
rect 10134 5284 10140 5296
rect 1820 5256 10140 5284
rect 1820 5244 1826 5256
rect 10134 5244 10140 5256
rect 10192 5244 10198 5296
rect 18969 5287 19027 5293
rect 18969 5253 18981 5287
rect 19015 5284 19027 5287
rect 20806 5284 20812 5296
rect 19015 5256 20812 5284
rect 19015 5253 19027 5256
rect 18969 5247 19027 5253
rect 20806 5244 20812 5256
rect 20864 5284 20870 5296
rect 20990 5284 20996 5296
rect 20864 5256 20996 5284
rect 20864 5244 20870 5256
rect 20990 5244 20996 5256
rect 21048 5284 21054 5296
rect 21177 5287 21235 5293
rect 21177 5284 21189 5287
rect 21048 5256 21189 5284
rect 21048 5244 21054 5256
rect 21177 5253 21189 5256
rect 21223 5253 21235 5287
rect 21910 5284 21916 5296
rect 21871 5256 21916 5284
rect 21177 5247 21235 5253
rect 21910 5244 21916 5256
rect 21968 5244 21974 5296
rect 2130 5216 2136 5228
rect 2091 5188 2136 5216
rect 2130 5176 2136 5188
rect 2188 5176 2194 5228
rect 5537 5219 5595 5225
rect 5537 5216 5549 5219
rect 4724 5188 5549 5216
rect 3237 5151 3295 5157
rect 3237 5117 3249 5151
rect 3283 5148 3295 5151
rect 3602 5148 3608 5160
rect 3283 5120 3608 5148
rect 3283 5117 3295 5120
rect 3237 5111 3295 5117
rect 3602 5108 3608 5120
rect 3660 5148 3666 5160
rect 3697 5151 3755 5157
rect 3697 5148 3709 5151
rect 3660 5120 3709 5148
rect 3660 5108 3666 5120
rect 3697 5117 3709 5120
rect 3743 5117 3755 5151
rect 3697 5111 3755 5117
rect 4433 5151 4491 5157
rect 4433 5117 4445 5151
rect 4479 5148 4491 5151
rect 4614 5148 4620 5160
rect 4479 5120 4620 5148
rect 4479 5117 4491 5120
rect 4433 5111 4491 5117
rect 4614 5108 4620 5120
rect 4672 5108 4678 5160
rect 4724 5157 4752 5188
rect 5537 5185 5549 5188
rect 5583 5216 5595 5219
rect 5626 5216 5632 5228
rect 5583 5188 5632 5216
rect 5583 5185 5595 5188
rect 5537 5179 5595 5185
rect 5626 5176 5632 5188
rect 5684 5176 5690 5228
rect 6730 5176 6736 5228
rect 6788 5216 6794 5228
rect 6917 5219 6975 5225
rect 6917 5216 6929 5219
rect 6788 5188 6929 5216
rect 6788 5176 6794 5188
rect 6917 5185 6929 5188
rect 6963 5216 6975 5219
rect 7558 5216 7564 5228
rect 6963 5188 7564 5216
rect 6963 5185 6975 5188
rect 6917 5179 6975 5185
rect 7558 5176 7564 5188
rect 7616 5216 7622 5228
rect 8389 5219 8447 5225
rect 8389 5216 8401 5219
rect 7616 5188 8401 5216
rect 7616 5176 7622 5188
rect 8389 5185 8401 5188
rect 8435 5185 8447 5219
rect 14734 5216 14740 5228
rect 14695 5188 14740 5216
rect 8389 5179 8447 5185
rect 14734 5176 14740 5188
rect 14792 5176 14798 5228
rect 16758 5176 16764 5228
rect 16816 5216 16822 5228
rect 20530 5216 20536 5228
rect 16816 5188 16896 5216
rect 20491 5188 20536 5216
rect 16816 5176 16822 5188
rect 4709 5151 4767 5157
rect 4709 5117 4721 5151
rect 4755 5117 4767 5151
rect 4709 5111 4767 5117
rect 5077 5151 5135 5157
rect 5077 5117 5089 5151
rect 5123 5117 5135 5151
rect 5077 5111 5135 5117
rect 1486 5080 1492 5092
rect 1447 5052 1492 5080
rect 1486 5040 1492 5052
rect 1544 5040 1550 5092
rect 1581 5083 1639 5089
rect 1581 5049 1593 5083
rect 1627 5080 1639 5083
rect 1670 5080 1676 5092
rect 1627 5052 1676 5080
rect 1627 5049 1639 5052
rect 1581 5043 1639 5049
rect 1670 5040 1676 5052
rect 1728 5040 1734 5092
rect 2682 5040 2688 5092
rect 2740 5080 2746 5092
rect 3513 5083 3571 5089
rect 3513 5080 3525 5083
rect 2740 5052 3525 5080
rect 2740 5040 2746 5052
rect 3513 5049 3525 5052
rect 3559 5080 3571 5083
rect 5092 5080 5120 5111
rect 6178 5108 6184 5160
rect 6236 5148 6242 5160
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 6236 5120 6837 5148
rect 6236 5108 6242 5120
rect 6825 5117 6837 5120
rect 6871 5117 6883 5151
rect 7098 5148 7104 5160
rect 7059 5120 7104 5148
rect 6825 5111 6883 5117
rect 7098 5108 7104 5120
rect 7156 5148 7162 5160
rect 7466 5148 7472 5160
rect 7156 5120 7472 5148
rect 7156 5108 7162 5120
rect 7466 5108 7472 5120
rect 7524 5108 7530 5160
rect 7653 5151 7711 5157
rect 7653 5117 7665 5151
rect 7699 5148 7711 5151
rect 8297 5151 8355 5157
rect 8297 5148 8309 5151
rect 7699 5120 8309 5148
rect 7699 5117 7711 5120
rect 7653 5111 7711 5117
rect 8297 5117 8309 5120
rect 8343 5148 8355 5151
rect 8481 5151 8539 5157
rect 8481 5148 8493 5151
rect 8343 5120 8493 5148
rect 8343 5117 8355 5120
rect 8297 5111 8355 5117
rect 8481 5117 8493 5120
rect 8527 5117 8539 5151
rect 8481 5111 8539 5117
rect 9490 5108 9496 5160
rect 9548 5148 9554 5160
rect 10594 5148 10600 5160
rect 9548 5120 10600 5148
rect 9548 5108 9554 5120
rect 10594 5108 10600 5120
rect 10652 5148 10658 5160
rect 10873 5151 10931 5157
rect 10873 5148 10885 5151
rect 10652 5120 10885 5148
rect 10652 5108 10658 5120
rect 10873 5117 10885 5120
rect 10919 5117 10931 5151
rect 10873 5111 10931 5117
rect 12253 5151 12311 5157
rect 12253 5117 12265 5151
rect 12299 5148 12311 5151
rect 12710 5148 12716 5160
rect 12299 5120 12716 5148
rect 12299 5117 12311 5120
rect 12253 5111 12311 5117
rect 12710 5108 12716 5120
rect 12768 5108 12774 5160
rect 13909 5151 13967 5157
rect 13909 5117 13921 5151
rect 13955 5148 13967 5151
rect 13998 5148 14004 5160
rect 13955 5120 14004 5148
rect 13955 5117 13967 5120
rect 13909 5111 13967 5117
rect 13998 5108 14004 5120
rect 14056 5148 14062 5160
rect 14645 5151 14703 5157
rect 14645 5148 14657 5151
rect 14056 5120 14657 5148
rect 14056 5108 14062 5120
rect 14645 5117 14657 5120
rect 14691 5148 14703 5151
rect 15473 5151 15531 5157
rect 15473 5148 15485 5151
rect 14691 5120 15485 5148
rect 14691 5117 14703 5120
rect 14645 5111 14703 5117
rect 15473 5117 15485 5120
rect 15519 5148 15531 5151
rect 15562 5148 15568 5160
rect 15519 5120 15568 5148
rect 15519 5117 15531 5120
rect 15473 5111 15531 5117
rect 15562 5108 15568 5120
rect 15620 5108 15626 5160
rect 15654 5108 15660 5160
rect 15712 5148 15718 5160
rect 16022 5148 16028 5160
rect 15712 5120 16028 5148
rect 15712 5108 15718 5120
rect 16022 5108 16028 5120
rect 16080 5108 16086 5160
rect 16114 5108 16120 5160
rect 16172 5148 16178 5160
rect 16390 5148 16396 5160
rect 16172 5120 16396 5148
rect 16172 5108 16178 5120
rect 16390 5108 16396 5120
rect 16448 5108 16454 5160
rect 16868 5157 16896 5188
rect 20530 5176 20536 5188
rect 20588 5176 20594 5228
rect 16853 5151 16911 5157
rect 16853 5117 16865 5151
rect 16899 5117 16911 5151
rect 16853 5111 16911 5117
rect 17037 5151 17095 5157
rect 17037 5117 17049 5151
rect 17083 5148 17095 5151
rect 18046 5148 18052 5160
rect 17083 5120 18052 5148
rect 17083 5117 17095 5120
rect 17037 5111 17095 5117
rect 18046 5108 18052 5120
rect 18104 5108 18110 5160
rect 21428 5151 21486 5157
rect 21428 5117 21440 5151
rect 21474 5148 21486 5151
rect 21928 5148 21956 5244
rect 21474 5120 21956 5148
rect 21474 5117 21486 5120
rect 21428 5111 21486 5117
rect 7742 5080 7748 5092
rect 3559 5052 7748 5080
rect 3559 5049 3571 5052
rect 3513 5043 3571 5049
rect 7742 5040 7748 5052
rect 7800 5040 7806 5092
rect 8570 5040 8576 5092
rect 8628 5080 8634 5092
rect 9861 5083 9919 5089
rect 9861 5080 9873 5083
rect 8628 5052 9873 5080
rect 8628 5040 8634 5052
rect 9861 5049 9873 5052
rect 9907 5080 9919 5083
rect 10318 5080 10324 5092
rect 9907 5052 10324 5080
rect 9907 5049 9919 5052
rect 9861 5043 9919 5049
rect 10318 5040 10324 5052
rect 10376 5040 10382 5092
rect 10778 5080 10784 5092
rect 10739 5052 10784 5080
rect 10778 5040 10784 5052
rect 10836 5040 10842 5092
rect 12434 5080 12440 5092
rect 12395 5052 12440 5080
rect 12434 5040 12440 5052
rect 12492 5040 12498 5092
rect 13262 5040 13268 5092
rect 13320 5080 13326 5092
rect 13722 5080 13728 5092
rect 13320 5052 13728 5080
rect 13320 5040 13326 5052
rect 13722 5040 13728 5052
rect 13780 5040 13786 5092
rect 16482 5040 16488 5092
rect 16540 5080 16546 5092
rect 17405 5083 17463 5089
rect 17405 5080 17417 5083
rect 16540 5052 17417 5080
rect 16540 5040 16546 5052
rect 17405 5049 17417 5052
rect 17451 5080 17463 5083
rect 18230 5080 18236 5092
rect 17451 5052 18236 5080
rect 17451 5049 17463 5052
rect 17405 5043 17463 5049
rect 18230 5040 18236 5052
rect 18288 5040 18294 5092
rect 18370 5083 18428 5089
rect 18370 5049 18382 5083
rect 18416 5049 18428 5083
rect 19889 5083 19947 5089
rect 19889 5080 19901 5083
rect 18370 5043 18428 5049
rect 19352 5052 19901 5080
rect 1688 5012 1716 5040
rect 2409 5015 2467 5021
rect 2409 5012 2421 5015
rect 1688 4984 2421 5012
rect 2409 4981 2421 4984
rect 2455 4981 2467 5015
rect 3786 5012 3792 5024
rect 3747 4984 3792 5012
rect 2409 4975 2467 4981
rect 3786 4972 3792 4984
rect 3844 4972 3850 5024
rect 6365 5015 6423 5021
rect 6365 4981 6377 5015
rect 6411 5012 6423 5015
rect 7098 5012 7104 5024
rect 6411 4984 7104 5012
rect 6411 4981 6423 4984
rect 6365 4975 6423 4981
rect 7098 4972 7104 4984
rect 7156 4972 7162 5024
rect 7466 4972 7472 5024
rect 7524 5012 7530 5024
rect 7837 5015 7895 5021
rect 7837 5012 7849 5015
rect 7524 4984 7849 5012
rect 7524 4972 7530 4984
rect 7837 4981 7849 4984
rect 7883 5012 7895 5015
rect 7926 5012 7932 5024
rect 7883 4984 7932 5012
rect 7883 4981 7895 4984
rect 7837 4975 7895 4981
rect 7926 4972 7932 4984
rect 7984 5012 7990 5024
rect 8110 5012 8116 5024
rect 7984 4984 8116 5012
rect 7984 4972 7990 4984
rect 8110 4972 8116 4984
rect 8168 4972 8174 5024
rect 15102 5012 15108 5024
rect 15063 4984 15108 5012
rect 15102 4972 15108 4984
rect 15160 4972 15166 5024
rect 16206 4972 16212 5024
rect 16264 5012 16270 5024
rect 16758 5012 16764 5024
rect 16264 4984 16764 5012
rect 16264 4972 16270 4984
rect 16758 4972 16764 4984
rect 16816 4972 16822 5024
rect 17678 4972 17684 5024
rect 17736 5012 17742 5024
rect 18385 5012 18413 5043
rect 19352 5024 19380 5052
rect 19889 5049 19901 5052
rect 19935 5049 19947 5083
rect 19889 5043 19947 5049
rect 19981 5083 20039 5089
rect 19981 5049 19993 5083
rect 20027 5049 20039 5083
rect 19981 5043 20039 5049
rect 17736 4984 18413 5012
rect 17736 4972 17742 4984
rect 19334 4972 19340 5024
rect 19392 5012 19398 5024
rect 19702 5012 19708 5024
rect 19392 4984 19437 5012
rect 19663 4984 19708 5012
rect 19392 4972 19398 4984
rect 19702 4972 19708 4984
rect 19760 5012 19766 5024
rect 19996 5012 20024 5043
rect 19760 4984 20024 5012
rect 19760 4972 19766 4984
rect 21266 4972 21272 5024
rect 21324 5012 21330 5024
rect 21499 5015 21557 5021
rect 21499 5012 21511 5015
rect 21324 4984 21511 5012
rect 21324 4972 21330 4984
rect 21499 4981 21511 4984
rect 21545 4981 21557 5015
rect 21499 4975 21557 4981
rect 1104 4922 22816 4944
rect 1104 4870 8982 4922
rect 9034 4870 9046 4922
rect 9098 4870 9110 4922
rect 9162 4870 9174 4922
rect 9226 4870 16982 4922
rect 17034 4870 17046 4922
rect 17098 4870 17110 4922
rect 17162 4870 17174 4922
rect 17226 4870 22816 4922
rect 1104 4848 22816 4870
rect 1210 4768 1216 4820
rect 1268 4808 1274 4820
rect 1673 4811 1731 4817
rect 1673 4808 1685 4811
rect 1268 4780 1685 4808
rect 1268 4768 1274 4780
rect 1673 4777 1685 4780
rect 1719 4808 1731 4811
rect 1854 4808 1860 4820
rect 1719 4780 1860 4808
rect 1719 4777 1731 4780
rect 1673 4771 1731 4777
rect 1854 4768 1860 4780
rect 1912 4768 1918 4820
rect 2406 4808 2412 4820
rect 1964 4780 2412 4808
rect 1964 4749 1992 4780
rect 2406 4768 2412 4780
rect 2464 4768 2470 4820
rect 3421 4811 3479 4817
rect 3421 4777 3433 4811
rect 3467 4808 3479 4811
rect 5718 4808 5724 4820
rect 3467 4780 5724 4808
rect 3467 4777 3479 4780
rect 3421 4771 3479 4777
rect 5718 4768 5724 4780
rect 5776 4768 5782 4820
rect 6178 4808 6184 4820
rect 6139 4780 6184 4808
rect 6178 4768 6184 4780
rect 6236 4768 6242 4820
rect 7282 4768 7288 4820
rect 7340 4808 7346 4820
rect 7558 4808 7564 4820
rect 7340 4780 7564 4808
rect 7340 4768 7346 4780
rect 7558 4768 7564 4780
rect 7616 4768 7622 4820
rect 9674 4768 9680 4820
rect 9732 4808 9738 4820
rect 9769 4811 9827 4817
rect 9769 4808 9781 4811
rect 9732 4780 9781 4808
rect 9732 4768 9738 4780
rect 9769 4777 9781 4780
rect 9815 4777 9827 4811
rect 9769 4771 9827 4777
rect 11882 4768 11888 4820
rect 11940 4808 11946 4820
rect 12069 4811 12127 4817
rect 12069 4808 12081 4811
rect 11940 4780 12081 4808
rect 11940 4768 11946 4780
rect 12069 4777 12081 4780
rect 12115 4777 12127 4811
rect 13814 4808 13820 4820
rect 12069 4771 12127 4777
rect 12360 4780 13820 4808
rect 1949 4743 2007 4749
rect 1949 4709 1961 4743
rect 1995 4709 2007 4743
rect 1949 4703 2007 4709
rect 4338 4700 4344 4752
rect 4396 4740 4402 4752
rect 4433 4743 4491 4749
rect 4433 4740 4445 4743
rect 4396 4712 4445 4740
rect 4396 4700 4402 4712
rect 4433 4709 4445 4712
rect 4479 4709 4491 4743
rect 4433 4703 4491 4709
rect 6196 4672 6224 4768
rect 6549 4743 6607 4749
rect 6549 4709 6561 4743
rect 6595 4740 6607 4743
rect 6822 4740 6828 4752
rect 6595 4712 6828 4740
rect 6595 4709 6607 4712
rect 6549 4703 6607 4709
rect 6822 4700 6828 4712
rect 6880 4740 6886 4752
rect 12360 4740 12388 4780
rect 13814 4768 13820 4780
rect 13872 4808 13878 4820
rect 14185 4811 14243 4817
rect 14185 4808 14197 4811
rect 13872 4780 14197 4808
rect 13872 4768 13878 4780
rect 14185 4777 14197 4780
rect 14231 4808 14243 4811
rect 14734 4808 14740 4820
rect 14231 4780 14740 4808
rect 14231 4777 14243 4780
rect 14185 4771 14243 4777
rect 14734 4768 14740 4780
rect 14792 4768 14798 4820
rect 17497 4811 17555 4817
rect 17497 4777 17509 4811
rect 17543 4808 17555 4811
rect 17678 4808 17684 4820
rect 17543 4780 17684 4808
rect 17543 4777 17555 4780
rect 17497 4771 17555 4777
rect 17678 4768 17684 4780
rect 17736 4768 17742 4820
rect 18046 4768 18052 4820
rect 18104 4808 18110 4820
rect 18325 4811 18383 4817
rect 18325 4808 18337 4811
rect 18104 4780 18337 4808
rect 18104 4768 18110 4780
rect 18325 4777 18337 4780
rect 18371 4777 18383 4811
rect 18325 4771 18383 4777
rect 13262 4740 13268 4752
rect 6880 4712 6960 4740
rect 6880 4700 6886 4712
rect 6454 4672 6460 4684
rect 6196 4644 6460 4672
rect 6454 4632 6460 4644
rect 6512 4672 6518 4684
rect 6932 4681 6960 4712
rect 9968 4712 12388 4740
rect 6641 4675 6699 4681
rect 6641 4672 6653 4675
rect 6512 4644 6653 4672
rect 6512 4632 6518 4644
rect 6641 4641 6653 4644
rect 6687 4641 6699 4675
rect 6641 4635 6699 4641
rect 6917 4675 6975 4681
rect 6917 4641 6929 4675
rect 6963 4641 6975 4675
rect 6917 4635 6975 4641
rect 8113 4675 8171 4681
rect 8113 4641 8125 4675
rect 8159 4672 8171 4675
rect 8294 4672 8300 4684
rect 8159 4644 8300 4672
rect 8159 4641 8171 4644
rect 8113 4635 8171 4641
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 8757 4675 8815 4681
rect 8757 4641 8769 4675
rect 8803 4672 8815 4675
rect 9398 4672 9404 4684
rect 8803 4644 9404 4672
rect 8803 4641 8815 4644
rect 8757 4635 8815 4641
rect 9398 4632 9404 4644
rect 9456 4672 9462 4684
rect 9968 4681 9996 4712
rect 9953 4675 10011 4681
rect 9953 4672 9965 4675
rect 9456 4644 9965 4672
rect 9456 4632 9462 4644
rect 9953 4641 9965 4644
rect 9999 4641 10011 4675
rect 10410 4672 10416 4684
rect 10371 4644 10416 4672
rect 9953 4635 10011 4641
rect 10410 4632 10416 4644
rect 10468 4632 10474 4684
rect 10686 4672 10692 4684
rect 10647 4644 10692 4672
rect 10686 4632 10692 4644
rect 10744 4632 10750 4684
rect 10873 4675 10931 4681
rect 10873 4641 10885 4675
rect 10919 4672 10931 4675
rect 11793 4675 11851 4681
rect 11793 4672 11805 4675
rect 10919 4644 11805 4672
rect 10919 4641 10931 4644
rect 10873 4635 10931 4641
rect 1857 4607 1915 4613
rect 1857 4573 1869 4607
rect 1903 4604 1915 4607
rect 1946 4604 1952 4616
rect 1903 4576 1952 4604
rect 1903 4573 1915 4576
rect 1857 4567 1915 4573
rect 1946 4564 1952 4576
rect 2004 4564 2010 4616
rect 2130 4604 2136 4616
rect 2091 4576 2136 4604
rect 2130 4564 2136 4576
rect 2188 4564 2194 4616
rect 4341 4607 4399 4613
rect 4341 4573 4353 4607
rect 4387 4604 4399 4607
rect 4522 4604 4528 4616
rect 4387 4576 4528 4604
rect 4387 4573 4399 4576
rect 4341 4567 4399 4573
rect 4522 4564 4528 4576
rect 4580 4564 4586 4616
rect 4706 4604 4712 4616
rect 4667 4576 4712 4604
rect 4706 4564 4712 4576
rect 4764 4564 4770 4616
rect 6730 4604 6736 4616
rect 6691 4576 6736 4604
rect 6730 4564 6736 4576
rect 6788 4564 6794 4616
rect 7374 4604 7380 4616
rect 7335 4576 7380 4604
rect 7374 4564 7380 4576
rect 7432 4564 7438 4616
rect 10778 4604 10784 4616
rect 7668 4576 10784 4604
rect 5718 4496 5724 4548
rect 5776 4536 5782 4548
rect 7668 4536 7696 4576
rect 10778 4564 10784 4576
rect 10836 4604 10842 4616
rect 10888 4604 10916 4635
rect 10836 4576 10916 4604
rect 10836 4564 10842 4576
rect 5776 4508 7696 4536
rect 8021 4539 8079 4545
rect 5776 4496 5782 4508
rect 8021 4505 8033 4539
rect 8067 4536 8079 4539
rect 8202 4536 8208 4548
rect 8067 4508 8208 4536
rect 8067 4505 8079 4508
rect 8021 4499 8079 4505
rect 8202 4496 8208 4508
rect 8260 4496 8266 4548
rect 11532 4536 11560 4644
rect 11793 4641 11805 4644
rect 11839 4641 11851 4675
rect 12250 4672 12256 4684
rect 12163 4644 12256 4672
rect 11793 4635 11851 4641
rect 12250 4632 12256 4644
rect 12308 4672 12314 4684
rect 12360 4672 12388 4712
rect 12728 4712 13268 4740
rect 12728 4681 12756 4712
rect 13262 4700 13268 4712
rect 13320 4700 13326 4752
rect 16298 4700 16304 4752
rect 16356 4740 16362 4752
rect 17037 4743 17095 4749
rect 16356 4712 16804 4740
rect 16356 4700 16362 4712
rect 12308 4644 12388 4672
rect 12713 4675 12771 4681
rect 12308 4632 12314 4644
rect 12713 4641 12725 4675
rect 12759 4641 12771 4675
rect 12713 4635 12771 4641
rect 12805 4675 12863 4681
rect 12805 4641 12817 4675
rect 12851 4641 12863 4675
rect 13170 4672 13176 4684
rect 13131 4644 13176 4672
rect 12805 4635 12863 4641
rect 11606 4564 11612 4616
rect 11664 4604 11670 4616
rect 12820 4604 12848 4635
rect 13170 4632 13176 4644
rect 13228 4672 13234 4684
rect 15013 4675 15071 4681
rect 15013 4672 15025 4675
rect 13228 4644 15025 4672
rect 13228 4632 13234 4644
rect 15013 4641 15025 4644
rect 15059 4641 15071 4675
rect 15013 4635 15071 4641
rect 15562 4632 15568 4684
rect 15620 4672 15626 4684
rect 15841 4675 15899 4681
rect 15841 4672 15853 4675
rect 15620 4644 15853 4672
rect 15620 4632 15626 4644
rect 15841 4641 15853 4644
rect 15887 4641 15899 4675
rect 16022 4672 16028 4684
rect 15983 4644 16028 4672
rect 15841 4635 15899 4641
rect 13725 4607 13783 4613
rect 13725 4604 13737 4607
rect 11664 4576 13737 4604
rect 11664 4564 11670 4576
rect 13725 4573 13737 4576
rect 13771 4604 13783 4607
rect 14182 4604 14188 4616
rect 13771 4576 14188 4604
rect 13771 4573 13783 4576
rect 13725 4567 13783 4573
rect 14182 4564 14188 4576
rect 14240 4604 14246 4616
rect 14366 4604 14372 4616
rect 14240 4576 14372 4604
rect 14240 4564 14246 4576
rect 14366 4564 14372 4576
rect 14424 4564 14430 4616
rect 15856 4604 15884 4635
rect 16022 4632 16028 4644
rect 16080 4632 16086 4684
rect 16390 4672 16396 4684
rect 16351 4644 16396 4672
rect 16390 4632 16396 4644
rect 16448 4632 16454 4684
rect 16776 4681 16804 4712
rect 17037 4709 17049 4743
rect 17083 4740 17095 4743
rect 17310 4740 17316 4752
rect 17083 4712 17316 4740
rect 17083 4709 17095 4712
rect 17037 4703 17095 4709
rect 17310 4700 17316 4712
rect 17368 4700 17374 4752
rect 19337 4743 19395 4749
rect 19337 4709 19349 4743
rect 19383 4740 19395 4743
rect 19702 4740 19708 4752
rect 19383 4712 19708 4740
rect 19383 4709 19395 4712
rect 19337 4703 19395 4709
rect 19702 4700 19708 4712
rect 19760 4700 19766 4752
rect 19886 4740 19892 4752
rect 19847 4712 19892 4740
rect 19886 4700 19892 4712
rect 19944 4700 19950 4752
rect 20622 4700 20628 4752
rect 20680 4740 20686 4752
rect 20901 4743 20959 4749
rect 20901 4740 20913 4743
rect 20680 4712 20913 4740
rect 20680 4700 20686 4712
rect 20901 4709 20913 4712
rect 20947 4709 20959 4743
rect 20901 4703 20959 4709
rect 16761 4675 16819 4681
rect 16761 4641 16773 4675
rect 16807 4641 16819 4675
rect 16761 4635 16819 4641
rect 17932 4675 17990 4681
rect 17932 4641 17944 4675
rect 17978 4672 17990 4675
rect 18322 4672 18328 4684
rect 17978 4644 18328 4672
rect 17978 4641 17990 4644
rect 17932 4635 17990 4641
rect 18322 4632 18328 4644
rect 18380 4672 18386 4684
rect 18690 4672 18696 4684
rect 18380 4644 18696 4672
rect 18380 4632 18386 4644
rect 18690 4632 18696 4644
rect 18748 4632 18754 4684
rect 20990 4672 20996 4684
rect 20951 4644 20996 4672
rect 20990 4632 20996 4644
rect 21048 4632 21054 4684
rect 16206 4604 16212 4616
rect 15856 4576 16212 4604
rect 16206 4564 16212 4576
rect 16264 4564 16270 4616
rect 19242 4604 19248 4616
rect 19203 4576 19248 4604
rect 19242 4564 19248 4576
rect 19300 4564 19306 4616
rect 13170 4536 13176 4548
rect 11532 4508 13176 4536
rect 13170 4496 13176 4508
rect 13228 4496 13234 4548
rect 3602 4428 3608 4480
rect 3660 4468 3666 4480
rect 3697 4471 3755 4477
rect 3697 4468 3709 4471
rect 3660 4440 3709 4468
rect 3660 4428 3666 4440
rect 3697 4437 3709 4440
rect 3743 4437 3755 4471
rect 3697 4431 3755 4437
rect 8110 4428 8116 4480
rect 8168 4468 8174 4480
rect 8343 4471 8401 4477
rect 8343 4468 8355 4471
rect 8168 4440 8355 4468
rect 8168 4428 8174 4440
rect 8343 4437 8355 4440
rect 8389 4437 8401 4471
rect 8343 4431 8401 4437
rect 14090 4428 14096 4480
rect 14148 4468 14154 4480
rect 18003 4471 18061 4477
rect 18003 4468 18015 4471
rect 14148 4440 18015 4468
rect 14148 4428 14154 4440
rect 18003 4437 18015 4440
rect 18049 4437 18061 4471
rect 18003 4431 18061 4437
rect 1104 4378 22816 4400
rect 1104 4326 4982 4378
rect 5034 4326 5046 4378
rect 5098 4326 5110 4378
rect 5162 4326 5174 4378
rect 5226 4326 12982 4378
rect 13034 4326 13046 4378
rect 13098 4326 13110 4378
rect 13162 4326 13174 4378
rect 13226 4326 20982 4378
rect 21034 4326 21046 4378
rect 21098 4326 21110 4378
rect 21162 4326 21174 4378
rect 21226 4326 22816 4378
rect 1104 4304 22816 4326
rect 2317 4267 2375 4273
rect 2317 4233 2329 4267
rect 2363 4264 2375 4267
rect 2406 4264 2412 4276
rect 2363 4236 2412 4264
rect 2363 4233 2375 4236
rect 2317 4227 2375 4233
rect 2406 4224 2412 4236
rect 2464 4224 2470 4276
rect 4522 4224 4528 4276
rect 4580 4264 4586 4276
rect 5445 4267 5503 4273
rect 5445 4264 5457 4267
rect 4580 4236 5457 4264
rect 4580 4224 4586 4236
rect 5445 4233 5457 4236
rect 5491 4264 5503 4267
rect 5767 4267 5825 4273
rect 5767 4264 5779 4267
rect 5491 4236 5779 4264
rect 5491 4233 5503 4236
rect 5445 4227 5503 4233
rect 5767 4233 5779 4236
rect 5813 4233 5825 4267
rect 5767 4227 5825 4233
rect 6641 4267 6699 4273
rect 6641 4233 6653 4267
rect 6687 4264 6699 4267
rect 6822 4264 6828 4276
rect 6687 4236 6828 4264
rect 6687 4233 6699 4236
rect 6641 4227 6699 4233
rect 6822 4224 6828 4236
rect 6880 4224 6886 4276
rect 7282 4224 7288 4276
rect 7340 4264 7346 4276
rect 7466 4264 7472 4276
rect 7340 4236 7472 4264
rect 7340 4224 7346 4236
rect 7466 4224 7472 4236
rect 7524 4224 7530 4276
rect 8754 4224 8760 4276
rect 8812 4264 8818 4276
rect 8812 4236 9536 4264
rect 8812 4224 8818 4236
rect 1854 4156 1860 4208
rect 1912 4196 1918 4208
rect 3605 4199 3663 4205
rect 3605 4196 3617 4199
rect 1912 4168 3617 4196
rect 1912 4156 1918 4168
rect 3605 4165 3617 4168
rect 3651 4196 3663 4199
rect 3697 4199 3755 4205
rect 3697 4196 3709 4199
rect 3651 4168 3709 4196
rect 3651 4165 3663 4168
rect 3605 4159 3663 4165
rect 3697 4165 3709 4168
rect 3743 4165 3755 4199
rect 7742 4196 7748 4208
rect 7703 4168 7748 4196
rect 3697 4159 3755 4165
rect 7742 4156 7748 4168
rect 7800 4156 7806 4208
rect 9398 4196 9404 4208
rect 8128 4168 9404 4196
rect 1946 4088 1952 4140
rect 2004 4128 2010 4140
rect 2593 4131 2651 4137
rect 2593 4128 2605 4131
rect 2004 4100 2605 4128
rect 2004 4088 2010 4100
rect 2593 4097 2605 4100
rect 2639 4128 2651 4131
rect 4706 4128 4712 4140
rect 2639 4100 4712 4128
rect 2639 4097 2651 4100
rect 2593 4091 2651 4097
rect 4706 4088 4712 4100
rect 4764 4088 4770 4140
rect 3421 4063 3479 4069
rect 3421 4029 3433 4063
rect 3467 4060 3479 4063
rect 3786 4060 3792 4072
rect 3467 4032 3792 4060
rect 3467 4029 3479 4032
rect 3421 4023 3479 4029
rect 3786 4020 3792 4032
rect 3844 4060 3850 4072
rect 3881 4063 3939 4069
rect 3881 4060 3893 4063
rect 3844 4032 3893 4060
rect 3844 4020 3850 4032
rect 3881 4029 3893 4032
rect 3927 4029 3939 4063
rect 3881 4023 3939 4029
rect 5534 4020 5540 4072
rect 5592 4060 5598 4072
rect 5664 4063 5722 4069
rect 5664 4060 5676 4063
rect 5592 4032 5676 4060
rect 5592 4020 5598 4032
rect 5664 4029 5676 4032
rect 5710 4060 5722 4063
rect 6089 4063 6147 4069
rect 6089 4060 6101 4063
rect 5710 4032 6101 4060
rect 5710 4029 5722 4032
rect 5664 4023 5722 4029
rect 6089 4029 6101 4032
rect 6135 4029 6147 4063
rect 6089 4023 6147 4029
rect 6984 4063 7042 4069
rect 6984 4029 6996 4063
rect 7030 4060 7042 4063
rect 7282 4060 7288 4072
rect 7030 4032 7288 4060
rect 7030 4029 7042 4032
rect 6984 4023 7042 4029
rect 7282 4020 7288 4032
rect 7340 4020 7346 4072
rect 8128 4069 8156 4168
rect 9398 4156 9404 4168
rect 9456 4156 9462 4208
rect 9508 4196 9536 4236
rect 10778 4224 10784 4276
rect 10836 4264 10842 4276
rect 11241 4267 11299 4273
rect 11241 4264 11253 4267
rect 10836 4236 11253 4264
rect 10836 4224 10842 4236
rect 11241 4233 11253 4236
rect 11287 4233 11299 4267
rect 11241 4227 11299 4233
rect 16390 4224 16396 4276
rect 16448 4264 16454 4276
rect 17221 4267 17279 4273
rect 17221 4264 17233 4267
rect 16448 4236 17233 4264
rect 16448 4224 16454 4236
rect 17221 4233 17233 4236
rect 17267 4233 17279 4267
rect 18322 4264 18328 4276
rect 18283 4236 18328 4264
rect 17221 4227 17279 4233
rect 18322 4224 18328 4236
rect 18380 4224 18386 4276
rect 18874 4264 18880 4276
rect 18835 4236 18880 4264
rect 18874 4224 18880 4236
rect 18932 4224 18938 4276
rect 20806 4224 20812 4276
rect 20864 4264 20870 4276
rect 20901 4267 20959 4273
rect 20901 4264 20913 4267
rect 20864 4236 20913 4264
rect 20864 4224 20870 4236
rect 20901 4233 20913 4236
rect 20947 4233 20959 4267
rect 20901 4227 20959 4233
rect 10137 4199 10195 4205
rect 10137 4196 10149 4199
rect 9508 4168 10149 4196
rect 10137 4165 10149 4168
rect 10183 4196 10195 4199
rect 10686 4196 10692 4208
rect 10183 4168 10692 4196
rect 10183 4165 10195 4168
rect 10137 4159 10195 4165
rect 10686 4156 10692 4168
rect 10744 4156 10750 4208
rect 15657 4199 15715 4205
rect 15657 4165 15669 4199
rect 15703 4196 15715 4199
rect 16298 4196 16304 4208
rect 15703 4168 16304 4196
rect 15703 4165 15715 4168
rect 15657 4159 15715 4165
rect 9582 4128 9588 4140
rect 8404 4100 9588 4128
rect 8113 4063 8171 4069
rect 8113 4029 8125 4063
rect 8159 4029 8171 4063
rect 8113 4023 8171 4029
rect 8202 4020 8208 4072
rect 8260 4060 8266 4072
rect 8404 4069 8432 4100
rect 9582 4088 9588 4100
rect 9640 4088 9646 4140
rect 11606 4128 11612 4140
rect 10428 4100 11612 4128
rect 8389 4063 8447 4069
rect 8389 4060 8401 4063
rect 8260 4032 8401 4060
rect 8260 4020 8266 4032
rect 8389 4029 8401 4032
rect 8435 4029 8447 4063
rect 8754 4060 8760 4072
rect 8715 4032 8760 4060
rect 8389 4023 8447 4029
rect 8754 4020 8760 4032
rect 8812 4020 8818 4072
rect 9309 4063 9367 4069
rect 9309 4029 9321 4063
rect 9355 4060 9367 4063
rect 9490 4060 9496 4072
rect 9355 4032 9496 4060
rect 9355 4029 9367 4032
rect 9309 4023 9367 4029
rect 9490 4020 9496 4032
rect 9548 4020 9554 4072
rect 10428 4060 10456 4100
rect 11606 4088 11612 4100
rect 11664 4088 11670 4140
rect 13449 4131 13507 4137
rect 13449 4097 13461 4131
rect 13495 4128 13507 4131
rect 13495 4100 14964 4128
rect 13495 4097 13507 4100
rect 13449 4091 13507 4097
rect 10594 4060 10600 4072
rect 9646 4032 10456 4060
rect 10555 4032 10600 4060
rect 1397 3995 1455 4001
rect 1397 3961 1409 3995
rect 1443 3992 1455 3995
rect 1486 3992 1492 4004
rect 1443 3964 1492 3992
rect 1443 3961 1455 3964
rect 1397 3955 1455 3961
rect 1486 3952 1492 3964
rect 1544 3992 1550 4004
rect 1857 3995 1915 4001
rect 1857 3992 1869 3995
rect 1544 3964 1869 3992
rect 1544 3952 1550 3964
rect 1857 3961 1869 3964
rect 1903 3961 1915 3995
rect 1857 3955 1915 3961
rect 3605 3995 3663 4001
rect 3605 3961 3617 3995
rect 3651 3992 3663 3995
rect 4202 3995 4260 4001
rect 4202 3992 4214 3995
rect 3651 3964 4214 3992
rect 3651 3961 3663 3964
rect 3605 3955 3663 3961
rect 4202 3961 4214 3964
rect 4248 3992 4260 3995
rect 6546 3992 6552 4004
rect 4248 3964 6552 3992
rect 4248 3961 4260 3964
rect 4202 3955 4260 3961
rect 6546 3952 6552 3964
rect 6604 3952 6610 4004
rect 7374 3952 7380 4004
rect 7432 3992 7438 4004
rect 9646 3992 9674 4032
rect 10594 4020 10600 4032
rect 10652 4020 10658 4072
rect 12504 4063 12562 4069
rect 12504 4029 12516 4063
rect 12550 4060 12562 4063
rect 13354 4060 13360 4072
rect 12550 4032 13360 4060
rect 12550 4029 12562 4032
rect 12504 4023 12562 4029
rect 13354 4020 13360 4032
rect 13412 4020 13418 4072
rect 13814 4020 13820 4072
rect 13872 4060 13878 4072
rect 14185 4063 14243 4069
rect 13872 4032 13917 4060
rect 13872 4020 13878 4032
rect 14185 4029 14197 4063
rect 14231 4029 14243 4063
rect 14366 4060 14372 4072
rect 14327 4032 14372 4060
rect 14185 4023 14243 4029
rect 7432 3964 9674 3992
rect 7432 3952 7438 3964
rect 9766 3952 9772 4004
rect 9824 3992 9830 4004
rect 10229 3995 10287 4001
rect 10229 3992 10241 3995
rect 9824 3964 10241 3992
rect 9824 3952 9830 3964
rect 10229 3961 10241 3964
rect 10275 3961 10287 3995
rect 12989 3995 13047 4001
rect 12989 3992 13001 3995
rect 10229 3955 10287 3961
rect 11992 3964 13001 3992
rect 4338 3884 4344 3936
rect 4396 3924 4402 3936
rect 4798 3924 4804 3936
rect 4396 3896 4804 3924
rect 4396 3884 4402 3896
rect 4798 3884 4804 3896
rect 4856 3924 4862 3936
rect 5077 3927 5135 3933
rect 5077 3924 5089 3927
rect 4856 3896 5089 3924
rect 4856 3884 4862 3896
rect 5077 3893 5089 3896
rect 5123 3893 5135 3927
rect 5077 3887 5135 3893
rect 7055 3927 7113 3933
rect 7055 3893 7067 3927
rect 7101 3924 7113 3927
rect 7282 3924 7288 3936
rect 7101 3896 7288 3924
rect 7101 3893 7113 3896
rect 7055 3887 7113 3893
rect 7282 3884 7288 3896
rect 7340 3884 7346 3936
rect 8018 3924 8024 3936
rect 7979 3896 8024 3924
rect 8018 3884 8024 3896
rect 8076 3884 8082 3936
rect 9582 3884 9588 3936
rect 9640 3924 9646 3936
rect 9677 3927 9735 3933
rect 9677 3924 9689 3927
rect 9640 3896 9689 3924
rect 9640 3884 9646 3896
rect 9677 3893 9689 3896
rect 9723 3924 9735 3927
rect 10410 3924 10416 3936
rect 9723 3896 10416 3924
rect 9723 3893 9735 3896
rect 9677 3887 9735 3893
rect 10410 3884 10416 3896
rect 10468 3924 10474 3936
rect 11992 3933 12020 3964
rect 12989 3961 13001 3964
rect 13035 3992 13047 3995
rect 13262 3992 13268 4004
rect 13035 3964 13268 3992
rect 13035 3961 13047 3964
rect 12989 3955 13047 3961
rect 13262 3952 13268 3964
rect 13320 3992 13326 4004
rect 14200 3992 14228 4023
rect 14366 4020 14372 4032
rect 14424 4020 14430 4072
rect 14936 4069 14964 4100
rect 14921 4063 14979 4069
rect 14921 4029 14933 4063
rect 14967 4060 14979 4063
rect 15672 4060 15700 4159
rect 16298 4156 16304 4168
rect 16356 4156 16362 4208
rect 15933 4131 15991 4137
rect 15933 4097 15945 4131
rect 15979 4128 15991 4131
rect 16574 4128 16580 4140
rect 15979 4100 16580 4128
rect 15979 4097 15991 4100
rect 15933 4091 15991 4097
rect 16574 4088 16580 4100
rect 16632 4128 16638 4140
rect 17589 4131 17647 4137
rect 17589 4128 17601 4131
rect 16632 4100 17601 4128
rect 16632 4088 16638 4100
rect 17589 4097 17601 4100
rect 17635 4097 17647 4131
rect 17589 4091 17647 4097
rect 14967 4032 15700 4060
rect 14967 4029 14979 4032
rect 14921 4023 14979 4029
rect 18874 4020 18880 4072
rect 18932 4060 18938 4072
rect 19061 4063 19119 4069
rect 19061 4060 19073 4063
rect 18932 4032 19073 4060
rect 18932 4020 18938 4032
rect 19061 4029 19073 4032
rect 19107 4029 19119 4063
rect 19061 4023 19119 4029
rect 16025 3995 16083 4001
rect 13320 3964 14964 3992
rect 13320 3952 13326 3964
rect 11977 3927 12035 3933
rect 11977 3924 11989 3927
rect 10468 3896 11989 3924
rect 10468 3884 10474 3896
rect 11977 3893 11989 3896
rect 12023 3893 12035 3927
rect 11977 3887 12035 3893
rect 12066 3884 12072 3936
rect 12124 3924 12130 3936
rect 12575 3927 12633 3933
rect 12575 3924 12587 3927
rect 12124 3896 12587 3924
rect 12124 3884 12130 3896
rect 12575 3893 12587 3896
rect 12621 3893 12633 3927
rect 14734 3924 14740 3936
rect 14695 3896 14740 3924
rect 12575 3887 12633 3893
rect 14734 3884 14740 3896
rect 14792 3884 14798 3936
rect 14936 3924 14964 3964
rect 16025 3961 16037 3995
rect 16071 3992 16083 3995
rect 16390 3992 16396 4004
rect 16071 3964 16396 3992
rect 16071 3961 16083 3964
rect 16025 3955 16083 3961
rect 16390 3952 16396 3964
rect 16448 3952 16454 4004
rect 16574 3992 16580 4004
rect 16535 3964 16580 3992
rect 16574 3952 16580 3964
rect 16632 3952 16638 4004
rect 19702 3992 19708 4004
rect 19615 3964 19708 3992
rect 19702 3952 19708 3964
rect 19760 3992 19766 4004
rect 19981 3995 20039 4001
rect 19981 3992 19993 3995
rect 19760 3964 19993 3992
rect 19760 3952 19766 3964
rect 19981 3961 19993 3964
rect 20027 3961 20039 3995
rect 19981 3955 20039 3961
rect 16114 3924 16120 3936
rect 14936 3896 16120 3924
rect 16114 3884 16120 3896
rect 16172 3924 16178 3936
rect 16945 3927 17003 3933
rect 16945 3924 16957 3927
rect 16172 3896 16957 3924
rect 16172 3884 16178 3896
rect 16945 3893 16957 3896
rect 16991 3924 17003 3927
rect 17310 3924 17316 3936
rect 16991 3896 17316 3924
rect 16991 3893 17003 3896
rect 16945 3887 17003 3893
rect 17310 3884 17316 3896
rect 17368 3884 17374 3936
rect 1104 3834 22816 3856
rect 1104 3782 8982 3834
rect 9034 3782 9046 3834
rect 9098 3782 9110 3834
rect 9162 3782 9174 3834
rect 9226 3782 16982 3834
rect 17034 3782 17046 3834
rect 17098 3782 17110 3834
rect 17162 3782 17174 3834
rect 17226 3782 22816 3834
rect 1104 3760 22816 3782
rect 6730 3720 6736 3732
rect 6691 3692 6736 3720
rect 6730 3680 6736 3692
rect 6788 3680 6794 3732
rect 8665 3723 8723 3729
rect 8665 3689 8677 3723
rect 8711 3720 8723 3723
rect 8754 3720 8760 3732
rect 8711 3692 8760 3720
rect 8711 3689 8723 3692
rect 8665 3683 8723 3689
rect 8754 3680 8760 3692
rect 8812 3680 8818 3732
rect 9398 3720 9404 3732
rect 9359 3692 9404 3720
rect 9398 3680 9404 3692
rect 9456 3680 9462 3732
rect 11701 3723 11759 3729
rect 11701 3689 11713 3723
rect 11747 3720 11759 3723
rect 12250 3720 12256 3732
rect 11747 3692 12256 3720
rect 11747 3689 11759 3692
rect 11701 3683 11759 3689
rect 12250 3680 12256 3692
rect 12308 3680 12314 3732
rect 12710 3720 12716 3732
rect 12671 3692 12716 3720
rect 12710 3680 12716 3692
rect 12768 3680 12774 3732
rect 13354 3720 13360 3732
rect 13315 3692 13360 3720
rect 13354 3680 13360 3692
rect 13412 3680 13418 3732
rect 14734 3720 14740 3732
rect 14695 3692 14740 3720
rect 14734 3680 14740 3692
rect 14792 3680 14798 3732
rect 15010 3720 15016 3732
rect 14971 3692 15016 3720
rect 15010 3680 15016 3692
rect 15068 3680 15074 3732
rect 16206 3680 16212 3732
rect 16264 3720 16270 3732
rect 16301 3723 16359 3729
rect 16301 3720 16313 3723
rect 16264 3692 16313 3720
rect 16264 3680 16270 3692
rect 16301 3689 16313 3692
rect 16347 3689 16359 3723
rect 16301 3683 16359 3689
rect 16390 3680 16396 3732
rect 16448 3720 16454 3732
rect 16669 3723 16727 3729
rect 16669 3720 16681 3723
rect 16448 3692 16681 3720
rect 16448 3680 16454 3692
rect 16669 3689 16681 3692
rect 16715 3689 16727 3723
rect 16669 3683 16727 3689
rect 17494 3680 17500 3732
rect 17552 3720 17558 3732
rect 18095 3723 18153 3729
rect 18095 3720 18107 3723
rect 17552 3692 18107 3720
rect 17552 3680 17558 3692
rect 18095 3689 18107 3692
rect 18141 3689 18153 3723
rect 19242 3720 19248 3732
rect 19203 3692 19248 3720
rect 18095 3683 18153 3689
rect 19242 3680 19248 3692
rect 19300 3680 19306 3732
rect 19334 3680 19340 3732
rect 19392 3720 19398 3732
rect 19429 3723 19487 3729
rect 19429 3720 19441 3723
rect 19392 3692 19441 3720
rect 19392 3680 19398 3692
rect 19429 3689 19441 3692
rect 19475 3689 19487 3723
rect 19429 3683 19487 3689
rect 20254 3680 20260 3732
rect 20312 3720 20318 3732
rect 21039 3723 21097 3729
rect 21039 3720 21051 3723
rect 20312 3692 21051 3720
rect 20312 3680 20318 3692
rect 21039 3689 21051 3692
rect 21085 3689 21097 3723
rect 21039 3683 21097 3689
rect 7374 3652 7380 3664
rect 7335 3624 7380 3652
rect 7374 3612 7380 3624
rect 7432 3612 7438 3664
rect 7742 3612 7748 3664
rect 7800 3652 7806 3664
rect 9490 3652 9496 3664
rect 7800 3624 9496 3652
rect 7800 3612 7806 3624
rect 9490 3612 9496 3624
rect 9548 3612 9554 3664
rect 9950 3652 9956 3664
rect 9911 3624 9956 3652
rect 9950 3612 9956 3624
rect 10008 3612 10014 3664
rect 11790 3612 11796 3664
rect 11848 3652 11854 3664
rect 12114 3655 12172 3661
rect 12114 3652 12126 3655
rect 11848 3624 12126 3652
rect 11848 3612 11854 3624
rect 12114 3621 12126 3624
rect 12160 3621 12172 3655
rect 15028 3652 15056 3680
rect 15381 3655 15439 3661
rect 15381 3652 15393 3655
rect 15028 3624 15393 3652
rect 12114 3615 12172 3621
rect 15381 3621 15393 3624
rect 15427 3621 15439 3655
rect 15381 3615 15439 3621
rect 15470 3612 15476 3664
rect 15528 3652 15534 3664
rect 16408 3652 16436 3680
rect 15528 3624 16436 3652
rect 15528 3612 15534 3624
rect 4798 3584 4804 3596
rect 4759 3556 4804 3584
rect 4798 3544 4804 3556
rect 4856 3544 4862 3596
rect 5721 3587 5779 3593
rect 5721 3553 5733 3587
rect 5767 3584 5779 3587
rect 5810 3584 5816 3596
rect 5767 3556 5816 3584
rect 5767 3553 5779 3556
rect 5721 3547 5779 3553
rect 5810 3544 5816 3556
rect 5868 3544 5874 3596
rect 8294 3584 8300 3596
rect 8207 3556 8300 3584
rect 8294 3544 8300 3556
rect 8352 3584 8358 3596
rect 13446 3584 13452 3596
rect 8352 3556 13452 3584
rect 8352 3544 8358 3556
rect 13446 3544 13452 3556
rect 13504 3544 13510 3596
rect 14274 3584 14280 3596
rect 14235 3556 14280 3584
rect 14274 3544 14280 3556
rect 14332 3544 14338 3596
rect 16850 3584 16856 3596
rect 16811 3556 16856 3584
rect 16850 3544 16856 3556
rect 16908 3544 16914 3596
rect 18024 3587 18082 3593
rect 18024 3553 18036 3587
rect 18070 3584 18082 3587
rect 18230 3584 18236 3596
rect 18070 3556 18236 3584
rect 18070 3553 18082 3556
rect 18024 3547 18082 3553
rect 18230 3544 18236 3556
rect 18288 3584 18294 3596
rect 18598 3584 18604 3596
rect 18288 3556 18604 3584
rect 18288 3544 18294 3556
rect 18598 3544 18604 3556
rect 18656 3544 18662 3596
rect 20968 3587 21026 3593
rect 20968 3553 20980 3587
rect 21014 3584 21026 3587
rect 21450 3584 21456 3596
rect 21014 3556 21456 3584
rect 21014 3553 21026 3556
rect 20968 3547 21026 3553
rect 21450 3544 21456 3556
rect 21508 3544 21514 3596
rect 7282 3516 7288 3528
rect 7243 3488 7288 3516
rect 7282 3476 7288 3488
rect 7340 3476 7346 3528
rect 9674 3516 9680 3528
rect 9635 3488 9680 3516
rect 9674 3476 9680 3488
rect 9732 3476 9738 3528
rect 11793 3519 11851 3525
rect 11793 3485 11805 3519
rect 11839 3516 11851 3519
rect 11882 3516 11888 3528
rect 11839 3488 11888 3516
rect 11839 3485 11851 3488
rect 11793 3479 11851 3485
rect 11882 3476 11888 3488
rect 11940 3476 11946 3528
rect 14369 3519 14427 3525
rect 14369 3485 14381 3519
rect 14415 3516 14427 3519
rect 15654 3516 15660 3528
rect 14415 3488 15660 3516
rect 14415 3485 14427 3488
rect 14369 3479 14427 3485
rect 15654 3476 15660 3488
rect 15712 3476 15718 3528
rect 7834 3448 7840 3460
rect 7795 3420 7840 3448
rect 7834 3408 7840 3420
rect 7892 3408 7898 3460
rect 12618 3408 12624 3460
rect 12676 3448 12682 3460
rect 13081 3451 13139 3457
rect 13081 3448 13093 3451
rect 12676 3420 13093 3448
rect 12676 3408 12682 3420
rect 13081 3417 13093 3420
rect 13127 3448 13139 3451
rect 15562 3448 15568 3460
rect 13127 3420 15568 3448
rect 13127 3417 13139 3420
rect 13081 3411 13139 3417
rect 15562 3408 15568 3420
rect 15620 3408 15626 3460
rect 15930 3448 15936 3460
rect 15891 3420 15936 3448
rect 15930 3408 15936 3420
rect 15988 3408 15994 3460
rect 16022 3408 16028 3460
rect 16080 3448 16086 3460
rect 17037 3451 17095 3457
rect 17037 3448 17049 3451
rect 16080 3420 17049 3448
rect 16080 3408 16086 3420
rect 17037 3417 17049 3420
rect 17083 3417 17095 3451
rect 17037 3411 17095 3417
rect 4430 3380 4436 3392
rect 4391 3352 4436 3380
rect 4430 3340 4436 3352
rect 4488 3340 4494 3392
rect 4522 3340 4528 3392
rect 4580 3380 4586 3392
rect 5261 3383 5319 3389
rect 5261 3380 5273 3383
rect 4580 3352 5273 3380
rect 4580 3340 4586 3352
rect 5261 3349 5273 3352
rect 5307 3380 5319 3383
rect 5859 3383 5917 3389
rect 5859 3380 5871 3383
rect 5307 3352 5871 3380
rect 5307 3349 5319 3352
rect 5261 3343 5319 3349
rect 5859 3349 5871 3352
rect 5905 3349 5917 3383
rect 5859 3343 5917 3349
rect 6178 3340 6184 3392
rect 6236 3380 6242 3392
rect 6454 3380 6460 3392
rect 6236 3352 6460 3380
rect 6236 3340 6242 3352
rect 6454 3340 6460 3352
rect 6512 3380 6518 3392
rect 7009 3383 7067 3389
rect 7009 3380 7021 3383
rect 6512 3352 7021 3380
rect 6512 3340 6518 3352
rect 7009 3349 7021 3352
rect 7055 3349 7067 3383
rect 10594 3380 10600 3392
rect 10555 3352 10600 3380
rect 7009 3343 7067 3349
rect 10594 3340 10600 3352
rect 10652 3380 10658 3392
rect 10873 3383 10931 3389
rect 10873 3380 10885 3383
rect 10652 3352 10885 3380
rect 10652 3340 10658 3352
rect 10873 3349 10885 3352
rect 10919 3349 10931 3383
rect 10873 3343 10931 3349
rect 11146 3340 11152 3392
rect 11204 3380 11210 3392
rect 11241 3383 11299 3389
rect 11241 3380 11253 3383
rect 11204 3352 11253 3380
rect 11204 3340 11210 3352
rect 11241 3349 11253 3352
rect 11287 3349 11299 3383
rect 11241 3343 11299 3349
rect 1104 3290 22816 3312
rect 1104 3238 4982 3290
rect 5034 3238 5046 3290
rect 5098 3238 5110 3290
rect 5162 3238 5174 3290
rect 5226 3238 12982 3290
rect 13034 3238 13046 3290
rect 13098 3238 13110 3290
rect 13162 3238 13174 3290
rect 13226 3238 20982 3290
rect 21034 3238 21046 3290
rect 21098 3238 21110 3290
rect 21162 3238 21174 3290
rect 21226 3238 22816 3290
rect 1104 3216 22816 3238
rect 1578 3176 1584 3188
rect 1539 3148 1584 3176
rect 1578 3136 1584 3148
rect 1636 3136 1642 3188
rect 3329 3179 3387 3185
rect 3329 3145 3341 3179
rect 3375 3176 3387 3179
rect 4246 3176 4252 3188
rect 3375 3148 4252 3176
rect 3375 3145 3387 3148
rect 3329 3139 3387 3145
rect 4246 3136 4252 3148
rect 4304 3136 4310 3188
rect 4341 3179 4399 3185
rect 4341 3145 4353 3179
rect 4387 3176 4399 3179
rect 4430 3176 4436 3188
rect 4387 3148 4436 3176
rect 4387 3145 4399 3148
rect 4341 3139 4399 3145
rect 4430 3136 4436 3148
rect 4488 3136 4494 3188
rect 6546 3176 6552 3188
rect 6507 3148 6552 3176
rect 6546 3136 6552 3148
rect 6604 3136 6610 3188
rect 7282 3136 7288 3188
rect 7340 3176 7346 3188
rect 8389 3179 8447 3185
rect 8389 3176 8401 3179
rect 7340 3148 8401 3176
rect 7340 3136 7346 3148
rect 8389 3145 8401 3148
rect 8435 3145 8447 3179
rect 8389 3139 8447 3145
rect 9674 3136 9680 3188
rect 9732 3176 9738 3188
rect 10965 3179 11023 3185
rect 10965 3176 10977 3179
rect 9732 3148 10977 3176
rect 9732 3136 9738 3148
rect 10965 3145 10977 3148
rect 11011 3145 11023 3179
rect 10965 3139 11023 3145
rect 13633 3179 13691 3185
rect 13633 3145 13645 3179
rect 13679 3176 13691 3179
rect 14274 3176 14280 3188
rect 13679 3148 14280 3176
rect 13679 3145 13691 3148
rect 13633 3139 13691 3145
rect 14274 3136 14280 3148
rect 14332 3176 14338 3188
rect 15013 3179 15071 3185
rect 15013 3176 15025 3179
rect 14332 3148 15025 3176
rect 14332 3136 14338 3148
rect 15013 3145 15025 3148
rect 15059 3176 15071 3179
rect 15381 3179 15439 3185
rect 15381 3176 15393 3179
rect 15059 3148 15393 3176
rect 15059 3145 15071 3148
rect 15013 3139 15071 3145
rect 15381 3145 15393 3148
rect 15427 3176 15439 3179
rect 15470 3176 15476 3188
rect 15427 3148 15476 3176
rect 15427 3145 15439 3148
rect 15381 3139 15439 3145
rect 15470 3136 15476 3148
rect 15528 3136 15534 3188
rect 15654 3176 15660 3188
rect 15615 3148 15660 3176
rect 15654 3136 15660 3148
rect 15712 3136 15718 3188
rect 16850 3176 16856 3188
rect 16811 3148 16856 3176
rect 16850 3136 16856 3148
rect 16908 3136 16914 3188
rect 19242 3136 19248 3188
rect 19300 3176 19306 3188
rect 19337 3179 19395 3185
rect 19337 3176 19349 3179
rect 19300 3148 19349 3176
rect 19300 3136 19306 3148
rect 19337 3145 19349 3148
rect 19383 3145 19395 3179
rect 19337 3139 19395 3145
rect 20806 3136 20812 3188
rect 20864 3176 20870 3188
rect 21039 3179 21097 3185
rect 21039 3176 21051 3179
rect 20864 3148 21051 3176
rect 20864 3136 20870 3148
rect 21039 3145 21051 3148
rect 21085 3145 21097 3179
rect 21450 3176 21456 3188
rect 21411 3148 21456 3176
rect 21039 3139 21097 3145
rect 21450 3136 21456 3148
rect 21508 3136 21514 3188
rect 3559 3111 3617 3117
rect 3559 3077 3571 3111
rect 3605 3108 3617 3111
rect 8478 3108 8484 3120
rect 3605 3080 8484 3108
rect 3605 3077 3617 3080
rect 3559 3071 3617 3077
rect 8478 3068 8484 3080
rect 8536 3068 8542 3120
rect 9582 3068 9588 3120
rect 9640 3108 9646 3120
rect 11333 3111 11391 3117
rect 11333 3108 11345 3111
rect 9640 3080 11345 3108
rect 9640 3068 9646 3080
rect 11333 3077 11345 3080
rect 11379 3077 11391 3111
rect 11333 3071 11391 3077
rect 14001 3111 14059 3117
rect 14001 3077 14013 3111
rect 14047 3108 14059 3111
rect 14458 3108 14464 3120
rect 14047 3080 14464 3108
rect 14047 3077 14059 3080
rect 14001 3071 14059 3077
rect 14458 3068 14464 3080
rect 14516 3108 14522 3120
rect 17678 3108 17684 3120
rect 14516 3080 17684 3108
rect 14516 3068 14522 3080
rect 17678 3068 17684 3080
rect 17736 3068 17742 3120
rect 4522 3040 4528 3052
rect 4483 3012 4528 3040
rect 4522 3000 4528 3012
rect 4580 3000 4586 3052
rect 4706 3000 4712 3052
rect 4764 3040 4770 3052
rect 4801 3043 4859 3049
rect 4801 3040 4813 3043
rect 4764 3012 4813 3040
rect 4764 3000 4770 3012
rect 4801 3009 4813 3012
rect 4847 3009 4859 3043
rect 4801 3003 4859 3009
rect 6273 3043 6331 3049
rect 6273 3009 6285 3043
rect 6319 3040 6331 3043
rect 6825 3043 6883 3049
rect 6825 3040 6837 3043
rect 6319 3012 6837 3040
rect 6319 3009 6331 3012
rect 6273 3003 6331 3009
rect 6825 3009 6837 3012
rect 6871 3040 6883 3043
rect 8018 3040 8024 3052
rect 6871 3012 8024 3040
rect 6871 3009 6883 3012
rect 6825 3003 6883 3009
rect 8018 3000 8024 3012
rect 8076 3000 8082 3052
rect 8573 3043 8631 3049
rect 8573 3009 8585 3043
rect 8619 3040 8631 3043
rect 9677 3043 9735 3049
rect 9677 3040 9689 3043
rect 8619 3012 9689 3040
rect 8619 3009 8631 3012
rect 8573 3003 8631 3009
rect 9677 3009 9689 3012
rect 9723 3040 9735 3043
rect 10597 3043 10655 3049
rect 10597 3040 10609 3043
rect 9723 3012 10609 3040
rect 9723 3009 9735 3012
rect 9677 3003 9735 3009
rect 10597 3009 10609 3012
rect 10643 3009 10655 3043
rect 12618 3040 12624 3052
rect 12579 3012 12624 3040
rect 10597 3003 10655 3009
rect 12618 3000 12624 3012
rect 12676 3000 12682 3052
rect 13265 3043 13323 3049
rect 13265 3009 13277 3043
rect 13311 3040 13323 3043
rect 13354 3040 13360 3052
rect 13311 3012 13360 3040
rect 13311 3009 13323 3012
rect 13265 3003 13323 3009
rect 13354 3000 13360 3012
rect 13412 3000 13418 3052
rect 14093 3043 14151 3049
rect 14093 3009 14105 3043
rect 14139 3040 14151 3043
rect 14734 3040 14740 3052
rect 14139 3012 14740 3040
rect 14139 3009 14151 3012
rect 14093 3003 14151 3009
rect 14734 3000 14740 3012
rect 14792 3000 14798 3052
rect 15562 3000 15568 3052
rect 15620 3040 15626 3052
rect 16209 3043 16267 3049
rect 16209 3040 16221 3043
rect 15620 3012 16221 3040
rect 15620 3000 15626 3012
rect 16209 3009 16221 3012
rect 16255 3040 16267 3043
rect 16574 3040 16580 3052
rect 16255 3012 16580 3040
rect 16255 3009 16267 3012
rect 16209 3003 16267 3009
rect 16574 3000 16580 3012
rect 16632 3000 16638 3052
rect 1397 2975 1455 2981
rect 1397 2941 1409 2975
rect 1443 2972 1455 2975
rect 3488 2975 3546 2981
rect 1443 2944 2084 2972
rect 1443 2941 1455 2944
rect 1397 2935 1455 2941
rect 2056 2848 2084 2944
rect 3488 2941 3500 2975
rect 3534 2972 3546 2975
rect 3881 2975 3939 2981
rect 3881 2972 3893 2975
rect 3534 2944 3893 2972
rect 3534 2941 3546 2944
rect 3488 2935 3546 2941
rect 3881 2941 3893 2944
rect 3927 2972 3939 2975
rect 4246 2972 4252 2984
rect 3927 2944 4252 2972
rect 3927 2941 3939 2944
rect 3881 2935 3939 2941
rect 4246 2932 4252 2944
rect 4304 2932 4310 2984
rect 6546 2932 6552 2984
rect 6604 2972 6610 2984
rect 7374 2972 7380 2984
rect 6604 2944 7380 2972
rect 6604 2932 6610 2944
rect 7374 2932 7380 2944
rect 7432 2972 7438 2984
rect 7745 2975 7803 2981
rect 7745 2972 7757 2975
rect 7432 2944 7757 2972
rect 7432 2932 7438 2944
rect 7745 2941 7757 2944
rect 7791 2972 7803 2975
rect 8113 2975 8171 2981
rect 8113 2972 8125 2975
rect 7791 2944 8125 2972
rect 7791 2941 7803 2944
rect 7745 2935 7803 2941
rect 8113 2941 8125 2944
rect 8159 2941 8171 2975
rect 11146 2972 11152 2984
rect 11107 2944 11152 2972
rect 8113 2935 8171 2941
rect 11146 2932 11152 2944
rect 11204 2932 11210 2984
rect 19128 2975 19186 2981
rect 19128 2941 19140 2975
rect 19174 2972 19186 2975
rect 19242 2972 19248 2984
rect 19174 2944 19248 2972
rect 19174 2941 19186 2944
rect 19128 2935 19186 2941
rect 19242 2932 19248 2944
rect 19300 2972 19306 2984
rect 19521 2975 19579 2981
rect 19521 2972 19533 2975
rect 19300 2944 19533 2972
rect 19300 2932 19306 2944
rect 19521 2941 19533 2944
rect 19567 2941 19579 2975
rect 19521 2935 19579 2941
rect 20968 2975 21026 2981
rect 20968 2941 20980 2975
rect 21014 2972 21026 2975
rect 21014 2944 21864 2972
rect 21014 2941 21026 2944
rect 20968 2935 21026 2941
rect 4617 2907 4675 2913
rect 4617 2873 4629 2907
rect 4663 2873 4675 2907
rect 4617 2867 4675 2873
rect 2038 2836 2044 2848
rect 1999 2808 2044 2836
rect 2038 2796 2044 2808
rect 2096 2796 2102 2848
rect 4430 2796 4436 2848
rect 4488 2836 4494 2848
rect 4632 2836 4660 2867
rect 6638 2864 6644 2916
rect 6696 2904 6702 2916
rect 7146 2907 7204 2913
rect 7146 2904 7158 2907
rect 6696 2876 7158 2904
rect 6696 2864 6702 2876
rect 7146 2873 7158 2876
rect 7192 2873 7204 2907
rect 7146 2867 7204 2873
rect 9125 2907 9183 2913
rect 9125 2873 9137 2907
rect 9171 2904 9183 2907
rect 9766 2904 9772 2916
rect 9171 2876 9772 2904
rect 9171 2873 9183 2876
rect 9125 2867 9183 2873
rect 5810 2836 5816 2848
rect 4488 2808 4660 2836
rect 5771 2808 5816 2836
rect 4488 2796 4494 2808
rect 5810 2796 5816 2808
rect 5868 2796 5874 2848
rect 7161 2836 7189 2867
rect 9766 2864 9772 2876
rect 9824 2864 9830 2916
rect 10318 2904 10324 2916
rect 10279 2876 10324 2904
rect 10318 2864 10324 2876
rect 10376 2864 10382 2916
rect 12253 2907 12311 2913
rect 12253 2873 12265 2907
rect 12299 2904 12311 2907
rect 12710 2904 12716 2916
rect 12299 2876 12716 2904
rect 12299 2873 12311 2876
rect 12253 2867 12311 2873
rect 12710 2864 12716 2876
rect 12768 2864 12774 2916
rect 14918 2864 14924 2916
rect 14976 2904 14982 2916
rect 15746 2904 15752 2916
rect 14976 2876 15752 2904
rect 14976 2864 14982 2876
rect 15746 2864 15752 2876
rect 15804 2904 15810 2916
rect 15933 2907 15991 2913
rect 15933 2904 15945 2907
rect 15804 2876 15945 2904
rect 15804 2864 15810 2876
rect 15933 2873 15945 2876
rect 15979 2873 15991 2907
rect 15933 2867 15991 2873
rect 16025 2907 16083 2913
rect 16025 2873 16037 2907
rect 16071 2873 16083 2907
rect 16025 2867 16083 2873
rect 9401 2839 9459 2845
rect 9401 2836 9413 2839
rect 7161 2808 9413 2836
rect 9401 2805 9413 2808
rect 9447 2836 9459 2839
rect 9950 2836 9956 2848
rect 9447 2808 9956 2836
rect 9447 2805 9459 2808
rect 9401 2799 9459 2805
rect 9950 2796 9956 2808
rect 10008 2836 10014 2848
rect 11790 2836 11796 2848
rect 10008 2808 11796 2836
rect 10008 2796 10014 2808
rect 11790 2796 11796 2808
rect 11848 2796 11854 2848
rect 14458 2836 14464 2848
rect 14419 2808 14464 2836
rect 14458 2796 14464 2808
rect 14516 2796 14522 2848
rect 15654 2796 15660 2848
rect 15712 2836 15718 2848
rect 16040 2836 16068 2867
rect 18046 2836 18052 2848
rect 15712 2808 16068 2836
rect 18007 2808 18052 2836
rect 15712 2796 15718 2808
rect 18046 2796 18052 2808
rect 18104 2796 18110 2848
rect 18598 2836 18604 2848
rect 18559 2808 18604 2836
rect 18598 2796 18604 2808
rect 18656 2796 18662 2848
rect 21836 2845 21864 2944
rect 21821 2839 21879 2845
rect 21821 2805 21833 2839
rect 21867 2836 21879 2839
rect 22278 2836 22284 2848
rect 21867 2808 22284 2836
rect 21867 2805 21879 2808
rect 21821 2799 21879 2805
rect 22278 2796 22284 2808
rect 22336 2796 22342 2848
rect 1104 2746 22816 2768
rect 1104 2694 8982 2746
rect 9034 2694 9046 2746
rect 9098 2694 9110 2746
rect 9162 2694 9174 2746
rect 9226 2694 16982 2746
rect 17034 2694 17046 2746
rect 17098 2694 17110 2746
rect 17162 2694 17174 2746
rect 17226 2694 22816 2746
rect 1104 2672 22816 2694
rect 1535 2635 1593 2641
rect 1535 2601 1547 2635
rect 1581 2632 1593 2635
rect 1762 2632 1768 2644
rect 1581 2604 1768 2632
rect 1581 2601 1593 2604
rect 1535 2595 1593 2601
rect 1762 2592 1768 2604
rect 1820 2592 1826 2644
rect 3510 2592 3516 2644
rect 3568 2632 3574 2644
rect 4203 2635 4261 2641
rect 4203 2632 4215 2635
rect 3568 2604 4215 2632
rect 3568 2592 3574 2604
rect 4203 2601 4215 2604
rect 4249 2601 4261 2635
rect 4203 2595 4261 2601
rect 8803 2635 8861 2641
rect 8803 2601 8815 2635
rect 8849 2632 8861 2635
rect 11146 2632 11152 2644
rect 8849 2604 11152 2632
rect 8849 2601 8861 2604
rect 8803 2595 8861 2601
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 11882 2632 11888 2644
rect 11843 2604 11888 2632
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 12434 2632 12440 2644
rect 12395 2604 12440 2632
rect 12434 2592 12440 2604
rect 12492 2632 12498 2644
rect 12492 2604 12848 2632
rect 12492 2592 12498 2604
rect 3145 2567 3203 2573
rect 3145 2533 3157 2567
rect 3191 2564 3203 2567
rect 6178 2564 6184 2576
rect 3191 2536 6184 2564
rect 3191 2533 3203 2536
rect 3145 2527 3203 2533
rect 6178 2524 6184 2536
rect 6236 2524 6242 2576
rect 7285 2567 7343 2573
rect 7285 2564 7297 2567
rect 6656 2536 7297 2564
rect 1118 2456 1124 2508
rect 1176 2496 1182 2508
rect 1432 2499 1490 2505
rect 1432 2496 1444 2499
rect 1176 2468 1444 2496
rect 1176 2456 1182 2468
rect 1432 2465 1444 2468
rect 1478 2496 1490 2499
rect 1857 2499 1915 2505
rect 1857 2496 1869 2499
rect 1478 2468 1869 2496
rect 1478 2465 1490 2468
rect 1432 2459 1490 2465
rect 1857 2465 1869 2468
rect 1903 2465 1915 2499
rect 2501 2499 2559 2505
rect 2501 2496 2513 2499
rect 1857 2459 1915 2465
rect 2240 2468 2513 2496
rect 842 2252 848 2304
rect 900 2292 906 2304
rect 2240 2301 2268 2468
rect 2501 2465 2513 2468
rect 2547 2465 2559 2499
rect 2501 2459 2559 2465
rect 4132 2499 4190 2505
rect 4132 2465 4144 2499
rect 4178 2496 4190 2499
rect 5169 2499 5227 2505
rect 4178 2468 4660 2496
rect 4178 2465 4190 2468
rect 4132 2459 4190 2465
rect 4632 2301 4660 2468
rect 5169 2465 5181 2499
rect 5215 2496 5227 2499
rect 5353 2499 5411 2505
rect 5353 2496 5365 2499
rect 5215 2468 5365 2496
rect 5215 2465 5227 2468
rect 5169 2459 5227 2465
rect 5353 2465 5365 2468
rect 5399 2496 5411 2499
rect 6546 2496 6552 2508
rect 5399 2468 6552 2496
rect 5399 2465 5411 2468
rect 5353 2459 5411 2465
rect 6546 2456 6552 2468
rect 6604 2456 6610 2508
rect 6656 2437 6684 2536
rect 7285 2533 7297 2536
rect 7331 2533 7343 2567
rect 7834 2564 7840 2576
rect 7795 2536 7840 2564
rect 7285 2527 7343 2533
rect 7834 2524 7840 2536
rect 7892 2564 7898 2576
rect 9125 2567 9183 2573
rect 9125 2564 9137 2567
rect 7892 2536 9137 2564
rect 7892 2524 7898 2536
rect 9125 2533 9137 2536
rect 9171 2533 9183 2567
rect 9125 2527 9183 2533
rect 9585 2567 9643 2573
rect 9585 2533 9597 2567
rect 9631 2564 9643 2567
rect 9953 2567 10011 2573
rect 9953 2564 9965 2567
rect 9631 2536 9965 2564
rect 9631 2533 9643 2536
rect 9585 2527 9643 2533
rect 9953 2533 9965 2536
rect 9999 2564 10011 2567
rect 10594 2564 10600 2576
rect 9999 2536 10600 2564
rect 9999 2533 10011 2536
rect 9953 2527 10011 2533
rect 8700 2499 8758 2505
rect 8700 2465 8712 2499
rect 8746 2465 8758 2499
rect 8700 2459 8758 2465
rect 5997 2431 6055 2437
rect 5997 2397 6009 2431
rect 6043 2428 6055 2431
rect 6641 2431 6699 2437
rect 6641 2428 6653 2431
rect 6043 2400 6653 2428
rect 6043 2397 6055 2400
rect 5997 2391 6055 2397
rect 6641 2397 6653 2400
rect 6687 2397 6699 2431
rect 6641 2391 6699 2397
rect 7193 2431 7251 2437
rect 7193 2397 7205 2431
rect 7239 2428 7251 2431
rect 8110 2428 8116 2440
rect 7239 2400 8116 2428
rect 7239 2397 7251 2400
rect 7193 2391 7251 2397
rect 6365 2363 6423 2369
rect 6365 2329 6377 2363
rect 6411 2360 6423 2363
rect 7208 2360 7236 2391
rect 8110 2388 8116 2400
rect 8168 2388 8174 2440
rect 6411 2332 7236 2360
rect 8573 2363 8631 2369
rect 6411 2329 6423 2332
rect 6365 2323 6423 2329
rect 8573 2329 8585 2363
rect 8619 2360 8631 2363
rect 8715 2360 8743 2459
rect 9140 2428 9168 2527
rect 10594 2524 10600 2536
rect 10652 2524 10658 2576
rect 11241 2567 11299 2573
rect 11241 2533 11253 2567
rect 11287 2564 11299 2567
rect 12066 2564 12072 2576
rect 11287 2536 12072 2564
rect 11287 2533 11299 2536
rect 11241 2527 11299 2533
rect 11348 2505 11376 2536
rect 12066 2524 12072 2536
rect 12124 2524 12130 2576
rect 12820 2573 12848 2604
rect 13262 2592 13268 2644
rect 13320 2632 13326 2644
rect 14369 2635 14427 2641
rect 14369 2632 14381 2635
rect 13320 2604 14381 2632
rect 13320 2592 13326 2604
rect 14369 2601 14381 2604
rect 14415 2601 14427 2635
rect 14369 2595 14427 2601
rect 15746 2592 15752 2644
rect 15804 2632 15810 2644
rect 16485 2635 16543 2641
rect 16485 2632 16497 2635
rect 15804 2604 16497 2632
rect 15804 2592 15810 2604
rect 16485 2601 16497 2604
rect 16531 2601 16543 2635
rect 16485 2595 16543 2601
rect 19794 2592 19800 2644
rect 19852 2632 19858 2644
rect 20073 2635 20131 2641
rect 20073 2632 20085 2635
rect 19852 2604 20085 2632
rect 19852 2592 19858 2604
rect 20073 2601 20085 2604
rect 20119 2601 20131 2635
rect 20073 2595 20131 2601
rect 12805 2567 12863 2573
rect 12805 2533 12817 2567
rect 12851 2533 12863 2567
rect 13354 2564 13360 2576
rect 13315 2536 13360 2564
rect 12805 2527 12863 2533
rect 13354 2524 13360 2536
rect 13412 2524 13418 2576
rect 15654 2573 15660 2576
rect 15289 2567 15347 2573
rect 15289 2533 15301 2567
rect 15335 2564 15347 2567
rect 15634 2567 15660 2573
rect 15634 2564 15646 2567
rect 15335 2536 15646 2564
rect 15335 2533 15347 2536
rect 15289 2527 15347 2533
rect 15634 2533 15646 2536
rect 15634 2527 15660 2533
rect 15654 2524 15660 2527
rect 15712 2524 15718 2576
rect 11333 2499 11391 2505
rect 11333 2496 11345 2499
rect 11311 2468 11345 2496
rect 11333 2465 11345 2468
rect 11379 2465 11391 2499
rect 14090 2496 14096 2508
rect 14051 2468 14096 2496
rect 11333 2459 11391 2465
rect 14090 2456 14096 2468
rect 14148 2456 14154 2508
rect 16666 2456 16672 2508
rect 16724 2496 16730 2508
rect 17037 2499 17095 2505
rect 17037 2496 17049 2499
rect 16724 2468 17049 2496
rect 16724 2456 16730 2468
rect 17037 2465 17049 2468
rect 17083 2496 17095 2499
rect 17589 2499 17647 2505
rect 17589 2496 17601 2499
rect 17083 2468 17601 2496
rect 17083 2465 17095 2468
rect 17037 2459 17095 2465
rect 17589 2465 17601 2468
rect 17635 2465 17647 2499
rect 17589 2459 17647 2465
rect 18325 2499 18383 2505
rect 18325 2465 18337 2499
rect 18371 2465 18383 2499
rect 18325 2459 18383 2465
rect 19521 2499 19579 2505
rect 19521 2465 19533 2499
rect 19567 2496 19579 2499
rect 19812 2496 19840 2592
rect 19567 2468 19840 2496
rect 21244 2499 21302 2505
rect 19567 2465 19579 2468
rect 19521 2459 19579 2465
rect 21244 2465 21256 2499
rect 21290 2496 21302 2499
rect 21290 2468 21772 2496
rect 21290 2465 21302 2468
rect 21244 2459 21302 2465
rect 9861 2431 9919 2437
rect 9861 2428 9873 2431
rect 9140 2400 9873 2428
rect 9861 2397 9873 2400
rect 9907 2397 9919 2431
rect 10318 2428 10324 2440
rect 10279 2400 10324 2428
rect 9861 2391 9919 2397
rect 10318 2388 10324 2400
rect 10376 2388 10382 2440
rect 12713 2431 12771 2437
rect 12713 2397 12725 2431
rect 12759 2428 12771 2431
rect 13633 2431 13691 2437
rect 13633 2428 13645 2431
rect 12759 2400 13645 2428
rect 12759 2397 12771 2400
rect 12713 2391 12771 2397
rect 13633 2397 13645 2400
rect 13679 2428 13691 2431
rect 14921 2431 14979 2437
rect 13679 2400 13814 2428
rect 13679 2397 13691 2400
rect 13633 2391 13691 2397
rect 10336 2360 10364 2388
rect 8619 2332 10364 2360
rect 8619 2329 8631 2332
rect 8573 2323 8631 2329
rect 10502 2320 10508 2372
rect 10560 2360 10566 2372
rect 11517 2363 11575 2369
rect 11517 2360 11529 2363
rect 10560 2332 11529 2360
rect 10560 2320 10566 2332
rect 11517 2329 11529 2332
rect 11563 2329 11575 2363
rect 13786 2360 13814 2400
rect 14921 2397 14933 2431
rect 14967 2428 14979 2431
rect 15565 2431 15623 2437
rect 15565 2428 15577 2431
rect 14967 2400 15577 2428
rect 14967 2397 14979 2400
rect 14921 2391 14979 2397
rect 15565 2397 15577 2400
rect 15611 2428 15623 2431
rect 18046 2428 18052 2440
rect 15611 2400 18052 2428
rect 15611 2397 15623 2400
rect 15565 2391 15623 2397
rect 18046 2388 18052 2400
rect 18104 2388 18110 2440
rect 18340 2428 18368 2459
rect 18598 2428 18604 2440
rect 18340 2400 18604 2428
rect 18598 2388 18604 2400
rect 18656 2428 18662 2440
rect 18969 2431 19027 2437
rect 18969 2428 18981 2431
rect 18656 2400 18981 2428
rect 18656 2388 18662 2400
rect 18969 2397 18981 2400
rect 19015 2428 19027 2431
rect 19610 2428 19616 2440
rect 19015 2400 19616 2428
rect 19015 2397 19027 2400
rect 18969 2391 19027 2397
rect 19610 2388 19616 2400
rect 19668 2388 19674 2440
rect 15930 2360 15936 2372
rect 13786 2332 15936 2360
rect 11517 2323 11575 2329
rect 15930 2320 15936 2332
rect 15988 2360 15994 2372
rect 16117 2363 16175 2369
rect 16117 2360 16129 2363
rect 15988 2332 16129 2360
rect 15988 2320 15994 2332
rect 16117 2329 16129 2332
rect 16163 2329 16175 2363
rect 16117 2323 16175 2329
rect 19705 2363 19763 2369
rect 19705 2329 19717 2363
rect 19751 2360 19763 2363
rect 20438 2360 20444 2372
rect 19751 2332 20444 2360
rect 19751 2329 19763 2332
rect 19705 2323 19763 2329
rect 20438 2320 20444 2332
rect 20496 2320 20502 2372
rect 2225 2295 2283 2301
rect 2225 2292 2237 2295
rect 900 2264 2237 2292
rect 900 2252 906 2264
rect 2225 2261 2237 2264
rect 2271 2261 2283 2295
rect 2225 2255 2283 2261
rect 4617 2295 4675 2301
rect 4617 2261 4629 2295
rect 4663 2292 4675 2295
rect 4798 2292 4804 2304
rect 4663 2264 4804 2292
rect 4663 2261 4675 2264
rect 4617 2255 4675 2261
rect 4798 2252 4804 2264
rect 4856 2252 4862 2304
rect 16942 2252 16948 2304
rect 17000 2292 17006 2304
rect 17221 2295 17279 2301
rect 17221 2292 17233 2295
rect 17000 2264 17233 2292
rect 17000 2252 17006 2264
rect 17221 2261 17233 2264
rect 17267 2261 17279 2295
rect 17221 2255 17279 2261
rect 18230 2252 18236 2304
rect 18288 2292 18294 2304
rect 18509 2295 18567 2301
rect 18509 2292 18521 2295
rect 18288 2264 18521 2292
rect 18288 2252 18294 2264
rect 18509 2261 18521 2264
rect 18555 2261 18567 2295
rect 18509 2255 18567 2261
rect 18966 2252 18972 2304
rect 19024 2292 19030 2304
rect 21744 2301 21772 2468
rect 21315 2295 21373 2301
rect 21315 2292 21327 2295
rect 19024 2264 21327 2292
rect 19024 2252 19030 2264
rect 21315 2261 21327 2264
rect 21361 2261 21373 2295
rect 21315 2255 21373 2261
rect 21729 2295 21787 2301
rect 21729 2261 21741 2295
rect 21775 2292 21787 2295
rect 23198 2292 23204 2304
rect 21775 2264 23204 2292
rect 21775 2261 21787 2264
rect 21729 2255 21787 2261
rect 23198 2252 23204 2264
rect 23256 2252 23262 2304
rect 1104 2202 22816 2224
rect 1104 2150 4982 2202
rect 5034 2150 5046 2202
rect 5098 2150 5110 2202
rect 5162 2150 5174 2202
rect 5226 2150 12982 2202
rect 13034 2150 13046 2202
rect 13098 2150 13110 2202
rect 13162 2150 13174 2202
rect 13226 2150 20982 2202
rect 21034 2150 21046 2202
rect 21098 2150 21110 2202
rect 21162 2150 21174 2202
rect 21226 2150 22816 2202
rect 1104 2128 22816 2150
rect 5810 2048 5816 2100
rect 5868 2088 5874 2100
rect 12158 2088 12164 2100
rect 5868 2060 12164 2088
rect 5868 2048 5874 2060
rect 12158 2048 12164 2060
rect 12216 2048 12222 2100
rect 11514 76 11520 128
rect 11572 116 11578 128
rect 13262 116 13268 128
rect 11572 88 13268 116
rect 11572 76 11578 88
rect 13262 76 13268 88
rect 13320 76 13326 128
<< via1 >>
rect 20 23536 72 23588
rect 572 23536 624 23588
rect 4982 21734 5034 21786
rect 5046 21734 5098 21786
rect 5110 21734 5162 21786
rect 5174 21734 5226 21786
rect 12982 21734 13034 21786
rect 13046 21734 13098 21786
rect 13110 21734 13162 21786
rect 13174 21734 13226 21786
rect 20982 21734 21034 21786
rect 21046 21734 21098 21786
rect 21110 21734 21162 21786
rect 21174 21734 21226 21786
rect 20076 21675 20128 21684
rect 20076 21641 20085 21675
rect 20085 21641 20119 21675
rect 20119 21641 20128 21675
rect 20076 21632 20128 21641
rect 8392 21292 8444 21344
rect 20076 21428 20128 21480
rect 10048 21292 10100 21344
rect 19340 21292 19392 21344
rect 8982 21190 9034 21242
rect 9046 21190 9098 21242
rect 9110 21190 9162 21242
rect 9174 21190 9226 21242
rect 16982 21190 17034 21242
rect 17046 21190 17098 21242
rect 17110 21190 17162 21242
rect 17174 21190 17226 21242
rect 9312 21088 9364 21140
rect 13268 21088 13320 21140
rect 19248 21088 19300 21140
rect 12348 20995 12400 21004
rect 12348 20961 12357 20995
rect 12357 20961 12391 20995
rect 12391 20961 12400 20995
rect 12348 20952 12400 20961
rect 18052 20995 18104 21004
rect 18052 20961 18061 20995
rect 18061 20961 18095 20995
rect 18095 20961 18104 20995
rect 18052 20952 18104 20961
rect 19984 20952 20036 21004
rect 19524 20748 19576 20800
rect 4982 20646 5034 20698
rect 5046 20646 5098 20698
rect 5110 20646 5162 20698
rect 5174 20646 5226 20698
rect 12982 20646 13034 20698
rect 13046 20646 13098 20698
rect 13110 20646 13162 20698
rect 13174 20646 13226 20698
rect 20982 20646 21034 20698
rect 21046 20646 21098 20698
rect 21110 20646 21162 20698
rect 21174 20646 21226 20698
rect 2780 20544 2832 20596
rect 4528 20587 4580 20596
rect 4528 20553 4537 20587
rect 4537 20553 4571 20587
rect 4571 20553 4580 20587
rect 4528 20544 4580 20553
rect 7932 20587 7984 20596
rect 7932 20553 7941 20587
rect 7941 20553 7975 20587
rect 7975 20553 7984 20587
rect 7932 20544 7984 20553
rect 8392 20587 8444 20596
rect 8392 20553 8401 20587
rect 8401 20553 8435 20587
rect 8435 20553 8444 20587
rect 8392 20544 8444 20553
rect 14188 20587 14240 20596
rect 14188 20553 14197 20587
rect 14197 20553 14231 20587
rect 14231 20553 14240 20587
rect 14188 20544 14240 20553
rect 12256 20408 12308 20460
rect 4528 20340 4580 20392
rect 8392 20340 8444 20392
rect 13912 20340 13964 20392
rect 17868 20544 17920 20596
rect 20444 20544 20496 20596
rect 21732 20544 21784 20596
rect 19984 20519 20036 20528
rect 19984 20485 19993 20519
rect 19993 20485 20027 20519
rect 20027 20485 20036 20519
rect 19984 20476 20036 20485
rect 18972 20383 19024 20392
rect 18972 20349 18981 20383
rect 18981 20349 19015 20383
rect 19015 20349 19024 20383
rect 18972 20340 19024 20349
rect 19892 20340 19944 20392
rect 9404 20315 9456 20324
rect 9404 20281 9413 20315
rect 9413 20281 9447 20315
rect 9447 20281 9456 20315
rect 9404 20272 9456 20281
rect 10048 20315 10100 20324
rect 2412 20204 2464 20256
rect 8852 20204 8904 20256
rect 9312 20204 9364 20256
rect 10048 20281 10057 20315
rect 10057 20281 10091 20315
rect 10091 20281 10100 20315
rect 10048 20272 10100 20281
rect 12532 20315 12584 20324
rect 12532 20281 12541 20315
rect 12541 20281 12575 20315
rect 12575 20281 12584 20315
rect 12532 20272 12584 20281
rect 12624 20315 12676 20324
rect 12624 20281 12633 20315
rect 12633 20281 12667 20315
rect 12667 20281 12676 20315
rect 12624 20272 12676 20281
rect 16396 20272 16448 20324
rect 18052 20272 18104 20324
rect 11612 20204 11664 20256
rect 12348 20204 12400 20256
rect 14740 20204 14792 20256
rect 8982 20102 9034 20154
rect 9046 20102 9098 20154
rect 9110 20102 9162 20154
rect 9174 20102 9226 20154
rect 16982 20102 17034 20154
rect 17046 20102 17098 20154
rect 17110 20102 17162 20154
rect 17174 20102 17226 20154
rect 18880 20000 18932 20052
rect 9772 19932 9824 19984
rect 11704 19975 11756 19984
rect 11704 19941 11713 19975
rect 11713 19941 11747 19975
rect 11747 19941 11756 19975
rect 11704 19932 11756 19941
rect 12624 19932 12676 19984
rect 13360 19932 13412 19984
rect 17500 19932 17552 19984
rect 19340 19975 19392 19984
rect 19340 19941 19349 19975
rect 19349 19941 19383 19975
rect 19383 19941 19392 19975
rect 19340 19932 19392 19941
rect 1584 19864 1636 19916
rect 8024 19864 8076 19916
rect 15844 19907 15896 19916
rect 15844 19873 15853 19907
rect 15853 19873 15887 19907
rect 15887 19873 15896 19907
rect 15844 19864 15896 19873
rect 20812 19864 20864 19916
rect 23020 19864 23072 19916
rect 10048 19839 10100 19848
rect 10048 19805 10057 19839
rect 10057 19805 10091 19839
rect 10091 19805 10100 19839
rect 10048 19796 10100 19805
rect 11612 19839 11664 19848
rect 11612 19805 11621 19839
rect 11621 19805 11655 19839
rect 11655 19805 11664 19839
rect 11612 19796 11664 19805
rect 13544 19796 13596 19848
rect 17224 19839 17276 19848
rect 17224 19805 17233 19839
rect 17233 19805 17267 19839
rect 17267 19805 17276 19839
rect 17224 19796 17276 19805
rect 19064 19796 19116 19848
rect 19984 19839 20036 19848
rect 19984 19805 19993 19839
rect 19993 19805 20027 19839
rect 20027 19805 20036 19839
rect 19984 19796 20036 19805
rect 10140 19728 10192 19780
rect 2872 19660 2924 19712
rect 9404 19703 9456 19712
rect 9404 19669 9413 19703
rect 9413 19669 9447 19703
rect 9447 19669 9456 19703
rect 9404 19660 9456 19669
rect 12256 19660 12308 19712
rect 16304 19660 16356 19712
rect 16580 19660 16632 19712
rect 20720 19660 20772 19712
rect 4982 19558 5034 19610
rect 5046 19558 5098 19610
rect 5110 19558 5162 19610
rect 5174 19558 5226 19610
rect 12982 19558 13034 19610
rect 13046 19558 13098 19610
rect 13110 19558 13162 19610
rect 13174 19558 13226 19610
rect 20982 19558 21034 19610
rect 21046 19558 21098 19610
rect 21110 19558 21162 19610
rect 21174 19558 21226 19610
rect 1584 19499 1636 19508
rect 1584 19465 1593 19499
rect 1593 19465 1627 19499
rect 1627 19465 1636 19499
rect 1584 19456 1636 19465
rect 8024 19499 8076 19508
rect 8024 19465 8033 19499
rect 8033 19465 8067 19499
rect 8067 19465 8076 19499
rect 8024 19456 8076 19465
rect 9312 19456 9364 19508
rect 9772 19499 9824 19508
rect 9772 19465 9781 19499
rect 9781 19465 9815 19499
rect 9815 19465 9824 19499
rect 9772 19456 9824 19465
rect 10140 19499 10192 19508
rect 10140 19465 10149 19499
rect 10149 19465 10183 19499
rect 10183 19465 10192 19499
rect 10140 19456 10192 19465
rect 11612 19456 11664 19508
rect 13360 19499 13412 19508
rect 11704 19320 11756 19372
rect 8576 19252 8628 19304
rect 10692 19295 10744 19304
rect 10692 19261 10701 19295
rect 10701 19261 10735 19295
rect 10735 19261 10744 19295
rect 10692 19252 10744 19261
rect 11612 19252 11664 19304
rect 13360 19465 13369 19499
rect 13369 19465 13403 19499
rect 13403 19465 13412 19499
rect 13360 19456 13412 19465
rect 13912 19499 13964 19508
rect 13912 19465 13921 19499
rect 13921 19465 13955 19499
rect 13955 19465 13964 19499
rect 13912 19456 13964 19465
rect 19340 19456 19392 19508
rect 20812 19456 20864 19508
rect 21640 19499 21692 19508
rect 21640 19465 21649 19499
rect 21649 19465 21683 19499
rect 21683 19465 21692 19499
rect 21640 19456 21692 19465
rect 12532 19388 12584 19440
rect 14740 19388 14792 19440
rect 19984 19388 20036 19440
rect 16212 19320 16264 19372
rect 17224 19320 17276 19372
rect 9680 19184 9732 19236
rect 14004 19252 14056 19304
rect 15660 19252 15712 19304
rect 17684 19252 17736 19304
rect 13544 19184 13596 19236
rect 16488 19227 16540 19236
rect 16488 19193 16497 19227
rect 16497 19193 16531 19227
rect 16531 19193 16540 19227
rect 16488 19184 16540 19193
rect 16580 19227 16632 19236
rect 16580 19193 16589 19227
rect 16589 19193 16623 19227
rect 16623 19193 16632 19227
rect 17500 19227 17552 19236
rect 16580 19184 16632 19193
rect 17500 19193 17509 19227
rect 17509 19193 17543 19227
rect 17543 19193 17552 19227
rect 21640 19252 21692 19304
rect 17500 19184 17552 19193
rect 12808 19116 12860 19168
rect 15844 19116 15896 19168
rect 18236 19116 18288 19168
rect 18788 19116 18840 19168
rect 18880 19116 18932 19168
rect 8982 19014 9034 19066
rect 9046 19014 9098 19066
rect 9110 19014 9162 19066
rect 9174 19014 9226 19066
rect 16982 19014 17034 19066
rect 17046 19014 17098 19066
rect 17110 19014 17162 19066
rect 17174 19014 17226 19066
rect 10692 18955 10744 18964
rect 10692 18921 10701 18955
rect 10701 18921 10735 18955
rect 10735 18921 10744 18955
rect 10692 18912 10744 18921
rect 13544 18955 13596 18964
rect 13544 18921 13553 18955
rect 13553 18921 13587 18955
rect 13587 18921 13596 18955
rect 13544 18912 13596 18921
rect 16212 18912 16264 18964
rect 16488 18955 16540 18964
rect 16488 18921 16497 18955
rect 16497 18921 16531 18955
rect 16531 18921 16540 18955
rect 16488 18912 16540 18921
rect 9680 18844 9732 18896
rect 11612 18844 11664 18896
rect 12256 18887 12308 18896
rect 12256 18853 12265 18887
rect 12265 18853 12299 18887
rect 12299 18853 12308 18887
rect 12256 18844 12308 18853
rect 15476 18844 15528 18896
rect 16304 18844 16356 18896
rect 17132 18887 17184 18896
rect 17132 18853 17141 18887
rect 17141 18853 17175 18887
rect 17175 18853 17184 18887
rect 17132 18844 17184 18853
rect 17500 18844 17552 18896
rect 18880 18887 18932 18896
rect 18880 18853 18889 18887
rect 18889 18853 18923 18887
rect 18923 18853 18932 18887
rect 18880 18844 18932 18853
rect 1308 18776 1360 18828
rect 12716 18776 12768 18828
rect 14096 18776 14148 18828
rect 9772 18751 9824 18760
rect 9772 18717 9781 18751
rect 9781 18717 9815 18751
rect 9815 18717 9824 18751
rect 9772 18708 9824 18717
rect 11244 18708 11296 18760
rect 15844 18708 15896 18760
rect 18788 18751 18840 18760
rect 18788 18717 18797 18751
rect 18797 18717 18831 18751
rect 18831 18717 18840 18751
rect 18788 18708 18840 18717
rect 19064 18751 19116 18760
rect 19064 18717 19073 18751
rect 19073 18717 19107 18751
rect 19107 18717 19116 18751
rect 19064 18708 19116 18717
rect 17500 18640 17552 18692
rect 17684 18683 17736 18692
rect 17684 18649 17693 18683
rect 17693 18649 17727 18683
rect 17727 18649 17736 18683
rect 17684 18640 17736 18649
rect 7656 18572 7708 18624
rect 8576 18615 8628 18624
rect 8576 18581 8585 18615
rect 8585 18581 8619 18615
rect 8619 18581 8628 18615
rect 8576 18572 8628 18581
rect 19708 18615 19760 18624
rect 19708 18581 19717 18615
rect 19717 18581 19751 18615
rect 19751 18581 19760 18615
rect 19708 18572 19760 18581
rect 4982 18470 5034 18522
rect 5046 18470 5098 18522
rect 5110 18470 5162 18522
rect 5174 18470 5226 18522
rect 12982 18470 13034 18522
rect 13046 18470 13098 18522
rect 13110 18470 13162 18522
rect 13174 18470 13226 18522
rect 20982 18470 21034 18522
rect 21046 18470 21098 18522
rect 21110 18470 21162 18522
rect 21174 18470 21226 18522
rect 1308 18368 1360 18420
rect 7656 18411 7708 18420
rect 7656 18377 7665 18411
rect 7665 18377 7699 18411
rect 7699 18377 7708 18411
rect 7656 18368 7708 18377
rect 9312 18411 9364 18420
rect 9312 18377 9321 18411
rect 9321 18377 9355 18411
rect 9355 18377 9364 18411
rect 9312 18368 9364 18377
rect 9772 18368 9824 18420
rect 11244 18411 11296 18420
rect 11244 18377 11253 18411
rect 11253 18377 11287 18411
rect 11287 18377 11296 18411
rect 11244 18368 11296 18377
rect 11612 18368 11664 18420
rect 16580 18368 16632 18420
rect 17132 18368 17184 18420
rect 18788 18368 18840 18420
rect 21272 18368 21324 18420
rect 2872 18232 2924 18284
rect 8392 18300 8444 18352
rect 10324 18300 10376 18352
rect 11980 18300 12032 18352
rect 2228 18207 2280 18216
rect 2228 18173 2237 18207
rect 2237 18173 2271 18207
rect 2271 18173 2280 18207
rect 2228 18164 2280 18173
rect 11152 18232 11204 18284
rect 16396 18300 16448 18352
rect 17500 18300 17552 18352
rect 1768 18028 1820 18080
rect 8392 18139 8444 18148
rect 8392 18105 8401 18139
rect 8401 18105 8435 18139
rect 8435 18105 8444 18139
rect 8392 18096 8444 18105
rect 8760 18096 8812 18148
rect 9680 18071 9732 18080
rect 9680 18037 9689 18071
rect 9689 18037 9723 18071
rect 9723 18037 9732 18071
rect 9680 18028 9732 18037
rect 9956 18139 10008 18148
rect 9956 18105 9965 18139
rect 9965 18105 9999 18139
rect 9999 18105 10008 18139
rect 9956 18096 10008 18105
rect 11244 18028 11296 18080
rect 12808 18164 12860 18216
rect 13452 18096 13504 18148
rect 14188 18164 14240 18216
rect 14096 18096 14148 18148
rect 18880 18232 18932 18284
rect 19524 18275 19576 18284
rect 19524 18241 19533 18275
rect 19533 18241 19567 18275
rect 19567 18241 19576 18275
rect 19524 18232 19576 18241
rect 19984 18275 20036 18284
rect 19984 18241 19993 18275
rect 19993 18241 20027 18275
rect 20027 18241 20036 18275
rect 19984 18232 20036 18241
rect 15568 18164 15620 18216
rect 11980 18028 12032 18080
rect 12256 18028 12308 18080
rect 12716 18028 12768 18080
rect 13728 18071 13780 18080
rect 13728 18037 13737 18071
rect 13737 18037 13771 18071
rect 13771 18037 13780 18071
rect 14832 18096 14884 18148
rect 15476 18139 15528 18148
rect 15476 18105 15485 18139
rect 15485 18105 15519 18139
rect 15519 18105 15528 18139
rect 15476 18096 15528 18105
rect 13728 18028 13780 18037
rect 15108 18028 15160 18080
rect 15844 18071 15896 18080
rect 15844 18037 15853 18071
rect 15853 18037 15887 18071
rect 15887 18037 15896 18071
rect 15844 18028 15896 18037
rect 16856 18028 16908 18080
rect 18788 18028 18840 18080
rect 19708 18096 19760 18148
rect 19156 18028 19208 18080
rect 8982 17926 9034 17978
rect 9046 17926 9098 17978
rect 9110 17926 9162 17978
rect 9174 17926 9226 17978
rect 16982 17926 17034 17978
rect 17046 17926 17098 17978
rect 17110 17926 17162 17978
rect 17174 17926 17226 17978
rect 1768 17824 1820 17876
rect 2320 17824 2372 17876
rect 9680 17824 9732 17876
rect 10232 17824 10284 17876
rect 13728 17824 13780 17876
rect 9956 17799 10008 17808
rect 9956 17765 9965 17799
rect 9965 17765 9999 17799
rect 9999 17765 10008 17799
rect 11704 17799 11756 17808
rect 9956 17756 10008 17765
rect 11704 17765 11713 17799
rect 11713 17765 11747 17799
rect 11747 17765 11756 17799
rect 11704 17756 11756 17765
rect 15844 17756 15896 17808
rect 16856 17799 16908 17808
rect 16856 17765 16865 17799
rect 16865 17765 16899 17799
rect 16899 17765 16908 17799
rect 16856 17756 16908 17765
rect 16948 17799 17000 17808
rect 16948 17765 16957 17799
rect 16957 17765 16991 17799
rect 16991 17765 17000 17799
rect 16948 17756 17000 17765
rect 18788 17756 18840 17808
rect 19524 17824 19576 17876
rect 21732 17824 21784 17876
rect 19248 17756 19300 17808
rect 19708 17756 19760 17808
rect 4804 17688 4856 17740
rect 5540 17688 5592 17740
rect 6644 17688 6696 17740
rect 10324 17731 10376 17740
rect 10324 17697 10333 17731
rect 10333 17697 10367 17731
rect 10367 17697 10376 17731
rect 10324 17688 10376 17697
rect 13360 17688 13412 17740
rect 5448 17663 5500 17672
rect 5448 17629 5457 17663
rect 5457 17629 5491 17663
rect 5491 17629 5500 17663
rect 5448 17620 5500 17629
rect 10784 17620 10836 17672
rect 11888 17663 11940 17672
rect 112 17552 164 17604
rect 11888 17629 11897 17663
rect 11897 17629 11931 17663
rect 11931 17629 11940 17663
rect 11888 17620 11940 17629
rect 12256 17552 12308 17604
rect 6920 17484 6972 17536
rect 8484 17527 8536 17536
rect 8484 17493 8493 17527
rect 8493 17493 8527 17527
rect 8527 17493 8536 17527
rect 8484 17484 8536 17493
rect 12164 17484 12216 17536
rect 13912 17484 13964 17536
rect 15200 17688 15252 17740
rect 19800 17688 19852 17740
rect 21732 17688 21784 17740
rect 18328 17663 18380 17672
rect 18328 17629 18337 17663
rect 18337 17629 18371 17663
rect 18371 17629 18380 17663
rect 18328 17620 18380 17629
rect 19064 17620 19116 17672
rect 17684 17552 17736 17604
rect 18696 17552 18748 17604
rect 14188 17484 14240 17536
rect 14924 17484 14976 17536
rect 15752 17527 15804 17536
rect 15752 17493 15761 17527
rect 15761 17493 15795 17527
rect 15795 17493 15804 17527
rect 15752 17484 15804 17493
rect 4982 17382 5034 17434
rect 5046 17382 5098 17434
rect 5110 17382 5162 17434
rect 5174 17382 5226 17434
rect 12982 17382 13034 17434
rect 13046 17382 13098 17434
rect 13110 17382 13162 17434
rect 13174 17382 13226 17434
rect 20982 17382 21034 17434
rect 21046 17382 21098 17434
rect 21110 17382 21162 17434
rect 21174 17382 21226 17434
rect 3148 17212 3200 17264
rect 4804 17280 4856 17332
rect 10324 17323 10376 17332
rect 10324 17289 10333 17323
rect 10333 17289 10367 17323
rect 10367 17289 10376 17323
rect 10324 17280 10376 17289
rect 12256 17280 12308 17332
rect 14832 17323 14884 17332
rect 14832 17289 14841 17323
rect 14841 17289 14875 17323
rect 14875 17289 14884 17323
rect 14832 17280 14884 17289
rect 15200 17323 15252 17332
rect 15200 17289 15209 17323
rect 15209 17289 15243 17323
rect 15243 17289 15252 17323
rect 15200 17280 15252 17289
rect 16856 17280 16908 17332
rect 18788 17280 18840 17332
rect 21456 17323 21508 17332
rect 21456 17289 21465 17323
rect 21465 17289 21499 17323
rect 21499 17289 21508 17323
rect 21456 17280 21508 17289
rect 21732 17323 21784 17332
rect 21732 17289 21741 17323
rect 21741 17289 21775 17323
rect 21775 17289 21784 17323
rect 21732 17280 21784 17289
rect 6184 17212 6236 17264
rect 13268 17255 13320 17264
rect 2320 17187 2372 17196
rect 2320 17153 2329 17187
rect 2329 17153 2363 17187
rect 2363 17153 2372 17187
rect 2320 17144 2372 17153
rect 2504 17144 2556 17196
rect 4620 17187 4672 17196
rect 4620 17153 4629 17187
rect 4629 17153 4663 17187
rect 4663 17153 4672 17187
rect 4620 17144 4672 17153
rect 7196 17144 7248 17196
rect 13268 17221 13277 17255
rect 13277 17221 13311 17255
rect 13311 17221 13320 17255
rect 13268 17212 13320 17221
rect 10784 17187 10836 17196
rect 10784 17153 10793 17187
rect 10793 17153 10827 17187
rect 10827 17153 10836 17187
rect 10784 17144 10836 17153
rect 11888 17144 11940 17196
rect 8484 17076 8536 17128
rect 12164 17076 12216 17128
rect 19248 17255 19300 17264
rect 14188 17187 14240 17196
rect 14188 17153 14197 17187
rect 14197 17153 14231 17187
rect 14231 17153 14240 17187
rect 14188 17144 14240 17153
rect 15752 17144 15804 17196
rect 19248 17221 19257 17255
rect 19257 17221 19291 17255
rect 19291 17221 19300 17255
rect 19248 17212 19300 17221
rect 16948 17144 17000 17196
rect 18328 17187 18380 17196
rect 18328 17153 18337 17187
rect 18337 17153 18371 17187
rect 18371 17153 18380 17187
rect 18328 17144 18380 17153
rect 13912 17119 13964 17128
rect 13912 17085 13921 17119
rect 13921 17085 13955 17119
rect 13955 17085 13964 17119
rect 13912 17076 13964 17085
rect 21456 17076 21508 17128
rect 3976 17008 4028 17060
rect 3700 16940 3752 16992
rect 7012 17051 7064 17060
rect 7012 17017 7021 17051
rect 7021 17017 7055 17051
rect 7055 17017 7064 17051
rect 7564 17051 7616 17060
rect 7012 17008 7064 17017
rect 7564 17017 7573 17051
rect 7573 17017 7607 17051
rect 7607 17017 7616 17051
rect 7564 17008 7616 17017
rect 5540 16983 5592 16992
rect 5540 16949 5549 16983
rect 5549 16949 5583 16983
rect 5583 16949 5592 16983
rect 5540 16940 5592 16949
rect 6644 16983 6696 16992
rect 6644 16949 6653 16983
rect 6653 16949 6687 16983
rect 6687 16949 6696 16983
rect 6644 16940 6696 16949
rect 8484 16983 8536 16992
rect 8484 16949 8493 16983
rect 8493 16949 8527 16983
rect 8527 16949 8536 16983
rect 8484 16940 8536 16949
rect 8760 16940 8812 16992
rect 9864 16940 9916 16992
rect 13360 17008 13412 17060
rect 14832 17008 14884 17060
rect 16028 17008 16080 17060
rect 11704 16983 11756 16992
rect 11704 16949 11713 16983
rect 11713 16949 11747 16983
rect 11747 16949 11756 16983
rect 11704 16940 11756 16949
rect 12808 16940 12860 16992
rect 17868 16983 17920 16992
rect 17868 16949 17877 16983
rect 17877 16949 17911 16983
rect 17911 16949 17920 16983
rect 19064 17008 19116 17060
rect 17868 16940 17920 16949
rect 19340 16940 19392 16992
rect 8982 16838 9034 16890
rect 9046 16838 9098 16890
rect 9110 16838 9162 16890
rect 9174 16838 9226 16890
rect 16982 16838 17034 16890
rect 17046 16838 17098 16890
rect 17110 16838 17162 16890
rect 17174 16838 17226 16890
rect 8760 16779 8812 16788
rect 8760 16745 8769 16779
rect 8769 16745 8803 16779
rect 8803 16745 8812 16779
rect 8760 16736 8812 16745
rect 10232 16736 10284 16788
rect 3976 16668 4028 16720
rect 5632 16668 5684 16720
rect 7932 16668 7984 16720
rect 15752 16736 15804 16788
rect 17408 16736 17460 16788
rect 17868 16779 17920 16788
rect 17868 16745 17877 16779
rect 17877 16745 17911 16779
rect 17911 16745 17920 16779
rect 17868 16736 17920 16745
rect 21732 16736 21784 16788
rect 11888 16711 11940 16720
rect 11888 16677 11897 16711
rect 11897 16677 11931 16711
rect 11931 16677 11940 16711
rect 11888 16668 11940 16677
rect 18880 16711 18932 16720
rect 18880 16677 18889 16711
rect 18889 16677 18923 16711
rect 18923 16677 18932 16711
rect 18880 16668 18932 16677
rect 5448 16643 5500 16652
rect 5448 16609 5457 16643
rect 5457 16609 5491 16643
rect 5491 16609 5500 16643
rect 5448 16600 5500 16609
rect 8484 16532 8536 16584
rect 4436 16464 4488 16516
rect 10876 16600 10928 16652
rect 13544 16600 13596 16652
rect 13912 16600 13964 16652
rect 15292 16643 15344 16652
rect 15292 16609 15301 16643
rect 15301 16609 15335 16643
rect 15335 16609 15344 16643
rect 15292 16600 15344 16609
rect 15752 16643 15804 16652
rect 15752 16609 15761 16643
rect 15761 16609 15795 16643
rect 15795 16609 15804 16643
rect 15752 16600 15804 16609
rect 20904 16643 20956 16652
rect 20904 16609 20913 16643
rect 20913 16609 20947 16643
rect 20947 16609 20956 16643
rect 20904 16600 20956 16609
rect 21272 16600 21324 16652
rect 9772 16532 9824 16584
rect 11796 16575 11848 16584
rect 11796 16541 11805 16575
rect 11805 16541 11839 16575
rect 11839 16541 11848 16575
rect 11796 16532 11848 16541
rect 12164 16575 12216 16584
rect 12164 16541 12173 16575
rect 12173 16541 12207 16575
rect 12207 16541 12216 16575
rect 12164 16532 12216 16541
rect 14372 16575 14424 16584
rect 14372 16541 14381 16575
rect 14381 16541 14415 16575
rect 14415 16541 14424 16575
rect 14372 16532 14424 16541
rect 16948 16575 17000 16584
rect 16948 16541 16957 16575
rect 16957 16541 16991 16575
rect 16991 16541 17000 16575
rect 16948 16532 17000 16541
rect 17776 16532 17828 16584
rect 18788 16575 18840 16584
rect 18788 16541 18797 16575
rect 18797 16541 18831 16575
rect 18831 16541 18840 16575
rect 18788 16532 18840 16541
rect 19064 16575 19116 16584
rect 19064 16541 19073 16575
rect 19073 16541 19107 16575
rect 19107 16541 19116 16575
rect 19064 16532 19116 16541
rect 3148 16396 3200 16448
rect 6368 16439 6420 16448
rect 6368 16405 6377 16439
rect 6377 16405 6411 16439
rect 6411 16405 6420 16439
rect 6368 16396 6420 16405
rect 7012 16396 7064 16448
rect 13452 16439 13504 16448
rect 13452 16405 13461 16439
rect 13461 16405 13495 16439
rect 13495 16405 13504 16439
rect 13452 16396 13504 16405
rect 13912 16396 13964 16448
rect 4982 16294 5034 16346
rect 5046 16294 5098 16346
rect 5110 16294 5162 16346
rect 5174 16294 5226 16346
rect 12982 16294 13034 16346
rect 13046 16294 13098 16346
rect 13110 16294 13162 16346
rect 13174 16294 13226 16346
rect 20982 16294 21034 16346
rect 21046 16294 21098 16346
rect 21110 16294 21162 16346
rect 21174 16294 21226 16346
rect 5448 16192 5500 16244
rect 7932 16235 7984 16244
rect 7932 16201 7941 16235
rect 7941 16201 7975 16235
rect 7975 16201 7984 16235
rect 7932 16192 7984 16201
rect 8484 16192 8536 16244
rect 10232 16192 10284 16244
rect 11888 16235 11940 16244
rect 11888 16201 11897 16235
rect 11897 16201 11931 16235
rect 11931 16201 11940 16235
rect 11888 16192 11940 16201
rect 13452 16192 13504 16244
rect 15292 16235 15344 16244
rect 15292 16201 15301 16235
rect 15301 16201 15335 16235
rect 15335 16201 15344 16235
rect 15292 16192 15344 16201
rect 16028 16235 16080 16244
rect 16028 16201 16037 16235
rect 16037 16201 16071 16235
rect 16071 16201 16080 16235
rect 16028 16192 16080 16201
rect 18880 16192 18932 16244
rect 21272 16192 21324 16244
rect 112 16124 164 16176
rect 1584 15988 1636 16040
rect 4344 16124 4396 16176
rect 4436 16056 4488 16108
rect 3148 15988 3200 16040
rect 4252 15988 4304 16040
rect 4160 15920 4212 15972
rect 5632 16056 5684 16108
rect 6920 16099 6972 16108
rect 6920 16065 6929 16099
rect 6929 16065 6963 16099
rect 6963 16065 6972 16099
rect 6920 16056 6972 16065
rect 7196 16099 7248 16108
rect 7196 16065 7205 16099
rect 7205 16065 7239 16099
rect 7239 16065 7248 16099
rect 7196 16056 7248 16065
rect 11244 16056 11296 16108
rect 11796 16124 11848 16176
rect 14372 16124 14424 16176
rect 9496 16031 9548 16040
rect 9496 15997 9505 16031
rect 9505 15997 9539 16031
rect 9539 15997 9548 16031
rect 9496 15988 9548 15997
rect 12808 15988 12860 16040
rect 9772 15963 9824 15972
rect 4988 15895 5040 15904
rect 4988 15861 4997 15895
rect 4997 15861 5031 15895
rect 5031 15861 5040 15895
rect 4988 15852 5040 15861
rect 6368 15852 6420 15904
rect 9772 15929 9781 15963
rect 9781 15929 9815 15963
rect 9815 15929 9824 15963
rect 9772 15920 9824 15929
rect 10600 15920 10652 15972
rect 13452 15920 13504 15972
rect 16948 16056 17000 16108
rect 19064 16124 19116 16176
rect 19984 16056 20036 16108
rect 14648 16031 14700 16040
rect 14648 15997 14657 16031
rect 14657 15997 14691 16031
rect 14691 15997 14700 16031
rect 14648 15988 14700 15997
rect 15752 15988 15804 16040
rect 16212 16031 16264 16040
rect 16212 15997 16221 16031
rect 16221 15997 16255 16031
rect 16255 15997 16264 16031
rect 16212 15988 16264 15997
rect 16028 15920 16080 15972
rect 17408 15963 17460 15972
rect 17408 15929 17417 15963
rect 17417 15929 17451 15963
rect 17451 15929 17460 15963
rect 17408 15920 17460 15929
rect 13544 15852 13596 15904
rect 14004 15895 14056 15904
rect 14004 15861 14013 15895
rect 14013 15861 14047 15895
rect 14047 15861 14056 15895
rect 14004 15852 14056 15861
rect 8982 15750 9034 15802
rect 9046 15750 9098 15802
rect 9110 15750 9162 15802
rect 9174 15750 9226 15802
rect 16982 15750 17034 15802
rect 17046 15750 17098 15802
rect 17110 15750 17162 15802
rect 17174 15750 17226 15802
rect 4252 15691 4304 15700
rect 4252 15657 4261 15691
rect 4261 15657 4295 15691
rect 4295 15657 4304 15691
rect 4252 15648 4304 15657
rect 8392 15691 8444 15700
rect 8392 15657 8401 15691
rect 8401 15657 8435 15691
rect 8435 15657 8444 15691
rect 8392 15648 8444 15657
rect 8852 15648 8904 15700
rect 9496 15648 9548 15700
rect 9772 15648 9824 15700
rect 11244 15648 11296 15700
rect 16580 15691 16632 15700
rect 16580 15657 16589 15691
rect 16589 15657 16623 15691
rect 16623 15657 16632 15691
rect 16580 15648 16632 15657
rect 17776 15691 17828 15700
rect 17776 15657 17785 15691
rect 17785 15657 17819 15691
rect 17819 15657 17828 15691
rect 17776 15648 17828 15657
rect 18788 15691 18840 15700
rect 18788 15657 18797 15691
rect 18797 15657 18831 15691
rect 18831 15657 18840 15691
rect 18788 15648 18840 15657
rect 19984 15648 20036 15700
rect 2596 15623 2648 15632
rect 2596 15589 2605 15623
rect 2605 15589 2639 15623
rect 2639 15589 2648 15623
rect 2596 15580 2648 15589
rect 4068 15580 4120 15632
rect 4988 15580 5040 15632
rect 6552 15623 6604 15632
rect 6552 15589 6561 15623
rect 6561 15589 6595 15623
rect 6595 15589 6604 15623
rect 6552 15580 6604 15589
rect 11612 15623 11664 15632
rect 9680 15555 9732 15564
rect 1584 15444 1636 15496
rect 9680 15521 9689 15555
rect 9689 15521 9723 15555
rect 9723 15521 9732 15555
rect 9680 15512 9732 15521
rect 11612 15589 11621 15623
rect 11621 15589 11655 15623
rect 11655 15589 11664 15623
rect 11612 15580 11664 15589
rect 16212 15623 16264 15632
rect 16212 15589 16221 15623
rect 16221 15589 16255 15623
rect 16255 15589 16264 15623
rect 16212 15580 16264 15589
rect 16856 15580 16908 15632
rect 13636 15555 13688 15564
rect 13636 15521 13645 15555
rect 13645 15521 13679 15555
rect 13679 15521 13688 15555
rect 13636 15512 13688 15521
rect 14188 15555 14240 15564
rect 14188 15521 14197 15555
rect 14197 15521 14231 15555
rect 14231 15521 14240 15555
rect 14648 15555 14700 15564
rect 14188 15512 14240 15521
rect 14648 15521 14657 15555
rect 14657 15521 14691 15555
rect 14691 15521 14700 15555
rect 14648 15512 14700 15521
rect 15752 15512 15804 15564
rect 18328 15555 18380 15564
rect 18328 15521 18337 15555
rect 18337 15521 18371 15555
rect 18371 15521 18380 15555
rect 18328 15512 18380 15521
rect 19064 15512 19116 15564
rect 2504 15487 2556 15496
rect 2504 15453 2513 15487
rect 2513 15453 2547 15487
rect 2547 15453 2556 15487
rect 2504 15444 2556 15453
rect 4620 15487 4672 15496
rect 4620 15453 4629 15487
rect 4629 15453 4663 15487
rect 4663 15453 4672 15487
rect 4620 15444 4672 15453
rect 6460 15487 6512 15496
rect 4804 15376 4856 15428
rect 6460 15453 6469 15487
rect 6469 15453 6503 15487
rect 6503 15453 6512 15487
rect 6460 15444 6512 15453
rect 10416 15487 10468 15496
rect 10416 15453 10425 15487
rect 10425 15453 10459 15487
rect 10459 15453 10468 15487
rect 10416 15444 10468 15453
rect 11152 15444 11204 15496
rect 11796 15444 11848 15496
rect 12164 15487 12216 15496
rect 12164 15453 12173 15487
rect 12173 15453 12207 15487
rect 12207 15453 12216 15487
rect 12164 15444 12216 15453
rect 1860 15351 1912 15360
rect 1860 15317 1869 15351
rect 1869 15317 1903 15351
rect 1903 15317 1912 15351
rect 1860 15308 1912 15317
rect 4620 15308 4672 15360
rect 7196 15376 7248 15428
rect 12532 15351 12584 15360
rect 12532 15317 12541 15351
rect 12541 15317 12575 15351
rect 12575 15317 12584 15351
rect 12532 15308 12584 15317
rect 16488 15308 16540 15360
rect 17316 15487 17368 15496
rect 17316 15453 17325 15487
rect 17325 15453 17359 15487
rect 17359 15453 17368 15487
rect 17316 15444 17368 15453
rect 16856 15308 16908 15360
rect 19800 15308 19852 15360
rect 4982 15206 5034 15258
rect 5046 15206 5098 15258
rect 5110 15206 5162 15258
rect 5174 15206 5226 15258
rect 12982 15206 13034 15258
rect 13046 15206 13098 15258
rect 13110 15206 13162 15258
rect 13174 15206 13226 15258
rect 20982 15206 21034 15258
rect 21046 15206 21098 15258
rect 21110 15206 21162 15258
rect 21174 15206 21226 15258
rect 2596 15104 2648 15156
rect 4068 15147 4120 15156
rect 4068 15113 4077 15147
rect 4077 15113 4111 15147
rect 4111 15113 4120 15147
rect 4068 15104 4120 15113
rect 6460 15147 6512 15156
rect 2504 15036 2556 15088
rect 1860 14968 1912 15020
rect 5356 15036 5408 15088
rect 6460 15113 6469 15147
rect 6469 15113 6503 15147
rect 6503 15113 6512 15147
rect 6460 15104 6512 15113
rect 10232 15104 10284 15156
rect 11612 15104 11664 15156
rect 11796 15147 11848 15156
rect 11796 15113 11805 15147
rect 11805 15113 11839 15147
rect 11839 15113 11848 15147
rect 11796 15104 11848 15113
rect 14188 15104 14240 15156
rect 15752 15147 15804 15156
rect 15752 15113 15761 15147
rect 15761 15113 15795 15147
rect 15795 15113 15804 15147
rect 15752 15104 15804 15113
rect 18328 15147 18380 15156
rect 18328 15113 18337 15147
rect 18337 15113 18371 15147
rect 18371 15113 18380 15147
rect 18328 15104 18380 15113
rect 19064 15104 19116 15156
rect 21456 15147 21508 15156
rect 21456 15113 21465 15147
rect 21465 15113 21499 15147
rect 21499 15113 21508 15147
rect 21456 15104 21508 15113
rect 7564 15036 7616 15088
rect 4804 14968 4856 15020
rect 7196 14968 7248 15020
rect 12164 14968 12216 15020
rect 8852 14943 8904 14952
rect 1768 14832 1820 14884
rect 6552 14832 6604 14884
rect 7012 14875 7064 14884
rect 7012 14841 7021 14875
rect 7021 14841 7055 14875
rect 7055 14841 7064 14875
rect 7012 14832 7064 14841
rect 8208 14875 8260 14884
rect 8208 14841 8217 14875
rect 8217 14841 8251 14875
rect 8251 14841 8260 14875
rect 8852 14909 8861 14943
rect 8861 14909 8895 14943
rect 8895 14909 8904 14943
rect 8852 14900 8904 14909
rect 9956 14943 10008 14952
rect 9956 14909 9965 14943
rect 9965 14909 9999 14943
rect 9999 14909 10008 14943
rect 9956 14900 10008 14909
rect 14372 14968 14424 15020
rect 15292 14968 15344 15020
rect 14464 14943 14516 14952
rect 14464 14909 14473 14943
rect 14473 14909 14507 14943
rect 14507 14909 14516 14943
rect 14464 14900 14516 14909
rect 12532 14875 12584 14884
rect 8208 14832 8260 14841
rect 12532 14841 12541 14875
rect 12541 14841 12575 14875
rect 12575 14841 12584 14875
rect 12532 14832 12584 14841
rect 14740 14875 14792 14884
rect 4988 14764 5040 14816
rect 5356 14764 5408 14816
rect 6828 14764 6880 14816
rect 7748 14764 7800 14816
rect 9680 14764 9732 14816
rect 10232 14764 10284 14816
rect 12164 14807 12216 14816
rect 12164 14773 12173 14807
rect 12173 14773 12207 14807
rect 12207 14773 12216 14807
rect 14740 14841 14749 14875
rect 14749 14841 14783 14875
rect 14783 14841 14792 14875
rect 14740 14832 14792 14841
rect 16580 15036 16632 15088
rect 16396 14968 16448 15020
rect 21456 14900 21508 14952
rect 13636 14807 13688 14816
rect 12164 14764 12216 14773
rect 13636 14773 13645 14807
rect 13645 14773 13679 14807
rect 13679 14773 13688 14807
rect 13636 14764 13688 14773
rect 16212 14807 16264 14816
rect 16212 14773 16221 14807
rect 16221 14773 16255 14807
rect 16255 14773 16264 14807
rect 16212 14764 16264 14773
rect 16764 14764 16816 14816
rect 18236 14764 18288 14816
rect 19064 14807 19116 14816
rect 19064 14773 19073 14807
rect 19073 14773 19107 14807
rect 19107 14773 19116 14807
rect 19064 14764 19116 14773
rect 20720 14764 20772 14816
rect 8982 14662 9034 14714
rect 9046 14662 9098 14714
rect 9110 14662 9162 14714
rect 9174 14662 9226 14714
rect 16982 14662 17034 14714
rect 17046 14662 17098 14714
rect 17110 14662 17162 14714
rect 17174 14662 17226 14714
rect 1860 14560 1912 14612
rect 4988 14603 5040 14612
rect 4988 14569 4997 14603
rect 4997 14569 5031 14603
rect 5031 14569 5040 14603
rect 4988 14560 5040 14569
rect 8024 14603 8076 14612
rect 8024 14569 8033 14603
rect 8033 14569 8067 14603
rect 8067 14569 8076 14603
rect 8024 14560 8076 14569
rect 8852 14560 8904 14612
rect 9956 14560 10008 14612
rect 12164 14560 12216 14612
rect 14372 14603 14424 14612
rect 14372 14569 14381 14603
rect 14381 14569 14415 14603
rect 14415 14569 14424 14603
rect 14372 14560 14424 14569
rect 15016 14560 15068 14612
rect 16212 14603 16264 14612
rect 16212 14569 16221 14603
rect 16221 14569 16255 14603
rect 16255 14569 16264 14603
rect 16212 14560 16264 14569
rect 16856 14603 16908 14612
rect 16856 14569 16865 14603
rect 16865 14569 16899 14603
rect 16899 14569 16908 14603
rect 16856 14560 16908 14569
rect 18236 14560 18288 14612
rect 3792 14492 3844 14544
rect 4160 14492 4212 14544
rect 4620 14492 4672 14544
rect 6368 14492 6420 14544
rect 1952 14467 2004 14476
rect 1952 14433 1961 14467
rect 1961 14433 1995 14467
rect 1995 14433 2004 14467
rect 1952 14424 2004 14433
rect 3516 14424 3568 14476
rect 7840 14424 7892 14476
rect 8116 14424 8168 14476
rect 8300 14467 8352 14476
rect 8300 14433 8309 14467
rect 8309 14433 8343 14467
rect 8343 14433 8352 14467
rect 10324 14492 10376 14544
rect 19064 14492 19116 14544
rect 19616 14492 19668 14544
rect 8300 14424 8352 14433
rect 10416 14424 10468 14476
rect 13268 14424 13320 14476
rect 4068 14399 4120 14408
rect 4068 14365 4077 14399
rect 4077 14365 4111 14399
rect 4111 14365 4120 14399
rect 4068 14356 4120 14365
rect 6828 14399 6880 14408
rect 6828 14365 6837 14399
rect 6837 14365 6871 14399
rect 6871 14365 6880 14399
rect 6828 14356 6880 14365
rect 10876 14356 10928 14408
rect 9680 14288 9732 14340
rect 13636 14288 13688 14340
rect 14740 14424 14792 14476
rect 15660 14424 15712 14476
rect 14096 14399 14148 14408
rect 14096 14365 14105 14399
rect 14105 14365 14139 14399
rect 14139 14365 14148 14399
rect 14096 14356 14148 14365
rect 16488 14356 16540 14408
rect 17592 14356 17644 14408
rect 18880 14356 18932 14408
rect 14464 14288 14516 14340
rect 16304 14288 16356 14340
rect 19248 14288 19300 14340
rect 2688 14263 2740 14272
rect 2688 14229 2697 14263
rect 2697 14229 2731 14263
rect 2731 14229 2740 14263
rect 2688 14220 2740 14229
rect 3884 14263 3936 14272
rect 3884 14229 3893 14263
rect 3893 14229 3927 14263
rect 3927 14229 3936 14263
rect 3884 14220 3936 14229
rect 5908 14263 5960 14272
rect 5908 14229 5917 14263
rect 5917 14229 5951 14263
rect 5951 14229 5960 14263
rect 5908 14220 5960 14229
rect 7012 14220 7064 14272
rect 12532 14263 12584 14272
rect 12532 14229 12541 14263
rect 12541 14229 12575 14263
rect 12575 14229 12584 14263
rect 12532 14220 12584 14229
rect 14740 14263 14792 14272
rect 14740 14229 14749 14263
rect 14749 14229 14783 14263
rect 14783 14229 14792 14263
rect 14740 14220 14792 14229
rect 4982 14118 5034 14170
rect 5046 14118 5098 14170
rect 5110 14118 5162 14170
rect 5174 14118 5226 14170
rect 12982 14118 13034 14170
rect 13046 14118 13098 14170
rect 13110 14118 13162 14170
rect 13174 14118 13226 14170
rect 20982 14118 21034 14170
rect 21046 14118 21098 14170
rect 21110 14118 21162 14170
rect 21174 14118 21226 14170
rect 1768 14059 1820 14068
rect 1768 14025 1777 14059
rect 1777 14025 1811 14059
rect 1811 14025 1820 14059
rect 1768 14016 1820 14025
rect 2136 14016 2188 14068
rect 3792 14059 3844 14068
rect 3792 14025 3801 14059
rect 3801 14025 3835 14059
rect 3835 14025 3844 14059
rect 3792 14016 3844 14025
rect 4068 14016 4120 14068
rect 6368 14059 6420 14068
rect 6368 14025 6377 14059
rect 6377 14025 6411 14059
rect 6411 14025 6420 14059
rect 6368 14016 6420 14025
rect 10232 14059 10284 14068
rect 10232 14025 10241 14059
rect 10241 14025 10275 14059
rect 10275 14025 10284 14059
rect 10232 14016 10284 14025
rect 10600 14016 10652 14068
rect 12624 14016 12676 14068
rect 15660 14059 15712 14068
rect 15660 14025 15669 14059
rect 15669 14025 15703 14059
rect 15703 14025 15712 14059
rect 15660 14016 15712 14025
rect 16212 14059 16264 14068
rect 16212 14025 16221 14059
rect 16221 14025 16255 14059
rect 16255 14025 16264 14059
rect 16212 14016 16264 14025
rect 16580 14016 16632 14068
rect 17592 14016 17644 14068
rect 19064 14016 19116 14068
rect 2228 13880 2280 13932
rect 2688 13880 2740 13932
rect 3884 13880 3936 13932
rect 9864 13991 9916 14000
rect 5356 13880 5408 13932
rect 8024 13923 8076 13932
rect 2136 13787 2188 13796
rect 2136 13753 2145 13787
rect 2145 13753 2179 13787
rect 2179 13753 2188 13787
rect 2136 13744 2188 13753
rect 3700 13744 3752 13796
rect 1952 13676 2004 13728
rect 3148 13719 3200 13728
rect 3148 13685 3157 13719
rect 3157 13685 3191 13719
rect 3191 13685 3200 13719
rect 3148 13676 3200 13685
rect 3516 13719 3568 13728
rect 3516 13685 3525 13719
rect 3525 13685 3559 13719
rect 3559 13685 3568 13719
rect 3516 13676 3568 13685
rect 3884 13676 3936 13728
rect 8024 13889 8033 13923
rect 8033 13889 8067 13923
rect 8067 13889 8076 13923
rect 8024 13880 8076 13889
rect 6460 13812 6512 13864
rect 9864 13957 9873 13991
rect 9873 13957 9907 13991
rect 9907 13957 9916 13991
rect 9864 13948 9916 13957
rect 11520 13948 11572 14000
rect 12440 13948 12492 14000
rect 13268 13948 13320 14000
rect 16764 13948 16816 14000
rect 10508 13923 10560 13932
rect 10508 13889 10517 13923
rect 10517 13889 10551 13923
rect 10551 13889 10560 13923
rect 10508 13880 10560 13889
rect 11796 13880 11848 13932
rect 14096 13923 14148 13932
rect 14096 13889 14105 13923
rect 14105 13889 14139 13923
rect 14139 13889 14148 13923
rect 14096 13880 14148 13889
rect 17316 13880 17368 13932
rect 9404 13744 9456 13796
rect 12532 13787 12584 13796
rect 12532 13753 12541 13787
rect 12541 13753 12575 13787
rect 12575 13753 12584 13787
rect 12532 13744 12584 13753
rect 12624 13787 12676 13796
rect 12624 13753 12633 13787
rect 12633 13753 12667 13787
rect 12667 13753 12676 13787
rect 12624 13744 12676 13753
rect 6092 13676 6144 13728
rect 6736 13676 6788 13728
rect 8392 13719 8444 13728
rect 8392 13685 8401 13719
rect 8401 13685 8435 13719
rect 8435 13685 8444 13719
rect 8392 13676 8444 13685
rect 10232 13676 10284 13728
rect 16488 13787 16540 13796
rect 16488 13753 16497 13787
rect 16497 13753 16531 13787
rect 16531 13753 16540 13787
rect 16488 13744 16540 13753
rect 16580 13787 16632 13796
rect 16580 13753 16589 13787
rect 16589 13753 16623 13787
rect 16623 13753 16632 13787
rect 16580 13744 16632 13753
rect 15016 13676 15068 13728
rect 15292 13719 15344 13728
rect 15292 13685 15301 13719
rect 15301 13685 15335 13719
rect 15335 13685 15344 13719
rect 15292 13676 15344 13685
rect 15384 13676 15436 13728
rect 18788 13812 18840 13864
rect 19432 13787 19484 13796
rect 19432 13753 19441 13787
rect 19441 13753 19475 13787
rect 19475 13753 19484 13787
rect 19432 13744 19484 13753
rect 20076 13787 20128 13796
rect 19340 13676 19392 13728
rect 20076 13753 20085 13787
rect 20085 13753 20119 13787
rect 20119 13753 20128 13787
rect 20076 13744 20128 13753
rect 20536 13744 20588 13796
rect 20812 13744 20864 13796
rect 21732 13744 21784 13796
rect 19616 13676 19668 13728
rect 20444 13676 20496 13728
rect 8982 13574 9034 13626
rect 9046 13574 9098 13626
rect 9110 13574 9162 13626
rect 9174 13574 9226 13626
rect 16982 13574 17034 13626
rect 17046 13574 17098 13626
rect 17110 13574 17162 13626
rect 17174 13574 17226 13626
rect 4068 13472 4120 13524
rect 7012 13472 7064 13524
rect 7840 13515 7892 13524
rect 7840 13481 7849 13515
rect 7849 13481 7883 13515
rect 7883 13481 7892 13515
rect 7840 13472 7892 13481
rect 8208 13472 8260 13524
rect 10600 13515 10652 13524
rect 2228 13447 2280 13456
rect 2228 13413 2237 13447
rect 2237 13413 2271 13447
rect 2271 13413 2280 13447
rect 2228 13404 2280 13413
rect 6552 13404 6604 13456
rect 8392 13404 8444 13456
rect 10048 13404 10100 13456
rect 10600 13481 10609 13515
rect 10609 13481 10643 13515
rect 10643 13481 10652 13515
rect 10600 13472 10652 13481
rect 10876 13515 10928 13524
rect 10876 13481 10885 13515
rect 10885 13481 10919 13515
rect 10919 13481 10928 13515
rect 10876 13472 10928 13481
rect 11888 13472 11940 13524
rect 13544 13472 13596 13524
rect 14096 13515 14148 13524
rect 14096 13481 14105 13515
rect 14105 13481 14139 13515
rect 14139 13481 14148 13515
rect 14096 13472 14148 13481
rect 17408 13472 17460 13524
rect 18144 13472 18196 13524
rect 19616 13515 19668 13524
rect 11796 13404 11848 13456
rect 12440 13404 12492 13456
rect 16856 13447 16908 13456
rect 16856 13413 16865 13447
rect 16865 13413 16899 13447
rect 16899 13413 16908 13447
rect 16856 13404 16908 13413
rect 19064 13404 19116 13456
rect 19616 13481 19625 13515
rect 19625 13481 19659 13515
rect 19659 13481 19668 13515
rect 19616 13472 19668 13481
rect 20076 13472 20128 13524
rect 20812 13404 20864 13456
rect 1860 13336 1912 13388
rect 2504 13336 2556 13388
rect 4160 13379 4212 13388
rect 4160 13345 4169 13379
rect 4169 13345 4203 13379
rect 4203 13345 4212 13379
rect 4620 13379 4672 13388
rect 4160 13336 4212 13345
rect 4620 13345 4629 13379
rect 4629 13345 4663 13379
rect 4663 13345 4672 13379
rect 4620 13336 4672 13345
rect 8484 13336 8536 13388
rect 10508 13336 10560 13388
rect 15568 13336 15620 13388
rect 9680 13311 9732 13320
rect 2320 13200 2372 13252
rect 1860 13132 1912 13184
rect 3792 13175 3844 13184
rect 3792 13141 3801 13175
rect 3801 13141 3835 13175
rect 3835 13141 3844 13175
rect 3792 13132 3844 13141
rect 5724 13175 5776 13184
rect 5724 13141 5733 13175
rect 5733 13141 5767 13175
rect 5767 13141 5776 13175
rect 9680 13277 9689 13311
rect 9689 13277 9723 13311
rect 9723 13277 9732 13311
rect 9680 13268 9732 13277
rect 11612 13311 11664 13320
rect 11612 13277 11621 13311
rect 11621 13277 11655 13311
rect 11655 13277 11664 13311
rect 11612 13268 11664 13277
rect 16948 13268 17000 13320
rect 17408 13311 17460 13320
rect 17408 13277 17417 13311
rect 17417 13277 17451 13311
rect 17451 13277 17460 13311
rect 17408 13268 17460 13277
rect 18420 13268 18472 13320
rect 18788 13268 18840 13320
rect 21456 13200 21508 13252
rect 5724 13132 5776 13141
rect 8300 13132 8352 13184
rect 9404 13132 9456 13184
rect 14096 13132 14148 13184
rect 14740 13132 14792 13184
rect 16488 13175 16540 13184
rect 16488 13141 16497 13175
rect 16497 13141 16531 13175
rect 16531 13141 16540 13175
rect 16488 13132 16540 13141
rect 17592 13132 17644 13184
rect 19432 13132 19484 13184
rect 20076 13132 20128 13184
rect 4982 13030 5034 13082
rect 5046 13030 5098 13082
rect 5110 13030 5162 13082
rect 5174 13030 5226 13082
rect 12982 13030 13034 13082
rect 13046 13030 13098 13082
rect 13110 13030 13162 13082
rect 13174 13030 13226 13082
rect 20982 13030 21034 13082
rect 21046 13030 21098 13082
rect 21110 13030 21162 13082
rect 21174 13030 21226 13082
rect 3148 12971 3200 12980
rect 3148 12937 3157 12971
rect 3157 12937 3191 12971
rect 3191 12937 3200 12971
rect 3148 12928 3200 12937
rect 4160 12928 4212 12980
rect 5908 12928 5960 12980
rect 20 12860 72 12912
rect 1860 12860 1912 12912
rect 4896 12860 4948 12912
rect 5632 12860 5684 12912
rect 6552 12903 6604 12912
rect 6552 12869 6561 12903
rect 6561 12869 6595 12903
rect 6595 12869 6604 12903
rect 6552 12860 6604 12869
rect 6828 12860 6880 12912
rect 4528 12835 4580 12844
rect 4528 12801 4537 12835
rect 4537 12801 4571 12835
rect 4571 12801 4580 12835
rect 4528 12792 4580 12801
rect 5356 12792 5408 12844
rect 6736 12792 6788 12844
rect 1676 12767 1728 12776
rect 1676 12733 1685 12767
rect 1685 12733 1719 12767
rect 1719 12733 1728 12767
rect 1676 12724 1728 12733
rect 2320 12724 2372 12776
rect 3792 12767 3844 12776
rect 3792 12733 3801 12767
rect 3801 12733 3835 12767
rect 3835 12733 3844 12767
rect 3792 12724 3844 12733
rect 3976 12724 4028 12776
rect 8484 12928 8536 12980
rect 8760 12928 8812 12980
rect 10600 12971 10652 12980
rect 10600 12937 10609 12971
rect 10609 12937 10643 12971
rect 10643 12937 10652 12971
rect 10600 12928 10652 12937
rect 11612 12928 11664 12980
rect 13544 12928 13596 12980
rect 16856 12928 16908 12980
rect 16948 12928 17000 12980
rect 18880 12928 18932 12980
rect 11796 12903 11848 12912
rect 11796 12869 11805 12903
rect 11805 12869 11839 12903
rect 11839 12869 11848 12903
rect 11796 12860 11848 12869
rect 18236 12860 18288 12912
rect 9680 12792 9732 12844
rect 11520 12835 11572 12844
rect 11520 12801 11529 12835
rect 11529 12801 11563 12835
rect 11563 12801 11572 12835
rect 11520 12792 11572 12801
rect 18144 12835 18196 12844
rect 18144 12801 18153 12835
rect 18153 12801 18187 12835
rect 18187 12801 18196 12835
rect 18144 12792 18196 12801
rect 18420 12835 18472 12844
rect 18420 12801 18429 12835
rect 18429 12801 18463 12835
rect 18463 12801 18472 12835
rect 18420 12792 18472 12801
rect 3516 12656 3568 12708
rect 4620 12656 4672 12708
rect 2688 12631 2740 12640
rect 2688 12597 2697 12631
rect 2697 12597 2731 12631
rect 2731 12597 2740 12631
rect 2688 12588 2740 12597
rect 3700 12631 3752 12640
rect 3700 12597 3709 12631
rect 3709 12597 3743 12631
rect 3743 12597 3752 12631
rect 3700 12588 3752 12597
rect 4068 12588 4120 12640
rect 4896 12631 4948 12640
rect 4896 12597 4905 12631
rect 4905 12597 4939 12631
rect 4939 12597 4948 12631
rect 4896 12588 4948 12597
rect 9404 12767 9456 12776
rect 7012 12699 7064 12708
rect 7012 12665 7021 12699
rect 7021 12665 7055 12699
rect 7055 12665 7064 12699
rect 9404 12733 9413 12767
rect 9413 12733 9447 12767
rect 9447 12733 9456 12767
rect 9404 12724 9456 12733
rect 13360 12724 13412 12776
rect 13544 12767 13596 12776
rect 13544 12733 13553 12767
rect 13553 12733 13587 12767
rect 13587 12733 13596 12767
rect 13544 12724 13596 12733
rect 14096 12767 14148 12776
rect 14096 12733 14105 12767
rect 14105 12733 14139 12767
rect 14139 12733 14148 12767
rect 14096 12724 14148 12733
rect 17408 12724 17460 12776
rect 19064 12724 19116 12776
rect 20812 12928 20864 12980
rect 21456 12928 21508 12980
rect 20260 12903 20312 12912
rect 20260 12869 20269 12903
rect 20269 12869 20303 12903
rect 20303 12869 20312 12903
rect 20260 12860 20312 12869
rect 21364 12903 21416 12912
rect 21364 12869 21373 12903
rect 21373 12869 21407 12903
rect 21407 12869 21416 12903
rect 21364 12860 21416 12869
rect 20444 12792 20496 12844
rect 7012 12656 7064 12665
rect 10508 12656 10560 12708
rect 10876 12699 10928 12708
rect 10876 12665 10885 12699
rect 10885 12665 10919 12699
rect 10919 12665 10928 12699
rect 10876 12656 10928 12665
rect 5816 12588 5868 12640
rect 6000 12588 6052 12640
rect 10232 12588 10284 12640
rect 10416 12588 10468 12640
rect 10600 12588 10652 12640
rect 15292 12656 15344 12708
rect 16028 12656 16080 12708
rect 18236 12699 18288 12708
rect 18236 12665 18245 12699
rect 18245 12665 18279 12699
rect 18279 12665 18288 12699
rect 20812 12724 20864 12776
rect 18236 12656 18288 12665
rect 15568 12588 15620 12640
rect 16764 12588 16816 12640
rect 8982 12486 9034 12538
rect 9046 12486 9098 12538
rect 9110 12486 9162 12538
rect 9174 12486 9226 12538
rect 16982 12486 17034 12538
rect 17046 12486 17098 12538
rect 17110 12486 17162 12538
rect 17174 12486 17226 12538
rect 1860 12384 1912 12436
rect 3976 12384 4028 12436
rect 4160 12384 4212 12436
rect 5724 12427 5776 12436
rect 5724 12393 5733 12427
rect 5733 12393 5767 12427
rect 5767 12393 5776 12427
rect 5724 12384 5776 12393
rect 1676 12316 1728 12368
rect 2688 12316 2740 12368
rect 1860 12291 1912 12300
rect 1860 12257 1869 12291
rect 1869 12257 1903 12291
rect 1903 12257 1912 12291
rect 2044 12291 2096 12300
rect 1860 12248 1912 12257
rect 2044 12257 2053 12291
rect 2053 12257 2087 12291
rect 2087 12257 2096 12291
rect 2044 12248 2096 12257
rect 2504 12291 2556 12300
rect 2504 12257 2513 12291
rect 2513 12257 2547 12291
rect 2547 12257 2556 12291
rect 5632 12316 5684 12368
rect 4160 12291 4212 12300
rect 2504 12248 2556 12257
rect 4160 12257 4169 12291
rect 4169 12257 4203 12291
rect 4203 12257 4212 12291
rect 4160 12248 4212 12257
rect 4896 12248 4948 12300
rect 5724 12248 5776 12300
rect 10876 12427 10928 12436
rect 10876 12393 10885 12427
rect 10885 12393 10919 12427
rect 10919 12393 10928 12427
rect 10876 12384 10928 12393
rect 16856 12384 16908 12436
rect 17408 12384 17460 12436
rect 18788 12427 18840 12436
rect 18788 12393 18797 12427
rect 18797 12393 18831 12427
rect 18831 12393 18840 12427
rect 18788 12384 18840 12393
rect 20444 12384 20496 12436
rect 12440 12316 12492 12368
rect 12808 12316 12860 12368
rect 16028 12316 16080 12368
rect 18144 12316 18196 12368
rect 20720 12316 20772 12368
rect 21272 12316 21324 12368
rect 6184 12291 6236 12300
rect 6184 12257 6193 12291
rect 6193 12257 6227 12291
rect 6227 12257 6236 12291
rect 6184 12248 6236 12257
rect 7288 12248 7340 12300
rect 7840 12248 7892 12300
rect 8024 12248 8076 12300
rect 10600 12248 10652 12300
rect 11888 12291 11940 12300
rect 11888 12257 11897 12291
rect 11897 12257 11931 12291
rect 11931 12257 11940 12291
rect 11888 12248 11940 12257
rect 12072 12291 12124 12300
rect 12072 12257 12081 12291
rect 12081 12257 12115 12291
rect 12115 12257 12124 12291
rect 12072 12248 12124 12257
rect 13636 12291 13688 12300
rect 13636 12257 13645 12291
rect 13645 12257 13679 12291
rect 13679 12257 13688 12291
rect 13636 12248 13688 12257
rect 14096 12248 14148 12300
rect 14464 12248 14516 12300
rect 19064 12248 19116 12300
rect 19340 12248 19392 12300
rect 19708 12291 19760 12300
rect 19708 12257 19717 12291
rect 19717 12257 19751 12291
rect 19751 12257 19760 12291
rect 19708 12248 19760 12257
rect 3976 12180 4028 12232
rect 12164 12223 12216 12232
rect 12164 12189 12173 12223
rect 12173 12189 12207 12223
rect 12207 12189 12216 12223
rect 12164 12180 12216 12189
rect 12808 12180 12860 12232
rect 15752 12180 15804 12232
rect 16948 12180 17000 12232
rect 21640 12223 21692 12232
rect 21640 12189 21649 12223
rect 21649 12189 21683 12223
rect 21683 12189 21692 12223
rect 21640 12180 21692 12189
rect 8208 12112 8260 12164
rect 19892 12155 19944 12164
rect 19892 12121 19901 12155
rect 19901 12121 19935 12155
rect 19935 12121 19944 12155
rect 19892 12112 19944 12121
rect 6920 12044 6972 12096
rect 9128 12087 9180 12096
rect 9128 12053 9137 12087
rect 9137 12053 9171 12087
rect 9171 12053 9180 12087
rect 9128 12044 9180 12053
rect 12716 12044 12768 12096
rect 16488 12044 16540 12096
rect 19984 12044 20036 12096
rect 23572 12044 23624 12096
rect 4982 11942 5034 11994
rect 5046 11942 5098 11994
rect 5110 11942 5162 11994
rect 5174 11942 5226 11994
rect 12982 11942 13034 11994
rect 13046 11942 13098 11994
rect 13110 11942 13162 11994
rect 13174 11942 13226 11994
rect 20982 11942 21034 11994
rect 21046 11942 21098 11994
rect 21110 11942 21162 11994
rect 21174 11942 21226 11994
rect 3700 11883 3752 11892
rect 3700 11849 3709 11883
rect 3709 11849 3743 11883
rect 3743 11849 3752 11883
rect 3700 11840 3752 11849
rect 4252 11840 4304 11892
rect 5724 11883 5776 11892
rect 5724 11849 5733 11883
rect 5733 11849 5767 11883
rect 5767 11849 5776 11883
rect 5724 11840 5776 11849
rect 5816 11840 5868 11892
rect 2044 11636 2096 11688
rect 3976 11815 4028 11824
rect 3976 11781 3985 11815
rect 3985 11781 4019 11815
rect 4019 11781 4028 11815
rect 3976 11772 4028 11781
rect 4160 11772 4212 11824
rect 6184 11772 6236 11824
rect 6920 11815 6972 11824
rect 6920 11781 6929 11815
rect 6929 11781 6963 11815
rect 6963 11781 6972 11815
rect 6920 11772 6972 11781
rect 2688 11747 2740 11756
rect 2688 11713 2697 11747
rect 2697 11713 2731 11747
rect 2731 11713 2740 11747
rect 2688 11704 2740 11713
rect 3700 11636 3752 11688
rect 2320 11611 2372 11620
rect 2320 11577 2329 11611
rect 2329 11577 2363 11611
rect 2363 11577 2372 11611
rect 2320 11568 2372 11577
rect 4068 11704 4120 11756
rect 6828 11679 6880 11688
rect 6828 11645 6837 11679
rect 6837 11645 6871 11679
rect 6871 11645 6880 11679
rect 6828 11636 6880 11645
rect 7288 11636 7340 11688
rect 11888 11840 11940 11892
rect 13636 11883 13688 11892
rect 13636 11849 13645 11883
rect 13645 11849 13679 11883
rect 13679 11849 13688 11883
rect 13636 11840 13688 11849
rect 15752 11883 15804 11892
rect 15752 11849 15761 11883
rect 15761 11849 15795 11883
rect 15795 11849 15804 11883
rect 15752 11840 15804 11849
rect 19708 11883 19760 11892
rect 19708 11849 19717 11883
rect 19717 11849 19751 11883
rect 19751 11849 19760 11883
rect 19708 11840 19760 11849
rect 20720 11840 20772 11892
rect 11060 11772 11112 11824
rect 12072 11772 12124 11824
rect 12624 11772 12676 11824
rect 12716 11704 12768 11756
rect 16028 11772 16080 11824
rect 16948 11704 17000 11756
rect 17408 11704 17460 11756
rect 19984 11772 20036 11824
rect 21272 11772 21324 11824
rect 7840 11636 7892 11688
rect 8116 11636 8168 11688
rect 9128 11636 9180 11688
rect 9588 11679 9640 11688
rect 6184 11568 6236 11620
rect 7656 11568 7708 11620
rect 9588 11645 9597 11679
rect 9597 11645 9631 11679
rect 9631 11645 9640 11679
rect 9588 11636 9640 11645
rect 9956 11679 10008 11688
rect 9956 11645 9965 11679
rect 9965 11645 9999 11679
rect 9999 11645 10008 11679
rect 9956 11636 10008 11645
rect 11336 11636 11388 11688
rect 11888 11636 11940 11688
rect 14464 11679 14516 11688
rect 10508 11568 10560 11620
rect 1768 11500 1820 11552
rect 2688 11500 2740 11552
rect 4344 11543 4396 11552
rect 4344 11509 4353 11543
rect 4353 11509 4387 11543
rect 4387 11509 4396 11543
rect 4344 11500 4396 11509
rect 6828 11500 6880 11552
rect 8024 11500 8076 11552
rect 8208 11543 8260 11552
rect 8208 11509 8217 11543
rect 8217 11509 8251 11543
rect 8251 11509 8260 11543
rect 8208 11500 8260 11509
rect 9312 11500 9364 11552
rect 10600 11543 10652 11552
rect 10600 11509 10609 11543
rect 10609 11509 10643 11543
rect 10643 11509 10652 11543
rect 10600 11500 10652 11509
rect 11244 11500 11296 11552
rect 11888 11543 11940 11552
rect 11888 11509 11897 11543
rect 11897 11509 11931 11543
rect 11931 11509 11940 11543
rect 11888 11500 11940 11509
rect 12808 11568 12860 11620
rect 14464 11645 14473 11679
rect 14473 11645 14507 11679
rect 14507 11645 14516 11679
rect 14464 11636 14516 11645
rect 16488 11611 16540 11620
rect 16488 11577 16497 11611
rect 16497 11577 16531 11611
rect 16531 11577 16540 11611
rect 16488 11568 16540 11577
rect 16580 11611 16632 11620
rect 16580 11577 16589 11611
rect 16589 11577 16623 11611
rect 16623 11577 16632 11611
rect 16580 11568 16632 11577
rect 13452 11500 13504 11552
rect 14004 11500 14056 11552
rect 16304 11543 16356 11552
rect 16304 11509 16313 11543
rect 16313 11509 16347 11543
rect 16347 11509 16356 11543
rect 16304 11500 16356 11509
rect 18144 11500 18196 11552
rect 18972 11543 19024 11552
rect 18972 11509 18981 11543
rect 18981 11509 19015 11543
rect 19015 11509 19024 11543
rect 18972 11500 19024 11509
rect 20168 11611 20220 11620
rect 20168 11577 20177 11611
rect 20177 11577 20211 11611
rect 20211 11577 20220 11611
rect 20720 11611 20772 11620
rect 20168 11568 20220 11577
rect 20720 11577 20729 11611
rect 20729 11577 20763 11611
rect 20763 11577 20772 11611
rect 20720 11568 20772 11577
rect 20628 11500 20680 11552
rect 21548 11500 21600 11552
rect 8982 11398 9034 11450
rect 9046 11398 9098 11450
rect 9110 11398 9162 11450
rect 9174 11398 9226 11450
rect 16982 11398 17034 11450
rect 17046 11398 17098 11450
rect 17110 11398 17162 11450
rect 17174 11398 17226 11450
rect 1768 11339 1820 11348
rect 1768 11305 1777 11339
rect 1777 11305 1811 11339
rect 1811 11305 1820 11339
rect 1768 11296 1820 11305
rect 2412 11296 2464 11348
rect 6552 11296 6604 11348
rect 2504 11228 2556 11280
rect 3792 11228 3844 11280
rect 2044 11203 2096 11212
rect 2044 11169 2053 11203
rect 2053 11169 2087 11203
rect 2087 11169 2096 11203
rect 2044 11160 2096 11169
rect 4712 11203 4764 11212
rect 4712 11169 4721 11203
rect 4721 11169 4755 11203
rect 4755 11169 4764 11203
rect 4712 11160 4764 11169
rect 8852 11296 8904 11348
rect 9588 11296 9640 11348
rect 12348 11296 12400 11348
rect 12808 11296 12860 11348
rect 14004 11339 14056 11348
rect 14004 11305 14013 11339
rect 14013 11305 14047 11339
rect 14047 11305 14056 11339
rect 14004 11296 14056 11305
rect 16028 11339 16080 11348
rect 16028 11305 16037 11339
rect 16037 11305 16071 11339
rect 16071 11305 16080 11339
rect 16028 11296 16080 11305
rect 16304 11296 16356 11348
rect 16580 11339 16632 11348
rect 16580 11305 16589 11339
rect 16589 11305 16623 11339
rect 16623 11305 16632 11339
rect 16580 11296 16632 11305
rect 9404 11228 9456 11280
rect 10416 11228 10468 11280
rect 12256 11228 12308 11280
rect 12164 11203 12216 11212
rect 1860 11092 1912 11144
rect 5908 11092 5960 11144
rect 12164 11169 12173 11203
rect 12173 11169 12207 11203
rect 12207 11169 12216 11203
rect 12164 11160 12216 11169
rect 17868 11160 17920 11212
rect 20168 11228 20220 11280
rect 21272 11228 21324 11280
rect 21640 11271 21692 11280
rect 21640 11237 21649 11271
rect 21649 11237 21683 11271
rect 21683 11237 21692 11271
rect 21640 11228 21692 11237
rect 19984 11203 20036 11212
rect 19984 11169 19993 11203
rect 19993 11169 20027 11203
rect 20027 11169 20036 11203
rect 19984 11160 20036 11169
rect 10876 11092 10928 11144
rect 15660 11135 15712 11144
rect 15660 11101 15669 11135
rect 15669 11101 15703 11135
rect 15703 11101 15712 11135
rect 15660 11092 15712 11101
rect 21456 11092 21508 11144
rect 8024 11024 8076 11076
rect 8208 11024 8260 11076
rect 14464 11067 14516 11076
rect 14464 11033 14473 11067
rect 14473 11033 14507 11067
rect 14507 11033 14516 11067
rect 14464 11024 14516 11033
rect 15844 11024 15896 11076
rect 3240 10956 3292 11008
rect 3700 10956 3752 11008
rect 5724 10956 5776 11008
rect 7380 10956 7432 11008
rect 7932 10956 7984 11008
rect 12808 10956 12860 11008
rect 15936 10956 15988 11008
rect 18144 10999 18196 11008
rect 18144 10965 18153 10999
rect 18153 10965 18187 10999
rect 18187 10965 18196 10999
rect 18144 10956 18196 10965
rect 18512 10956 18564 11008
rect 20628 10999 20680 11008
rect 20628 10965 20637 10999
rect 20637 10965 20671 10999
rect 20671 10965 20680 10999
rect 20628 10956 20680 10965
rect 4982 10854 5034 10906
rect 5046 10854 5098 10906
rect 5110 10854 5162 10906
rect 5174 10854 5226 10906
rect 12982 10854 13034 10906
rect 13046 10854 13098 10906
rect 13110 10854 13162 10906
rect 13174 10854 13226 10906
rect 20982 10854 21034 10906
rect 21046 10854 21098 10906
rect 21110 10854 21162 10906
rect 21174 10854 21226 10906
rect 1584 10795 1636 10804
rect 1584 10761 1593 10795
rect 1593 10761 1627 10795
rect 1627 10761 1636 10795
rect 1584 10752 1636 10761
rect 2504 10752 2556 10804
rect 4344 10752 4396 10804
rect 5908 10795 5960 10804
rect 4068 10684 4120 10736
rect 2412 10616 2464 10668
rect 2964 10659 3016 10668
rect 2964 10625 2973 10659
rect 2973 10625 3007 10659
rect 3007 10625 3016 10659
rect 2964 10616 3016 10625
rect 5908 10761 5917 10795
rect 5917 10761 5951 10795
rect 5951 10761 5960 10795
rect 5908 10752 5960 10761
rect 6552 10752 6604 10804
rect 10416 10795 10468 10804
rect 10416 10761 10425 10795
rect 10425 10761 10459 10795
rect 10459 10761 10468 10795
rect 10416 10752 10468 10761
rect 12164 10752 12216 10804
rect 20168 10752 20220 10804
rect 21272 10795 21324 10804
rect 21272 10761 21281 10795
rect 21281 10761 21315 10795
rect 21315 10761 21324 10795
rect 21272 10752 21324 10761
rect 21548 10795 21600 10804
rect 21548 10761 21557 10795
rect 21557 10761 21591 10795
rect 21591 10761 21600 10795
rect 21548 10752 21600 10761
rect 9956 10684 10008 10736
rect 10600 10684 10652 10736
rect 19984 10727 20036 10736
rect 10324 10616 10376 10668
rect 19984 10693 19993 10727
rect 19993 10693 20027 10727
rect 20027 10693 20036 10727
rect 19984 10684 20036 10693
rect 18972 10616 19024 10668
rect 20260 10659 20312 10668
rect 20260 10625 20269 10659
rect 20269 10625 20303 10659
rect 20303 10625 20312 10659
rect 20260 10616 20312 10625
rect 20720 10659 20772 10668
rect 20720 10625 20729 10659
rect 20729 10625 20763 10659
rect 20763 10625 20772 10659
rect 20720 10616 20772 10625
rect 2780 10523 2832 10532
rect 2780 10489 2789 10523
rect 2789 10489 2823 10523
rect 2823 10489 2832 10523
rect 2780 10480 2832 10489
rect 7564 10548 7616 10600
rect 8116 10591 8168 10600
rect 8116 10557 8125 10591
rect 8125 10557 8159 10591
rect 8159 10557 8168 10591
rect 8116 10548 8168 10557
rect 8208 10548 8260 10600
rect 8852 10548 8904 10600
rect 9312 10591 9364 10600
rect 9312 10557 9321 10591
rect 9321 10557 9355 10591
rect 9355 10557 9364 10591
rect 9312 10548 9364 10557
rect 10508 10591 10560 10600
rect 10508 10557 10517 10591
rect 10517 10557 10551 10591
rect 10551 10557 10560 10591
rect 10508 10548 10560 10557
rect 11060 10591 11112 10600
rect 11060 10557 11069 10591
rect 11069 10557 11103 10591
rect 11103 10557 11112 10591
rect 11060 10548 11112 10557
rect 15016 10548 15068 10600
rect 15936 10591 15988 10600
rect 3792 10455 3844 10464
rect 3792 10421 3801 10455
rect 3801 10421 3835 10455
rect 3835 10421 3844 10455
rect 3792 10412 3844 10421
rect 5448 10480 5500 10532
rect 9496 10480 9548 10532
rect 12624 10480 12676 10532
rect 12900 10523 12952 10532
rect 12900 10489 12909 10523
rect 12909 10489 12943 10523
rect 12943 10489 12952 10523
rect 13452 10523 13504 10532
rect 12900 10480 12952 10489
rect 13452 10489 13461 10523
rect 13461 10489 13495 10523
rect 13495 10489 13504 10523
rect 13452 10480 13504 10489
rect 13912 10480 13964 10532
rect 14004 10480 14056 10532
rect 15936 10557 15945 10591
rect 15945 10557 15979 10591
rect 15979 10557 15988 10591
rect 15936 10548 15988 10557
rect 16304 10591 16356 10600
rect 16304 10557 16313 10591
rect 16313 10557 16347 10591
rect 16347 10557 16356 10591
rect 16304 10548 16356 10557
rect 15660 10480 15712 10532
rect 17868 10523 17920 10532
rect 17868 10489 17877 10523
rect 17877 10489 17911 10523
rect 17911 10489 17920 10523
rect 17868 10480 17920 10489
rect 19984 10480 20036 10532
rect 8024 10455 8076 10464
rect 8024 10421 8033 10455
rect 8033 10421 8067 10455
rect 8067 10421 8076 10455
rect 8024 10412 8076 10421
rect 8576 10412 8628 10464
rect 10876 10412 10928 10464
rect 12256 10455 12308 10464
rect 12256 10421 12265 10455
rect 12265 10421 12299 10455
rect 12299 10421 12308 10455
rect 12256 10412 12308 10421
rect 18144 10412 18196 10464
rect 8982 10310 9034 10362
rect 9046 10310 9098 10362
rect 9110 10310 9162 10362
rect 9174 10310 9226 10362
rect 16982 10310 17034 10362
rect 17046 10310 17098 10362
rect 17110 10310 17162 10362
rect 17174 10310 17226 10362
rect 4712 10251 4764 10260
rect 2136 10140 2188 10192
rect 4712 10217 4721 10251
rect 4721 10217 4755 10251
rect 4755 10217 4764 10251
rect 4712 10208 4764 10217
rect 8852 10208 8904 10260
rect 10508 10251 10560 10260
rect 10508 10217 10517 10251
rect 10517 10217 10551 10251
rect 10551 10217 10560 10251
rect 10508 10208 10560 10217
rect 10876 10251 10928 10260
rect 10876 10217 10885 10251
rect 10885 10217 10919 10251
rect 10919 10217 10928 10251
rect 10876 10208 10928 10217
rect 12808 10251 12860 10260
rect 12808 10217 12817 10251
rect 12817 10217 12851 10251
rect 12851 10217 12860 10251
rect 12808 10208 12860 10217
rect 15660 10208 15712 10260
rect 16028 10208 16080 10260
rect 18144 10208 18196 10260
rect 20628 10208 20680 10260
rect 21364 10208 21416 10260
rect 2780 10140 2832 10192
rect 3976 10140 4028 10192
rect 5816 10183 5868 10192
rect 5816 10149 5819 10183
rect 5819 10149 5853 10183
rect 5853 10149 5868 10183
rect 5816 10140 5868 10149
rect 6552 10140 6604 10192
rect 7380 10183 7432 10192
rect 7380 10149 7389 10183
rect 7389 10149 7423 10183
rect 7423 10149 7432 10183
rect 7380 10140 7432 10149
rect 11428 10183 11480 10192
rect 11428 10149 11437 10183
rect 11437 10149 11471 10183
rect 11471 10149 11480 10183
rect 11428 10140 11480 10149
rect 14188 10140 14240 10192
rect 17500 10140 17552 10192
rect 20260 10183 20312 10192
rect 20260 10149 20269 10183
rect 20269 10149 20303 10183
rect 20303 10149 20312 10183
rect 20260 10140 20312 10149
rect 1768 10072 1820 10124
rect 4068 10072 4120 10124
rect 7012 10072 7064 10124
rect 13268 10115 13320 10124
rect 13268 10081 13277 10115
rect 13277 10081 13311 10115
rect 13311 10081 13320 10115
rect 13268 10072 13320 10081
rect 13544 10115 13596 10124
rect 13544 10081 13553 10115
rect 13553 10081 13587 10115
rect 13587 10081 13596 10115
rect 13544 10072 13596 10081
rect 15476 10115 15528 10124
rect 15476 10081 15485 10115
rect 15485 10081 15519 10115
rect 15519 10081 15528 10115
rect 15476 10072 15528 10081
rect 15844 10115 15896 10124
rect 15844 10081 15853 10115
rect 15853 10081 15887 10115
rect 15887 10081 15896 10115
rect 15844 10072 15896 10081
rect 16856 10115 16908 10124
rect 16856 10081 16865 10115
rect 16865 10081 16899 10115
rect 16899 10081 16908 10115
rect 16856 10072 16908 10081
rect 19156 10072 19208 10124
rect 19524 10072 19576 10124
rect 20904 10115 20956 10124
rect 20904 10081 20913 10115
rect 20913 10081 20947 10115
rect 20947 10081 20956 10115
rect 20904 10072 20956 10081
rect 21548 10072 21600 10124
rect 5448 10047 5500 10056
rect 5448 10013 5457 10047
rect 5457 10013 5491 10047
rect 5491 10013 5500 10047
rect 5448 10004 5500 10013
rect 7104 10004 7156 10056
rect 7564 10047 7616 10056
rect 7564 10013 7573 10047
rect 7573 10013 7607 10047
rect 7607 10013 7616 10047
rect 7564 10004 7616 10013
rect 11336 10047 11388 10056
rect 11336 10013 11345 10047
rect 11345 10013 11379 10047
rect 11379 10013 11388 10047
rect 11336 10004 11388 10013
rect 11612 10047 11664 10056
rect 11612 10013 11621 10047
rect 11621 10013 11655 10047
rect 11655 10013 11664 10047
rect 11612 10004 11664 10013
rect 12624 10004 12676 10056
rect 17960 10047 18012 10056
rect 17960 10013 17969 10047
rect 17969 10013 18003 10047
rect 18003 10013 18012 10047
rect 17960 10004 18012 10013
rect 18788 10004 18840 10056
rect 3700 9936 3752 9988
rect 13912 9936 13964 9988
rect 3608 9911 3660 9920
rect 3608 9877 3617 9911
rect 3617 9877 3651 9911
rect 3651 9877 3660 9911
rect 3608 9868 3660 9877
rect 3884 9868 3936 9920
rect 4712 9868 4764 9920
rect 7104 9911 7156 9920
rect 7104 9877 7113 9911
rect 7113 9877 7147 9911
rect 7147 9877 7156 9911
rect 7104 9868 7156 9877
rect 8208 9911 8260 9920
rect 8208 9877 8217 9911
rect 8217 9877 8251 9911
rect 8251 9877 8260 9911
rect 8208 9868 8260 9877
rect 9312 9868 9364 9920
rect 14832 9868 14884 9920
rect 18144 9868 18196 9920
rect 4982 9766 5034 9818
rect 5046 9766 5098 9818
rect 5110 9766 5162 9818
rect 5174 9766 5226 9818
rect 12982 9766 13034 9818
rect 13046 9766 13098 9818
rect 13110 9766 13162 9818
rect 13174 9766 13226 9818
rect 20982 9766 21034 9818
rect 21046 9766 21098 9818
rect 21110 9766 21162 9818
rect 21174 9766 21226 9818
rect 2136 9664 2188 9716
rect 3608 9664 3660 9716
rect 5448 9664 5500 9716
rect 7380 9664 7432 9716
rect 7748 9664 7800 9716
rect 8852 9664 8904 9716
rect 11428 9664 11480 9716
rect 16856 9707 16908 9716
rect 16856 9673 16865 9707
rect 16865 9673 16899 9707
rect 16899 9673 16908 9707
rect 16856 9664 16908 9673
rect 21548 9707 21600 9716
rect 21548 9673 21557 9707
rect 21557 9673 21591 9707
rect 21591 9673 21600 9707
rect 21548 9664 21600 9673
rect 2964 9596 3016 9648
rect 8024 9596 8076 9648
rect 13544 9596 13596 9648
rect 14556 9639 14608 9648
rect 14556 9605 14565 9639
rect 14565 9605 14599 9639
rect 14599 9605 14608 9639
rect 14556 9596 14608 9605
rect 14832 9596 14884 9648
rect 3700 9528 3752 9580
rect 4436 9528 4488 9580
rect 5540 9528 5592 9580
rect 11612 9528 11664 9580
rect 15384 9528 15436 9580
rect 4068 9503 4120 9512
rect 4068 9469 4077 9503
rect 4077 9469 4111 9503
rect 4111 9469 4120 9503
rect 4068 9460 4120 9469
rect 7656 9460 7708 9512
rect 9496 9503 9548 9512
rect 9496 9469 9505 9503
rect 9505 9469 9539 9503
rect 9539 9469 9548 9503
rect 9496 9460 9548 9469
rect 12440 9503 12492 9512
rect 12440 9469 12449 9503
rect 12449 9469 12483 9503
rect 12483 9469 12492 9503
rect 12440 9460 12492 9469
rect 12900 9503 12952 9512
rect 12900 9469 12909 9503
rect 12909 9469 12943 9503
rect 12943 9469 12952 9503
rect 12900 9460 12952 9469
rect 14556 9460 14608 9512
rect 15016 9503 15068 9512
rect 15016 9469 15025 9503
rect 15025 9469 15059 9503
rect 15059 9469 15068 9503
rect 15016 9460 15068 9469
rect 3516 9435 3568 9444
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 2044 9324 2096 9376
rect 3516 9401 3525 9435
rect 3525 9401 3559 9435
rect 3559 9401 3568 9435
rect 3516 9392 3568 9401
rect 3976 9392 4028 9444
rect 4436 9435 4488 9444
rect 3148 9324 3200 9376
rect 4436 9401 4445 9435
rect 4445 9401 4479 9435
rect 4479 9401 4488 9435
rect 4436 9392 4488 9401
rect 6736 9392 6788 9444
rect 6920 9435 6972 9444
rect 6920 9401 6929 9435
rect 6929 9401 6963 9435
rect 6963 9401 6972 9435
rect 6920 9392 6972 9401
rect 7012 9435 7064 9444
rect 7012 9401 7021 9435
rect 7021 9401 7055 9435
rect 7055 9401 7064 9435
rect 7564 9435 7616 9444
rect 7012 9392 7064 9401
rect 7564 9401 7573 9435
rect 7573 9401 7607 9435
rect 7607 9401 7616 9435
rect 7564 9392 7616 9401
rect 9680 9435 9732 9444
rect 9680 9401 9689 9435
rect 9689 9401 9723 9435
rect 9723 9401 9732 9435
rect 9680 9392 9732 9401
rect 10692 9435 10744 9444
rect 10692 9401 10701 9435
rect 10701 9401 10735 9435
rect 10735 9401 10744 9435
rect 10692 9392 10744 9401
rect 5816 9324 5868 9376
rect 8116 9324 8168 9376
rect 8484 9367 8536 9376
rect 8484 9333 8493 9367
rect 8493 9333 8527 9367
rect 8527 9333 8536 9367
rect 8484 9324 8536 9333
rect 10232 9324 10284 9376
rect 11336 9392 11388 9444
rect 12716 9367 12768 9376
rect 12716 9333 12725 9367
rect 12725 9333 12759 9367
rect 12759 9333 12768 9367
rect 12716 9324 12768 9333
rect 13820 9367 13872 9376
rect 13820 9333 13829 9367
rect 13829 9333 13863 9367
rect 13863 9333 13872 9367
rect 13820 9324 13872 9333
rect 15108 9324 15160 9376
rect 15936 9460 15988 9512
rect 17960 9596 18012 9648
rect 18144 9571 18196 9580
rect 18144 9537 18153 9571
rect 18153 9537 18187 9571
rect 18187 9537 18196 9571
rect 18144 9528 18196 9537
rect 20720 9528 20772 9580
rect 16488 9460 16540 9512
rect 18788 9435 18840 9444
rect 16028 9324 16080 9376
rect 17500 9367 17552 9376
rect 17500 9333 17509 9367
rect 17509 9333 17543 9367
rect 17543 9333 17552 9367
rect 17500 9324 17552 9333
rect 17868 9367 17920 9376
rect 17868 9333 17877 9367
rect 17877 9333 17911 9367
rect 17911 9333 17920 9367
rect 18788 9401 18797 9435
rect 18797 9401 18831 9435
rect 18831 9401 18840 9435
rect 18788 9392 18840 9401
rect 20812 9392 20864 9444
rect 21272 9435 21324 9444
rect 21272 9401 21281 9435
rect 21281 9401 21315 9435
rect 21315 9401 21324 9435
rect 21272 9392 21324 9401
rect 17868 9324 17920 9333
rect 19524 9324 19576 9376
rect 8982 9222 9034 9274
rect 9046 9222 9098 9274
rect 9110 9222 9162 9274
rect 9174 9222 9226 9274
rect 16982 9222 17034 9274
rect 17046 9222 17098 9274
rect 17110 9222 17162 9274
rect 17174 9222 17226 9274
rect 3148 9163 3200 9172
rect 3148 9129 3157 9163
rect 3157 9129 3191 9163
rect 3191 9129 3200 9163
rect 3148 9120 3200 9129
rect 3700 9120 3752 9172
rect 4436 9120 4488 9172
rect 7012 9120 7064 9172
rect 8576 9120 8628 9172
rect 9496 9120 9548 9172
rect 10416 9120 10468 9172
rect 10692 9120 10744 9172
rect 14740 9163 14792 9172
rect 14740 9129 14749 9163
rect 14749 9129 14783 9163
rect 14783 9129 14792 9163
rect 14740 9120 14792 9129
rect 15016 9120 15068 9172
rect 15476 9163 15528 9172
rect 15476 9129 15485 9163
rect 15485 9129 15519 9163
rect 15519 9129 15528 9163
rect 15476 9120 15528 9129
rect 17500 9120 17552 9172
rect 5816 9052 5868 9104
rect 2044 9027 2096 9036
rect 2044 8993 2053 9027
rect 2053 8993 2087 9027
rect 2087 8993 2096 9027
rect 2044 8984 2096 8993
rect 2320 9027 2372 9036
rect 2320 8993 2329 9027
rect 2329 8993 2363 9027
rect 2363 8993 2372 9027
rect 2320 8984 2372 8993
rect 3884 8984 3936 9036
rect 4436 8984 4488 9036
rect 6000 8984 6052 9036
rect 6644 9052 6696 9104
rect 11336 9095 11388 9104
rect 11336 9061 11345 9095
rect 11345 9061 11379 9095
rect 11379 9061 11388 9095
rect 11336 9052 11388 9061
rect 12256 9052 12308 9104
rect 16212 9052 16264 9104
rect 18512 9095 18564 9104
rect 18512 9061 18521 9095
rect 18521 9061 18555 9095
rect 18555 9061 18564 9095
rect 18512 9052 18564 9061
rect 20720 9120 20772 9172
rect 19248 9052 19300 9104
rect 21640 9120 21692 9172
rect 21088 9095 21140 9104
rect 21088 9061 21097 9095
rect 21097 9061 21131 9095
rect 21131 9061 21140 9095
rect 21088 9052 21140 9061
rect 9680 9027 9732 9036
rect 9680 8993 9689 9027
rect 9689 8993 9723 9027
rect 9723 8993 9732 9027
rect 9680 8984 9732 8993
rect 11244 8984 11296 9036
rect 12716 9027 12768 9036
rect 12716 8993 12725 9027
rect 12725 8993 12759 9027
rect 12759 8993 12768 9027
rect 12716 8984 12768 8993
rect 1860 8916 1912 8968
rect 1952 8780 2004 8832
rect 3792 8916 3844 8968
rect 5356 8959 5408 8968
rect 5356 8925 5365 8959
rect 5365 8925 5399 8959
rect 5399 8925 5408 8959
rect 5356 8916 5408 8925
rect 6736 8916 6788 8968
rect 7380 8916 7432 8968
rect 7564 8959 7616 8968
rect 7564 8925 7573 8959
rect 7573 8925 7607 8959
rect 7607 8925 7616 8959
rect 7564 8916 7616 8925
rect 11060 8916 11112 8968
rect 12900 8916 12952 8968
rect 13268 8916 13320 8968
rect 15016 8959 15068 8968
rect 15016 8925 15025 8959
rect 15025 8925 15059 8959
rect 15059 8925 15068 8959
rect 15016 8916 15068 8925
rect 16028 8959 16080 8968
rect 16028 8925 16037 8959
rect 16037 8925 16071 8959
rect 16071 8925 16080 8959
rect 16028 8916 16080 8925
rect 18972 8959 19024 8968
rect 18972 8925 18981 8959
rect 18981 8925 19015 8959
rect 19015 8925 19024 8959
rect 18972 8916 19024 8925
rect 21272 8959 21324 8968
rect 21272 8925 21281 8959
rect 21281 8925 21315 8959
rect 21315 8925 21324 8959
rect 21272 8916 21324 8925
rect 10692 8848 10744 8900
rect 20720 8848 20772 8900
rect 21088 8848 21140 8900
rect 4712 8823 4764 8832
rect 4712 8789 4721 8823
rect 4721 8789 4755 8823
rect 4755 8789 4764 8823
rect 4712 8780 4764 8789
rect 4804 8780 4856 8832
rect 10232 8780 10284 8832
rect 13636 8823 13688 8832
rect 13636 8789 13645 8823
rect 13645 8789 13679 8823
rect 13679 8789 13688 8823
rect 13636 8780 13688 8789
rect 15844 8823 15896 8832
rect 15844 8789 15853 8823
rect 15853 8789 15887 8823
rect 15887 8789 15896 8823
rect 15844 8780 15896 8789
rect 18236 8823 18288 8832
rect 18236 8789 18245 8823
rect 18245 8789 18279 8823
rect 18279 8789 18288 8823
rect 18236 8780 18288 8789
rect 4982 8678 5034 8730
rect 5046 8678 5098 8730
rect 5110 8678 5162 8730
rect 5174 8678 5226 8730
rect 12982 8678 13034 8730
rect 13046 8678 13098 8730
rect 13110 8678 13162 8730
rect 13174 8678 13226 8730
rect 20982 8678 21034 8730
rect 21046 8678 21098 8730
rect 21110 8678 21162 8730
rect 21174 8678 21226 8730
rect 2320 8576 2372 8628
rect 2044 8508 2096 8560
rect 3240 8551 3292 8560
rect 3240 8517 3249 8551
rect 3249 8517 3283 8551
rect 3283 8517 3292 8551
rect 3240 8508 3292 8517
rect 1860 8440 1912 8492
rect 1676 8415 1728 8424
rect 1676 8381 1685 8415
rect 1685 8381 1719 8415
rect 1719 8381 1728 8415
rect 1676 8372 1728 8381
rect 1952 8415 2004 8424
rect 1952 8381 1961 8415
rect 1961 8381 1995 8415
rect 1995 8381 2004 8415
rect 1952 8372 2004 8381
rect 6092 8576 6144 8628
rect 6644 8619 6696 8628
rect 6644 8585 6653 8619
rect 6653 8585 6687 8619
rect 6687 8585 6696 8619
rect 6644 8576 6696 8585
rect 10324 8576 10376 8628
rect 11428 8576 11480 8628
rect 12716 8576 12768 8628
rect 4528 8508 4580 8560
rect 5356 8483 5408 8492
rect 5356 8449 5365 8483
rect 5365 8449 5399 8483
rect 5399 8449 5408 8483
rect 5356 8440 5408 8449
rect 4712 8415 4764 8424
rect 4712 8381 4721 8415
rect 4721 8381 4755 8415
rect 4755 8381 4764 8415
rect 4712 8372 4764 8381
rect 4804 8372 4856 8424
rect 5816 8372 5868 8424
rect 11244 8440 11296 8492
rect 12256 8440 12308 8492
rect 13544 8508 13596 8560
rect 13452 8483 13504 8492
rect 13452 8449 13461 8483
rect 13461 8449 13495 8483
rect 13495 8449 13504 8483
rect 13452 8440 13504 8449
rect 16028 8576 16080 8628
rect 20720 8576 20772 8628
rect 21640 8576 21692 8628
rect 17500 8508 17552 8560
rect 16212 8440 16264 8492
rect 18236 8483 18288 8492
rect 1768 8279 1820 8288
rect 1768 8245 1777 8279
rect 1777 8245 1811 8279
rect 1811 8245 1820 8279
rect 1768 8236 1820 8245
rect 3884 8236 3936 8288
rect 4436 8279 4488 8288
rect 4436 8245 4445 8279
rect 4445 8245 4479 8279
rect 4479 8245 4488 8279
rect 4436 8236 4488 8245
rect 6736 8236 6788 8288
rect 8576 8415 8628 8424
rect 8576 8381 8585 8415
rect 8585 8381 8619 8415
rect 8619 8381 8628 8415
rect 8576 8372 8628 8381
rect 7564 8236 7616 8288
rect 10416 8304 10468 8356
rect 13636 8304 13688 8356
rect 18236 8449 18245 8483
rect 18245 8449 18279 8483
rect 18279 8449 18288 8483
rect 18236 8440 18288 8449
rect 19616 8440 19668 8492
rect 19248 8415 19300 8424
rect 19248 8381 19257 8415
rect 19257 8381 19291 8415
rect 19291 8381 19300 8415
rect 19248 8372 19300 8381
rect 21272 8372 21324 8424
rect 17684 8304 17736 8356
rect 17868 8347 17920 8356
rect 17868 8313 17877 8347
rect 17877 8313 17911 8347
rect 17911 8313 17920 8347
rect 17868 8304 17920 8313
rect 15384 8236 15436 8288
rect 18972 8304 19024 8356
rect 19156 8236 19208 8288
rect 8982 8134 9034 8186
rect 9046 8134 9098 8186
rect 9110 8134 9162 8186
rect 9174 8134 9226 8186
rect 16982 8134 17034 8186
rect 17046 8134 17098 8186
rect 17110 8134 17162 8186
rect 17174 8134 17226 8186
rect 1676 8075 1728 8084
rect 1676 8041 1685 8075
rect 1685 8041 1719 8075
rect 1719 8041 1728 8075
rect 1676 8032 1728 8041
rect 2136 8075 2188 8084
rect 2136 8041 2145 8075
rect 2145 8041 2179 8075
rect 2179 8041 2188 8075
rect 2136 8032 2188 8041
rect 4712 8032 4764 8084
rect 3884 7964 3936 8016
rect 4252 8007 4304 8016
rect 4252 7973 4261 8007
rect 4261 7973 4295 8007
rect 4295 7973 4304 8007
rect 4252 7964 4304 7973
rect 6736 8007 6788 8016
rect 6736 7973 6745 8007
rect 6745 7973 6779 8007
rect 6779 7973 6788 8007
rect 6736 7964 6788 7973
rect 6828 8007 6880 8016
rect 6828 7973 6837 8007
rect 6837 7973 6871 8007
rect 6871 7973 6880 8007
rect 7380 8032 7432 8084
rect 8576 8032 8628 8084
rect 9680 8032 9732 8084
rect 15384 8075 15436 8084
rect 15384 8041 15393 8075
rect 15393 8041 15427 8075
rect 15427 8041 15436 8075
rect 15384 8032 15436 8041
rect 18512 8032 18564 8084
rect 19616 8075 19668 8084
rect 19616 8041 19625 8075
rect 19625 8041 19659 8075
rect 19659 8041 19668 8075
rect 19616 8032 19668 8041
rect 6828 7964 6880 7973
rect 7840 7964 7892 8016
rect 6460 7896 6512 7948
rect 12256 7964 12308 8016
rect 12624 7964 12676 8016
rect 18236 8007 18288 8016
rect 18236 7973 18245 8007
rect 18245 7973 18279 8007
rect 18279 7973 18288 8007
rect 18236 7964 18288 7973
rect 20812 7964 20864 8016
rect 1768 7871 1820 7880
rect 1768 7837 1777 7871
rect 1777 7837 1811 7871
rect 1811 7837 1820 7871
rect 1768 7828 1820 7837
rect 3516 7828 3568 7880
rect 7104 7828 7156 7880
rect 10508 7828 10560 7880
rect 11060 7896 11112 7948
rect 15292 7939 15344 7948
rect 15292 7905 15301 7939
rect 15301 7905 15335 7939
rect 15335 7905 15344 7939
rect 15292 7896 15344 7905
rect 15752 7939 15804 7948
rect 15752 7905 15761 7939
rect 15761 7905 15795 7939
rect 15795 7905 15804 7939
rect 15752 7896 15804 7905
rect 15936 7896 15988 7948
rect 16304 7896 16356 7948
rect 20720 7896 20772 7948
rect 11428 7828 11480 7880
rect 11796 7828 11848 7880
rect 18788 7828 18840 7880
rect 13268 7803 13320 7812
rect 13268 7769 13277 7803
rect 13277 7769 13311 7803
rect 13311 7769 13320 7803
rect 13268 7760 13320 7769
rect 18696 7803 18748 7812
rect 18696 7769 18705 7803
rect 18705 7769 18739 7803
rect 18739 7769 18748 7803
rect 18696 7760 18748 7769
rect 6920 7692 6972 7744
rect 8484 7692 8536 7744
rect 9404 7692 9456 7744
rect 13544 7735 13596 7744
rect 13544 7701 13553 7735
rect 13553 7701 13587 7735
rect 13587 7701 13596 7735
rect 13544 7692 13596 7701
rect 4982 7590 5034 7642
rect 5046 7590 5098 7642
rect 5110 7590 5162 7642
rect 5174 7590 5226 7642
rect 12982 7590 13034 7642
rect 13046 7590 13098 7642
rect 13110 7590 13162 7642
rect 13174 7590 13226 7642
rect 20982 7590 21034 7642
rect 21046 7590 21098 7642
rect 21110 7590 21162 7642
rect 21174 7590 21226 7642
rect 1768 7488 1820 7540
rect 6460 7488 6512 7540
rect 7656 7488 7708 7540
rect 1860 7420 1912 7472
rect 2136 7352 2188 7404
rect 2964 7352 3016 7404
rect 6920 7395 6972 7404
rect 6920 7361 6929 7395
rect 6929 7361 6963 7395
rect 6963 7361 6972 7395
rect 6920 7352 6972 7361
rect 7380 7395 7432 7404
rect 7380 7361 7389 7395
rect 7389 7361 7423 7395
rect 7423 7361 7432 7395
rect 7380 7352 7432 7361
rect 4712 7284 4764 7336
rect 1952 7259 2004 7268
rect 1952 7225 1961 7259
rect 1961 7225 1995 7259
rect 1995 7225 2004 7259
rect 1952 7216 2004 7225
rect 2044 7259 2096 7268
rect 2044 7225 2053 7259
rect 2053 7225 2087 7259
rect 2087 7225 2096 7259
rect 3516 7259 3568 7268
rect 2044 7216 2096 7225
rect 3516 7225 3525 7259
rect 3525 7225 3559 7259
rect 3559 7225 3568 7259
rect 3516 7216 3568 7225
rect 3332 7191 3384 7200
rect 3332 7157 3341 7191
rect 3341 7157 3375 7191
rect 3375 7157 3384 7191
rect 5816 7216 5868 7268
rect 3332 7148 3384 7157
rect 4252 7148 4304 7200
rect 7564 7284 7616 7336
rect 8852 7488 8904 7540
rect 11060 7488 11112 7540
rect 11428 7531 11480 7540
rect 11428 7497 11437 7531
rect 11437 7497 11471 7531
rect 11471 7497 11480 7531
rect 11428 7488 11480 7497
rect 11796 7531 11848 7540
rect 11796 7497 11805 7531
rect 11805 7497 11839 7531
rect 11839 7497 11848 7531
rect 11796 7488 11848 7497
rect 12624 7531 12676 7540
rect 12624 7497 12633 7531
rect 12633 7497 12667 7531
rect 12667 7497 12676 7531
rect 12624 7488 12676 7497
rect 15936 7488 15988 7540
rect 17960 7488 18012 7540
rect 21272 7488 21324 7540
rect 13452 7463 13504 7472
rect 13452 7429 13461 7463
rect 13461 7429 13495 7463
rect 13495 7429 13504 7463
rect 13452 7420 13504 7429
rect 16304 7420 16356 7472
rect 18236 7420 18288 7472
rect 19064 7420 19116 7472
rect 20720 7420 20772 7472
rect 10508 7395 10560 7404
rect 10508 7361 10517 7395
rect 10517 7361 10551 7395
rect 10551 7361 10560 7395
rect 10508 7352 10560 7361
rect 10968 7395 11020 7404
rect 10968 7361 10977 7395
rect 10977 7361 11011 7395
rect 11011 7361 11020 7395
rect 10968 7352 11020 7361
rect 13268 7352 13320 7404
rect 14556 7352 14608 7404
rect 8852 7327 8904 7336
rect 8852 7293 8861 7327
rect 8861 7293 8895 7327
rect 8895 7293 8904 7327
rect 8852 7284 8904 7293
rect 9404 7284 9456 7336
rect 10232 7284 10284 7336
rect 14832 7284 14884 7336
rect 15292 7284 15344 7336
rect 18972 7352 19024 7404
rect 6736 7148 6788 7200
rect 8668 7216 8720 7268
rect 12900 7259 12952 7268
rect 12900 7225 12909 7259
rect 12909 7225 12943 7259
rect 12943 7225 12952 7259
rect 12900 7216 12952 7225
rect 13268 7216 13320 7268
rect 18420 7259 18472 7268
rect 18420 7225 18429 7259
rect 18429 7225 18463 7259
rect 18463 7225 18472 7259
rect 18420 7216 18472 7225
rect 18696 7216 18748 7268
rect 20812 7148 20864 7200
rect 8982 7046 9034 7098
rect 9046 7046 9098 7098
rect 9110 7046 9162 7098
rect 9174 7046 9226 7098
rect 16982 7046 17034 7098
rect 17046 7046 17098 7098
rect 17110 7046 17162 7098
rect 17174 7046 17226 7098
rect 1584 6987 1636 6996
rect 1584 6953 1593 6987
rect 1593 6953 1627 6987
rect 1627 6953 1636 6987
rect 1584 6944 1636 6953
rect 1952 6987 2004 6996
rect 1952 6953 1961 6987
rect 1961 6953 1995 6987
rect 1995 6953 2004 6987
rect 1952 6944 2004 6953
rect 3884 6987 3936 6996
rect 3884 6953 3893 6987
rect 3893 6953 3927 6987
rect 3927 6953 3936 6987
rect 3884 6944 3936 6953
rect 4252 6987 4304 6996
rect 4252 6953 4261 6987
rect 4261 6953 4295 6987
rect 4295 6953 4304 6987
rect 4252 6944 4304 6953
rect 4712 6987 4764 6996
rect 4712 6953 4721 6987
rect 4721 6953 4755 6987
rect 4755 6953 4764 6987
rect 4712 6944 4764 6953
rect 6920 6944 6972 6996
rect 14832 6944 14884 6996
rect 15752 6944 15804 6996
rect 2044 6876 2096 6928
rect 3332 6876 3384 6928
rect 6736 6919 6788 6928
rect 6736 6885 6745 6919
rect 6745 6885 6779 6919
rect 6779 6885 6788 6919
rect 6736 6876 6788 6885
rect 2872 6808 2924 6860
rect 4528 6851 4580 6860
rect 4528 6817 4537 6851
rect 4537 6817 4571 6851
rect 4571 6817 4580 6851
rect 4528 6808 4580 6817
rect 4804 6808 4856 6860
rect 5632 6808 5684 6860
rect 8760 6876 8812 6928
rect 10324 6919 10376 6928
rect 10324 6885 10333 6919
rect 10333 6885 10367 6919
rect 10367 6885 10376 6919
rect 10324 6876 10376 6885
rect 12348 6919 12400 6928
rect 12348 6885 12357 6919
rect 12357 6885 12391 6919
rect 12391 6885 12400 6919
rect 12348 6876 12400 6885
rect 14004 6808 14056 6860
rect 15292 6851 15344 6860
rect 15292 6817 15301 6851
rect 15301 6817 15335 6851
rect 15335 6817 15344 6851
rect 15292 6808 15344 6817
rect 18236 6944 18288 6996
rect 18788 6987 18840 6996
rect 18788 6953 18797 6987
rect 18797 6953 18831 6987
rect 18831 6953 18840 6987
rect 18788 6944 18840 6953
rect 17684 6876 17736 6928
rect 20536 6876 20588 6928
rect 21456 6876 21508 6928
rect 15936 6808 15988 6860
rect 16488 6851 16540 6860
rect 16488 6817 16497 6851
rect 16497 6817 16531 6851
rect 16531 6817 16540 6851
rect 16488 6808 16540 6817
rect 19708 6851 19760 6860
rect 19708 6817 19717 6851
rect 19717 6817 19751 6851
rect 19751 6817 19760 6851
rect 19708 6808 19760 6817
rect 6644 6783 6696 6792
rect 6644 6749 6653 6783
rect 6653 6749 6687 6783
rect 6687 6749 6696 6783
rect 6644 6740 6696 6749
rect 7012 6783 7064 6792
rect 7012 6749 7021 6783
rect 7021 6749 7055 6783
rect 7055 6749 7064 6783
rect 7012 6740 7064 6749
rect 11060 6740 11112 6792
rect 12256 6783 12308 6792
rect 12256 6749 12265 6783
rect 12265 6749 12299 6783
rect 12299 6749 12308 6783
rect 12256 6740 12308 6749
rect 16764 6783 16816 6792
rect 16764 6749 16773 6783
rect 16773 6749 16807 6783
rect 16807 6749 16816 6783
rect 16764 6740 16816 6749
rect 21272 6783 21324 6792
rect 21272 6749 21281 6783
rect 21281 6749 21315 6783
rect 21315 6749 21324 6783
rect 21272 6740 21324 6749
rect 10784 6715 10836 6724
rect 10784 6681 10793 6715
rect 10793 6681 10827 6715
rect 10827 6681 10836 6715
rect 10784 6672 10836 6681
rect 12900 6672 12952 6724
rect 14556 6672 14608 6724
rect 19524 6672 19576 6724
rect 3516 6647 3568 6656
rect 3516 6613 3525 6647
rect 3525 6613 3559 6647
rect 3559 6613 3568 6647
rect 3516 6604 3568 6613
rect 5356 6604 5408 6656
rect 14188 6647 14240 6656
rect 14188 6613 14197 6647
rect 14197 6613 14231 6647
rect 14231 6613 14240 6647
rect 14188 6604 14240 6613
rect 16396 6604 16448 6656
rect 4982 6502 5034 6554
rect 5046 6502 5098 6554
rect 5110 6502 5162 6554
rect 5174 6502 5226 6554
rect 12982 6502 13034 6554
rect 13046 6502 13098 6554
rect 13110 6502 13162 6554
rect 13174 6502 13226 6554
rect 20982 6502 21034 6554
rect 21046 6502 21098 6554
rect 21110 6502 21162 6554
rect 21174 6502 21226 6554
rect 3608 6400 3660 6452
rect 4528 6400 4580 6452
rect 4712 6400 4764 6452
rect 4804 6332 4856 6384
rect 2872 6307 2924 6316
rect 2872 6273 2881 6307
rect 2881 6273 2915 6307
rect 2915 6273 2924 6307
rect 2872 6264 2924 6273
rect 2136 6196 2188 6248
rect 2688 6128 2740 6180
rect 6552 6332 6604 6384
rect 8668 6443 8720 6452
rect 8668 6409 8677 6443
rect 8677 6409 8711 6443
rect 8711 6409 8720 6443
rect 8668 6400 8720 6409
rect 8760 6400 8812 6452
rect 10324 6400 10376 6452
rect 11060 6443 11112 6452
rect 11060 6409 11069 6443
rect 11069 6409 11103 6443
rect 11103 6409 11112 6443
rect 11060 6400 11112 6409
rect 12348 6400 12400 6452
rect 14004 6400 14056 6452
rect 15752 6400 15804 6452
rect 16764 6443 16816 6452
rect 16764 6409 16773 6443
rect 16773 6409 16807 6443
rect 16807 6409 16816 6443
rect 16764 6400 16816 6409
rect 17684 6400 17736 6452
rect 18420 6400 18472 6452
rect 19064 6443 19116 6452
rect 19064 6409 19073 6443
rect 19073 6409 19107 6443
rect 19107 6409 19116 6443
rect 19064 6400 19116 6409
rect 20536 6400 20588 6452
rect 14832 6332 14884 6384
rect 16488 6332 16540 6384
rect 19708 6332 19760 6384
rect 21364 6332 21416 6384
rect 21456 6375 21508 6384
rect 21456 6341 21465 6375
rect 21465 6341 21499 6375
rect 21499 6341 21508 6375
rect 21456 6332 21508 6341
rect 5356 6264 5408 6316
rect 5632 6264 5684 6316
rect 10784 6307 10836 6316
rect 10784 6273 10793 6307
rect 10793 6273 10827 6307
rect 10827 6273 10836 6307
rect 10784 6264 10836 6273
rect 10968 6264 11020 6316
rect 13544 6264 13596 6316
rect 13636 6264 13688 6316
rect 6920 6196 6972 6248
rect 7104 6239 7156 6248
rect 7104 6205 7113 6239
rect 7113 6205 7147 6239
rect 7147 6205 7156 6239
rect 7104 6196 7156 6205
rect 8024 6196 8076 6248
rect 7564 6128 7616 6180
rect 14188 6196 14240 6248
rect 15936 6264 15988 6316
rect 16764 6264 16816 6316
rect 20536 6307 20588 6316
rect 20536 6273 20545 6307
rect 20545 6273 20579 6307
rect 20579 6273 20588 6307
rect 20536 6264 20588 6273
rect 21272 6264 21324 6316
rect 10140 6171 10192 6180
rect 10140 6137 10149 6171
rect 10149 6137 10183 6171
rect 10183 6137 10192 6171
rect 10140 6128 10192 6137
rect 10232 6171 10284 6180
rect 10232 6137 10241 6171
rect 10241 6137 10275 6171
rect 10275 6137 10284 6171
rect 12624 6171 12676 6180
rect 10232 6128 10284 6137
rect 12624 6137 12633 6171
rect 12633 6137 12667 6171
rect 12667 6137 12676 6171
rect 12624 6128 12676 6137
rect 1676 6103 1728 6112
rect 1676 6069 1685 6103
rect 1685 6069 1719 6103
rect 1719 6069 1728 6103
rect 1676 6060 1728 6069
rect 2412 6103 2464 6112
rect 2412 6069 2421 6103
rect 2421 6069 2455 6103
rect 2455 6069 2464 6103
rect 2412 6060 2464 6069
rect 5448 6060 5500 6112
rect 6368 6060 6420 6112
rect 7104 6060 7156 6112
rect 8208 6103 8260 6112
rect 8208 6069 8217 6103
rect 8217 6069 8251 6103
rect 8251 6069 8260 6103
rect 8208 6060 8260 6069
rect 12348 6060 12400 6112
rect 14004 6103 14056 6112
rect 14004 6069 14013 6103
rect 14013 6069 14047 6103
rect 14047 6069 14056 6103
rect 15844 6196 15896 6248
rect 16580 6196 16632 6248
rect 19064 6196 19116 6248
rect 15292 6103 15344 6112
rect 14004 6060 14056 6069
rect 15292 6069 15301 6103
rect 15301 6069 15335 6103
rect 15335 6069 15344 6103
rect 15292 6060 15344 6069
rect 17316 6060 17368 6112
rect 20628 6171 20680 6180
rect 20628 6137 20637 6171
rect 20637 6137 20671 6171
rect 20671 6137 20680 6171
rect 20628 6128 20680 6137
rect 20812 6128 20864 6180
rect 21272 6128 21324 6180
rect 23480 6060 23532 6112
rect 8982 5958 9034 6010
rect 9046 5958 9098 6010
rect 9110 5958 9162 6010
rect 9174 5958 9226 6010
rect 16982 5958 17034 6010
rect 17046 5958 17098 6010
rect 17110 5958 17162 6010
rect 17174 5958 17226 6010
rect 5356 5856 5408 5908
rect 1860 5831 1912 5840
rect 1860 5797 1863 5831
rect 1863 5797 1897 5831
rect 1897 5797 1912 5831
rect 1860 5788 1912 5797
rect 2872 5788 2924 5840
rect 2412 5763 2464 5772
rect 2412 5729 2421 5763
rect 2421 5729 2455 5763
rect 2455 5729 2464 5763
rect 2412 5720 2464 5729
rect 3608 5720 3660 5772
rect 4528 5720 4580 5772
rect 4712 5763 4764 5772
rect 4712 5729 4721 5763
rect 4721 5729 4755 5763
rect 4755 5729 4764 5763
rect 4712 5720 4764 5729
rect 5724 5720 5776 5772
rect 6184 5720 6236 5772
rect 10232 5856 10284 5908
rect 12256 5899 12308 5908
rect 12256 5865 12265 5899
rect 12265 5865 12299 5899
rect 12299 5865 12308 5899
rect 12256 5856 12308 5865
rect 17316 5856 17368 5908
rect 20536 5899 20588 5908
rect 10324 5788 10376 5840
rect 10968 5831 11020 5840
rect 10968 5797 10977 5831
rect 10977 5797 11011 5831
rect 11011 5797 11020 5831
rect 10968 5788 11020 5797
rect 17684 5831 17736 5840
rect 17684 5797 17693 5831
rect 17693 5797 17727 5831
rect 17727 5797 17736 5831
rect 17684 5788 17736 5797
rect 20536 5865 20545 5899
rect 20545 5865 20579 5899
rect 20579 5865 20588 5899
rect 20536 5856 20588 5865
rect 19432 5831 19484 5840
rect 19432 5797 19441 5831
rect 19441 5797 19475 5831
rect 19475 5797 19484 5831
rect 21456 5856 21508 5908
rect 19432 5788 19484 5797
rect 20812 5788 20864 5840
rect 6828 5720 6880 5772
rect 8116 5763 8168 5772
rect 8116 5729 8125 5763
rect 8125 5729 8159 5763
rect 8159 5729 8168 5763
rect 8116 5720 8168 5729
rect 15108 5720 15160 5772
rect 16488 5720 16540 5772
rect 5632 5652 5684 5704
rect 6920 5652 6972 5704
rect 8760 5652 8812 5704
rect 10324 5695 10376 5704
rect 10324 5661 10333 5695
rect 10333 5661 10367 5695
rect 10367 5661 10376 5695
rect 10324 5652 10376 5661
rect 21272 5695 21324 5704
rect 4528 5584 4580 5636
rect 6368 5584 6420 5636
rect 6552 5627 6604 5636
rect 6552 5593 6561 5627
rect 6561 5593 6595 5627
rect 6595 5593 6604 5627
rect 6552 5584 6604 5593
rect 14188 5584 14240 5636
rect 16120 5584 16172 5636
rect 4436 5516 4488 5568
rect 7012 5516 7064 5568
rect 7564 5559 7616 5568
rect 7564 5525 7573 5559
rect 7573 5525 7607 5559
rect 7607 5525 7616 5559
rect 7564 5516 7616 5525
rect 12624 5559 12676 5568
rect 12624 5525 12633 5559
rect 12633 5525 12667 5559
rect 12667 5525 12676 5559
rect 12624 5516 12676 5525
rect 15016 5516 15068 5568
rect 15660 5559 15712 5568
rect 15660 5525 15669 5559
rect 15669 5525 15703 5559
rect 15703 5525 15712 5559
rect 15660 5516 15712 5525
rect 16672 5516 16724 5568
rect 17316 5559 17368 5568
rect 17316 5525 17325 5559
rect 17325 5525 17359 5559
rect 17359 5525 17368 5559
rect 18880 5584 18932 5636
rect 19432 5584 19484 5636
rect 19892 5627 19944 5636
rect 19892 5593 19901 5627
rect 19901 5593 19935 5627
rect 19935 5593 19944 5627
rect 21272 5661 21281 5695
rect 21281 5661 21315 5695
rect 21315 5661 21324 5695
rect 21272 5652 21324 5661
rect 19892 5584 19944 5593
rect 21456 5584 21508 5636
rect 17316 5516 17368 5525
rect 4982 5414 5034 5466
rect 5046 5414 5098 5466
rect 5110 5414 5162 5466
rect 5174 5414 5226 5466
rect 12982 5414 13034 5466
rect 13046 5414 13098 5466
rect 13110 5414 13162 5466
rect 13174 5414 13226 5466
rect 20982 5414 21034 5466
rect 21046 5414 21098 5466
rect 21110 5414 21162 5466
rect 21174 5414 21226 5466
rect 2872 5355 2924 5364
rect 2872 5321 2881 5355
rect 2881 5321 2915 5355
rect 2915 5321 2924 5355
rect 2872 5312 2924 5321
rect 5448 5312 5500 5364
rect 6552 5355 6604 5364
rect 6552 5321 6561 5355
rect 6561 5321 6595 5355
rect 6595 5321 6604 5355
rect 6552 5312 6604 5321
rect 7748 5355 7800 5364
rect 7748 5321 7757 5355
rect 7757 5321 7791 5355
rect 7791 5321 7800 5355
rect 10232 5355 10284 5364
rect 7748 5312 7800 5321
rect 10232 5321 10241 5355
rect 10241 5321 10275 5355
rect 10275 5321 10284 5355
rect 10232 5312 10284 5321
rect 10600 5355 10652 5364
rect 10600 5321 10609 5355
rect 10609 5321 10643 5355
rect 10643 5321 10652 5355
rect 10600 5312 10652 5321
rect 17684 5312 17736 5364
rect 21364 5312 21416 5364
rect 21456 5312 21508 5364
rect 1768 5244 1820 5296
rect 10140 5244 10192 5296
rect 20812 5244 20864 5296
rect 20996 5244 21048 5296
rect 21916 5287 21968 5296
rect 21916 5253 21925 5287
rect 21925 5253 21959 5287
rect 21959 5253 21968 5287
rect 21916 5244 21968 5253
rect 2136 5219 2188 5228
rect 2136 5185 2145 5219
rect 2145 5185 2179 5219
rect 2179 5185 2188 5219
rect 2136 5176 2188 5185
rect 3608 5108 3660 5160
rect 4620 5108 4672 5160
rect 5632 5176 5684 5228
rect 6736 5176 6788 5228
rect 7564 5176 7616 5228
rect 14740 5219 14792 5228
rect 14740 5185 14749 5219
rect 14749 5185 14783 5219
rect 14783 5185 14792 5219
rect 14740 5176 14792 5185
rect 16764 5176 16816 5228
rect 20536 5219 20588 5228
rect 1492 5083 1544 5092
rect 1492 5049 1501 5083
rect 1501 5049 1535 5083
rect 1535 5049 1544 5083
rect 1492 5040 1544 5049
rect 1676 5040 1728 5092
rect 2688 5040 2740 5092
rect 6184 5108 6236 5160
rect 7104 5151 7156 5160
rect 7104 5117 7113 5151
rect 7113 5117 7147 5151
rect 7147 5117 7156 5151
rect 7104 5108 7156 5117
rect 7472 5108 7524 5160
rect 9496 5108 9548 5160
rect 10600 5108 10652 5160
rect 12716 5151 12768 5160
rect 12716 5117 12725 5151
rect 12725 5117 12759 5151
rect 12759 5117 12768 5151
rect 12716 5108 12768 5117
rect 14004 5108 14056 5160
rect 15568 5151 15620 5160
rect 15568 5117 15577 5151
rect 15577 5117 15611 5151
rect 15611 5117 15620 5151
rect 15568 5108 15620 5117
rect 15660 5108 15712 5160
rect 16028 5151 16080 5160
rect 16028 5117 16037 5151
rect 16037 5117 16071 5151
rect 16071 5117 16080 5151
rect 16028 5108 16080 5117
rect 16120 5108 16172 5160
rect 16396 5151 16448 5160
rect 16396 5117 16405 5151
rect 16405 5117 16439 5151
rect 16439 5117 16448 5151
rect 16396 5108 16448 5117
rect 20536 5185 20545 5219
rect 20545 5185 20579 5219
rect 20579 5185 20588 5219
rect 20536 5176 20588 5185
rect 18052 5151 18104 5160
rect 18052 5117 18061 5151
rect 18061 5117 18095 5151
rect 18095 5117 18104 5151
rect 18052 5108 18104 5117
rect 7748 5040 7800 5092
rect 8576 5040 8628 5092
rect 10324 5040 10376 5092
rect 10784 5083 10836 5092
rect 10784 5049 10793 5083
rect 10793 5049 10827 5083
rect 10827 5049 10836 5083
rect 10784 5040 10836 5049
rect 12440 5083 12492 5092
rect 12440 5049 12449 5083
rect 12449 5049 12483 5083
rect 12483 5049 12492 5083
rect 12440 5040 12492 5049
rect 13268 5040 13320 5092
rect 13728 5040 13780 5092
rect 16488 5040 16540 5092
rect 18236 5040 18288 5092
rect 3792 5015 3844 5024
rect 3792 4981 3801 5015
rect 3801 4981 3835 5015
rect 3835 4981 3844 5015
rect 3792 4972 3844 4981
rect 7104 4972 7156 5024
rect 7472 4972 7524 5024
rect 7932 4972 7984 5024
rect 8116 4972 8168 5024
rect 15108 5015 15160 5024
rect 15108 4981 15117 5015
rect 15117 4981 15151 5015
rect 15151 4981 15160 5015
rect 15108 4972 15160 4981
rect 16212 4972 16264 5024
rect 16764 4972 16816 5024
rect 17684 4972 17736 5024
rect 19340 5015 19392 5024
rect 19340 4981 19349 5015
rect 19349 4981 19383 5015
rect 19383 4981 19392 5015
rect 19708 5015 19760 5024
rect 19340 4972 19392 4981
rect 19708 4981 19717 5015
rect 19717 4981 19751 5015
rect 19751 4981 19760 5015
rect 19708 4972 19760 4981
rect 21272 4972 21324 5024
rect 8982 4870 9034 4922
rect 9046 4870 9098 4922
rect 9110 4870 9162 4922
rect 9174 4870 9226 4922
rect 16982 4870 17034 4922
rect 17046 4870 17098 4922
rect 17110 4870 17162 4922
rect 17174 4870 17226 4922
rect 1216 4768 1268 4820
rect 1860 4768 1912 4820
rect 2412 4768 2464 4820
rect 5724 4768 5776 4820
rect 6184 4811 6236 4820
rect 6184 4777 6193 4811
rect 6193 4777 6227 4811
rect 6227 4777 6236 4811
rect 6184 4768 6236 4777
rect 7288 4768 7340 4820
rect 7564 4768 7616 4820
rect 9680 4768 9732 4820
rect 11888 4768 11940 4820
rect 4344 4700 4396 4752
rect 6828 4700 6880 4752
rect 13820 4768 13872 4820
rect 14740 4768 14792 4820
rect 17684 4768 17736 4820
rect 18052 4768 18104 4820
rect 6460 4632 6512 4684
rect 8300 4632 8352 4684
rect 9404 4632 9456 4684
rect 10416 4675 10468 4684
rect 10416 4641 10425 4675
rect 10425 4641 10459 4675
rect 10459 4641 10468 4675
rect 10416 4632 10468 4641
rect 10692 4675 10744 4684
rect 10692 4641 10701 4675
rect 10701 4641 10735 4675
rect 10735 4641 10744 4675
rect 10692 4632 10744 4641
rect 1952 4564 2004 4616
rect 2136 4607 2188 4616
rect 2136 4573 2145 4607
rect 2145 4573 2179 4607
rect 2179 4573 2188 4607
rect 2136 4564 2188 4573
rect 4528 4564 4580 4616
rect 4712 4607 4764 4616
rect 4712 4573 4721 4607
rect 4721 4573 4755 4607
rect 4755 4573 4764 4607
rect 4712 4564 4764 4573
rect 6736 4607 6788 4616
rect 6736 4573 6745 4607
rect 6745 4573 6779 4607
rect 6779 4573 6788 4607
rect 6736 4564 6788 4573
rect 7380 4607 7432 4616
rect 7380 4573 7389 4607
rect 7389 4573 7423 4607
rect 7423 4573 7432 4607
rect 7380 4564 7432 4573
rect 5724 4496 5776 4548
rect 10784 4564 10836 4616
rect 8208 4496 8260 4548
rect 12256 4675 12308 4684
rect 12256 4641 12265 4675
rect 12265 4641 12299 4675
rect 12299 4641 12308 4675
rect 13268 4700 13320 4752
rect 16304 4700 16356 4752
rect 12256 4632 12308 4641
rect 13176 4675 13228 4684
rect 11612 4564 11664 4616
rect 13176 4641 13185 4675
rect 13185 4641 13219 4675
rect 13219 4641 13228 4675
rect 13176 4632 13228 4641
rect 15568 4632 15620 4684
rect 16028 4675 16080 4684
rect 14188 4564 14240 4616
rect 14372 4564 14424 4616
rect 16028 4641 16037 4675
rect 16037 4641 16071 4675
rect 16071 4641 16080 4675
rect 16028 4632 16080 4641
rect 16396 4675 16448 4684
rect 16396 4641 16405 4675
rect 16405 4641 16439 4675
rect 16439 4641 16448 4675
rect 16396 4632 16448 4641
rect 17316 4700 17368 4752
rect 19708 4700 19760 4752
rect 19892 4743 19944 4752
rect 19892 4709 19901 4743
rect 19901 4709 19935 4743
rect 19935 4709 19944 4743
rect 19892 4700 19944 4709
rect 20628 4700 20680 4752
rect 18328 4632 18380 4684
rect 18696 4632 18748 4684
rect 20996 4675 21048 4684
rect 20996 4641 21005 4675
rect 21005 4641 21039 4675
rect 21039 4641 21048 4675
rect 20996 4632 21048 4641
rect 16212 4564 16264 4616
rect 19248 4607 19300 4616
rect 19248 4573 19257 4607
rect 19257 4573 19291 4607
rect 19291 4573 19300 4607
rect 19248 4564 19300 4573
rect 13176 4496 13228 4548
rect 3608 4428 3660 4480
rect 8116 4428 8168 4480
rect 14096 4428 14148 4480
rect 4982 4326 5034 4378
rect 5046 4326 5098 4378
rect 5110 4326 5162 4378
rect 5174 4326 5226 4378
rect 12982 4326 13034 4378
rect 13046 4326 13098 4378
rect 13110 4326 13162 4378
rect 13174 4326 13226 4378
rect 20982 4326 21034 4378
rect 21046 4326 21098 4378
rect 21110 4326 21162 4378
rect 21174 4326 21226 4378
rect 2412 4224 2464 4276
rect 4528 4224 4580 4276
rect 6828 4224 6880 4276
rect 7288 4224 7340 4276
rect 7472 4267 7524 4276
rect 7472 4233 7481 4267
rect 7481 4233 7515 4267
rect 7515 4233 7524 4267
rect 7472 4224 7524 4233
rect 8760 4224 8812 4276
rect 1860 4156 1912 4208
rect 7748 4199 7800 4208
rect 7748 4165 7757 4199
rect 7757 4165 7791 4199
rect 7791 4165 7800 4199
rect 7748 4156 7800 4165
rect 1952 4088 2004 4140
rect 4712 4088 4764 4140
rect 3792 4020 3844 4072
rect 5540 4020 5592 4072
rect 7288 4020 7340 4072
rect 9404 4156 9456 4208
rect 10784 4224 10836 4276
rect 16396 4224 16448 4276
rect 18328 4267 18380 4276
rect 18328 4233 18337 4267
rect 18337 4233 18371 4267
rect 18371 4233 18380 4267
rect 18328 4224 18380 4233
rect 18880 4267 18932 4276
rect 18880 4233 18889 4267
rect 18889 4233 18923 4267
rect 18923 4233 18932 4267
rect 18880 4224 18932 4233
rect 20812 4224 20864 4276
rect 10692 4156 10744 4208
rect 8208 4020 8260 4072
rect 9588 4088 9640 4140
rect 11612 4131 11664 4140
rect 8760 4063 8812 4072
rect 8760 4029 8769 4063
rect 8769 4029 8803 4063
rect 8803 4029 8812 4063
rect 8760 4020 8812 4029
rect 9496 4020 9548 4072
rect 11612 4097 11621 4131
rect 11621 4097 11655 4131
rect 11655 4097 11664 4131
rect 11612 4088 11664 4097
rect 10600 4063 10652 4072
rect 1492 3952 1544 4004
rect 6552 3952 6604 4004
rect 7380 3952 7432 4004
rect 10600 4029 10609 4063
rect 10609 4029 10643 4063
rect 10643 4029 10652 4063
rect 10600 4020 10652 4029
rect 13360 4020 13412 4072
rect 13820 4063 13872 4072
rect 13820 4029 13829 4063
rect 13829 4029 13863 4063
rect 13863 4029 13872 4063
rect 13820 4020 13872 4029
rect 14372 4063 14424 4072
rect 9772 3952 9824 4004
rect 4344 3884 4396 3936
rect 4804 3927 4856 3936
rect 4804 3893 4813 3927
rect 4813 3893 4847 3927
rect 4847 3893 4856 3927
rect 4804 3884 4856 3893
rect 7288 3884 7340 3936
rect 8024 3927 8076 3936
rect 8024 3893 8033 3927
rect 8033 3893 8067 3927
rect 8067 3893 8076 3927
rect 8024 3884 8076 3893
rect 9588 3884 9640 3936
rect 10416 3884 10468 3936
rect 13268 3952 13320 4004
rect 14372 4029 14381 4063
rect 14381 4029 14415 4063
rect 14415 4029 14424 4063
rect 14372 4020 14424 4029
rect 16304 4156 16356 4208
rect 16580 4088 16632 4140
rect 18880 4020 18932 4072
rect 12072 3884 12124 3936
rect 14740 3927 14792 3936
rect 14740 3893 14749 3927
rect 14749 3893 14783 3927
rect 14783 3893 14792 3927
rect 14740 3884 14792 3893
rect 16396 3952 16448 4004
rect 16580 3995 16632 4004
rect 16580 3961 16589 3995
rect 16589 3961 16623 3995
rect 16623 3961 16632 3995
rect 16580 3952 16632 3961
rect 19708 3995 19760 4004
rect 19708 3961 19717 3995
rect 19717 3961 19751 3995
rect 19751 3961 19760 3995
rect 19708 3952 19760 3961
rect 16120 3884 16172 3936
rect 17316 3884 17368 3936
rect 8982 3782 9034 3834
rect 9046 3782 9098 3834
rect 9110 3782 9162 3834
rect 9174 3782 9226 3834
rect 16982 3782 17034 3834
rect 17046 3782 17098 3834
rect 17110 3782 17162 3834
rect 17174 3782 17226 3834
rect 6736 3723 6788 3732
rect 6736 3689 6745 3723
rect 6745 3689 6779 3723
rect 6779 3689 6788 3723
rect 6736 3680 6788 3689
rect 8760 3680 8812 3732
rect 9404 3723 9456 3732
rect 9404 3689 9413 3723
rect 9413 3689 9447 3723
rect 9447 3689 9456 3723
rect 9404 3680 9456 3689
rect 12256 3680 12308 3732
rect 12716 3723 12768 3732
rect 12716 3689 12725 3723
rect 12725 3689 12759 3723
rect 12759 3689 12768 3723
rect 12716 3680 12768 3689
rect 13360 3723 13412 3732
rect 13360 3689 13369 3723
rect 13369 3689 13403 3723
rect 13403 3689 13412 3723
rect 13360 3680 13412 3689
rect 14740 3723 14792 3732
rect 14740 3689 14749 3723
rect 14749 3689 14783 3723
rect 14783 3689 14792 3723
rect 14740 3680 14792 3689
rect 15016 3723 15068 3732
rect 15016 3689 15025 3723
rect 15025 3689 15059 3723
rect 15059 3689 15068 3723
rect 15016 3680 15068 3689
rect 16212 3680 16264 3732
rect 16396 3680 16448 3732
rect 17500 3680 17552 3732
rect 19248 3723 19300 3732
rect 19248 3689 19257 3723
rect 19257 3689 19291 3723
rect 19291 3689 19300 3723
rect 19248 3680 19300 3689
rect 19340 3680 19392 3732
rect 20260 3680 20312 3732
rect 7380 3655 7432 3664
rect 7380 3621 7389 3655
rect 7389 3621 7423 3655
rect 7423 3621 7432 3655
rect 7380 3612 7432 3621
rect 7748 3612 7800 3664
rect 9496 3612 9548 3664
rect 9956 3655 10008 3664
rect 9956 3621 9965 3655
rect 9965 3621 9999 3655
rect 9999 3621 10008 3655
rect 9956 3612 10008 3621
rect 11796 3612 11848 3664
rect 15476 3655 15528 3664
rect 15476 3621 15485 3655
rect 15485 3621 15519 3655
rect 15519 3621 15528 3655
rect 15476 3612 15528 3621
rect 4804 3587 4856 3596
rect 4804 3553 4813 3587
rect 4813 3553 4847 3587
rect 4847 3553 4856 3587
rect 4804 3544 4856 3553
rect 5816 3544 5868 3596
rect 8300 3587 8352 3596
rect 8300 3553 8309 3587
rect 8309 3553 8343 3587
rect 8343 3553 8352 3587
rect 8300 3544 8352 3553
rect 13452 3544 13504 3596
rect 14280 3587 14332 3596
rect 14280 3553 14289 3587
rect 14289 3553 14323 3587
rect 14323 3553 14332 3587
rect 14280 3544 14332 3553
rect 16856 3587 16908 3596
rect 16856 3553 16865 3587
rect 16865 3553 16899 3587
rect 16899 3553 16908 3587
rect 16856 3544 16908 3553
rect 18236 3544 18288 3596
rect 18604 3544 18656 3596
rect 21456 3544 21508 3596
rect 7288 3519 7340 3528
rect 7288 3485 7297 3519
rect 7297 3485 7331 3519
rect 7331 3485 7340 3519
rect 7288 3476 7340 3485
rect 9680 3519 9732 3528
rect 9680 3485 9689 3519
rect 9689 3485 9723 3519
rect 9723 3485 9732 3519
rect 9680 3476 9732 3485
rect 11888 3476 11940 3528
rect 15660 3476 15712 3528
rect 7840 3451 7892 3460
rect 7840 3417 7849 3451
rect 7849 3417 7883 3451
rect 7883 3417 7892 3451
rect 7840 3408 7892 3417
rect 12624 3408 12676 3460
rect 15568 3408 15620 3460
rect 15936 3451 15988 3460
rect 15936 3417 15945 3451
rect 15945 3417 15979 3451
rect 15979 3417 15988 3451
rect 15936 3408 15988 3417
rect 16028 3408 16080 3460
rect 4436 3383 4488 3392
rect 4436 3349 4445 3383
rect 4445 3349 4479 3383
rect 4479 3349 4488 3383
rect 4436 3340 4488 3349
rect 4528 3340 4580 3392
rect 6184 3340 6236 3392
rect 6460 3340 6512 3392
rect 10600 3383 10652 3392
rect 10600 3349 10609 3383
rect 10609 3349 10643 3383
rect 10643 3349 10652 3383
rect 10600 3340 10652 3349
rect 11152 3340 11204 3392
rect 4982 3238 5034 3290
rect 5046 3238 5098 3290
rect 5110 3238 5162 3290
rect 5174 3238 5226 3290
rect 12982 3238 13034 3290
rect 13046 3238 13098 3290
rect 13110 3238 13162 3290
rect 13174 3238 13226 3290
rect 20982 3238 21034 3290
rect 21046 3238 21098 3290
rect 21110 3238 21162 3290
rect 21174 3238 21226 3290
rect 1584 3179 1636 3188
rect 1584 3145 1593 3179
rect 1593 3145 1627 3179
rect 1627 3145 1636 3179
rect 1584 3136 1636 3145
rect 4252 3136 4304 3188
rect 4436 3136 4488 3188
rect 6552 3179 6604 3188
rect 6552 3145 6561 3179
rect 6561 3145 6595 3179
rect 6595 3145 6604 3179
rect 6552 3136 6604 3145
rect 7288 3136 7340 3188
rect 9680 3136 9732 3188
rect 14280 3136 14332 3188
rect 15476 3136 15528 3188
rect 15660 3179 15712 3188
rect 15660 3145 15669 3179
rect 15669 3145 15703 3179
rect 15703 3145 15712 3179
rect 15660 3136 15712 3145
rect 16856 3179 16908 3188
rect 16856 3145 16865 3179
rect 16865 3145 16899 3179
rect 16899 3145 16908 3179
rect 16856 3136 16908 3145
rect 19248 3136 19300 3188
rect 20812 3136 20864 3188
rect 21456 3179 21508 3188
rect 21456 3145 21465 3179
rect 21465 3145 21499 3179
rect 21499 3145 21508 3179
rect 21456 3136 21508 3145
rect 8484 3068 8536 3120
rect 9588 3068 9640 3120
rect 14464 3068 14516 3120
rect 17684 3068 17736 3120
rect 4528 3043 4580 3052
rect 4528 3009 4537 3043
rect 4537 3009 4571 3043
rect 4571 3009 4580 3043
rect 4528 3000 4580 3009
rect 4712 3000 4764 3052
rect 8024 3000 8076 3052
rect 12624 3043 12676 3052
rect 12624 3009 12633 3043
rect 12633 3009 12667 3043
rect 12667 3009 12676 3043
rect 12624 3000 12676 3009
rect 13360 3000 13412 3052
rect 14740 3000 14792 3052
rect 15568 3000 15620 3052
rect 16580 3000 16632 3052
rect 4252 2932 4304 2984
rect 6552 2932 6604 2984
rect 7380 2932 7432 2984
rect 11152 2975 11204 2984
rect 11152 2941 11161 2975
rect 11161 2941 11195 2975
rect 11195 2941 11204 2975
rect 11152 2932 11204 2941
rect 19248 2932 19300 2984
rect 2044 2839 2096 2848
rect 2044 2805 2053 2839
rect 2053 2805 2087 2839
rect 2087 2805 2096 2839
rect 2044 2796 2096 2805
rect 4436 2796 4488 2848
rect 6644 2864 6696 2916
rect 9772 2907 9824 2916
rect 5816 2839 5868 2848
rect 5816 2805 5825 2839
rect 5825 2805 5859 2839
rect 5859 2805 5868 2839
rect 5816 2796 5868 2805
rect 9772 2873 9781 2907
rect 9781 2873 9815 2907
rect 9815 2873 9824 2907
rect 9772 2864 9824 2873
rect 10324 2907 10376 2916
rect 10324 2873 10333 2907
rect 10333 2873 10367 2907
rect 10367 2873 10376 2907
rect 10324 2864 10376 2873
rect 12716 2907 12768 2916
rect 12716 2873 12725 2907
rect 12725 2873 12759 2907
rect 12759 2873 12768 2907
rect 12716 2864 12768 2873
rect 14924 2864 14976 2916
rect 15752 2864 15804 2916
rect 9956 2796 10008 2848
rect 11796 2839 11848 2848
rect 11796 2805 11805 2839
rect 11805 2805 11839 2839
rect 11839 2805 11848 2839
rect 11796 2796 11848 2805
rect 14464 2839 14516 2848
rect 14464 2805 14473 2839
rect 14473 2805 14507 2839
rect 14507 2805 14516 2839
rect 14464 2796 14516 2805
rect 15660 2796 15712 2848
rect 18052 2839 18104 2848
rect 18052 2805 18061 2839
rect 18061 2805 18095 2839
rect 18095 2805 18104 2839
rect 18052 2796 18104 2805
rect 18604 2839 18656 2848
rect 18604 2805 18613 2839
rect 18613 2805 18647 2839
rect 18647 2805 18656 2839
rect 18604 2796 18656 2805
rect 22284 2796 22336 2848
rect 8982 2694 9034 2746
rect 9046 2694 9098 2746
rect 9110 2694 9162 2746
rect 9174 2694 9226 2746
rect 16982 2694 17034 2746
rect 17046 2694 17098 2746
rect 17110 2694 17162 2746
rect 17174 2694 17226 2746
rect 1768 2592 1820 2644
rect 3516 2592 3568 2644
rect 11152 2592 11204 2644
rect 11888 2635 11940 2644
rect 11888 2601 11897 2635
rect 11897 2601 11931 2635
rect 11931 2601 11940 2635
rect 11888 2592 11940 2601
rect 12440 2635 12492 2644
rect 12440 2601 12449 2635
rect 12449 2601 12483 2635
rect 12483 2601 12492 2635
rect 12440 2592 12492 2601
rect 6184 2524 6236 2576
rect 1124 2456 1176 2508
rect 848 2252 900 2304
rect 6552 2456 6604 2508
rect 7840 2567 7892 2576
rect 7840 2533 7849 2567
rect 7849 2533 7883 2567
rect 7883 2533 7892 2567
rect 7840 2524 7892 2533
rect 8116 2388 8168 2440
rect 10600 2524 10652 2576
rect 12072 2524 12124 2576
rect 13268 2592 13320 2644
rect 15752 2592 15804 2644
rect 19800 2592 19852 2644
rect 13360 2567 13412 2576
rect 13360 2533 13369 2567
rect 13369 2533 13403 2567
rect 13403 2533 13412 2567
rect 13360 2524 13412 2533
rect 15660 2567 15712 2576
rect 15660 2533 15680 2567
rect 15680 2533 15712 2567
rect 15660 2524 15712 2533
rect 14096 2499 14148 2508
rect 14096 2465 14105 2499
rect 14105 2465 14139 2499
rect 14139 2465 14148 2499
rect 14096 2456 14148 2465
rect 16672 2456 16724 2508
rect 10324 2431 10376 2440
rect 10324 2397 10333 2431
rect 10333 2397 10367 2431
rect 10367 2397 10376 2431
rect 10324 2388 10376 2397
rect 10508 2320 10560 2372
rect 18052 2388 18104 2440
rect 18604 2388 18656 2440
rect 19616 2388 19668 2440
rect 15936 2320 15988 2372
rect 20444 2320 20496 2372
rect 4804 2252 4856 2304
rect 16948 2252 17000 2304
rect 18236 2252 18288 2304
rect 18972 2252 19024 2304
rect 23204 2252 23256 2304
rect 4982 2150 5034 2202
rect 5046 2150 5098 2202
rect 5110 2150 5162 2202
rect 5174 2150 5226 2202
rect 12982 2150 13034 2202
rect 13046 2150 13098 2202
rect 13110 2150 13162 2202
rect 13174 2150 13226 2202
rect 20982 2150 21034 2202
rect 21046 2150 21098 2202
rect 21110 2150 21162 2202
rect 21174 2150 21226 2202
rect 5816 2048 5868 2100
rect 12164 2048 12216 2100
rect 11520 76 11572 128
rect 13268 76 13320 128
<< metal2 >>
rect 20 23588 72 23594
rect 20 23530 72 23536
rect 570 23588 626 24000
rect 1766 23610 1822 24000
rect 3054 23610 3110 24000
rect 570 23536 572 23588
rect 624 23536 626 23588
rect 32 12918 60 23530
rect 570 23520 626 23536
rect 1688 23582 1822 23610
rect 584 23499 612 23520
rect 1306 22536 1362 22545
rect 1306 22471 1362 22480
rect 1320 18834 1348 22471
rect 1582 20768 1638 20777
rect 1582 20703 1638 20712
rect 1596 19922 1624 20703
rect 1584 19916 1636 19922
rect 1584 19858 1636 19864
rect 1596 19514 1624 19858
rect 1584 19508 1636 19514
rect 1584 19450 1636 19456
rect 1308 18828 1360 18834
rect 1308 18770 1360 18776
rect 1320 18426 1348 18770
rect 1308 18420 1360 18426
rect 1308 18362 1360 18368
rect 110 17912 166 17921
rect 110 17847 166 17856
rect 124 17610 152 17847
rect 112 17604 164 17610
rect 112 17546 164 17552
rect 110 16280 166 16289
rect 110 16215 166 16224
rect 124 16182 152 16215
rect 112 16176 164 16182
rect 112 16118 164 16124
rect 1584 16040 1636 16046
rect 1584 15982 1636 15988
rect 1596 15502 1624 15982
rect 1584 15496 1636 15502
rect 1584 15438 1636 15444
rect 1688 13814 1716 23582
rect 1766 23520 1822 23582
rect 2792 23582 3110 23610
rect 2792 20602 2820 23582
rect 3054 23520 3110 23582
rect 4342 23610 4398 24000
rect 5538 23610 5594 24000
rect 6826 23610 6882 24000
rect 8114 23610 8170 24000
rect 9402 23610 9458 24000
rect 4342 23582 4568 23610
rect 4342 23520 4398 23582
rect 4540 20602 4568 23582
rect 5538 23582 5856 23610
rect 5538 23520 5594 23582
rect 4956 21788 5252 21808
rect 5012 21786 5036 21788
rect 5092 21786 5116 21788
rect 5172 21786 5196 21788
rect 5034 21734 5036 21786
rect 5098 21734 5110 21786
rect 5172 21734 5174 21786
rect 5012 21732 5036 21734
rect 5092 21732 5116 21734
rect 5172 21732 5196 21734
rect 4956 21712 5252 21732
rect 4956 20700 5252 20720
rect 5012 20698 5036 20700
rect 5092 20698 5116 20700
rect 5172 20698 5196 20700
rect 5034 20646 5036 20698
rect 5098 20646 5110 20698
rect 5172 20646 5174 20698
rect 5012 20644 5036 20646
rect 5092 20644 5116 20646
rect 5172 20644 5196 20646
rect 4956 20624 5252 20644
rect 2780 20596 2832 20602
rect 2780 20538 2832 20544
rect 4528 20596 4580 20602
rect 4528 20538 4580 20544
rect 4540 20398 4568 20538
rect 4528 20392 4580 20398
rect 4528 20334 4580 20340
rect 2412 20256 2464 20262
rect 2412 20198 2464 20204
rect 2226 19272 2282 19281
rect 2226 19207 2282 19216
rect 2240 18222 2268 19207
rect 2228 18216 2280 18222
rect 2228 18158 2280 18164
rect 1768 18080 1820 18086
rect 1768 18022 1820 18028
rect 1780 17882 1808 18022
rect 1768 17876 1820 17882
rect 1768 17818 1820 17824
rect 2320 17876 2372 17882
rect 2320 17818 2372 17824
rect 2332 17202 2360 17818
rect 2320 17196 2372 17202
rect 2320 17138 2372 17144
rect 1860 15360 1912 15366
rect 1860 15302 1912 15308
rect 1872 15026 1900 15302
rect 1860 15020 1912 15026
rect 1860 14962 1912 14968
rect 1768 14884 1820 14890
rect 1768 14826 1820 14832
rect 1780 14074 1808 14826
rect 1872 14618 1900 14962
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 1952 14476 2004 14482
rect 1952 14418 2004 14424
rect 1768 14068 1820 14074
rect 1768 14010 1820 14016
rect 1688 13786 1808 13814
rect 20 12912 72 12918
rect 20 12854 72 12860
rect 1676 12776 1728 12782
rect 1676 12718 1728 12724
rect 1688 12374 1716 12718
rect 1676 12368 1728 12374
rect 1582 12336 1638 12345
rect 1676 12310 1728 12316
rect 1582 12271 1638 12280
rect 1596 10810 1624 12271
rect 1780 11558 1808 13786
rect 1964 13734 1992 14418
rect 2136 14068 2188 14074
rect 2136 14010 2188 14016
rect 2148 13802 2176 14010
rect 2228 13932 2280 13938
rect 2228 13874 2280 13880
rect 2136 13796 2188 13802
rect 2136 13738 2188 13744
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1860 13388 1912 13394
rect 1964 13376 1992 13670
rect 1912 13348 1992 13376
rect 1860 13330 1912 13336
rect 1860 13184 1912 13190
rect 1860 13126 1912 13132
rect 1872 12918 1900 13126
rect 1860 12912 1912 12918
rect 1860 12854 1912 12860
rect 1872 12442 1900 12854
rect 1860 12436 1912 12442
rect 1860 12378 1912 12384
rect 1872 12306 1900 12378
rect 1860 12300 1912 12306
rect 1860 12242 1912 12248
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 1768 11552 1820 11558
rect 1768 11494 1820 11500
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 1780 10130 1808 11290
rect 1872 11150 1900 12242
rect 2056 11694 2084 12242
rect 2044 11688 2096 11694
rect 2044 11630 2096 11636
rect 2044 11212 2096 11218
rect 2044 11154 2096 11160
rect 1860 11144 1912 11150
rect 1860 11086 1912 11092
rect 1768 10124 1820 10130
rect 1768 10066 1820 10072
rect 1674 9616 1730 9625
rect 1674 9551 1730 9560
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1596 9081 1624 9318
rect 1582 9072 1638 9081
rect 1582 9007 1638 9016
rect 110 8936 166 8945
rect 110 8871 166 8880
rect 124 2553 152 8871
rect 1688 8430 1716 9551
rect 1872 8974 1900 11086
rect 2056 9382 2084 11154
rect 2148 10198 2176 13738
rect 2240 13462 2268 13874
rect 2228 13456 2280 13462
rect 2228 13398 2280 13404
rect 2320 13252 2372 13258
rect 2320 13194 2372 13200
rect 2332 12782 2360 13194
rect 2320 12776 2372 12782
rect 2320 12718 2372 12724
rect 2332 11626 2360 12718
rect 2320 11620 2372 11626
rect 2320 11562 2372 11568
rect 2136 10192 2188 10198
rect 2136 10134 2188 10140
rect 2148 9722 2176 10134
rect 2136 9716 2188 9722
rect 2136 9658 2188 9664
rect 2044 9376 2096 9382
rect 1964 9336 2044 9364
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 1872 8498 1900 8910
rect 1964 8838 1992 9336
rect 2044 9318 2096 9324
rect 2044 9036 2096 9042
rect 2044 8978 2096 8984
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1964 8430 1992 8774
rect 2056 8566 2084 8978
rect 2044 8560 2096 8566
rect 2044 8502 2096 8508
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 1688 8090 1716 8366
rect 1768 8288 1820 8294
rect 1768 8230 1820 8236
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1780 7886 1808 8230
rect 2148 8090 2176 9658
rect 2332 9042 2360 11562
rect 2424 11354 2452 20198
rect 2872 19712 2924 19718
rect 2872 19654 2924 19660
rect 2884 18290 2912 19654
rect 4956 19612 5252 19632
rect 5012 19610 5036 19612
rect 5092 19610 5116 19612
rect 5172 19610 5196 19612
rect 5034 19558 5036 19610
rect 5098 19558 5110 19610
rect 5172 19558 5174 19610
rect 5012 19556 5036 19558
rect 5092 19556 5116 19558
rect 5172 19556 5196 19558
rect 4956 19536 5252 19556
rect 4956 18524 5252 18544
rect 5012 18522 5036 18524
rect 5092 18522 5116 18524
rect 5172 18522 5196 18524
rect 5034 18470 5036 18522
rect 5098 18470 5110 18522
rect 5172 18470 5174 18522
rect 5012 18468 5036 18470
rect 5092 18468 5116 18470
rect 5172 18468 5196 18470
rect 4956 18448 5252 18468
rect 5828 18329 5856 23582
rect 6826 23582 7144 23610
rect 6826 23520 6882 23582
rect 5814 18320 5870 18329
rect 2872 18284 2924 18290
rect 5814 18255 5870 18264
rect 2872 18226 2924 18232
rect 7116 18193 7144 23582
rect 7944 23582 8170 23610
rect 7944 20602 7972 23582
rect 8114 23520 8170 23582
rect 9324 23582 9458 23610
rect 8392 21344 8444 21350
rect 8392 21286 8444 21292
rect 8404 20602 8432 21286
rect 8956 21244 9252 21264
rect 9012 21242 9036 21244
rect 9092 21242 9116 21244
rect 9172 21242 9196 21244
rect 9034 21190 9036 21242
rect 9098 21190 9110 21242
rect 9172 21190 9174 21242
rect 9012 21188 9036 21190
rect 9092 21188 9116 21190
rect 9172 21188 9196 21190
rect 8956 21168 9252 21188
rect 9324 21146 9352 23582
rect 9402 23520 9458 23582
rect 10598 23610 10654 24000
rect 11886 23610 11942 24000
rect 13174 23610 13230 24000
rect 14462 23610 14518 24000
rect 15658 23610 15714 24000
rect 16946 23610 17002 24000
rect 18234 23610 18290 24000
rect 19522 23610 19578 24000
rect 20718 23610 20774 24000
rect 22006 23610 22062 24000
rect 23294 23610 23350 24000
rect 10598 23582 10916 23610
rect 10598 23520 10654 23582
rect 10048 21344 10100 21350
rect 10048 21286 10100 21292
rect 9312 21140 9364 21146
rect 9312 21082 9364 21088
rect 7932 20596 7984 20602
rect 7932 20538 7984 20544
rect 8392 20596 8444 20602
rect 8392 20538 8444 20544
rect 8404 20398 8432 20538
rect 8392 20392 8444 20398
rect 8392 20334 8444 20340
rect 10060 20330 10088 21286
rect 9404 20324 9456 20330
rect 9404 20266 9456 20272
rect 10048 20324 10100 20330
rect 10048 20266 10100 20272
rect 8852 20256 8904 20262
rect 8852 20198 8904 20204
rect 9312 20256 9364 20262
rect 9312 20198 9364 20204
rect 8024 19916 8076 19922
rect 8024 19858 8076 19864
rect 8036 19514 8064 19858
rect 8024 19508 8076 19514
rect 8024 19450 8076 19456
rect 8576 19304 8628 19310
rect 8576 19246 8628 19252
rect 8588 18630 8616 19246
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 7668 18426 7696 18566
rect 7656 18420 7708 18426
rect 7656 18362 7708 18368
rect 8392 18352 8444 18358
rect 8392 18294 8444 18300
rect 7102 18184 7158 18193
rect 8404 18154 8432 18294
rect 7102 18119 7158 18128
rect 8392 18148 8444 18154
rect 8392 18090 8444 18096
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 5540 17740 5592 17746
rect 5540 17682 5592 17688
rect 6644 17740 6696 17746
rect 6644 17682 6696 17688
rect 4816 17338 4844 17682
rect 5448 17672 5500 17678
rect 5448 17614 5500 17620
rect 4956 17436 5252 17456
rect 5012 17434 5036 17436
rect 5092 17434 5116 17436
rect 5172 17434 5196 17436
rect 5034 17382 5036 17434
rect 5098 17382 5110 17434
rect 5172 17382 5174 17434
rect 5012 17380 5036 17382
rect 5092 17380 5116 17382
rect 5172 17380 5196 17382
rect 4956 17360 5252 17380
rect 4804 17332 4856 17338
rect 4804 17274 4856 17280
rect 3148 17264 3200 17270
rect 3148 17206 3200 17212
rect 2504 17196 2556 17202
rect 2504 17138 2556 17144
rect 2516 15502 2544 17138
rect 3160 16454 3188 17206
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 3976 17060 4028 17066
rect 3976 17002 4028 17008
rect 3700 16992 3752 16998
rect 3700 16934 3752 16940
rect 3148 16448 3200 16454
rect 3148 16390 3200 16396
rect 3160 16046 3188 16390
rect 3148 16040 3200 16046
rect 3148 15982 3200 15988
rect 2596 15632 2648 15638
rect 2596 15574 2648 15580
rect 2504 15496 2556 15502
rect 2504 15438 2556 15444
rect 2516 15094 2544 15438
rect 2608 15162 2636 15574
rect 2596 15156 2648 15162
rect 2596 15098 2648 15104
rect 2504 15088 2556 15094
rect 2504 15030 2556 15036
rect 2688 14272 2740 14278
rect 2688 14214 2740 14220
rect 2700 13938 2728 14214
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 3160 13734 3188 15982
rect 3514 14784 3570 14793
rect 3514 14719 3570 14728
rect 3528 14482 3556 14719
rect 3516 14476 3568 14482
rect 3516 14418 3568 14424
rect 3528 13734 3556 14418
rect 3712 13802 3740 16934
rect 3988 16726 4016 17002
rect 3976 16720 4028 16726
rect 3976 16662 4028 16668
rect 4436 16516 4488 16522
rect 4436 16458 4488 16464
rect 4344 16176 4396 16182
rect 4344 16118 4396 16124
rect 4252 16040 4304 16046
rect 4252 15982 4304 15988
rect 4160 15972 4212 15978
rect 4160 15914 4212 15920
rect 4068 15632 4120 15638
rect 4068 15574 4120 15580
rect 4080 15162 4108 15574
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 4172 14550 4200 15914
rect 4264 15706 4292 15982
rect 4252 15700 4304 15706
rect 4252 15642 4304 15648
rect 3792 14544 3844 14550
rect 3792 14486 3844 14492
rect 4160 14544 4212 14550
rect 4160 14486 4212 14492
rect 3804 14074 3832 14486
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 3884 14272 3936 14278
rect 3884 14214 3936 14220
rect 3792 14068 3844 14074
rect 3792 14010 3844 14016
rect 3896 13938 3924 14214
rect 4080 14074 4108 14350
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 3700 13796 3752 13802
rect 3700 13738 3752 13744
rect 3148 13728 3200 13734
rect 3148 13670 3200 13676
rect 3516 13728 3568 13734
rect 3516 13670 3568 13676
rect 3884 13728 3936 13734
rect 3884 13670 3936 13676
rect 2504 13388 2556 13394
rect 2504 13330 2556 13336
rect 2516 12306 2544 13330
rect 3160 12986 3188 13670
rect 3792 13184 3844 13190
rect 3792 13126 3844 13132
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 3804 12782 3832 13126
rect 3792 12776 3844 12782
rect 3792 12718 3844 12724
rect 3516 12708 3568 12714
rect 3516 12650 3568 12656
rect 2688 12640 2740 12646
rect 2688 12582 2740 12588
rect 2700 12374 2728 12582
rect 2688 12368 2740 12374
rect 2688 12310 2740 12316
rect 2504 12300 2556 12306
rect 2504 12242 2556 12248
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2424 10674 2452 11290
rect 2516 11286 2544 12242
rect 2700 11762 2728 12310
rect 2688 11756 2740 11762
rect 2688 11698 2740 11704
rect 2688 11552 2740 11558
rect 2688 11494 2740 11500
rect 2504 11280 2556 11286
rect 2504 11222 2556 11228
rect 2516 10810 2544 11222
rect 2504 10804 2556 10810
rect 2504 10746 2556 10752
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 2320 9036 2372 9042
rect 2320 8978 2372 8984
rect 2332 8634 2360 8978
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 1780 7546 1808 7822
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 1860 7472 1912 7478
rect 1860 7414 1912 7420
rect 1582 7168 1638 7177
rect 1582 7103 1638 7112
rect 1596 7002 1624 7103
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1582 5400 1638 5409
rect 1582 5335 1638 5344
rect 1492 5092 1544 5098
rect 1492 5034 1544 5040
rect 1216 4820 1268 4826
rect 1216 4762 1268 4768
rect 110 2544 166 2553
rect 110 2479 166 2488
rect 1124 2508 1176 2514
rect 1124 2450 1176 2456
rect 848 2304 900 2310
rect 848 2246 900 2252
rect 478 82 534 480
rect 860 82 888 2246
rect 1136 1465 1164 2450
rect 1122 1456 1178 1465
rect 1122 1391 1178 1400
rect 478 54 888 82
rect 1228 82 1256 4762
rect 1504 4010 1532 5034
rect 1492 4004 1544 4010
rect 1492 3946 1544 3952
rect 1596 3194 1624 5335
rect 1688 5098 1716 6054
rect 1872 5846 1900 7414
rect 2148 7410 2176 8026
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 1952 7268 2004 7274
rect 1952 7210 2004 7216
rect 2044 7268 2096 7274
rect 2044 7210 2096 7216
rect 1964 7002 1992 7210
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 2056 6934 2084 7210
rect 2044 6928 2096 6934
rect 2044 6870 2096 6876
rect 2136 6248 2188 6254
rect 2136 6190 2188 6196
rect 1860 5840 1912 5846
rect 1860 5782 1912 5788
rect 1768 5296 1820 5302
rect 1768 5238 1820 5244
rect 1676 5092 1728 5098
rect 1676 5034 1728 5040
rect 1584 3188 1636 3194
rect 1584 3130 1636 3136
rect 1780 2650 1808 5238
rect 1872 4826 1900 5782
rect 2148 5234 2176 6190
rect 2700 6186 2728 11494
rect 3240 11008 3292 11014
rect 3240 10950 3292 10956
rect 2964 10668 3016 10674
rect 2964 10610 3016 10616
rect 2780 10532 2832 10538
rect 2780 10474 2832 10480
rect 2792 10198 2820 10474
rect 2780 10192 2832 10198
rect 2780 10134 2832 10140
rect 2976 9654 3004 10610
rect 2964 9648 3016 9654
rect 2964 9590 3016 9596
rect 2976 7410 3004 9590
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 3160 9178 3188 9318
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 3252 8566 3280 10950
rect 3528 9625 3556 12650
rect 3700 12640 3752 12646
rect 3700 12582 3752 12588
rect 3712 11898 3740 12582
rect 3700 11892 3752 11898
rect 3700 11834 3752 11840
rect 3700 11688 3752 11694
rect 3804 11676 3832 12718
rect 3752 11648 3832 11676
rect 3700 11630 3752 11636
rect 3712 11014 3740 11630
rect 3792 11280 3844 11286
rect 3792 11222 3844 11228
rect 3700 11008 3752 11014
rect 3700 10950 3752 10956
rect 3804 10470 3832 11222
rect 3792 10464 3844 10470
rect 3792 10406 3844 10412
rect 3700 9988 3752 9994
rect 3700 9930 3752 9936
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 3620 9722 3648 9862
rect 3608 9716 3660 9722
rect 3608 9658 3660 9664
rect 3514 9616 3570 9625
rect 3514 9551 3570 9560
rect 3516 9444 3568 9450
rect 3516 9386 3568 9392
rect 3240 8560 3292 8566
rect 3240 8502 3292 8508
rect 3528 7886 3556 9386
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 2964 7404 3016 7410
rect 2964 7346 3016 7352
rect 3516 7268 3568 7274
rect 3516 7210 3568 7216
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3344 6934 3372 7142
rect 3332 6928 3384 6934
rect 3332 6870 3384 6876
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 2884 6322 2912 6802
rect 3528 6662 3556 7210
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 2884 6225 2912 6258
rect 2870 6216 2926 6225
rect 2688 6180 2740 6186
rect 2870 6151 2926 6160
rect 2688 6122 2740 6128
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2424 5778 2452 6054
rect 2872 5840 2924 5846
rect 2872 5782 2924 5788
rect 2412 5772 2464 5778
rect 2412 5714 2464 5720
rect 2136 5228 2188 5234
rect 2136 5170 2188 5176
rect 1860 4820 1912 4826
rect 1860 4762 1912 4768
rect 1872 4214 1900 4762
rect 2148 4622 2176 5170
rect 2424 4826 2452 5714
rect 2884 5370 2912 5782
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 2688 5092 2740 5098
rect 2688 5034 2740 5040
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 2136 4616 2188 4622
rect 2136 4558 2188 4564
rect 1860 4208 1912 4214
rect 1860 4150 1912 4156
rect 1964 4146 1992 4558
rect 2424 4282 2452 4762
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 2044 2848 2096 2854
rect 2044 2790 2096 2796
rect 1768 2644 1820 2650
rect 1768 2586 1820 2592
rect 2056 1737 2084 2790
rect 2042 1728 2098 1737
rect 2042 1663 2098 1672
rect 1398 82 1454 480
rect 1228 54 1454 82
rect 478 0 534 54
rect 1398 0 1454 54
rect 2318 82 2374 480
rect 2700 82 2728 5034
rect 3528 2650 3556 6598
rect 3620 6458 3648 9658
rect 3712 9586 3740 9930
rect 3700 9580 3752 9586
rect 3700 9522 3752 9528
rect 3712 9178 3740 9522
rect 3700 9172 3752 9178
rect 3700 9114 3752 9120
rect 3804 8974 3832 10406
rect 3896 9926 3924 13670
rect 4080 13530 4108 14010
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 4160 13388 4212 13394
rect 4160 13330 4212 13336
rect 4172 12986 4200 13330
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 3976 12776 4028 12782
rect 3976 12718 4028 12724
rect 3988 12442 4016 12718
rect 4068 12640 4120 12646
rect 4068 12582 4120 12588
rect 3976 12436 4028 12442
rect 3976 12378 4028 12384
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 3988 11830 4016 12174
rect 3976 11824 4028 11830
rect 3976 11766 4028 11772
rect 4080 11762 4108 12582
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 4172 12306 4200 12378
rect 4160 12300 4212 12306
rect 4212 12260 4292 12288
rect 4160 12242 4212 12248
rect 4264 11898 4292 12260
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4160 11824 4212 11830
rect 4160 11766 4212 11772
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 4068 10736 4120 10742
rect 4068 10678 4120 10684
rect 3976 10192 4028 10198
rect 3976 10134 4028 10140
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3896 9042 3924 9862
rect 3988 9450 4016 10134
rect 4080 10130 4108 10678
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 4080 9518 4108 10066
rect 4172 9625 4200 11766
rect 4356 11558 4384 16118
rect 4448 16114 4476 16458
rect 4436 16108 4488 16114
rect 4436 16050 4488 16056
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4356 10810 4384 11494
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4158 9616 4214 9625
rect 4448 9586 4476 16050
rect 4632 15502 4660 17138
rect 5460 16658 5488 17614
rect 5552 16998 5580 17682
rect 6184 17264 6236 17270
rect 6184 17206 6236 17212
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 4956 16348 5252 16368
rect 5012 16346 5036 16348
rect 5092 16346 5116 16348
rect 5172 16346 5196 16348
rect 5034 16294 5036 16346
rect 5098 16294 5110 16346
rect 5172 16294 5174 16346
rect 5012 16292 5036 16294
rect 5092 16292 5116 16294
rect 5172 16292 5196 16294
rect 4956 16272 5252 16292
rect 5460 16250 5488 16594
rect 5448 16244 5500 16250
rect 5448 16186 5500 16192
rect 4988 15904 5040 15910
rect 4988 15846 5040 15852
rect 5000 15638 5028 15846
rect 4988 15632 5040 15638
rect 4988 15574 5040 15580
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4632 15366 4660 15438
rect 4804 15428 4856 15434
rect 4804 15370 4856 15376
rect 4620 15360 4672 15366
rect 4620 15302 4672 15308
rect 4632 14550 4660 15302
rect 4816 15026 4844 15370
rect 4956 15260 5252 15280
rect 5012 15258 5036 15260
rect 5092 15258 5116 15260
rect 5172 15258 5196 15260
rect 5034 15206 5036 15258
rect 5098 15206 5110 15258
rect 5172 15206 5174 15258
rect 5012 15204 5036 15206
rect 5092 15204 5116 15206
rect 5172 15204 5196 15206
rect 4956 15184 5252 15204
rect 5356 15088 5408 15094
rect 5356 15030 5408 15036
rect 4804 15020 4856 15026
rect 4804 14962 4856 14968
rect 5368 14822 5396 15030
rect 4988 14816 5040 14822
rect 4988 14758 5040 14764
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5000 14618 5028 14758
rect 4988 14612 5040 14618
rect 4988 14554 5040 14560
rect 4620 14544 4672 14550
rect 4620 14486 4672 14492
rect 4956 14172 5252 14192
rect 5012 14170 5036 14172
rect 5092 14170 5116 14172
rect 5172 14170 5196 14172
rect 5034 14118 5036 14170
rect 5098 14118 5110 14170
rect 5172 14118 5174 14170
rect 5012 14116 5036 14118
rect 5092 14116 5116 14118
rect 5172 14116 5196 14118
rect 4956 14096 5252 14116
rect 5368 13938 5396 14758
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 5552 13841 5580 16934
rect 5632 16720 5684 16726
rect 5632 16662 5684 16668
rect 5644 16114 5672 16662
rect 5632 16108 5684 16114
rect 5632 16050 5684 16056
rect 5908 14272 5960 14278
rect 5908 14214 5960 14220
rect 5354 13832 5410 13841
rect 5354 13767 5410 13776
rect 5538 13832 5594 13841
rect 5538 13767 5594 13776
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4528 12844 4580 12850
rect 4528 12786 4580 12792
rect 4158 9551 4214 9560
rect 4436 9580 4488 9586
rect 4436 9522 4488 9528
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 3976 9444 4028 9450
rect 3976 9386 4028 9392
rect 3884 9036 3936 9042
rect 3884 8978 3936 8984
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 4080 8537 4108 9454
rect 4436 9444 4488 9450
rect 4436 9386 4488 9392
rect 4448 9178 4476 9386
rect 4436 9172 4488 9178
rect 4436 9114 4488 9120
rect 4436 9036 4488 9042
rect 4436 8978 4488 8984
rect 4066 8528 4122 8537
rect 4066 8463 4122 8472
rect 4448 8294 4476 8978
rect 4540 8566 4568 12786
rect 4632 12714 4660 13330
rect 4956 13084 5252 13104
rect 5012 13082 5036 13084
rect 5092 13082 5116 13084
rect 5172 13082 5196 13084
rect 5034 13030 5036 13082
rect 5098 13030 5110 13082
rect 5172 13030 5174 13082
rect 5012 13028 5036 13030
rect 5092 13028 5116 13030
rect 5172 13028 5196 13030
rect 4956 13008 5252 13028
rect 4896 12912 4948 12918
rect 4896 12854 4948 12860
rect 4620 12708 4672 12714
rect 4620 12650 4672 12656
rect 4908 12646 4936 12854
rect 5368 12850 5396 13767
rect 5724 13184 5776 13190
rect 5724 13126 5776 13132
rect 5632 12912 5684 12918
rect 5632 12854 5684 12860
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 4908 12306 4936 12582
rect 5644 12374 5672 12854
rect 5736 12442 5764 13126
rect 5920 12986 5948 14214
rect 6092 13728 6144 13734
rect 6092 13670 6144 13676
rect 5908 12980 5960 12986
rect 5908 12922 5960 12928
rect 5816 12640 5868 12646
rect 5816 12582 5868 12588
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 5632 12368 5684 12374
rect 5632 12310 5684 12316
rect 4896 12300 4948 12306
rect 4896 12242 4948 12248
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 4956 11996 5252 12016
rect 5012 11994 5036 11996
rect 5092 11994 5116 11996
rect 5172 11994 5196 11996
rect 5034 11942 5036 11994
rect 5098 11942 5110 11994
rect 5172 11942 5174 11994
rect 5012 11940 5036 11942
rect 5092 11940 5116 11942
rect 5172 11940 5196 11942
rect 4956 11920 5252 11940
rect 5736 11898 5764 12242
rect 5828 11898 5856 12582
rect 5724 11892 5776 11898
rect 5724 11834 5776 11840
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4724 10266 4752 11154
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 5724 11008 5776 11014
rect 5724 10950 5776 10956
rect 4956 10908 5252 10928
rect 5012 10906 5036 10908
rect 5092 10906 5116 10908
rect 5172 10906 5196 10908
rect 5034 10854 5036 10906
rect 5098 10854 5110 10906
rect 5172 10854 5174 10906
rect 5012 10852 5036 10854
rect 5092 10852 5116 10854
rect 5172 10852 5196 10854
rect 4956 10832 5252 10852
rect 5448 10532 5500 10538
rect 5448 10474 5500 10480
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 4724 9926 4752 10202
rect 5460 10062 5488 10474
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4956 9820 5252 9840
rect 5012 9818 5036 9820
rect 5092 9818 5116 9820
rect 5172 9818 5196 9820
rect 5034 9766 5036 9818
rect 5098 9766 5110 9818
rect 5172 9766 5174 9818
rect 5012 9764 5036 9766
rect 5092 9764 5116 9766
rect 5172 9764 5196 9766
rect 4956 9744 5252 9764
rect 5460 9722 5488 9998
rect 5736 9761 5764 10950
rect 5920 10810 5948 11086
rect 5908 10804 5960 10810
rect 5908 10746 5960 10752
rect 5816 10192 5868 10198
rect 5816 10134 5868 10140
rect 5722 9752 5778 9761
rect 5448 9716 5500 9722
rect 5722 9687 5778 9696
rect 5448 9658 5500 9664
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4528 8560 4580 8566
rect 4528 8502 4580 8508
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 4436 8288 4488 8294
rect 4436 8230 4488 8236
rect 3896 8022 3924 8230
rect 3884 8016 3936 8022
rect 3884 7958 3936 7964
rect 4252 8016 4304 8022
rect 4252 7958 4304 7964
rect 3896 7002 3924 7958
rect 4264 7206 4292 7958
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4264 7002 4292 7142
rect 3884 6996 3936 7002
rect 3884 6938 3936 6944
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 3608 6452 3660 6458
rect 3608 6394 3660 6400
rect 3608 5772 3660 5778
rect 3608 5714 3660 5720
rect 3620 5166 3648 5714
rect 4448 5574 4476 8230
rect 4540 6866 4568 8502
rect 4724 8430 4752 8774
rect 4816 8430 4844 8774
rect 4956 8732 5252 8752
rect 5012 8730 5036 8732
rect 5092 8730 5116 8732
rect 5172 8730 5196 8732
rect 5034 8678 5036 8730
rect 5098 8678 5110 8730
rect 5172 8678 5174 8730
rect 5012 8676 5036 8678
rect 5092 8676 5116 8678
rect 5172 8676 5196 8678
rect 4956 8656 5252 8676
rect 5368 8498 5396 8910
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4804 8424 4856 8430
rect 4804 8366 4856 8372
rect 4724 8090 4752 8366
rect 4712 8084 4764 8090
rect 4712 8026 4764 8032
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4724 7002 4752 7278
rect 4712 6996 4764 7002
rect 4712 6938 4764 6944
rect 4816 6866 4844 8366
rect 4956 7644 5252 7664
rect 5012 7642 5036 7644
rect 5092 7642 5116 7644
rect 5172 7642 5196 7644
rect 5034 7590 5036 7642
rect 5098 7590 5110 7642
rect 5172 7590 5174 7642
rect 5012 7588 5036 7590
rect 5092 7588 5116 7590
rect 5172 7588 5196 7590
rect 4956 7568 5252 7588
rect 4528 6860 4580 6866
rect 4528 6802 4580 6808
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4540 6458 4568 6802
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4724 5778 4752 6394
rect 4816 6390 4844 6802
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 4956 6556 5252 6576
rect 5012 6554 5036 6556
rect 5092 6554 5116 6556
rect 5172 6554 5196 6556
rect 5034 6502 5036 6554
rect 5098 6502 5110 6554
rect 5172 6502 5174 6554
rect 5012 6500 5036 6502
rect 5092 6500 5116 6502
rect 5172 6500 5196 6502
rect 4956 6480 5252 6500
rect 4804 6384 4856 6390
rect 4804 6326 4856 6332
rect 5368 6322 5396 6598
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5368 5914 5396 6258
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 4540 5642 4568 5714
rect 4528 5636 4580 5642
rect 4528 5578 4580 5584
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 3608 5160 3660 5166
rect 3608 5102 3660 5108
rect 4620 5160 4672 5166
rect 4724 5148 4752 5714
rect 4956 5468 5252 5488
rect 5012 5466 5036 5468
rect 5092 5466 5116 5468
rect 5172 5466 5196 5468
rect 5034 5414 5036 5466
rect 5098 5414 5110 5466
rect 5172 5414 5174 5466
rect 5012 5412 5036 5414
rect 5092 5412 5116 5414
rect 5172 5412 5196 5414
rect 4956 5392 5252 5412
rect 5460 5370 5488 6054
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 4672 5120 4752 5148
rect 4620 5102 4672 5108
rect 3620 4486 3648 5102
rect 3792 5024 3844 5030
rect 3792 4966 3844 4972
rect 3608 4480 3660 4486
rect 3608 4422 3660 4428
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 2318 54 2728 82
rect 3238 82 3294 480
rect 3620 82 3648 4422
rect 3804 4078 3832 4966
rect 4344 4752 4396 4758
rect 4344 4694 4396 4700
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 4356 3942 4384 4694
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4540 4282 4568 4558
rect 4528 4276 4580 4282
rect 4528 4218 4580 4224
rect 4724 4146 4752 4558
rect 4956 4380 5252 4400
rect 5012 4378 5036 4380
rect 5092 4378 5116 4380
rect 5172 4378 5196 4380
rect 5034 4326 5036 4378
rect 5098 4326 5110 4378
rect 5172 4326 5174 4378
rect 5012 4324 5036 4326
rect 5092 4324 5116 4326
rect 5172 4324 5196 4326
rect 4956 4304 5252 4324
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 4252 3188 4304 3194
rect 4356 3176 4384 3878
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4528 3392 4580 3398
rect 4528 3334 4580 3340
rect 4448 3194 4476 3334
rect 4304 3148 4384 3176
rect 4436 3188 4488 3194
rect 4252 3130 4304 3136
rect 4436 3130 4488 3136
rect 4252 2984 4304 2990
rect 4252 2926 4304 2932
rect 3238 54 3648 82
rect 4158 82 4214 480
rect 4264 82 4292 2926
rect 4448 2854 4476 3130
rect 4540 3058 4568 3334
rect 4724 3058 4752 4082
rect 5552 4078 5580 9522
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5644 6322 5672 6802
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 5736 5778 5764 9687
rect 5828 9382 5856 10134
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5828 9110 5856 9318
rect 5816 9104 5868 9110
rect 5816 9046 5868 9052
rect 5828 8430 5856 9046
rect 6012 9042 6040 12582
rect 6000 9036 6052 9042
rect 6000 8978 6052 8984
rect 6104 8634 6132 13670
rect 6196 12306 6224 17206
rect 6656 17105 6684 17682
rect 6920 17536 6972 17542
rect 6920 17478 6972 17484
rect 8484 17536 8536 17542
rect 8484 17478 8536 17484
rect 6642 17096 6698 17105
rect 6642 17031 6698 17040
rect 6656 16998 6684 17031
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 6368 16448 6420 16454
rect 6368 16390 6420 16396
rect 6380 15910 6408 16390
rect 6932 16114 6960 17478
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 7012 17060 7064 17066
rect 7012 17002 7064 17008
rect 7024 16454 7052 17002
rect 7208 16561 7236 17138
rect 8496 17134 8524 17478
rect 8484 17128 8536 17134
rect 8404 17088 8484 17116
rect 7564 17060 7616 17066
rect 7564 17002 7616 17008
rect 7194 16552 7250 16561
rect 7194 16487 7250 16496
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 7196 16108 7248 16114
rect 7196 16050 7248 16056
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 6380 14550 6408 15846
rect 6552 15632 6604 15638
rect 6552 15574 6604 15580
rect 6460 15496 6512 15502
rect 6460 15438 6512 15444
rect 6472 15162 6500 15438
rect 6460 15156 6512 15162
rect 6460 15098 6512 15104
rect 6564 14890 6592 15574
rect 7208 15434 7236 16050
rect 7196 15428 7248 15434
rect 7196 15370 7248 15376
rect 7576 15094 7604 17002
rect 7932 16720 7984 16726
rect 7932 16662 7984 16668
rect 7944 16250 7972 16662
rect 7932 16244 7984 16250
rect 7932 16186 7984 16192
rect 8404 15706 8432 17088
rect 8484 17070 8536 17076
rect 8484 16992 8536 16998
rect 8484 16934 8536 16940
rect 8496 16590 8524 16934
rect 8484 16584 8536 16590
rect 8484 16526 8536 16532
rect 8496 16250 8524 16526
rect 8484 16244 8536 16250
rect 8484 16186 8536 16192
rect 8392 15700 8444 15706
rect 8392 15642 8444 15648
rect 8114 15464 8170 15473
rect 8114 15399 8170 15408
rect 7564 15088 7616 15094
rect 7564 15030 7616 15036
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 6552 14884 6604 14890
rect 6552 14826 6604 14832
rect 7012 14884 7064 14890
rect 7012 14826 7064 14832
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6368 14544 6420 14550
rect 6368 14486 6420 14492
rect 6380 14074 6408 14486
rect 6840 14414 6868 14758
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6460 13864 6512 13870
rect 6460 13806 6512 13812
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 6196 11830 6224 12242
rect 6184 11824 6236 11830
rect 6184 11766 6236 11772
rect 6196 11626 6224 11766
rect 6184 11620 6236 11626
rect 6184 11562 6236 11568
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 5816 8424 5868 8430
rect 5816 8366 5868 8372
rect 5828 7274 5856 8366
rect 5816 7268 5868 7274
rect 5816 7210 5868 7216
rect 5724 5772 5776 5778
rect 5724 5714 5776 5720
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5644 5409 5672 5646
rect 5630 5400 5686 5409
rect 5630 5335 5686 5344
rect 5644 5234 5672 5335
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5736 4826 5764 5714
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 5736 4554 5764 4762
rect 5724 4548 5776 4554
rect 5724 4490 5776 4496
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4816 3602 4844 3878
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 5816 3596 5868 3602
rect 5816 3538 5868 3544
rect 4956 3292 5252 3312
rect 5012 3290 5036 3292
rect 5092 3290 5116 3292
rect 5172 3290 5196 3292
rect 5034 3238 5036 3290
rect 5098 3238 5110 3290
rect 5172 3238 5174 3290
rect 5012 3236 5036 3238
rect 5092 3236 5116 3238
rect 5172 3236 5196 3238
rect 4956 3216 5252 3236
rect 4528 3052 4580 3058
rect 4528 2994 4580 3000
rect 4712 3052 4764 3058
rect 4712 2994 4764 3000
rect 5828 2854 5856 3538
rect 4436 2848 4488 2854
rect 4436 2790 4488 2796
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 4804 2304 4856 2310
rect 4804 2246 4856 2252
rect 4158 54 4292 82
rect 4816 82 4844 2246
rect 4956 2204 5252 2224
rect 5012 2202 5036 2204
rect 5092 2202 5116 2204
rect 5172 2202 5196 2204
rect 5034 2150 5036 2202
rect 5098 2150 5110 2202
rect 5172 2150 5174 2202
rect 5012 2148 5036 2150
rect 5092 2148 5116 2150
rect 5172 2148 5196 2150
rect 4956 2128 5252 2148
rect 5828 2106 5856 2790
rect 5816 2100 5868 2106
rect 5816 2042 5868 2048
rect 5078 82 5134 480
rect 4816 54 5134 82
rect 2318 0 2374 54
rect 3238 0 3294 54
rect 4158 0 4214 54
rect 5078 0 5134 54
rect 5998 82 6054 480
rect 6104 82 6132 8570
rect 6472 7954 6500 13806
rect 6736 13728 6788 13734
rect 6736 13670 6788 13676
rect 6552 13456 6604 13462
rect 6552 13398 6604 13404
rect 6564 12918 6592 13398
rect 6552 12912 6604 12918
rect 6552 12854 6604 12860
rect 6564 11354 6592 12854
rect 6748 12850 6776 13670
rect 6840 12918 6868 14350
rect 7024 14278 7052 14826
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 7024 13530 7052 14214
rect 7012 13524 7064 13530
rect 7012 13466 7064 13472
rect 6828 12912 6880 12918
rect 6828 12854 6880 12860
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 7024 12714 7052 13466
rect 7012 12708 7064 12714
rect 7012 12650 7064 12656
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6932 11830 6960 12038
rect 6920 11824 6972 11830
rect 6920 11766 6972 11772
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6840 11558 6868 11630
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 6564 10810 6592 11290
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6564 10198 6592 10746
rect 6552 10192 6604 10198
rect 6552 10134 6604 10140
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 7024 9450 7052 10066
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 7116 9926 7144 9998
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 6644 9104 6696 9110
rect 6644 9046 6696 9052
rect 6656 8634 6684 9046
rect 6748 8974 6776 9386
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6932 8786 6960 9386
rect 7024 9178 7052 9386
rect 7012 9172 7064 9178
rect 7012 9114 7064 9120
rect 6932 8758 7052 8786
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6736 8288 6788 8294
rect 6736 8230 6788 8236
rect 6748 8022 6776 8230
rect 6736 8016 6788 8022
rect 6736 7958 6788 7964
rect 6828 8016 6880 8022
rect 6828 7958 6880 7964
rect 6460 7948 6512 7954
rect 6460 7890 6512 7896
rect 6472 7546 6500 7890
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 6736 7200 6788 7206
rect 6840 7188 6868 7958
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6932 7410 6960 7686
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6788 7160 6868 7188
rect 6736 7142 6788 7148
rect 6748 6934 6776 7142
rect 6932 7002 6960 7346
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 6736 6928 6788 6934
rect 6736 6870 6788 6876
rect 7024 6798 7052 8758
rect 7116 7886 7144 9862
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 6552 6384 6604 6390
rect 6552 6326 6604 6332
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 6196 5166 6224 5714
rect 6380 5642 6408 6054
rect 6564 5642 6592 6326
rect 6368 5636 6420 5642
rect 6368 5578 6420 5584
rect 6552 5636 6604 5642
rect 6552 5578 6604 5584
rect 6564 5370 6592 5578
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 6656 5273 6684 6734
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 6828 5772 6880 5778
rect 6828 5714 6880 5720
rect 6642 5264 6698 5273
rect 6642 5199 6698 5208
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6184 5160 6236 5166
rect 6184 5102 6236 5108
rect 6196 4826 6224 5102
rect 6184 4820 6236 4826
rect 6184 4762 6236 4768
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6472 3398 6500 4626
rect 6748 4622 6776 5170
rect 6840 4758 6868 5714
rect 6932 5710 6960 6190
rect 7116 6118 7144 6190
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 6828 4752 6880 4758
rect 6828 4694 6880 4700
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6552 4004 6604 4010
rect 6552 3946 6604 3952
rect 6184 3392 6236 3398
rect 6184 3334 6236 3340
rect 6460 3392 6512 3398
rect 6460 3334 6512 3340
rect 6196 2582 6224 3334
rect 6564 3194 6592 3946
rect 6748 3738 6776 4558
rect 6840 4282 6868 4694
rect 6828 4276 6880 4282
rect 6828 4218 6880 4224
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6552 3188 6604 3194
rect 6604 3148 6684 3176
rect 6552 3130 6604 3136
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 6184 2576 6236 2582
rect 6184 2518 6236 2524
rect 6564 2514 6592 2926
rect 6656 2922 6684 3148
rect 6644 2916 6696 2922
rect 6644 2858 6696 2864
rect 6552 2508 6604 2514
rect 6552 2450 6604 2456
rect 5998 54 6132 82
rect 6918 82 6974 480
rect 7024 82 7052 5510
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 7116 5030 7144 5102
rect 7104 5024 7156 5030
rect 7104 4966 7156 4972
rect 7208 4154 7236 14962
rect 7748 14816 7800 14822
rect 7748 14758 7800 14764
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 7300 11694 7328 12242
rect 7288 11688 7340 11694
rect 7760 11676 7788 14758
rect 8024 14612 8076 14618
rect 8024 14554 8076 14560
rect 7840 14476 7892 14482
rect 7840 14418 7892 14424
rect 7852 13841 7880 14418
rect 8036 13938 8064 14554
rect 8128 14482 8156 15399
rect 8208 14884 8260 14890
rect 8208 14826 8260 14832
rect 8220 14793 8248 14826
rect 8206 14784 8262 14793
rect 8206 14719 8262 14728
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 8024 13932 8076 13938
rect 8024 13874 8076 13880
rect 7838 13832 7894 13841
rect 7838 13767 7894 13776
rect 7852 13530 7880 13767
rect 8220 13530 8248 14719
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 7840 13524 7892 13530
rect 7840 13466 7892 13472
rect 8208 13524 8260 13530
rect 8208 13466 8260 13472
rect 8312 13190 8340 14418
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 8404 13462 8432 13670
rect 8392 13456 8444 13462
rect 8392 13398 8444 13404
rect 8484 13388 8536 13394
rect 8484 13330 8536 13336
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 8496 12986 8524 13330
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 7840 12300 7892 12306
rect 8024 12300 8076 12306
rect 7892 12260 7972 12288
rect 7840 12242 7892 12248
rect 7840 11688 7892 11694
rect 7760 11648 7840 11676
rect 7288 11630 7340 11636
rect 7840 11630 7892 11636
rect 7300 4826 7328 11630
rect 7656 11620 7708 11626
rect 7656 11562 7708 11568
rect 7380 11008 7432 11014
rect 7380 10950 7432 10956
rect 7392 10198 7420 10950
rect 7564 10600 7616 10606
rect 7564 10542 7616 10548
rect 7380 10192 7432 10198
rect 7380 10134 7432 10140
rect 7392 9722 7420 10134
rect 7576 10062 7604 10542
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7380 9716 7432 9722
rect 7380 9658 7432 9664
rect 7576 9450 7604 9998
rect 7668 9518 7696 11562
rect 7748 9716 7800 9722
rect 7748 9658 7800 9664
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 7564 9444 7616 9450
rect 7564 9386 7616 9392
rect 7576 8974 7604 9386
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 7392 8090 7420 8910
rect 7564 8288 7616 8294
rect 7564 8230 7616 8236
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7392 7410 7420 8026
rect 7576 7993 7604 8230
rect 7562 7984 7618 7993
rect 7484 7942 7562 7970
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 7484 5556 7512 7942
rect 7562 7919 7618 7928
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7576 6186 7604 7278
rect 7564 6180 7616 6186
rect 7564 6122 7616 6128
rect 7392 5528 7512 5556
rect 7564 5568 7616 5574
rect 7288 4820 7340 4826
rect 7392 4808 7420 5528
rect 7564 5510 7616 5516
rect 7576 5234 7604 5510
rect 7564 5228 7616 5234
rect 7564 5170 7616 5176
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7484 5030 7512 5102
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7564 4820 7616 4826
rect 7392 4780 7512 4808
rect 7288 4762 7340 4768
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 7116 4126 7236 4154
rect 7116 1873 7144 4126
rect 7300 4078 7328 4218
rect 7288 4072 7340 4078
rect 7288 4014 7340 4020
rect 7392 4010 7420 4558
rect 7484 4282 7512 4780
rect 7564 4762 7616 4768
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7380 4004 7432 4010
rect 7380 3946 7432 3952
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7300 3534 7328 3878
rect 7380 3664 7432 3670
rect 7380 3606 7432 3612
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 7300 3194 7328 3470
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 7392 2990 7420 3606
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 7102 1864 7158 1873
rect 7102 1799 7158 1808
rect 7576 105 7604 4762
rect 6918 54 7052 82
rect 7562 96 7618 105
rect 5998 0 6054 54
rect 6918 0 6974 54
rect 7668 82 7696 7482
rect 7760 5409 7788 9658
rect 7852 8022 7880 11630
rect 7944 11014 7972 12260
rect 8024 12242 8076 12248
rect 8036 11558 8064 12242
rect 8208 12164 8260 12170
rect 8208 12106 8260 12112
rect 8116 11688 8168 11694
rect 8116 11630 8168 11636
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 8036 11082 8064 11494
rect 8024 11076 8076 11082
rect 8024 11018 8076 11024
rect 7932 11008 7984 11014
rect 7932 10950 7984 10956
rect 7944 9081 7972 10950
rect 8036 10470 8064 11018
rect 8128 10606 8156 11630
rect 8220 11558 8248 12106
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8220 11082 8248 11494
rect 8208 11076 8260 11082
rect 8208 11018 8260 11024
rect 8220 10606 8248 11018
rect 8116 10600 8168 10606
rect 8116 10542 8168 10548
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 8036 9654 8064 10406
rect 8024 9648 8076 9654
rect 8024 9590 8076 9596
rect 7930 9072 7986 9081
rect 7930 9007 7986 9016
rect 7840 8016 7892 8022
rect 7840 7958 7892 7964
rect 8036 6254 8064 9590
rect 8128 9382 8156 10542
rect 8220 9926 8248 10542
rect 8588 10470 8616 18566
rect 8760 18148 8812 18154
rect 8760 18090 8812 18096
rect 8666 17096 8722 17105
rect 8666 17031 8722 17040
rect 8576 10464 8628 10470
rect 8576 10406 8628 10412
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 8220 6118 8248 9862
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8496 7750 8524 9318
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 8588 8430 8616 9114
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8588 8090 8616 8366
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8680 7562 8708 17031
rect 8772 16998 8800 18090
rect 8760 16992 8812 16998
rect 8760 16934 8812 16940
rect 8772 16794 8800 16934
rect 8760 16788 8812 16794
rect 8760 16730 8812 16736
rect 8864 16017 8892 20198
rect 8956 20156 9252 20176
rect 9012 20154 9036 20156
rect 9092 20154 9116 20156
rect 9172 20154 9196 20156
rect 9034 20102 9036 20154
rect 9098 20102 9110 20154
rect 9172 20102 9174 20154
rect 9012 20100 9036 20102
rect 9092 20100 9116 20102
rect 9172 20100 9196 20102
rect 8956 20080 9252 20100
rect 9324 19514 9352 20198
rect 9416 19718 9444 20266
rect 9772 19984 9824 19990
rect 9772 19926 9824 19932
rect 9404 19712 9456 19718
rect 9404 19654 9456 19660
rect 9784 19514 9812 19926
rect 10060 19854 10088 20266
rect 10048 19848 10100 19854
rect 10048 19790 10100 19796
rect 10140 19780 10192 19786
rect 10140 19722 10192 19728
rect 10152 19514 10180 19722
rect 9312 19508 9364 19514
rect 9312 19450 9364 19456
rect 9772 19508 9824 19514
rect 9772 19450 9824 19456
rect 10140 19508 10192 19514
rect 10140 19450 10192 19456
rect 10692 19304 10744 19310
rect 10692 19246 10744 19252
rect 9680 19236 9732 19242
rect 9680 19178 9732 19184
rect 8956 19068 9252 19088
rect 9012 19066 9036 19068
rect 9092 19066 9116 19068
rect 9172 19066 9196 19068
rect 9034 19014 9036 19066
rect 9098 19014 9110 19066
rect 9172 19014 9174 19066
rect 9012 19012 9036 19014
rect 9092 19012 9116 19014
rect 9172 19012 9196 19014
rect 8956 18992 9252 19012
rect 9692 18902 9720 19178
rect 10704 18970 10732 19246
rect 10692 18964 10744 18970
rect 10692 18906 10744 18912
rect 9680 18896 9732 18902
rect 9680 18838 9732 18844
rect 9312 18420 9364 18426
rect 9312 18362 9364 18368
rect 8956 17980 9252 18000
rect 9012 17978 9036 17980
rect 9092 17978 9116 17980
rect 9172 17978 9196 17980
rect 9034 17926 9036 17978
rect 9098 17926 9110 17978
rect 9172 17926 9174 17978
rect 9012 17924 9036 17926
rect 9092 17924 9116 17926
rect 9172 17924 9196 17926
rect 8956 17904 9252 17924
rect 8956 16892 9252 16912
rect 9012 16890 9036 16892
rect 9092 16890 9116 16892
rect 9172 16890 9196 16892
rect 9034 16838 9036 16890
rect 9098 16838 9110 16890
rect 9172 16838 9174 16890
rect 9012 16836 9036 16838
rect 9092 16836 9116 16838
rect 9172 16836 9196 16838
rect 8956 16816 9252 16836
rect 8850 16008 8906 16017
rect 8850 15943 8906 15952
rect 8956 15804 9252 15824
rect 9012 15802 9036 15804
rect 9092 15802 9116 15804
rect 9172 15802 9196 15804
rect 9034 15750 9036 15802
rect 9098 15750 9110 15802
rect 9172 15750 9174 15802
rect 9012 15748 9036 15750
rect 9092 15748 9116 15750
rect 9172 15748 9196 15750
rect 8956 15728 9252 15748
rect 8852 15700 8904 15706
rect 8852 15642 8904 15648
rect 8864 14958 8892 15642
rect 8852 14952 8904 14958
rect 8852 14894 8904 14900
rect 8864 14618 8892 14894
rect 8956 14716 9252 14736
rect 9012 14714 9036 14716
rect 9092 14714 9116 14716
rect 9172 14714 9196 14716
rect 9034 14662 9036 14714
rect 9098 14662 9110 14714
rect 9172 14662 9174 14714
rect 9012 14660 9036 14662
rect 9092 14660 9116 14662
rect 9172 14660 9196 14662
rect 8956 14640 9252 14660
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8956 13628 9252 13648
rect 9012 13626 9036 13628
rect 9092 13626 9116 13628
rect 9172 13626 9196 13628
rect 9034 13574 9036 13626
rect 9098 13574 9110 13626
rect 9172 13574 9174 13626
rect 9012 13572 9036 13574
rect 9092 13572 9116 13574
rect 9172 13572 9196 13574
rect 8956 13552 9252 13572
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8312 7534 8708 7562
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 7746 5400 7802 5409
rect 7746 5335 7748 5344
rect 7800 5335 7802 5344
rect 7748 5306 7800 5312
rect 7760 5275 7788 5306
rect 7748 5092 7800 5098
rect 7748 5034 7800 5040
rect 7760 4214 7788 5034
rect 8128 5030 8156 5714
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 8116 5024 8168 5030
rect 8116 4966 8168 4972
rect 7748 4208 7800 4214
rect 7748 4150 7800 4156
rect 7760 3670 7788 4150
rect 7944 4049 7972 4966
rect 8220 4554 8248 6054
rect 8312 4690 8340 7534
rect 8668 7268 8720 7274
rect 8668 7210 8720 7216
rect 8680 6458 8708 7210
rect 8772 6934 8800 12922
rect 8956 12540 9252 12560
rect 9012 12538 9036 12540
rect 9092 12538 9116 12540
rect 9172 12538 9196 12540
rect 9034 12486 9036 12538
rect 9098 12486 9110 12538
rect 9172 12486 9174 12538
rect 9012 12484 9036 12486
rect 9092 12484 9116 12486
rect 9172 12484 9196 12486
rect 8956 12464 9252 12484
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 9140 11694 9168 12038
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9324 11558 9352 18362
rect 9692 18086 9720 18838
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 9784 18426 9812 18702
rect 9772 18420 9824 18426
rect 9772 18362 9824 18368
rect 10324 18352 10376 18358
rect 10324 18294 10376 18300
rect 9956 18148 10008 18154
rect 9956 18090 10008 18096
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9692 17882 9720 18022
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9968 17814 9996 18090
rect 10232 17876 10284 17882
rect 10232 17818 10284 17824
rect 9956 17808 10008 17814
rect 9956 17750 10008 17756
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9496 16040 9548 16046
rect 9496 15982 9548 15988
rect 9508 15706 9536 15982
rect 9784 15978 9812 16526
rect 9772 15972 9824 15978
rect 9772 15914 9824 15920
rect 9784 15706 9812 15914
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9692 14822 9720 15506
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9692 14346 9720 14758
rect 9680 14340 9732 14346
rect 9680 14282 9732 14288
rect 9876 14006 9904 16934
rect 10244 16794 10272 17818
rect 10336 17746 10364 18294
rect 10324 17740 10376 17746
rect 10324 17682 10376 17688
rect 10336 17338 10364 17682
rect 10784 17672 10836 17678
rect 10784 17614 10836 17620
rect 10324 17332 10376 17338
rect 10324 17274 10376 17280
rect 10796 17202 10824 17614
rect 10888 17241 10916 23582
rect 11886 23582 12020 23610
rect 11886 23520 11942 23582
rect 11612 20256 11664 20262
rect 11612 20198 11664 20204
rect 11624 19854 11652 20198
rect 11704 19984 11756 19990
rect 11704 19926 11756 19932
rect 11612 19848 11664 19854
rect 11612 19790 11664 19796
rect 11624 19514 11652 19790
rect 11612 19508 11664 19514
rect 11612 19450 11664 19456
rect 11716 19378 11744 19926
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11612 19304 11664 19310
rect 11612 19246 11664 19252
rect 11624 18902 11652 19246
rect 11612 18896 11664 18902
rect 11612 18838 11664 18844
rect 11244 18760 11296 18766
rect 11244 18702 11296 18708
rect 11256 18426 11284 18702
rect 11624 18426 11652 18838
rect 11244 18420 11296 18426
rect 11244 18362 11296 18368
rect 11612 18420 11664 18426
rect 11612 18362 11664 18368
rect 11992 18358 12020 23582
rect 13174 23582 13308 23610
rect 13174 23520 13230 23582
rect 12956 21788 13252 21808
rect 13012 21786 13036 21788
rect 13092 21786 13116 21788
rect 13172 21786 13196 21788
rect 13034 21734 13036 21786
rect 13098 21734 13110 21786
rect 13172 21734 13174 21786
rect 13012 21732 13036 21734
rect 13092 21732 13116 21734
rect 13172 21732 13196 21734
rect 12956 21712 13252 21732
rect 13280 21146 13308 23582
rect 14200 23582 14518 23610
rect 13268 21140 13320 21146
rect 13268 21082 13320 21088
rect 12348 21004 12400 21010
rect 12348 20946 12400 20952
rect 12256 20460 12308 20466
rect 12256 20402 12308 20408
rect 12268 19718 12296 20402
rect 12360 20262 12388 20946
rect 12956 20700 13252 20720
rect 13012 20698 13036 20700
rect 13092 20698 13116 20700
rect 13172 20698 13196 20700
rect 13034 20646 13036 20698
rect 13098 20646 13110 20698
rect 13172 20646 13174 20698
rect 13012 20644 13036 20646
rect 13092 20644 13116 20646
rect 13172 20644 13196 20646
rect 12956 20624 13252 20644
rect 14200 20602 14228 23582
rect 14462 23520 14518 23582
rect 15396 23582 15714 23610
rect 14188 20596 14240 20602
rect 14188 20538 14240 20544
rect 13912 20392 13964 20398
rect 13912 20334 13964 20340
rect 12532 20324 12584 20330
rect 12532 20266 12584 20272
rect 12624 20324 12676 20330
rect 12624 20266 12676 20272
rect 12348 20256 12400 20262
rect 12348 20198 12400 20204
rect 12256 19712 12308 19718
rect 12256 19654 12308 19660
rect 12268 18902 12296 19654
rect 12256 18896 12308 18902
rect 12256 18838 12308 18844
rect 11980 18352 12032 18358
rect 11980 18294 12032 18300
rect 11152 18284 11204 18290
rect 11152 18226 11204 18232
rect 10874 17232 10930 17241
rect 10784 17196 10836 17202
rect 10874 17167 10930 17176
rect 10784 17138 10836 17144
rect 10232 16788 10284 16794
rect 10232 16730 10284 16736
rect 10244 16250 10272 16730
rect 10888 16658 10916 17167
rect 10876 16652 10928 16658
rect 10876 16594 10928 16600
rect 10232 16244 10284 16250
rect 10232 16186 10284 16192
rect 10244 15162 10272 16186
rect 10600 15972 10652 15978
rect 10600 15914 10652 15920
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10232 15156 10284 15162
rect 10232 15098 10284 15104
rect 9956 14952 10008 14958
rect 9956 14894 10008 14900
rect 9968 14618 9996 14894
rect 10244 14822 10272 15098
rect 10232 14816 10284 14822
rect 10232 14758 10284 14764
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 10244 14532 10272 14758
rect 10324 14544 10376 14550
rect 10244 14504 10324 14532
rect 10244 14074 10272 14504
rect 10324 14486 10376 14492
rect 10428 14482 10456 15438
rect 10416 14476 10468 14482
rect 10416 14418 10468 14424
rect 10612 14074 10640 15914
rect 11164 15502 11192 18226
rect 11244 18080 11296 18086
rect 11244 18022 11296 18028
rect 11980 18080 12032 18086
rect 11980 18022 12032 18028
rect 12256 18080 12308 18086
rect 12256 18022 12308 18028
rect 11256 16114 11284 18022
rect 11704 17808 11756 17814
rect 11704 17750 11756 17756
rect 11716 16998 11744 17750
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 11900 17202 11928 17614
rect 11888 17196 11940 17202
rect 11808 17156 11888 17184
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 11244 16108 11296 16114
rect 11244 16050 11296 16056
rect 11256 15706 11284 16050
rect 11244 15700 11296 15706
rect 11244 15642 11296 15648
rect 11612 15632 11664 15638
rect 11612 15574 11664 15580
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 11624 15162 11652 15574
rect 11612 15156 11664 15162
rect 11612 15098 11664 15104
rect 10876 14408 10928 14414
rect 10876 14350 10928 14356
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 9864 14000 9916 14006
rect 9864 13942 9916 13948
rect 9404 13796 9456 13802
rect 9404 13738 9456 13744
rect 9416 13705 9444 13738
rect 10244 13734 10272 14010
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10232 13728 10284 13734
rect 9402 13696 9458 13705
rect 10232 13670 10284 13676
rect 9402 13631 9458 13640
rect 10048 13456 10100 13462
rect 10244 13444 10272 13670
rect 10100 13416 10272 13444
rect 10048 13398 10100 13404
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9416 12782 9444 13126
rect 9692 12850 9720 13262
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 8956 11452 9252 11472
rect 9012 11450 9036 11452
rect 9092 11450 9116 11452
rect 9172 11450 9196 11452
rect 9034 11398 9036 11450
rect 9098 11398 9110 11450
rect 9172 11398 9174 11450
rect 9012 11396 9036 11398
rect 9092 11396 9116 11398
rect 9172 11396 9196 11398
rect 8956 11376 9252 11396
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8864 10606 8892 11290
rect 9416 11286 9444 12718
rect 10244 12646 10272 13416
rect 10520 13394 10548 13874
rect 10612 13530 10640 14010
rect 10888 13530 10916 14350
rect 11520 14000 11572 14006
rect 11334 13968 11390 13977
rect 11520 13942 11572 13948
rect 11334 13903 11390 13912
rect 10600 13524 10652 13530
rect 10600 13466 10652 13472
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10508 13388 10560 13394
rect 10508 13330 10560 13336
rect 10612 12986 10640 13466
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 10508 12708 10560 12714
rect 10508 12650 10560 12656
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 10416 12640 10468 12646
rect 10416 12582 10468 12588
rect 9588 11688 9640 11694
rect 9588 11630 9640 11636
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 9600 11354 9628 11630
rect 9588 11348 9640 11354
rect 9588 11290 9640 11296
rect 9404 11280 9456 11286
rect 9404 11222 9456 11228
rect 9968 10742 9996 11630
rect 10428 11286 10456 12582
rect 10520 11626 10548 12650
rect 10612 12646 10640 12922
rect 10876 12708 10928 12714
rect 10876 12650 10928 12656
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10888 12442 10916 12650
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 10600 12300 10652 12306
rect 10600 12242 10652 12248
rect 10508 11620 10560 11626
rect 10508 11562 10560 11568
rect 10416 11280 10468 11286
rect 10416 11222 10468 11228
rect 10428 10810 10456 11222
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 9956 10736 10008 10742
rect 9956 10678 10008 10684
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 9312 10600 9364 10606
rect 10336 10577 10364 10610
rect 9312 10542 9364 10548
rect 10322 10568 10378 10577
rect 8864 10266 8892 10542
rect 8956 10364 9252 10384
rect 9012 10362 9036 10364
rect 9092 10362 9116 10364
rect 9172 10362 9196 10364
rect 9034 10310 9036 10362
rect 9098 10310 9110 10362
rect 9172 10310 9174 10362
rect 9012 10308 9036 10310
rect 9092 10308 9116 10310
rect 9172 10308 9196 10310
rect 8956 10288 9252 10308
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 8864 9722 8892 10202
rect 9324 9926 9352 10542
rect 9496 10532 9548 10538
rect 10322 10503 10378 10512
rect 9496 10474 9548 10480
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9324 9761 9352 9862
rect 9310 9752 9366 9761
rect 8852 9716 8904 9722
rect 9310 9687 9366 9696
rect 8852 9658 8904 9664
rect 9324 9625 9352 9687
rect 9310 9616 9366 9625
rect 9310 9551 9366 9560
rect 9508 9518 9536 10474
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 8956 9276 9252 9296
rect 9012 9274 9036 9276
rect 9092 9274 9116 9276
rect 9172 9274 9196 9276
rect 9034 9222 9036 9274
rect 9098 9222 9110 9274
rect 9172 9222 9174 9274
rect 9012 9220 9036 9222
rect 9092 9220 9116 9222
rect 9172 9220 9196 9222
rect 8956 9200 9252 9220
rect 9508 9178 9536 9454
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 8850 9072 8906 9081
rect 9692 9042 9720 9386
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 8850 9007 8906 9016
rect 9680 9036 9732 9042
rect 8864 7546 8892 9007
rect 9680 8978 9732 8984
rect 8956 8188 9252 8208
rect 9012 8186 9036 8188
rect 9092 8186 9116 8188
rect 9172 8186 9196 8188
rect 9034 8134 9036 8186
rect 9098 8134 9110 8186
rect 9172 8134 9174 8186
rect 9012 8132 9036 8134
rect 9092 8132 9116 8134
rect 9172 8132 9196 8134
rect 8956 8112 9252 8132
rect 9692 8090 9720 8978
rect 10244 8838 10272 9318
rect 10428 9178 10456 10746
rect 10520 10606 10548 11562
rect 10612 11558 10640 12242
rect 11060 11824 11112 11830
rect 11060 11766 11112 11772
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10600 10736 10652 10742
rect 10600 10678 10652 10684
rect 10508 10600 10560 10606
rect 10508 10542 10560 10548
rect 10520 10266 10548 10542
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9404 7744 9456 7750
rect 9404 7686 9456 7692
rect 8852 7540 8904 7546
rect 8852 7482 8904 7488
rect 8850 7440 8906 7449
rect 8850 7375 8906 7384
rect 8864 7342 8892 7375
rect 9416 7342 9444 7686
rect 10244 7342 10272 8774
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 10232 7336 10284 7342
rect 10232 7278 10284 7284
rect 8956 7100 9252 7120
rect 9012 7098 9036 7100
rect 9092 7098 9116 7100
rect 9172 7098 9196 7100
rect 9034 7046 9036 7098
rect 9098 7046 9110 7098
rect 9172 7046 9174 7098
rect 9012 7044 9036 7046
rect 9092 7044 9116 7046
rect 9172 7044 9196 7046
rect 8956 7024 9252 7044
rect 8760 6928 8812 6934
rect 8760 6870 8812 6876
rect 8772 6458 8800 6870
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8760 6452 8812 6458
rect 8812 6412 8892 6440
rect 8760 6394 8812 6400
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8576 5092 8628 5098
rect 8496 5052 8576 5080
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8208 4548 8260 4554
rect 8208 4490 8260 4496
rect 8116 4480 8168 4486
rect 8116 4422 8168 4428
rect 7930 4040 7986 4049
rect 7930 3975 7986 3984
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 7748 3664 7800 3670
rect 7748 3606 7800 3612
rect 7840 3460 7892 3466
rect 7840 3402 7892 3408
rect 7852 2582 7880 3402
rect 8036 3058 8064 3878
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 7840 2576 7892 2582
rect 7840 2518 7892 2524
rect 8128 2446 8156 4422
rect 8220 4078 8248 4490
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 8312 3602 8340 4626
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8496 3126 8524 5052
rect 8576 5034 8628 5040
rect 8772 4282 8800 5646
rect 8760 4276 8812 4282
rect 8760 4218 8812 4224
rect 8772 4078 8800 4218
rect 8760 4072 8812 4078
rect 8760 4014 8812 4020
rect 8772 3738 8800 4014
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8484 3120 8536 3126
rect 8484 3062 8536 3068
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 7838 82 7894 480
rect 7668 54 7894 82
rect 7562 31 7618 40
rect 7838 0 7894 54
rect 8758 82 8814 480
rect 8864 82 8892 6412
rect 8956 6012 9252 6032
rect 9012 6010 9036 6012
rect 9092 6010 9116 6012
rect 9172 6010 9196 6012
rect 9034 5958 9036 6010
rect 9098 5958 9110 6010
rect 9172 5958 9174 6010
rect 9012 5956 9036 5958
rect 9092 5956 9116 5958
rect 9172 5956 9196 5958
rect 8956 5936 9252 5956
rect 8956 4924 9252 4944
rect 9012 4922 9036 4924
rect 9092 4922 9116 4924
rect 9172 4922 9196 4924
rect 9034 4870 9036 4922
rect 9098 4870 9110 4922
rect 9172 4870 9174 4922
rect 9012 4868 9036 4870
rect 9092 4868 9116 4870
rect 9172 4868 9196 4870
rect 8956 4848 9252 4868
rect 9416 4690 9444 7278
rect 10244 6186 10272 7278
rect 10336 6934 10364 8570
rect 10428 8362 10456 9114
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10520 7410 10548 7822
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10324 6928 10376 6934
rect 10324 6870 10376 6876
rect 10336 6458 10364 6870
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10140 6180 10192 6186
rect 10140 6122 10192 6128
rect 10232 6180 10284 6186
rect 10232 6122 10284 6128
rect 10152 5302 10180 6122
rect 10244 5914 10272 6122
rect 10232 5908 10284 5914
rect 10232 5850 10284 5856
rect 10336 5846 10364 6394
rect 10324 5840 10376 5846
rect 10244 5788 10324 5794
rect 10244 5782 10376 5788
rect 10244 5766 10364 5782
rect 10244 5370 10272 5766
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 10140 5296 10192 5302
rect 10140 5238 10192 5244
rect 9496 5160 9548 5166
rect 9496 5102 9548 5108
rect 9404 4684 9456 4690
rect 9404 4626 9456 4632
rect 9416 4214 9444 4626
rect 9404 4208 9456 4214
rect 9404 4150 9456 4156
rect 8956 3836 9252 3856
rect 9012 3834 9036 3836
rect 9092 3834 9116 3836
rect 9172 3834 9196 3836
rect 9034 3782 9036 3834
rect 9098 3782 9110 3834
rect 9172 3782 9174 3834
rect 9012 3780 9036 3782
rect 9092 3780 9116 3782
rect 9172 3780 9196 3782
rect 8956 3760 9252 3780
rect 9416 3738 9444 4150
rect 9508 4078 9536 5102
rect 10336 5098 10364 5646
rect 10612 5370 10640 10678
rect 10888 10470 10916 11086
rect 11072 10606 11100 11766
rect 11348 11694 11376 13903
rect 11532 12850 11560 13942
rect 11716 13814 11744 16934
rect 11808 16590 11836 17156
rect 11888 17138 11940 17144
rect 11888 16720 11940 16726
rect 11888 16662 11940 16668
rect 11796 16584 11848 16590
rect 11796 16526 11848 16532
rect 11808 16182 11836 16526
rect 11900 16250 11928 16662
rect 11888 16244 11940 16250
rect 11888 16186 11940 16192
rect 11796 16176 11848 16182
rect 11796 16118 11848 16124
rect 11796 15496 11848 15502
rect 11796 15438 11848 15444
rect 11808 15162 11836 15438
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 11808 13938 11836 15098
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 11716 13786 11836 13814
rect 11808 13705 11836 13786
rect 11794 13696 11850 13705
rect 11794 13631 11850 13640
rect 11808 13462 11836 13631
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11796 13456 11848 13462
rect 11796 13398 11848 13404
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 11624 12986 11652 13262
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11808 12918 11836 13398
rect 11796 12912 11848 12918
rect 11796 12854 11848 12860
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 11900 12306 11928 13466
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 11900 11898 11928 12242
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11336 11688 11388 11694
rect 11888 11688 11940 11694
rect 11336 11630 11388 11636
rect 11886 11656 11888 11665
rect 11940 11656 11942 11665
rect 11886 11591 11942 11600
rect 11900 11558 11928 11591
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 11888 11552 11940 11558
rect 11888 11494 11940 11500
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 10888 10266 10916 10406
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10692 9444 10744 9450
rect 10692 9386 10744 9392
rect 10704 9178 10732 9386
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 11072 8974 11100 10542
rect 11256 9042 11284 11494
rect 11992 11121 12020 18022
rect 12268 17610 12296 18022
rect 12256 17604 12308 17610
rect 12256 17546 12308 17552
rect 12164 17536 12216 17542
rect 12164 17478 12216 17484
rect 12176 17134 12204 17478
rect 12268 17338 12296 17546
rect 12256 17332 12308 17338
rect 12256 17274 12308 17280
rect 12164 17128 12216 17134
rect 12164 17070 12216 17076
rect 12176 16590 12204 17070
rect 12164 16584 12216 16590
rect 12164 16526 12216 16532
rect 12176 15502 12204 16526
rect 12360 15609 12388 20198
rect 12544 19446 12572 20266
rect 12636 19990 12664 20266
rect 12624 19984 12676 19990
rect 12624 19926 12676 19932
rect 13360 19984 13412 19990
rect 13360 19926 13412 19932
rect 12956 19612 13252 19632
rect 13012 19610 13036 19612
rect 13092 19610 13116 19612
rect 13172 19610 13196 19612
rect 13034 19558 13036 19610
rect 13098 19558 13110 19610
rect 13172 19558 13174 19610
rect 13012 19556 13036 19558
rect 13092 19556 13116 19558
rect 13172 19556 13196 19558
rect 12956 19536 13252 19556
rect 13372 19514 13400 19926
rect 13544 19848 13596 19854
rect 13544 19790 13596 19796
rect 13360 19508 13412 19514
rect 13360 19450 13412 19456
rect 12532 19440 12584 19446
rect 12532 19382 12584 19388
rect 13556 19242 13584 19790
rect 13924 19514 13952 20334
rect 14740 20256 14792 20262
rect 14740 20198 14792 20204
rect 13912 19508 13964 19514
rect 13912 19450 13964 19456
rect 14752 19446 14780 20198
rect 14740 19440 14792 19446
rect 14740 19382 14792 19388
rect 14004 19304 14056 19310
rect 14004 19246 14056 19252
rect 13544 19236 13596 19242
rect 13544 19178 13596 19184
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 12716 18828 12768 18834
rect 12716 18770 12768 18776
rect 12728 18086 12756 18770
rect 12820 18222 12848 19110
rect 13556 18970 13584 19178
rect 13544 18964 13596 18970
rect 13544 18906 13596 18912
rect 12956 18524 13252 18544
rect 13012 18522 13036 18524
rect 13092 18522 13116 18524
rect 13172 18522 13196 18524
rect 13034 18470 13036 18522
rect 13098 18470 13110 18522
rect 13172 18470 13174 18522
rect 13012 18468 13036 18470
rect 13092 18468 13116 18470
rect 13172 18468 13196 18470
rect 12956 18448 13252 18468
rect 12808 18216 12860 18222
rect 12808 18158 12860 18164
rect 13452 18148 13504 18154
rect 13452 18090 13504 18096
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12346 15600 12402 15609
rect 12346 15535 12402 15544
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12176 15026 12204 15438
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12164 15020 12216 15026
rect 12164 14962 12216 14968
rect 12544 14890 12572 15302
rect 12532 14884 12584 14890
rect 12452 14844 12532 14872
rect 12164 14816 12216 14822
rect 12164 14758 12216 14764
rect 12176 14618 12204 14758
rect 12164 14612 12216 14618
rect 12164 14554 12216 14560
rect 12452 14006 12480 14844
rect 12532 14826 12584 14832
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12440 14000 12492 14006
rect 12440 13942 12492 13948
rect 12452 13462 12480 13942
rect 12544 13802 12572 14214
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12636 13802 12664 14010
rect 12728 13977 12756 18022
rect 13360 17740 13412 17746
rect 13360 17682 13412 17688
rect 12956 17436 13252 17456
rect 13012 17434 13036 17436
rect 13092 17434 13116 17436
rect 13172 17434 13196 17436
rect 13034 17382 13036 17434
rect 13098 17382 13110 17434
rect 13172 17382 13174 17434
rect 13012 17380 13036 17382
rect 13092 17380 13116 17382
rect 13172 17380 13196 17382
rect 12956 17360 13252 17380
rect 13268 17264 13320 17270
rect 13268 17206 13320 17212
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 12820 16153 12848 16934
rect 12956 16348 13252 16368
rect 13012 16346 13036 16348
rect 13092 16346 13116 16348
rect 13172 16346 13196 16348
rect 13034 16294 13036 16346
rect 13098 16294 13110 16346
rect 13172 16294 13174 16346
rect 13012 16292 13036 16294
rect 13092 16292 13116 16294
rect 13172 16292 13196 16294
rect 12956 16272 13252 16292
rect 12806 16144 12862 16153
rect 12806 16079 12862 16088
rect 12808 16040 12860 16046
rect 12808 15982 12860 15988
rect 12820 14521 12848 15982
rect 12956 15260 13252 15280
rect 13012 15258 13036 15260
rect 13092 15258 13116 15260
rect 13172 15258 13196 15260
rect 13034 15206 13036 15258
rect 13098 15206 13110 15258
rect 13172 15206 13174 15258
rect 13012 15204 13036 15206
rect 13092 15204 13116 15206
rect 13172 15204 13196 15206
rect 12956 15184 13252 15204
rect 12806 14512 12862 14521
rect 13280 14482 13308 17206
rect 13372 17066 13400 17682
rect 13464 17377 13492 18090
rect 13728 18080 13780 18086
rect 13728 18022 13780 18028
rect 13740 17882 13768 18022
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13912 17536 13964 17542
rect 13912 17478 13964 17484
rect 13450 17368 13506 17377
rect 13450 17303 13506 17312
rect 13924 17134 13952 17478
rect 13912 17128 13964 17134
rect 13912 17070 13964 17076
rect 13360 17060 13412 17066
rect 13360 17002 13412 17008
rect 12806 14447 12862 14456
rect 13268 14476 13320 14482
rect 12714 13968 12770 13977
rect 12714 13903 12770 13912
rect 12532 13796 12584 13802
rect 12532 13738 12584 13744
rect 12624 13796 12676 13802
rect 12624 13738 12676 13744
rect 12440 13456 12492 13462
rect 12440 13398 12492 13404
rect 12440 12368 12492 12374
rect 12440 12310 12492 12316
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 12084 11830 12112 12242
rect 12164 12232 12216 12238
rect 12164 12174 12216 12180
rect 12072 11824 12124 11830
rect 12072 11766 12124 11772
rect 12176 11218 12204 12174
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 12256 11280 12308 11286
rect 12256 11222 12308 11228
rect 12164 11212 12216 11218
rect 12164 11154 12216 11160
rect 11978 11112 12034 11121
rect 11978 11047 12034 11056
rect 12176 10810 12204 11154
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12268 10470 12296 11222
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 11428 10192 11480 10198
rect 11428 10134 11480 10140
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11348 9450 11376 9998
rect 11440 9722 11468 10134
rect 11612 10056 11664 10062
rect 11612 9998 11664 10004
rect 11428 9716 11480 9722
rect 11428 9658 11480 9664
rect 11336 9444 11388 9450
rect 11336 9386 11388 9392
rect 11348 9110 11376 9386
rect 11336 9104 11388 9110
rect 11336 9046 11388 9052
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 11060 8968 11112 8974
rect 11256 8945 11284 8978
rect 11060 8910 11112 8916
rect 11242 8936 11298 8945
rect 10692 8900 10744 8906
rect 10692 8842 10744 8848
rect 10600 5364 10652 5370
rect 10600 5306 10652 5312
rect 10612 5166 10640 5306
rect 10600 5160 10652 5166
rect 10600 5102 10652 5108
rect 10324 5092 10376 5098
rect 10324 5034 10376 5040
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 9508 3670 9536 4014
rect 9600 3942 9628 4082
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 9496 3664 9548 3670
rect 9496 3606 9548 3612
rect 9692 3534 9720 4762
rect 10704 4690 10732 8842
rect 11072 7954 11100 8910
rect 11242 8871 11298 8880
rect 11256 8498 11284 8871
rect 11440 8634 11468 9658
rect 11624 9586 11652 9998
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 12268 9110 12296 10406
rect 12256 9104 12308 9110
rect 12256 9046 12308 9052
rect 11428 8628 11480 8634
rect 11428 8570 11480 8576
rect 12268 8498 12296 9046
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 12268 8022 12296 8434
rect 12256 8016 12308 8022
rect 12256 7958 12308 7964
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 11072 7546 11100 7890
rect 11428 7880 11480 7886
rect 11428 7822 11480 7828
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11440 7546 11468 7822
rect 11808 7546 11836 7822
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 11428 7540 11480 7546
rect 11428 7482 11480 7488
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10784 6724 10836 6730
rect 10784 6666 10836 6672
rect 10796 6322 10824 6666
rect 10980 6322 11008 7346
rect 12360 6934 12388 11290
rect 12452 9518 12480 12310
rect 12544 9908 12572 13738
rect 12820 12374 12848 14447
rect 13268 14418 13320 14424
rect 12956 14172 13252 14192
rect 13012 14170 13036 14172
rect 13092 14170 13116 14172
rect 13172 14170 13196 14172
rect 13034 14118 13036 14170
rect 13098 14118 13110 14170
rect 13172 14118 13174 14170
rect 13012 14116 13036 14118
rect 13092 14116 13116 14118
rect 13172 14116 13196 14118
rect 12956 14096 13252 14116
rect 13280 14006 13308 14418
rect 13268 14000 13320 14006
rect 13268 13942 13320 13948
rect 13372 13814 13400 17002
rect 13924 16658 13952 17070
rect 13544 16652 13596 16658
rect 13544 16594 13596 16600
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 13464 16250 13492 16390
rect 13452 16244 13504 16250
rect 13452 16186 13504 16192
rect 13464 15978 13492 16186
rect 13452 15972 13504 15978
rect 13452 15914 13504 15920
rect 13556 15910 13584 16594
rect 13924 16454 13952 16594
rect 13912 16448 13964 16454
rect 13912 16390 13964 16396
rect 14016 16266 14044 19246
rect 14096 18828 14148 18834
rect 14096 18770 14148 18776
rect 14108 18154 14136 18770
rect 14188 18216 14240 18222
rect 14188 18158 14240 18164
rect 14096 18148 14148 18154
rect 14096 18090 14148 18096
rect 14200 17542 14228 18158
rect 14832 18148 14884 18154
rect 14832 18090 14884 18096
rect 14188 17536 14240 17542
rect 14188 17478 14240 17484
rect 14200 17202 14228 17478
rect 14844 17338 14872 18090
rect 15108 18080 15160 18086
rect 15160 18040 15240 18068
rect 15108 18022 15160 18028
rect 15212 17746 15240 18040
rect 15200 17740 15252 17746
rect 15200 17682 15252 17688
rect 14924 17536 14976 17542
rect 14924 17478 14976 17484
rect 14832 17332 14884 17338
rect 14832 17274 14884 17280
rect 14188 17196 14240 17202
rect 14188 17138 14240 17144
rect 14844 17066 14872 17274
rect 14832 17060 14884 17066
rect 14832 17002 14884 17008
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 13924 16238 14044 16266
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13372 13786 13492 13814
rect 12956 13084 13252 13104
rect 13012 13082 13036 13084
rect 13092 13082 13116 13084
rect 13172 13082 13196 13084
rect 13034 13030 13036 13082
rect 13098 13030 13110 13082
rect 13172 13030 13174 13082
rect 13012 13028 13036 13030
rect 13092 13028 13116 13030
rect 13172 13028 13196 13030
rect 12956 13008 13252 13028
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 12808 12368 12860 12374
rect 12808 12310 12860 12316
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12624 11824 12676 11830
rect 12624 11766 12676 11772
rect 12636 10538 12664 11766
rect 12728 11762 12756 12038
rect 12716 11756 12768 11762
rect 12716 11698 12768 11704
rect 12820 11626 12848 12174
rect 12956 11996 13252 12016
rect 13012 11994 13036 11996
rect 13092 11994 13116 11996
rect 13172 11994 13196 11996
rect 13034 11942 13036 11994
rect 13098 11942 13110 11994
rect 13172 11942 13174 11994
rect 13012 11940 13036 11942
rect 13092 11940 13116 11942
rect 13172 11940 13196 11942
rect 12956 11920 13252 11940
rect 12808 11620 12860 11626
rect 12808 11562 12860 11568
rect 12820 11354 12848 11562
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12820 10520 12848 10950
rect 12956 10908 13252 10928
rect 13012 10906 13036 10908
rect 13092 10906 13116 10908
rect 13172 10906 13196 10908
rect 13034 10854 13036 10906
rect 13098 10854 13110 10906
rect 13172 10854 13174 10906
rect 13012 10852 13036 10854
rect 13092 10852 13116 10854
rect 13172 10852 13196 10854
rect 12956 10832 13252 10852
rect 12900 10532 12952 10538
rect 12820 10492 12900 10520
rect 12636 10062 12664 10474
rect 12820 10266 12848 10492
rect 12900 10474 12952 10480
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12544 9880 12848 9908
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12728 9042 12756 9318
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12728 8634 12756 8978
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 12636 7546 12664 7958
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12348 6928 12400 6934
rect 12348 6870 12400 6876
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 11072 6458 11100 6734
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 10980 5846 11008 6258
rect 12268 5914 12296 6734
rect 12360 6458 12388 6870
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 12360 6118 12388 6394
rect 12624 6180 12676 6186
rect 12624 6122 12676 6128
rect 12348 6112 12400 6118
rect 12348 6054 12400 6060
rect 12256 5908 12308 5914
rect 12256 5850 12308 5856
rect 10968 5840 11020 5846
rect 10968 5782 11020 5788
rect 12636 5574 12664 6122
rect 12624 5568 12676 5574
rect 12624 5510 12676 5516
rect 12636 5137 12664 5510
rect 12716 5160 12768 5166
rect 12622 5128 12678 5137
rect 10784 5092 10836 5098
rect 10784 5034 10836 5040
rect 12440 5092 12492 5098
rect 12716 5102 12768 5108
rect 12622 5063 12678 5072
rect 12440 5034 12492 5040
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 10692 4684 10744 4690
rect 10692 4626 10744 4632
rect 9772 4004 9824 4010
rect 9772 3946 9824 3952
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9692 3194 9720 3470
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9588 3120 9640 3126
rect 9588 3062 9640 3068
rect 8956 2748 9252 2768
rect 9012 2746 9036 2748
rect 9092 2746 9116 2748
rect 9172 2746 9196 2748
rect 9034 2694 9036 2746
rect 9098 2694 9110 2746
rect 9172 2694 9174 2746
rect 9012 2692 9036 2694
rect 9092 2692 9116 2694
rect 9172 2692 9196 2694
rect 8956 2672 9252 2692
rect 8758 54 8892 82
rect 9600 82 9628 3062
rect 9784 2922 9812 3946
rect 10428 3942 10456 4626
rect 10704 4214 10732 4626
rect 10796 4622 10824 5034
rect 11888 4820 11940 4826
rect 11888 4762 11940 4768
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 10796 4282 10824 4558
rect 10784 4276 10836 4282
rect 10784 4218 10836 4224
rect 10692 4208 10744 4214
rect 10692 4150 10744 4156
rect 11624 4146 11652 4558
rect 11612 4140 11664 4146
rect 11612 4082 11664 4088
rect 10600 4072 10652 4078
rect 10600 4014 10652 4020
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 9772 2916 9824 2922
rect 9772 2858 9824 2864
rect 9968 2854 9996 3606
rect 10612 3398 10640 4014
rect 11796 3664 11848 3670
rect 11796 3606 11848 3612
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 10324 2916 10376 2922
rect 10324 2858 10376 2864
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 10336 2446 10364 2858
rect 10612 2582 10640 3334
rect 11164 2990 11192 3334
rect 11152 2984 11204 2990
rect 11152 2926 11204 2932
rect 11164 2650 11192 2926
rect 11808 2854 11836 3606
rect 11900 3534 11928 4762
rect 12256 4684 12308 4690
rect 12256 4626 12308 4632
rect 12072 3936 12124 3942
rect 12072 3878 12124 3884
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11796 2848 11848 2854
rect 11796 2790 11848 2796
rect 11900 2650 11928 3470
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 12084 2582 12112 3878
rect 12268 3738 12296 4626
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 12452 2650 12480 5034
rect 12728 3738 12756 5102
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 12624 3460 12676 3466
rect 12624 3402 12676 3408
rect 12636 3058 12664 3402
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 12728 2922 12756 3674
rect 12820 3641 12848 9880
rect 12956 9820 13252 9840
rect 13012 9818 13036 9820
rect 13092 9818 13116 9820
rect 13172 9818 13196 9820
rect 13034 9766 13036 9818
rect 13098 9766 13110 9818
rect 13172 9766 13174 9818
rect 13012 9764 13036 9766
rect 13092 9764 13116 9766
rect 13172 9764 13196 9766
rect 12956 9744 13252 9764
rect 12900 9512 12952 9518
rect 12900 9454 12952 9460
rect 12912 8974 12940 9454
rect 13280 8974 13308 10066
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 12956 8732 13252 8752
rect 13012 8730 13036 8732
rect 13092 8730 13116 8732
rect 13172 8730 13196 8732
rect 13034 8678 13036 8730
rect 13098 8678 13110 8730
rect 13172 8678 13174 8730
rect 13012 8676 13036 8678
rect 13092 8676 13116 8678
rect 13172 8676 13196 8678
rect 12956 8656 13252 8676
rect 13268 7812 13320 7818
rect 13268 7754 13320 7760
rect 12956 7644 13252 7664
rect 13012 7642 13036 7644
rect 13092 7642 13116 7644
rect 13172 7642 13196 7644
rect 13034 7590 13036 7642
rect 13098 7590 13110 7642
rect 13172 7590 13174 7642
rect 13012 7588 13036 7590
rect 13092 7588 13116 7590
rect 13172 7588 13196 7590
rect 12956 7568 13252 7588
rect 13280 7410 13308 7754
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 13280 7274 13308 7346
rect 13372 7313 13400 12718
rect 13464 11558 13492 13786
rect 13556 13530 13584 15846
rect 13636 15564 13688 15570
rect 13636 15506 13688 15512
rect 13648 14822 13676 15506
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 13648 14346 13676 14758
rect 13636 14340 13688 14346
rect 13636 14282 13688 14288
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13556 12986 13584 13466
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13556 12782 13584 12922
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 13648 12306 13676 14282
rect 13636 12300 13688 12306
rect 13636 12242 13688 12248
rect 13648 11898 13676 12242
rect 13636 11892 13688 11898
rect 13636 11834 13688 11840
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13924 10538 13952 16238
rect 14384 16182 14412 16526
rect 14372 16176 14424 16182
rect 14372 16118 14424 16124
rect 14648 16040 14700 16046
rect 14648 15982 14700 15988
rect 14004 15904 14056 15910
rect 14004 15846 14056 15852
rect 14016 14521 14044 15846
rect 14554 15600 14610 15609
rect 14188 15564 14240 15570
rect 14660 15570 14688 15982
rect 14554 15535 14610 15544
rect 14648 15564 14700 15570
rect 14188 15506 14240 15512
rect 14200 15162 14228 15506
rect 14370 15464 14426 15473
rect 14370 15399 14426 15408
rect 14188 15156 14240 15162
rect 14188 15098 14240 15104
rect 14002 14512 14058 14521
rect 14002 14447 14058 14456
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 14108 13938 14136 14350
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 14108 13530 14136 13874
rect 14096 13524 14148 13530
rect 14096 13466 14148 13472
rect 14096 13184 14148 13190
rect 14096 13126 14148 13132
rect 14108 12782 14136 13126
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14108 12306 14136 12718
rect 14096 12300 14148 12306
rect 14096 12242 14148 12248
rect 14004 11552 14056 11558
rect 14004 11494 14056 11500
rect 14016 11354 14044 11494
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 13452 10532 13504 10538
rect 13452 10474 13504 10480
rect 13912 10532 13964 10538
rect 13912 10474 13964 10480
rect 14004 10532 14056 10538
rect 14004 10474 14056 10480
rect 13464 8498 13492 10474
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13556 9654 13584 10066
rect 13912 9988 13964 9994
rect 14016 9976 14044 10474
rect 14200 10198 14228 15098
rect 14384 15026 14412 15399
rect 14372 15020 14424 15026
rect 14372 14962 14424 14968
rect 14384 14618 14412 14962
rect 14464 14952 14516 14958
rect 14464 14894 14516 14900
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 14476 14346 14504 14894
rect 14464 14340 14516 14346
rect 14464 14282 14516 14288
rect 14464 12300 14516 12306
rect 14464 12242 14516 12248
rect 14476 11694 14504 12242
rect 14464 11688 14516 11694
rect 14464 11630 14516 11636
rect 14476 11082 14504 11630
rect 14464 11076 14516 11082
rect 14464 11018 14516 11024
rect 14188 10192 14240 10198
rect 14188 10134 14240 10140
rect 13964 9948 14044 9976
rect 13912 9930 13964 9936
rect 13544 9648 13596 9654
rect 13544 9590 13596 9596
rect 13556 8922 13584 9590
rect 13820 9376 13872 9382
rect 13924 9364 13952 9930
rect 14568 9654 14596 15535
rect 14648 15506 14700 15512
rect 14740 14884 14792 14890
rect 14740 14826 14792 14832
rect 14752 14482 14780 14826
rect 14740 14476 14792 14482
rect 14740 14418 14792 14424
rect 14740 14272 14792 14278
rect 14740 14214 14792 14220
rect 14752 13190 14780 14214
rect 14740 13184 14792 13190
rect 14740 13126 14792 13132
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 14844 9654 14872 9862
rect 14556 9648 14608 9654
rect 14832 9648 14884 9654
rect 14556 9590 14608 9596
rect 14830 9616 14832 9625
rect 14884 9616 14886 9625
rect 14568 9518 14596 9590
rect 14830 9551 14886 9560
rect 14844 9525 14872 9551
rect 14556 9512 14608 9518
rect 14556 9454 14608 9460
rect 13872 9336 13952 9364
rect 13820 9318 13872 9324
rect 13556 8894 13768 8922
rect 13636 8832 13688 8838
rect 13636 8774 13688 8780
rect 13544 8560 13596 8566
rect 13544 8502 13596 8508
rect 13452 8492 13504 8498
rect 13452 8434 13504 8440
rect 13464 7478 13492 8434
rect 13556 7750 13584 8502
rect 13648 8362 13676 8774
rect 13636 8356 13688 8362
rect 13636 8298 13688 8304
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13452 7472 13504 7478
rect 13452 7414 13504 7420
rect 13358 7304 13414 7313
rect 12900 7268 12952 7274
rect 12900 7210 12952 7216
rect 13268 7268 13320 7274
rect 13358 7239 13414 7248
rect 13268 7210 13320 7216
rect 12912 6730 12940 7210
rect 12900 6724 12952 6730
rect 12900 6666 12952 6672
rect 12956 6556 13252 6576
rect 13012 6554 13036 6556
rect 13092 6554 13116 6556
rect 13172 6554 13196 6556
rect 13034 6502 13036 6554
rect 13098 6502 13110 6554
rect 13172 6502 13174 6554
rect 13012 6500 13036 6502
rect 13092 6500 13116 6502
rect 13172 6500 13196 6502
rect 12956 6480 13252 6500
rect 13556 6322 13584 7686
rect 13740 6610 13768 8894
rect 13648 6582 13768 6610
rect 13648 6322 13676 6582
rect 13832 6474 13860 9318
rect 14568 7410 14596 9454
rect 14740 9172 14792 9178
rect 14740 9114 14792 9120
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 14002 7304 14058 7313
rect 14002 7239 14058 7248
rect 14016 6866 14044 7239
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 13740 6446 13860 6474
rect 14016 6458 14044 6802
rect 14556 6724 14608 6730
rect 14556 6666 14608 6672
rect 14188 6656 14240 6662
rect 14188 6598 14240 6604
rect 14004 6452 14056 6458
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 12956 5468 13252 5488
rect 13012 5466 13036 5468
rect 13092 5466 13116 5468
rect 13172 5466 13196 5468
rect 13034 5414 13036 5466
rect 13098 5414 13110 5466
rect 13172 5414 13174 5466
rect 13012 5412 13036 5414
rect 13092 5412 13116 5414
rect 13172 5412 13196 5414
rect 12956 5392 13252 5412
rect 13740 5098 13768 6446
rect 14004 6394 14056 6400
rect 14200 6254 14228 6598
rect 14188 6248 14240 6254
rect 14188 6190 14240 6196
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 14016 5166 14044 6054
rect 14200 5642 14228 6190
rect 14188 5636 14240 5642
rect 14188 5578 14240 5584
rect 14004 5160 14056 5166
rect 14004 5102 14056 5108
rect 13268 5092 13320 5098
rect 13268 5034 13320 5040
rect 13728 5092 13780 5098
rect 13728 5034 13780 5040
rect 13280 4758 13308 5034
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13268 4752 13320 4758
rect 13268 4694 13320 4700
rect 13176 4684 13228 4690
rect 13176 4626 13228 4632
rect 13188 4554 13216 4626
rect 13176 4548 13228 4554
rect 13176 4490 13228 4496
rect 12956 4380 13252 4400
rect 13012 4378 13036 4380
rect 13092 4378 13116 4380
rect 13172 4378 13196 4380
rect 13034 4326 13036 4378
rect 13098 4326 13110 4378
rect 13172 4326 13174 4378
rect 13012 4324 13036 4326
rect 13092 4324 13116 4326
rect 13172 4324 13196 4326
rect 12956 4304 13252 4324
rect 13280 4010 13308 4694
rect 13832 4078 13860 4762
rect 14200 4622 14228 5578
rect 14188 4616 14240 4622
rect 14188 4558 14240 4564
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 14096 4480 14148 4486
rect 14096 4422 14148 4428
rect 13360 4072 13412 4078
rect 13360 4014 13412 4020
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 13268 4004 13320 4010
rect 13268 3946 13320 3952
rect 13372 3738 13400 4014
rect 13360 3732 13412 3738
rect 13360 3674 13412 3680
rect 12806 3632 12862 3641
rect 12806 3567 12862 3576
rect 12956 3292 13252 3312
rect 13012 3290 13036 3292
rect 13092 3290 13116 3292
rect 13172 3290 13196 3292
rect 13034 3238 13036 3290
rect 13098 3238 13110 3290
rect 13172 3238 13174 3290
rect 13012 3236 13036 3238
rect 13092 3236 13116 3238
rect 13172 3236 13196 3238
rect 12956 3216 13252 3236
rect 13372 3058 13400 3674
rect 13452 3596 13504 3602
rect 13452 3538 13504 3544
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 12716 2916 12768 2922
rect 12716 2858 12768 2864
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 10600 2576 10652 2582
rect 10600 2518 10652 2524
rect 12072 2576 12124 2582
rect 12072 2518 12124 2524
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10508 2372 10560 2378
rect 10508 2314 10560 2320
rect 9678 82 9734 480
rect 9600 54 9734 82
rect 10520 82 10548 2314
rect 12956 2204 13252 2224
rect 13012 2202 13036 2204
rect 13092 2202 13116 2204
rect 13172 2202 13196 2204
rect 13034 2150 13036 2202
rect 13098 2150 13110 2202
rect 13172 2150 13174 2202
rect 13012 2148 13036 2150
rect 13092 2148 13116 2150
rect 13172 2148 13196 2150
rect 12956 2128 13252 2148
rect 12164 2100 12216 2106
rect 12164 2042 12216 2048
rect 10598 82 10654 480
rect 10520 54 10654 82
rect 8758 0 8814 54
rect 9678 0 9734 54
rect 10598 0 10654 54
rect 11518 128 11574 480
rect 11518 76 11520 128
rect 11572 76 11574 128
rect 11518 0 11574 76
rect 12176 82 12204 2042
rect 12438 82 12494 480
rect 13280 134 13308 2586
rect 13372 2582 13400 2994
rect 13360 2576 13412 2582
rect 13360 2518 13412 2524
rect 12176 54 12494 82
rect 13268 128 13320 134
rect 13268 70 13320 76
rect 13358 82 13414 480
rect 13464 82 13492 3538
rect 14108 2514 14136 4422
rect 14384 4078 14412 4558
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14280 3596 14332 3602
rect 14280 3538 14332 3544
rect 14292 3194 14320 3538
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14464 3120 14516 3126
rect 14464 3062 14516 3068
rect 14476 2854 14504 3062
rect 14464 2848 14516 2854
rect 14464 2790 14516 2796
rect 14096 2508 14148 2514
rect 14096 2450 14148 2456
rect 12438 0 12494 54
rect 13358 54 13492 82
rect 14278 82 14334 480
rect 14568 82 14596 6666
rect 14752 5234 14780 9114
rect 14830 7440 14886 7449
rect 14830 7375 14886 7384
rect 14844 7342 14872 7375
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 14844 7002 14872 7278
rect 14832 6996 14884 7002
rect 14832 6938 14884 6944
rect 14844 6390 14872 6938
rect 14832 6384 14884 6390
rect 14832 6326 14884 6332
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 14752 4826 14780 5170
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 14752 3738 14780 3878
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 14752 3058 14780 3674
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 14936 2922 14964 17478
rect 15212 17338 15240 17682
rect 15200 17332 15252 17338
rect 15200 17274 15252 17280
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 15304 16250 15332 16594
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 15304 15026 15332 16186
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 15016 14612 15068 14618
rect 15016 14554 15068 14560
rect 15028 13734 15056 14554
rect 15396 13734 15424 23582
rect 15658 23520 15714 23582
rect 16684 23582 17002 23610
rect 16396 20324 16448 20330
rect 16396 20266 16448 20272
rect 15844 19916 15896 19922
rect 15844 19858 15896 19864
rect 15660 19304 15712 19310
rect 15660 19246 15712 19252
rect 15476 18896 15528 18902
rect 15476 18838 15528 18844
rect 15488 18154 15516 18838
rect 15568 18216 15620 18222
rect 15672 18193 15700 19246
rect 15856 19174 15884 19858
rect 16304 19712 16356 19718
rect 16304 19654 16356 19660
rect 16212 19372 16264 19378
rect 16212 19314 16264 19320
rect 15844 19168 15896 19174
rect 15764 19128 15844 19156
rect 15764 18329 15792 19128
rect 15844 19110 15896 19116
rect 16224 18970 16252 19314
rect 16212 18964 16264 18970
rect 16212 18906 16264 18912
rect 16316 18902 16344 19654
rect 16304 18896 16356 18902
rect 16304 18838 16356 18844
rect 15844 18760 15896 18766
rect 15844 18702 15896 18708
rect 15750 18320 15806 18329
rect 15750 18255 15806 18264
rect 15568 18158 15620 18164
rect 15658 18184 15714 18193
rect 15476 18148 15528 18154
rect 15476 18090 15528 18096
rect 15016 13728 15068 13734
rect 15016 13670 15068 13676
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 15384 13728 15436 13734
rect 15384 13670 15436 13676
rect 15304 12714 15332 13670
rect 15580 13394 15608 18158
rect 15658 18119 15714 18128
rect 15672 15552 15700 18119
rect 15856 18086 15884 18702
rect 16408 18358 16436 20266
rect 16580 19712 16632 19718
rect 16580 19654 16632 19660
rect 16592 19242 16620 19654
rect 16488 19236 16540 19242
rect 16488 19178 16540 19184
rect 16580 19236 16632 19242
rect 16580 19178 16632 19184
rect 16500 18970 16528 19178
rect 16488 18964 16540 18970
rect 16488 18906 16540 18912
rect 16592 18426 16620 19178
rect 16580 18420 16632 18426
rect 16580 18362 16632 18368
rect 16396 18352 16448 18358
rect 16396 18294 16448 18300
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 15856 17814 15884 18022
rect 15844 17808 15896 17814
rect 15844 17750 15896 17756
rect 15752 17536 15804 17542
rect 15752 17478 15804 17484
rect 15764 17202 15792 17478
rect 15752 17196 15804 17202
rect 15752 17138 15804 17144
rect 15764 16794 15792 17138
rect 16028 17060 16080 17066
rect 16028 17002 16080 17008
rect 15752 16788 15804 16794
rect 15752 16730 15804 16736
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 15764 16046 15792 16594
rect 16040 16250 16068 17002
rect 16028 16244 16080 16250
rect 16028 16186 16080 16192
rect 15752 16040 15804 16046
rect 15752 15982 15804 15988
rect 16040 15978 16068 16186
rect 16212 16040 16264 16046
rect 16212 15982 16264 15988
rect 16578 16008 16634 16017
rect 16028 15972 16080 15978
rect 16028 15914 16080 15920
rect 16224 15638 16252 15982
rect 16578 15943 16634 15952
rect 16592 15706 16620 15943
rect 16580 15700 16632 15706
rect 16580 15642 16632 15648
rect 16212 15632 16264 15638
rect 16212 15574 16264 15580
rect 15752 15564 15804 15570
rect 15672 15524 15752 15552
rect 15752 15506 15804 15512
rect 15764 15162 15792 15506
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 16396 15020 16448 15026
rect 16316 14980 16396 15008
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 16224 14618 16252 14758
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15672 14074 15700 14418
rect 16224 14074 16252 14554
rect 16316 14346 16344 14980
rect 16396 14962 16448 14968
rect 16500 14414 16528 15302
rect 16592 15094 16620 15642
rect 16580 15088 16632 15094
rect 16580 15030 16632 15036
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 16304 14340 16356 14346
rect 16304 14282 16356 14288
rect 15660 14068 15712 14074
rect 15660 14010 15712 14016
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 15568 13388 15620 13394
rect 15568 13330 15620 13336
rect 15292 12708 15344 12714
rect 15292 12650 15344 12656
rect 15580 12646 15608 13330
rect 16028 12708 16080 12714
rect 16028 12650 16080 12656
rect 15568 12640 15620 12646
rect 15568 12582 15620 12588
rect 15016 10600 15068 10606
rect 15016 10542 15068 10548
rect 15028 9518 15056 10542
rect 15476 10124 15528 10130
rect 15476 10066 15528 10072
rect 15384 9580 15436 9586
rect 15488 9568 15516 10066
rect 15436 9540 15516 9568
rect 15384 9522 15436 9528
rect 15016 9512 15068 9518
rect 15016 9454 15068 9460
rect 15028 9178 15056 9454
rect 15108 9376 15160 9382
rect 15108 9318 15160 9324
rect 15016 9172 15068 9178
rect 15016 9114 15068 9120
rect 15014 9072 15070 9081
rect 15120 9058 15148 9318
rect 15488 9178 15516 9540
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 15580 9058 15608 12582
rect 16040 12374 16068 12650
rect 16028 12368 16080 12374
rect 16028 12310 16080 12316
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15764 11898 15792 12174
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 16040 11830 16068 12310
rect 16316 12084 16344 14282
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16592 13802 16620 14010
rect 16488 13796 16540 13802
rect 16488 13738 16540 13744
rect 16580 13796 16632 13802
rect 16580 13738 16632 13744
rect 16500 13190 16528 13738
rect 16488 13184 16540 13190
rect 16488 13126 16540 13132
rect 16488 12096 16540 12102
rect 16316 12056 16488 12084
rect 16488 12038 16540 12044
rect 16028 11824 16080 11830
rect 16028 11766 16080 11772
rect 16040 11354 16068 11766
rect 16500 11626 16528 12038
rect 16488 11620 16540 11626
rect 16488 11562 16540 11568
rect 16580 11620 16632 11626
rect 16580 11562 16632 11568
rect 16304 11552 16356 11558
rect 16304 11494 16356 11500
rect 16316 11354 16344 11494
rect 16592 11354 16620 11562
rect 16028 11348 16080 11354
rect 16028 11290 16080 11296
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16580 11348 16632 11354
rect 16580 11290 16632 11296
rect 15660 11144 15712 11150
rect 15660 11086 15712 11092
rect 15672 10538 15700 11086
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 15660 10532 15712 10538
rect 15660 10474 15712 10480
rect 15672 10266 15700 10474
rect 15660 10260 15712 10266
rect 15660 10202 15712 10208
rect 15856 10130 15884 11018
rect 15936 11008 15988 11014
rect 15936 10950 15988 10956
rect 15948 10606 15976 10950
rect 15936 10600 15988 10606
rect 15936 10542 15988 10548
rect 15844 10124 15896 10130
rect 15844 10066 15896 10072
rect 15070 9030 15148 9058
rect 15488 9030 15608 9058
rect 15014 9007 15070 9016
rect 15028 8974 15056 9007
rect 15016 8968 15068 8974
rect 15016 8910 15068 8916
rect 15384 8288 15436 8294
rect 15384 8230 15436 8236
rect 15396 8090 15424 8230
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 15304 7342 15332 7890
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15304 6866 15332 7278
rect 15292 6860 15344 6866
rect 15292 6802 15344 6808
rect 15304 6118 15332 6802
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 15016 5568 15068 5574
rect 15016 5510 15068 5516
rect 15028 3738 15056 5510
rect 15120 5030 15148 5714
rect 15108 5024 15160 5030
rect 15108 4966 15160 4972
rect 15016 3732 15068 3738
rect 15016 3674 15068 3680
rect 14924 2916 14976 2922
rect 14924 2858 14976 2864
rect 14278 54 14596 82
rect 15120 82 15148 4966
rect 15488 4185 15516 9030
rect 15856 8838 15884 10066
rect 15948 9518 15976 10542
rect 16040 10266 16068 11290
rect 16304 10600 16356 10606
rect 16304 10542 16356 10548
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 15936 9512 15988 9518
rect 15936 9454 15988 9460
rect 15844 8832 15896 8838
rect 15844 8774 15896 8780
rect 15752 7948 15804 7954
rect 15752 7890 15804 7896
rect 15764 7002 15792 7890
rect 15752 6996 15804 7002
rect 15752 6938 15804 6944
rect 15764 6458 15792 6938
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15856 6254 15884 8774
rect 15948 7954 15976 9454
rect 16028 9376 16080 9382
rect 16028 9318 16080 9324
rect 16040 8974 16068 9318
rect 16212 9104 16264 9110
rect 16212 9046 16264 9052
rect 16028 8968 16080 8974
rect 16028 8910 16080 8916
rect 16040 8634 16068 8910
rect 16028 8628 16080 8634
rect 16028 8570 16080 8576
rect 16224 8498 16252 9046
rect 16212 8492 16264 8498
rect 16212 8434 16264 8440
rect 16210 7984 16266 7993
rect 15936 7948 15988 7954
rect 16316 7954 16344 10542
rect 16488 9512 16540 9518
rect 16488 9454 16540 9460
rect 16210 7919 16266 7928
rect 16304 7948 16356 7954
rect 15936 7890 15988 7896
rect 15948 7546 15976 7890
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 15948 6866 15976 7482
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 15948 6322 15976 6802
rect 15936 6316 15988 6322
rect 15936 6258 15988 6264
rect 15844 6248 15896 6254
rect 15844 6190 15896 6196
rect 16120 5636 16172 5642
rect 16120 5578 16172 5584
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 15672 5166 15700 5510
rect 16132 5166 16160 5578
rect 15568 5160 15620 5166
rect 15568 5102 15620 5108
rect 15660 5160 15712 5166
rect 15660 5102 15712 5108
rect 16028 5160 16080 5166
rect 16028 5102 16080 5108
rect 16120 5160 16172 5166
rect 16120 5102 16172 5108
rect 15580 4690 15608 5102
rect 16040 4690 16068 5102
rect 16224 5030 16252 7919
rect 16304 7890 16356 7896
rect 16316 7478 16344 7890
rect 16304 7472 16356 7478
rect 16304 7414 16356 7420
rect 16212 5024 16264 5030
rect 16212 4966 16264 4972
rect 16316 4758 16344 7414
rect 16500 6866 16528 9454
rect 16578 8528 16634 8537
rect 16578 8463 16634 8472
rect 16488 6860 16540 6866
rect 16488 6802 16540 6808
rect 16396 6656 16448 6662
rect 16396 6598 16448 6604
rect 16408 5273 16436 6598
rect 16500 6390 16528 6802
rect 16488 6384 16540 6390
rect 16488 6326 16540 6332
rect 16592 6254 16620 8463
rect 16684 7993 16712 23582
rect 16946 23520 17002 23582
rect 17880 23582 18290 23610
rect 16956 21244 17252 21264
rect 17012 21242 17036 21244
rect 17092 21242 17116 21244
rect 17172 21242 17196 21244
rect 17034 21190 17036 21242
rect 17098 21190 17110 21242
rect 17172 21190 17174 21242
rect 17012 21188 17036 21190
rect 17092 21188 17116 21190
rect 17172 21188 17196 21190
rect 16956 21168 17252 21188
rect 17880 20602 17908 23582
rect 18234 23520 18290 23582
rect 19260 23582 19578 23610
rect 19260 21146 19288 23582
rect 19522 23520 19578 23582
rect 20456 23582 20774 23610
rect 20074 22808 20130 22817
rect 20074 22743 20130 22752
rect 19982 21992 20038 22001
rect 19982 21927 20038 21936
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19248 21140 19300 21146
rect 19248 21082 19300 21088
rect 18052 21004 18104 21010
rect 18052 20946 18104 20952
rect 17868 20596 17920 20602
rect 17868 20538 17920 20544
rect 18064 20330 18092 20946
rect 18972 20392 19024 20398
rect 18972 20334 19024 20340
rect 18052 20324 18104 20330
rect 18052 20266 18104 20272
rect 16956 20156 17252 20176
rect 17012 20154 17036 20156
rect 17092 20154 17116 20156
rect 17172 20154 17196 20156
rect 17034 20102 17036 20154
rect 17098 20102 17110 20154
rect 17172 20102 17174 20154
rect 17012 20100 17036 20102
rect 17092 20100 17116 20102
rect 17172 20100 17196 20102
rect 16956 20080 17252 20100
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 17500 19984 17552 19990
rect 17500 19926 17552 19932
rect 17224 19848 17276 19854
rect 17224 19790 17276 19796
rect 17236 19378 17264 19790
rect 17224 19372 17276 19378
rect 17224 19314 17276 19320
rect 17512 19242 17540 19926
rect 17684 19304 17736 19310
rect 17684 19246 17736 19252
rect 17500 19236 17552 19242
rect 17500 19178 17552 19184
rect 16956 19068 17252 19088
rect 17012 19066 17036 19068
rect 17092 19066 17116 19068
rect 17172 19066 17196 19068
rect 17034 19014 17036 19066
rect 17098 19014 17110 19066
rect 17172 19014 17174 19066
rect 17012 19012 17036 19014
rect 17092 19012 17116 19014
rect 17172 19012 17196 19014
rect 16956 18992 17252 19012
rect 17512 18902 17540 19178
rect 17132 18896 17184 18902
rect 17132 18838 17184 18844
rect 17500 18896 17552 18902
rect 17500 18838 17552 18844
rect 17144 18426 17172 18838
rect 17512 18698 17540 18838
rect 17696 18698 17724 19246
rect 18892 19174 18920 19994
rect 18236 19168 18288 19174
rect 18236 19110 18288 19116
rect 18788 19168 18840 19174
rect 18788 19110 18840 19116
rect 18880 19168 18932 19174
rect 18880 19110 18932 19116
rect 17500 18692 17552 18698
rect 17500 18634 17552 18640
rect 17684 18692 17736 18698
rect 17684 18634 17736 18640
rect 17132 18420 17184 18426
rect 17132 18362 17184 18368
rect 17512 18358 17540 18634
rect 17500 18352 17552 18358
rect 17500 18294 17552 18300
rect 16856 18080 16908 18086
rect 16856 18022 16908 18028
rect 16868 17814 16896 18022
rect 16956 17980 17252 18000
rect 17012 17978 17036 17980
rect 17092 17978 17116 17980
rect 17172 17978 17196 17980
rect 17034 17926 17036 17978
rect 17098 17926 17110 17978
rect 17172 17926 17174 17978
rect 17012 17924 17036 17926
rect 17092 17924 17116 17926
rect 17172 17924 17196 17926
rect 16956 17904 17252 17924
rect 16856 17808 16908 17814
rect 16856 17750 16908 17756
rect 16948 17808 17000 17814
rect 16948 17750 17000 17756
rect 16868 17338 16896 17750
rect 16856 17332 16908 17338
rect 16856 17274 16908 17280
rect 16960 17202 16988 17750
rect 17696 17610 17724 18634
rect 17684 17604 17736 17610
rect 17684 17546 17736 17552
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 17868 16992 17920 16998
rect 17868 16934 17920 16940
rect 16956 16892 17252 16912
rect 17012 16890 17036 16892
rect 17092 16890 17116 16892
rect 17172 16890 17196 16892
rect 17034 16838 17036 16890
rect 17098 16838 17110 16890
rect 17172 16838 17174 16890
rect 17012 16836 17036 16838
rect 17092 16836 17116 16838
rect 17172 16836 17196 16838
rect 16956 16816 17252 16836
rect 17880 16794 17908 16934
rect 17408 16788 17460 16794
rect 17408 16730 17460 16736
rect 17868 16788 17920 16794
rect 17868 16730 17920 16736
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 16960 16114 16988 16526
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 17420 15978 17448 16730
rect 17776 16584 17828 16590
rect 17776 16526 17828 16532
rect 17408 15972 17460 15978
rect 17408 15914 17460 15920
rect 16956 15804 17252 15824
rect 17012 15802 17036 15804
rect 17092 15802 17116 15804
rect 17172 15802 17196 15804
rect 17034 15750 17036 15802
rect 17098 15750 17110 15802
rect 17172 15750 17174 15802
rect 17012 15748 17036 15750
rect 17092 15748 17116 15750
rect 17172 15748 17196 15750
rect 16956 15728 17252 15748
rect 17788 15706 17816 16526
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 16856 15632 16908 15638
rect 16776 15592 16856 15620
rect 16776 14822 16804 15592
rect 16856 15574 16908 15580
rect 18248 15552 18276 19110
rect 18800 18766 18828 19110
rect 18892 18902 18920 19110
rect 18880 18896 18932 18902
rect 18880 18838 18932 18844
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18800 18426 18828 18702
rect 18788 18420 18840 18426
rect 18788 18362 18840 18368
rect 18892 18290 18920 18838
rect 18880 18284 18932 18290
rect 18880 18226 18932 18232
rect 18788 18080 18840 18086
rect 18788 18022 18840 18028
rect 18800 17814 18828 18022
rect 18788 17808 18840 17814
rect 18788 17750 18840 17756
rect 18328 17672 18380 17678
rect 18328 17614 18380 17620
rect 18340 17202 18368 17614
rect 18696 17604 18748 17610
rect 18696 17546 18748 17552
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 18708 16572 18736 17546
rect 18800 17338 18828 17750
rect 18788 17332 18840 17338
rect 18788 17274 18840 17280
rect 18984 17105 19012 20334
rect 19352 19990 19380 21286
rect 19996 21010 20024 21927
rect 20088 21690 20116 22743
rect 20076 21684 20128 21690
rect 20076 21626 20128 21632
rect 20088 21486 20116 21626
rect 20076 21480 20128 21486
rect 20076 21422 20128 21428
rect 19984 21004 20036 21010
rect 19984 20946 20036 20952
rect 19524 20800 19576 20806
rect 19524 20742 19576 20748
rect 19340 19984 19392 19990
rect 19340 19926 19392 19932
rect 19064 19848 19116 19854
rect 19064 19790 19116 19796
rect 19076 18766 19104 19790
rect 19352 19514 19380 19926
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 19064 18760 19116 18766
rect 19064 18702 19116 18708
rect 19076 17678 19104 18702
rect 19536 18290 19564 20742
rect 19996 20534 20024 20946
rect 20456 20602 20484 23582
rect 20718 23520 20774 23582
rect 21744 23582 22062 23610
rect 20956 21788 21252 21808
rect 21012 21786 21036 21788
rect 21092 21786 21116 21788
rect 21172 21786 21196 21788
rect 21034 21734 21036 21786
rect 21098 21734 21110 21786
rect 21172 21734 21174 21786
rect 21012 21732 21036 21734
rect 21092 21732 21116 21734
rect 21172 21732 21196 21734
rect 20956 21712 21252 21732
rect 21454 20904 21510 20913
rect 21454 20839 21510 20848
rect 20956 20700 21252 20720
rect 21012 20698 21036 20700
rect 21092 20698 21116 20700
rect 21172 20698 21196 20700
rect 21034 20646 21036 20698
rect 21098 20646 21110 20698
rect 21172 20646 21174 20698
rect 21012 20644 21036 20646
rect 21092 20644 21116 20646
rect 21172 20644 21196 20646
rect 20956 20624 21252 20644
rect 20444 20596 20496 20602
rect 20444 20538 20496 20544
rect 19984 20528 20036 20534
rect 19984 20470 20036 20476
rect 19892 20392 19944 20398
rect 19892 20334 19944 20340
rect 19708 18624 19760 18630
rect 19708 18566 19760 18572
rect 19524 18284 19576 18290
rect 19524 18226 19576 18232
rect 19156 18080 19208 18086
rect 19156 18022 19208 18028
rect 19064 17672 19116 17678
rect 19064 17614 19116 17620
rect 18970 17096 19026 17105
rect 18970 17031 19026 17040
rect 19064 17060 19116 17066
rect 19064 17002 19116 17008
rect 18880 16720 18932 16726
rect 18880 16662 18932 16668
rect 18788 16584 18840 16590
rect 18708 16544 18788 16572
rect 18788 16526 18840 16532
rect 18800 15706 18828 16526
rect 18892 16250 18920 16662
rect 19076 16590 19104 17002
rect 19064 16584 19116 16590
rect 19064 16526 19116 16532
rect 18880 16244 18932 16250
rect 18880 16186 18932 16192
rect 19076 16182 19104 16526
rect 19064 16176 19116 16182
rect 19064 16118 19116 16124
rect 18788 15700 18840 15706
rect 18788 15642 18840 15648
rect 19076 15570 19104 16118
rect 18328 15564 18380 15570
rect 18248 15524 18328 15552
rect 18328 15506 18380 15512
rect 19064 15564 19116 15570
rect 19064 15506 19116 15512
rect 17316 15496 17368 15502
rect 17316 15438 17368 15444
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16764 14816 16816 14822
rect 16764 14758 16816 14764
rect 16776 14006 16804 14758
rect 16868 14618 16896 15302
rect 16956 14716 17252 14736
rect 17012 14714 17036 14716
rect 17092 14714 17116 14716
rect 17172 14714 17196 14716
rect 17034 14662 17036 14714
rect 17098 14662 17110 14714
rect 17172 14662 17174 14714
rect 17012 14660 17036 14662
rect 17092 14660 17116 14662
rect 17172 14660 17196 14662
rect 16956 14640 17252 14660
rect 16856 14612 16908 14618
rect 16856 14554 16908 14560
rect 16764 14000 16816 14006
rect 16764 13942 16816 13948
rect 17328 13938 17356 15438
rect 18340 15162 18368 15506
rect 19076 15162 19104 15506
rect 18328 15156 18380 15162
rect 18328 15098 18380 15104
rect 19064 15156 19116 15162
rect 19064 15098 19116 15104
rect 18236 14816 18288 14822
rect 18236 14758 18288 14764
rect 19064 14816 19116 14822
rect 19064 14758 19116 14764
rect 18248 14618 18276 14758
rect 18236 14612 18288 14618
rect 18236 14554 18288 14560
rect 19076 14550 19104 14758
rect 19064 14544 19116 14550
rect 19064 14486 19116 14492
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 18880 14408 18932 14414
rect 18880 14350 18932 14356
rect 17604 14074 17632 14350
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 17328 13814 17356 13874
rect 18788 13864 18840 13870
rect 17328 13786 17448 13814
rect 18788 13806 18840 13812
rect 16956 13628 17252 13648
rect 17012 13626 17036 13628
rect 17092 13626 17116 13628
rect 17172 13626 17196 13628
rect 17034 13574 17036 13626
rect 17098 13574 17110 13626
rect 17172 13574 17174 13626
rect 17012 13572 17036 13574
rect 17092 13572 17116 13574
rect 17172 13572 17196 13574
rect 16956 13552 17252 13572
rect 17420 13530 17448 13786
rect 17408 13524 17460 13530
rect 17408 13466 17460 13472
rect 18144 13524 18196 13530
rect 18144 13466 18196 13472
rect 16856 13456 16908 13462
rect 16856 13398 16908 13404
rect 16868 12986 16896 13398
rect 16948 13320 17000 13326
rect 16948 13262 17000 13268
rect 17408 13320 17460 13326
rect 17408 13262 17460 13268
rect 16960 12986 16988 13262
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 16764 12640 16816 12646
rect 16764 12582 16816 12588
rect 16776 8378 16804 12582
rect 16868 12442 16896 12922
rect 17420 12782 17448 13262
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17408 12776 17460 12782
rect 17408 12718 17460 12724
rect 16956 12540 17252 12560
rect 17012 12538 17036 12540
rect 17092 12538 17116 12540
rect 17172 12538 17196 12540
rect 17034 12486 17036 12538
rect 17098 12486 17110 12538
rect 17172 12486 17174 12538
rect 17012 12484 17036 12486
rect 17092 12484 17116 12486
rect 17172 12484 17196 12486
rect 16956 12464 17252 12484
rect 17420 12442 17448 12718
rect 16856 12436 16908 12442
rect 16856 12378 16908 12384
rect 17408 12436 17460 12442
rect 17408 12378 17460 12384
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 16960 11762 16988 12174
rect 17420 11762 17448 12378
rect 16948 11756 17000 11762
rect 16948 11698 17000 11704
rect 17408 11756 17460 11762
rect 17408 11698 17460 11704
rect 16956 11452 17252 11472
rect 17012 11450 17036 11452
rect 17092 11450 17116 11452
rect 17172 11450 17196 11452
rect 17034 11398 17036 11450
rect 17098 11398 17110 11450
rect 17172 11398 17174 11450
rect 17012 11396 17036 11398
rect 17092 11396 17116 11398
rect 17172 11396 17196 11398
rect 16956 11376 17252 11396
rect 16854 11112 16910 11121
rect 16854 11047 16910 11056
rect 16868 10130 16896 11047
rect 16956 10364 17252 10384
rect 17012 10362 17036 10364
rect 17092 10362 17116 10364
rect 17172 10362 17196 10364
rect 17034 10310 17036 10362
rect 17098 10310 17110 10362
rect 17172 10310 17174 10362
rect 17012 10308 17036 10310
rect 17092 10308 17116 10310
rect 17172 10308 17196 10310
rect 16956 10288 17252 10308
rect 17500 10192 17552 10198
rect 17500 10134 17552 10140
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16868 9722 16896 10066
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 17512 9382 17540 10134
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 16956 9276 17252 9296
rect 17012 9274 17036 9276
rect 17092 9274 17116 9276
rect 17172 9274 17196 9276
rect 17034 9222 17036 9274
rect 17098 9222 17110 9274
rect 17172 9222 17174 9274
rect 17012 9220 17036 9222
rect 17092 9220 17116 9222
rect 17172 9220 17196 9222
rect 16956 9200 17252 9220
rect 17512 9178 17540 9318
rect 17500 9172 17552 9178
rect 17500 9114 17552 9120
rect 17512 8566 17540 9114
rect 17500 8560 17552 8566
rect 17500 8502 17552 8508
rect 16776 8350 16896 8378
rect 16670 7984 16726 7993
rect 16670 7919 16726 7928
rect 16764 6792 16816 6798
rect 16764 6734 16816 6740
rect 16776 6458 16804 6734
rect 16764 6452 16816 6458
rect 16764 6394 16816 6400
rect 16764 6316 16816 6322
rect 16764 6258 16816 6264
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 16488 5772 16540 5778
rect 16488 5714 16540 5720
rect 16394 5264 16450 5273
rect 16394 5199 16450 5208
rect 16396 5160 16448 5166
rect 16396 5102 16448 5108
rect 16304 4752 16356 4758
rect 16304 4694 16356 4700
rect 15568 4684 15620 4690
rect 15568 4626 15620 4632
rect 16028 4684 16080 4690
rect 16080 4644 16160 4672
rect 16028 4626 16080 4632
rect 15474 4176 15530 4185
rect 15474 4111 15530 4120
rect 16132 3942 16160 4644
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 16224 3738 16252 4558
rect 16316 4214 16344 4694
rect 16408 4690 16436 5102
rect 16500 5098 16528 5714
rect 16672 5568 16724 5574
rect 16592 5528 16672 5556
rect 16488 5092 16540 5098
rect 16488 5034 16540 5040
rect 16396 4684 16448 4690
rect 16396 4626 16448 4632
rect 16408 4282 16436 4626
rect 16396 4276 16448 4282
rect 16396 4218 16448 4224
rect 16304 4208 16356 4214
rect 16304 4150 16356 4156
rect 16592 4146 16620 5528
rect 16672 5510 16724 5516
rect 16776 5234 16804 6258
rect 16764 5228 16816 5234
rect 16764 5170 16816 5176
rect 16764 5024 16816 5030
rect 16764 4966 16816 4972
rect 16776 4154 16804 4966
rect 16580 4140 16632 4146
rect 16580 4082 16632 4088
rect 16684 4126 16804 4154
rect 16396 4004 16448 4010
rect 16396 3946 16448 3952
rect 16580 4004 16632 4010
rect 16580 3946 16632 3952
rect 16408 3738 16436 3946
rect 16212 3732 16264 3738
rect 16212 3674 16264 3680
rect 16396 3732 16448 3738
rect 16396 3674 16448 3680
rect 15476 3664 15528 3670
rect 15476 3606 15528 3612
rect 15488 3194 15516 3606
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 15568 3460 15620 3466
rect 15568 3402 15620 3408
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 15580 3058 15608 3402
rect 15672 3194 15700 3470
rect 15936 3460 15988 3466
rect 15936 3402 15988 3408
rect 16028 3460 16080 3466
rect 16028 3402 16080 3408
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 15568 3052 15620 3058
rect 15568 2994 15620 3000
rect 15672 2854 15700 3130
rect 15752 2916 15804 2922
rect 15752 2858 15804 2864
rect 15660 2848 15712 2854
rect 15660 2790 15712 2796
rect 15672 2582 15700 2790
rect 15764 2650 15792 2858
rect 15752 2644 15804 2650
rect 15752 2586 15804 2592
rect 15660 2576 15712 2582
rect 15660 2518 15712 2524
rect 15948 2378 15976 3402
rect 15936 2372 15988 2378
rect 15936 2314 15988 2320
rect 15198 82 15254 480
rect 15120 54 15254 82
rect 16040 82 16068 3402
rect 16592 3058 16620 3946
rect 16580 3052 16632 3058
rect 16580 2994 16632 3000
rect 16684 2514 16712 4126
rect 16868 3602 16896 8350
rect 16956 8188 17252 8208
rect 17012 8186 17036 8188
rect 17092 8186 17116 8188
rect 17172 8186 17196 8188
rect 17034 8134 17036 8186
rect 17098 8134 17110 8186
rect 17172 8134 17174 8186
rect 17012 8132 17036 8134
rect 17092 8132 17116 8134
rect 17172 8132 17196 8134
rect 16956 8112 17252 8132
rect 16956 7100 17252 7120
rect 17012 7098 17036 7100
rect 17092 7098 17116 7100
rect 17172 7098 17196 7100
rect 17034 7046 17036 7098
rect 17098 7046 17110 7098
rect 17172 7046 17174 7098
rect 17012 7044 17036 7046
rect 17092 7044 17116 7046
rect 17172 7044 17196 7046
rect 16956 7024 17252 7044
rect 17316 6112 17368 6118
rect 17316 6054 17368 6060
rect 16956 6012 17252 6032
rect 17012 6010 17036 6012
rect 17092 6010 17116 6012
rect 17172 6010 17196 6012
rect 17034 5958 17036 6010
rect 17098 5958 17110 6010
rect 17172 5958 17174 6010
rect 17012 5956 17036 5958
rect 17092 5956 17116 5958
rect 17172 5956 17196 5958
rect 16956 5936 17252 5956
rect 17328 5914 17356 6054
rect 17316 5908 17368 5914
rect 17316 5850 17368 5856
rect 17316 5568 17368 5574
rect 17316 5510 17368 5516
rect 16956 4924 17252 4944
rect 17012 4922 17036 4924
rect 17092 4922 17116 4924
rect 17172 4922 17196 4924
rect 17034 4870 17036 4922
rect 17098 4870 17110 4922
rect 17172 4870 17174 4922
rect 17012 4868 17036 4870
rect 17092 4868 17116 4870
rect 17172 4868 17196 4870
rect 16956 4848 17252 4868
rect 17328 4758 17356 5510
rect 17316 4752 17368 4758
rect 17316 4694 17368 4700
rect 17604 4154 17632 13126
rect 18156 12850 18184 13466
rect 18800 13326 18828 13806
rect 18892 13705 18920 14350
rect 19076 14074 19104 14486
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 18878 13696 18934 13705
rect 18878 13631 18934 13640
rect 18420 13320 18472 13326
rect 18420 13262 18472 13268
rect 18788 13320 18840 13326
rect 18788 13262 18840 13268
rect 18236 12912 18288 12918
rect 18236 12854 18288 12860
rect 18144 12844 18196 12850
rect 18144 12786 18196 12792
rect 18248 12714 18276 12854
rect 18432 12850 18460 13262
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 18236 12708 18288 12714
rect 18236 12650 18288 12656
rect 18800 12442 18828 13262
rect 18892 12986 18920 13631
rect 19064 13456 19116 13462
rect 19064 13398 19116 13404
rect 18880 12980 18932 12986
rect 18880 12922 18932 12928
rect 19076 12782 19104 13398
rect 19064 12776 19116 12782
rect 19064 12718 19116 12724
rect 18788 12436 18840 12442
rect 18788 12378 18840 12384
rect 18144 12368 18196 12374
rect 18144 12310 18196 12316
rect 18156 11558 18184 12310
rect 19076 12306 19104 12718
rect 19064 12300 19116 12306
rect 19064 12242 19116 12248
rect 18144 11552 18196 11558
rect 18144 11494 18196 11500
rect 18972 11552 19024 11558
rect 18972 11494 19024 11500
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17880 10538 17908 11154
rect 18156 11014 18184 11494
rect 18144 11008 18196 11014
rect 18144 10950 18196 10956
rect 18512 11008 18564 11014
rect 18512 10950 18564 10956
rect 17868 10532 17920 10538
rect 17868 10474 17920 10480
rect 17880 10441 17908 10474
rect 18156 10470 18184 10950
rect 18144 10464 18196 10470
rect 17866 10432 17922 10441
rect 18144 10406 18196 10412
rect 17866 10367 17922 10376
rect 18156 10266 18184 10406
rect 18144 10260 18196 10266
rect 18144 10202 18196 10208
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 17972 9654 18000 9998
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 17960 9648 18012 9654
rect 17960 9590 18012 9596
rect 17868 9376 17920 9382
rect 17868 9318 17920 9324
rect 17880 8362 17908 9318
rect 17684 8356 17736 8362
rect 17684 8298 17736 8304
rect 17868 8356 17920 8362
rect 17868 8298 17920 8304
rect 17696 6934 17724 8298
rect 17972 7546 18000 9590
rect 18156 9586 18184 9862
rect 18144 9580 18196 9586
rect 18144 9522 18196 9528
rect 18524 9110 18552 10950
rect 18984 10674 19012 11494
rect 18972 10668 19024 10674
rect 18972 10610 19024 10616
rect 19168 10130 19196 18022
rect 19536 17882 19564 18226
rect 19720 18154 19748 18566
rect 19708 18148 19760 18154
rect 19708 18090 19760 18096
rect 19524 17876 19576 17882
rect 19524 17818 19576 17824
rect 19720 17814 19748 18090
rect 19248 17808 19300 17814
rect 19248 17750 19300 17756
rect 19708 17808 19760 17814
rect 19708 17750 19760 17756
rect 19260 17270 19288 17750
rect 19800 17740 19852 17746
rect 19800 17682 19852 17688
rect 19248 17264 19300 17270
rect 19248 17206 19300 17212
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19352 16561 19380 16934
rect 19338 16552 19394 16561
rect 19338 16487 19394 16496
rect 19812 16153 19840 17682
rect 19904 17377 19932 20334
rect 20812 19916 20864 19922
rect 20812 19858 20864 19864
rect 19984 19848 20036 19854
rect 19984 19790 20036 19796
rect 19996 19446 20024 19790
rect 20720 19712 20772 19718
rect 20720 19654 20772 19660
rect 19984 19440 20036 19446
rect 19984 19382 20036 19388
rect 19996 18290 20024 19382
rect 19984 18284 20036 18290
rect 19984 18226 20036 18232
rect 19890 17368 19946 17377
rect 19890 17303 19946 17312
rect 19798 16144 19854 16153
rect 19798 16079 19854 16088
rect 19800 15360 19852 15366
rect 19800 15302 19852 15308
rect 19616 14544 19668 14550
rect 19616 14486 19668 14492
rect 19248 14340 19300 14346
rect 19248 14282 19300 14288
rect 19260 13433 19288 14282
rect 19432 13796 19484 13802
rect 19432 13738 19484 13744
rect 19340 13728 19392 13734
rect 19340 13670 19392 13676
rect 19246 13424 19302 13433
rect 19246 13359 19302 13368
rect 19352 12306 19380 13670
rect 19444 13190 19472 13738
rect 19628 13734 19656 14486
rect 19616 13728 19668 13734
rect 19616 13670 19668 13676
rect 19628 13530 19656 13670
rect 19616 13524 19668 13530
rect 19616 13466 19668 13472
rect 19432 13184 19484 13190
rect 19432 13126 19484 13132
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 19708 12300 19760 12306
rect 19708 12242 19760 12248
rect 19720 11898 19748 12242
rect 19708 11892 19760 11898
rect 19708 11834 19760 11840
rect 19156 10124 19208 10130
rect 19156 10066 19208 10072
rect 19524 10124 19576 10130
rect 19524 10066 19576 10072
rect 18788 10056 18840 10062
rect 18788 9998 18840 10004
rect 18800 9450 18828 9998
rect 18788 9444 18840 9450
rect 18788 9386 18840 9392
rect 18512 9104 18564 9110
rect 18512 9046 18564 9052
rect 18236 8832 18288 8838
rect 18236 8774 18288 8780
rect 18248 8498 18276 8774
rect 18236 8492 18288 8498
rect 18236 8434 18288 8440
rect 18524 8090 18552 9046
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 18236 8016 18288 8022
rect 18236 7958 18288 7964
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 18248 7478 18276 7958
rect 18800 7886 18828 9386
rect 19536 9382 19564 10066
rect 19524 9376 19576 9382
rect 19524 9318 19576 9324
rect 19248 9104 19300 9110
rect 19248 9046 19300 9052
rect 18972 8968 19024 8974
rect 18972 8910 19024 8916
rect 18984 8362 19012 8910
rect 19260 8430 19288 9046
rect 19248 8424 19300 8430
rect 19248 8366 19300 8372
rect 18972 8356 19024 8362
rect 18972 8298 19024 8304
rect 18788 7880 18840 7886
rect 18788 7822 18840 7828
rect 18696 7812 18748 7818
rect 18696 7754 18748 7760
rect 18236 7472 18288 7478
rect 18236 7414 18288 7420
rect 18248 7002 18276 7414
rect 18708 7274 18736 7754
rect 18420 7268 18472 7274
rect 18420 7210 18472 7216
rect 18696 7268 18748 7274
rect 18696 7210 18748 7216
rect 18236 6996 18288 7002
rect 18236 6938 18288 6944
rect 17684 6928 17736 6934
rect 17684 6870 17736 6876
rect 17696 6458 17724 6870
rect 18432 6458 18460 7210
rect 17684 6452 17736 6458
rect 17684 6394 17736 6400
rect 18420 6452 18472 6458
rect 18420 6394 18472 6400
rect 17696 5846 17724 6394
rect 17684 5840 17736 5846
rect 17684 5782 17736 5788
rect 17696 5370 17724 5782
rect 17684 5364 17736 5370
rect 17684 5306 17736 5312
rect 17696 5030 17724 5306
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 17684 5024 17736 5030
rect 17684 4966 17736 4972
rect 17696 4826 17724 4966
rect 18064 4826 18092 5102
rect 18236 5092 18288 5098
rect 18236 5034 18288 5040
rect 17684 4820 17736 4826
rect 17684 4762 17736 4768
rect 18052 4820 18104 4826
rect 18052 4762 18104 4768
rect 17512 4126 17632 4154
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 16956 3836 17252 3856
rect 17012 3834 17036 3836
rect 17092 3834 17116 3836
rect 17172 3834 17196 3836
rect 17034 3782 17036 3834
rect 17098 3782 17110 3834
rect 17172 3782 17174 3834
rect 17012 3780 17036 3782
rect 17092 3780 17116 3782
rect 17172 3780 17196 3782
rect 16956 3760 17252 3780
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 16868 3194 16896 3538
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 17328 2961 17356 3878
rect 17512 3738 17540 4126
rect 17500 3732 17552 3738
rect 17500 3674 17552 3680
rect 17696 3126 17724 4762
rect 18248 3602 18276 5034
rect 18708 4690 18736 7210
rect 18800 7002 18828 7822
rect 18984 7410 19012 8298
rect 19156 8288 19208 8294
rect 19156 8230 19208 8236
rect 19064 7472 19116 7478
rect 19064 7414 19116 7420
rect 18972 7404 19024 7410
rect 18972 7346 19024 7352
rect 18788 6996 18840 7002
rect 18788 6938 18840 6944
rect 19076 6458 19104 7414
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 19076 6254 19104 6394
rect 19064 6248 19116 6254
rect 19168 6225 19196 8230
rect 19536 6730 19564 9318
rect 19616 8492 19668 8498
rect 19616 8434 19668 8440
rect 19628 8090 19656 8434
rect 19616 8084 19668 8090
rect 19616 8026 19668 8032
rect 19708 6860 19760 6866
rect 19708 6802 19760 6808
rect 19524 6724 19576 6730
rect 19524 6666 19576 6672
rect 19720 6390 19748 6802
rect 19708 6384 19760 6390
rect 19708 6326 19760 6332
rect 19064 6190 19116 6196
rect 19154 6216 19210 6225
rect 19154 6151 19210 6160
rect 19432 5840 19484 5846
rect 19432 5782 19484 5788
rect 19444 5642 19472 5782
rect 18880 5636 18932 5642
rect 18880 5578 18932 5584
rect 19432 5636 19484 5642
rect 19432 5578 19484 5584
rect 18328 4684 18380 4690
rect 18328 4626 18380 4632
rect 18696 4684 18748 4690
rect 18696 4626 18748 4632
rect 18340 4282 18368 4626
rect 18892 4282 18920 5578
rect 19340 5024 19392 5030
rect 19340 4966 19392 4972
rect 19708 5024 19760 5030
rect 19708 4966 19760 4972
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 18328 4276 18380 4282
rect 18328 4218 18380 4224
rect 18880 4276 18932 4282
rect 18880 4218 18932 4224
rect 18892 4078 18920 4218
rect 18880 4072 18932 4078
rect 18880 4014 18932 4020
rect 19260 3738 19288 4558
rect 19352 3738 19380 4966
rect 19720 4758 19748 4966
rect 19708 4752 19760 4758
rect 19708 4694 19760 4700
rect 19720 4010 19748 4694
rect 19708 4004 19760 4010
rect 19708 3946 19760 3952
rect 19248 3732 19300 3738
rect 19248 3674 19300 3680
rect 19340 3732 19392 3738
rect 19340 3674 19392 3680
rect 18236 3596 18288 3602
rect 18236 3538 18288 3544
rect 18604 3596 18656 3602
rect 18604 3538 18656 3544
rect 17684 3120 17736 3126
rect 17684 3062 17736 3068
rect 17314 2952 17370 2961
rect 17314 2887 17370 2896
rect 18616 2854 18644 3538
rect 19260 3194 19288 3674
rect 19248 3188 19300 3194
rect 19248 3130 19300 3136
rect 19248 2984 19300 2990
rect 19248 2926 19300 2932
rect 18052 2848 18104 2854
rect 18052 2790 18104 2796
rect 18604 2848 18656 2854
rect 18604 2790 18656 2796
rect 16956 2748 17252 2768
rect 17012 2746 17036 2748
rect 17092 2746 17116 2748
rect 17172 2746 17196 2748
rect 17034 2694 17036 2746
rect 17098 2694 17110 2746
rect 17172 2694 17174 2746
rect 17012 2692 17036 2694
rect 17092 2692 17116 2694
rect 17172 2692 17196 2694
rect 16956 2672 17252 2692
rect 16672 2508 16724 2514
rect 16672 2450 16724 2456
rect 18064 2446 18092 2790
rect 18616 2446 18644 2790
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 18604 2440 18656 2446
rect 18604 2382 18656 2388
rect 16948 2304 17000 2310
rect 16948 2246 17000 2252
rect 18236 2304 18288 2310
rect 18236 2246 18288 2252
rect 18972 2304 19024 2310
rect 18972 2246 19024 2252
rect 16118 82 16174 480
rect 16040 54 16174 82
rect 16960 82 16988 2246
rect 17038 82 17094 480
rect 16960 54 17094 82
rect 13358 0 13414 54
rect 14278 0 14334 54
rect 15198 0 15254 54
rect 16118 0 16174 54
rect 17038 0 17094 54
rect 17958 82 18014 480
rect 18248 82 18276 2246
rect 18984 1873 19012 2246
rect 18970 1864 19026 1873
rect 18970 1799 19026 1808
rect 17958 54 18276 82
rect 18878 82 18934 480
rect 19260 82 19288 2926
rect 19812 2650 19840 15302
rect 19904 13814 19932 17303
rect 19996 16114 20024 18226
rect 20732 16776 20760 19654
rect 20824 19514 20852 19858
rect 20956 19612 21252 19632
rect 21012 19610 21036 19612
rect 21092 19610 21116 19612
rect 21172 19610 21196 19612
rect 21034 19558 21036 19610
rect 21098 19558 21110 19610
rect 21172 19558 21174 19610
rect 21012 19556 21036 19558
rect 21092 19556 21116 19558
rect 21172 19556 21196 19558
rect 20956 19536 21252 19556
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 21270 18864 21326 18873
rect 21270 18799 21326 18808
rect 20956 18524 21252 18544
rect 21012 18522 21036 18524
rect 21092 18522 21116 18524
rect 21172 18522 21196 18524
rect 21034 18470 21036 18522
rect 21098 18470 21110 18522
rect 21172 18470 21174 18522
rect 21012 18468 21036 18470
rect 21092 18468 21116 18470
rect 21172 18468 21196 18470
rect 20956 18448 21252 18468
rect 21284 18426 21312 18799
rect 21272 18420 21324 18426
rect 21272 18362 21324 18368
rect 20956 17436 21252 17456
rect 21012 17434 21036 17436
rect 21092 17434 21116 17436
rect 21172 17434 21196 17436
rect 21034 17382 21036 17434
rect 21098 17382 21110 17434
rect 21172 17382 21174 17434
rect 21012 17380 21036 17382
rect 21092 17380 21116 17382
rect 21172 17380 21196 17382
rect 20956 17360 21252 17380
rect 21468 17338 21496 20839
rect 21744 20602 21772 23582
rect 22006 23520 22062 23582
rect 23032 23582 23350 23610
rect 21732 20596 21784 20602
rect 21732 20538 21784 20544
rect 23032 19922 23060 23582
rect 23294 23520 23350 23582
rect 23020 19916 23072 19922
rect 23020 19858 23072 19864
rect 21638 19816 21694 19825
rect 21638 19751 21694 19760
rect 21652 19514 21680 19751
rect 21640 19508 21692 19514
rect 21640 19450 21692 19456
rect 21652 19310 21680 19450
rect 21640 19304 21692 19310
rect 21640 19246 21692 19252
rect 21730 18048 21786 18057
rect 21730 17983 21786 17992
rect 21744 17882 21772 17983
rect 21732 17876 21784 17882
rect 21732 17818 21784 17824
rect 21732 17740 21784 17746
rect 21732 17682 21784 17688
rect 21744 17338 21772 17682
rect 21456 17332 21508 17338
rect 21456 17274 21508 17280
rect 21732 17332 21784 17338
rect 21732 17274 21784 17280
rect 20902 17232 20958 17241
rect 20902 17167 20958 17176
rect 20732 16748 20852 16776
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 19996 15706 20024 16050
rect 19984 15700 20036 15706
rect 19984 15642 20036 15648
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 19904 13786 20024 13814
rect 19890 12472 19946 12481
rect 19890 12407 19946 12416
rect 19904 12170 19932 12407
rect 19892 12164 19944 12170
rect 19892 12106 19944 12112
rect 19996 12102 20024 13786
rect 20076 13796 20128 13802
rect 20076 13738 20128 13744
rect 20536 13796 20588 13802
rect 20536 13738 20588 13744
rect 20088 13705 20116 13738
rect 20444 13728 20496 13734
rect 20074 13696 20130 13705
rect 20444 13670 20496 13676
rect 20074 13631 20130 13640
rect 20088 13530 20116 13631
rect 20076 13524 20128 13530
rect 20076 13466 20128 13472
rect 20258 13424 20314 13433
rect 20258 13359 20314 13368
rect 20076 13184 20128 13190
rect 20076 13126 20128 13132
rect 19984 12096 20036 12102
rect 19984 12038 20036 12044
rect 19984 11824 20036 11830
rect 19984 11766 20036 11772
rect 19996 11218 20024 11766
rect 19984 11212 20036 11218
rect 19984 11154 20036 11160
rect 19996 10742 20024 11154
rect 19984 10736 20036 10742
rect 19984 10678 20036 10684
rect 19996 10538 20024 10678
rect 19984 10532 20036 10538
rect 19984 10474 20036 10480
rect 19892 5636 19944 5642
rect 19892 5578 19944 5584
rect 19904 4758 19932 5578
rect 19892 4752 19944 4758
rect 19892 4694 19944 4700
rect 20088 4154 20116 13126
rect 20272 12918 20300 13359
rect 20260 12912 20312 12918
rect 20260 12854 20312 12860
rect 20456 12850 20484 13670
rect 20444 12844 20496 12850
rect 20444 12786 20496 12792
rect 20456 12442 20484 12786
rect 20444 12436 20496 12442
rect 20444 12378 20496 12384
rect 20168 11620 20220 11626
rect 20168 11562 20220 11568
rect 20180 11286 20208 11562
rect 20168 11280 20220 11286
rect 20168 11222 20220 11228
rect 20180 10810 20208 11222
rect 20168 10804 20220 10810
rect 20168 10746 20220 10752
rect 20260 10668 20312 10674
rect 20260 10610 20312 10616
rect 20272 10198 20300 10610
rect 20260 10192 20312 10198
rect 20260 10134 20312 10140
rect 20548 6934 20576 13738
rect 20732 12374 20760 14758
rect 20824 13802 20852 16748
rect 20916 16658 20944 17167
rect 21468 17134 21496 17274
rect 21456 17128 21508 17134
rect 21456 17070 21508 17076
rect 21730 16960 21786 16969
rect 21730 16895 21786 16904
rect 21744 16794 21772 16895
rect 21732 16788 21784 16794
rect 21732 16730 21784 16736
rect 20904 16652 20956 16658
rect 20904 16594 20956 16600
rect 21272 16652 21324 16658
rect 21272 16594 21324 16600
rect 20956 16348 21252 16368
rect 21012 16346 21036 16348
rect 21092 16346 21116 16348
rect 21172 16346 21196 16348
rect 21034 16294 21036 16346
rect 21098 16294 21110 16346
rect 21172 16294 21174 16346
rect 21012 16292 21036 16294
rect 21092 16292 21116 16294
rect 21172 16292 21196 16294
rect 20956 16272 21252 16292
rect 21284 16250 21312 16594
rect 21272 16244 21324 16250
rect 21272 16186 21324 16192
rect 21454 15872 21510 15881
rect 21454 15807 21510 15816
rect 20956 15260 21252 15280
rect 21012 15258 21036 15260
rect 21092 15258 21116 15260
rect 21172 15258 21196 15260
rect 21034 15206 21036 15258
rect 21098 15206 21110 15258
rect 21172 15206 21174 15258
rect 21012 15204 21036 15206
rect 21092 15204 21116 15206
rect 21172 15204 21196 15206
rect 20956 15184 21252 15204
rect 21468 15162 21496 15807
rect 21456 15156 21508 15162
rect 21456 15098 21508 15104
rect 21468 14958 21496 15098
rect 21456 14952 21508 14958
rect 21456 14894 21508 14900
rect 23570 14376 23626 14385
rect 23492 14334 23570 14362
rect 20956 14172 21252 14192
rect 21012 14170 21036 14172
rect 21092 14170 21116 14172
rect 21172 14170 21196 14172
rect 21034 14118 21036 14170
rect 21098 14118 21110 14170
rect 21172 14118 21174 14170
rect 21012 14116 21036 14118
rect 21092 14116 21116 14118
rect 21172 14116 21196 14118
rect 20956 14096 21252 14116
rect 20812 13796 20864 13802
rect 20812 13738 20864 13744
rect 21732 13796 21784 13802
rect 21732 13738 21784 13744
rect 20812 13456 20864 13462
rect 20812 13398 20864 13404
rect 20824 12986 20852 13398
rect 21456 13252 21508 13258
rect 21456 13194 21508 13200
rect 20956 13084 21252 13104
rect 21012 13082 21036 13084
rect 21092 13082 21116 13084
rect 21172 13082 21196 13084
rect 21034 13030 21036 13082
rect 21098 13030 21110 13082
rect 21172 13030 21174 13082
rect 21012 13028 21036 13030
rect 21092 13028 21116 13030
rect 21172 13028 21196 13030
rect 20956 13008 21252 13028
rect 21362 13016 21418 13025
rect 20812 12980 20864 12986
rect 21468 12986 21496 13194
rect 21362 12951 21418 12960
rect 21456 12980 21508 12986
rect 20812 12922 20864 12928
rect 21376 12918 21404 12951
rect 21456 12922 21508 12928
rect 21364 12912 21416 12918
rect 21364 12854 21416 12860
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 20720 12368 20772 12374
rect 20720 12310 20772 12316
rect 20732 11898 20760 12310
rect 20720 11892 20772 11898
rect 20720 11834 20772 11840
rect 20824 11665 20852 12718
rect 21272 12368 21324 12374
rect 21272 12310 21324 12316
rect 20956 11996 21252 12016
rect 21012 11994 21036 11996
rect 21092 11994 21116 11996
rect 21172 11994 21196 11996
rect 21034 11942 21036 11994
rect 21098 11942 21110 11994
rect 21172 11942 21174 11994
rect 21012 11940 21036 11942
rect 21092 11940 21116 11942
rect 21172 11940 21196 11942
rect 20956 11920 21252 11940
rect 21284 11830 21312 12310
rect 21640 12232 21692 12238
rect 21640 12174 21692 12180
rect 21272 11824 21324 11830
rect 21272 11766 21324 11772
rect 20810 11656 20866 11665
rect 20720 11620 20772 11626
rect 20810 11591 20866 11600
rect 20720 11562 20772 11568
rect 20628 11552 20680 11558
rect 20628 11494 20680 11500
rect 20640 11014 20668 11494
rect 20628 11008 20680 11014
rect 20628 10950 20680 10956
rect 20640 10266 20668 10950
rect 20732 10674 20760 11562
rect 21548 11552 21600 11558
rect 21548 11494 21600 11500
rect 21272 11280 21324 11286
rect 21272 11222 21324 11228
rect 20956 10908 21252 10928
rect 21012 10906 21036 10908
rect 21092 10906 21116 10908
rect 21172 10906 21196 10908
rect 21034 10854 21036 10906
rect 21098 10854 21110 10906
rect 21172 10854 21174 10906
rect 21012 10852 21036 10854
rect 21092 10852 21116 10854
rect 21172 10852 21196 10854
rect 20956 10832 21252 10852
rect 21284 10810 21312 11222
rect 21456 11144 21508 11150
rect 21560 11132 21588 11494
rect 21652 11286 21680 12174
rect 21640 11280 21692 11286
rect 21640 11222 21692 11228
rect 21508 11104 21588 11132
rect 21456 11086 21508 11092
rect 21362 10840 21418 10849
rect 21272 10804 21324 10810
rect 21560 10810 21588 11104
rect 21362 10775 21418 10784
rect 21548 10804 21600 10810
rect 21272 10746 21324 10752
rect 20720 10668 20772 10674
rect 20720 10610 20772 10616
rect 20628 10260 20680 10266
rect 20628 10202 20680 10208
rect 20732 9586 20760 10610
rect 20902 10568 20958 10577
rect 20902 10503 20958 10512
rect 20916 10130 20944 10503
rect 21376 10266 21404 10775
rect 21548 10746 21600 10752
rect 21364 10260 21416 10266
rect 21364 10202 21416 10208
rect 20904 10124 20956 10130
rect 20904 10066 20956 10072
rect 21548 10124 21600 10130
rect 21548 10066 21600 10072
rect 20956 9820 21252 9840
rect 21012 9818 21036 9820
rect 21092 9818 21116 9820
rect 21172 9818 21196 9820
rect 21034 9766 21036 9818
rect 21098 9766 21110 9818
rect 21172 9766 21174 9818
rect 21012 9764 21036 9766
rect 21092 9764 21116 9766
rect 21172 9764 21196 9766
rect 20956 9744 21252 9764
rect 21560 9722 21588 10066
rect 21548 9716 21600 9722
rect 21548 9658 21600 9664
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20732 9178 20760 9522
rect 20812 9444 20864 9450
rect 20812 9386 20864 9392
rect 21272 9444 21324 9450
rect 21272 9386 21324 9392
rect 20720 9172 20772 9178
rect 20720 9114 20772 9120
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 20732 8634 20760 8842
rect 20720 8628 20772 8634
rect 20720 8570 20772 8576
rect 20732 7954 20760 8570
rect 20824 8022 20852 9386
rect 21088 9104 21140 9110
rect 21088 9046 21140 9052
rect 21100 8906 21128 9046
rect 21284 8974 21312 9386
rect 21652 9178 21680 11222
rect 21640 9172 21692 9178
rect 21640 9114 21692 9120
rect 21272 8968 21324 8974
rect 21272 8910 21324 8916
rect 21088 8900 21140 8906
rect 21088 8842 21140 8848
rect 20956 8732 21252 8752
rect 21012 8730 21036 8732
rect 21092 8730 21116 8732
rect 21172 8730 21196 8732
rect 21034 8678 21036 8730
rect 21098 8678 21110 8730
rect 21172 8678 21174 8730
rect 21012 8676 21036 8678
rect 21092 8676 21116 8678
rect 21172 8676 21196 8678
rect 20956 8656 21252 8676
rect 21284 8430 21312 8910
rect 21652 8634 21680 9114
rect 21640 8628 21692 8634
rect 21640 8570 21692 8576
rect 21272 8424 21324 8430
rect 21272 8366 21324 8372
rect 20812 8016 20864 8022
rect 20812 7958 20864 7964
rect 20720 7948 20772 7954
rect 20720 7890 20772 7896
rect 20732 7478 20760 7890
rect 21270 7848 21326 7857
rect 21270 7783 21326 7792
rect 20956 7644 21252 7664
rect 21012 7642 21036 7644
rect 21092 7642 21116 7644
rect 21172 7642 21196 7644
rect 21034 7590 21036 7642
rect 21098 7590 21110 7642
rect 21172 7590 21174 7642
rect 21012 7588 21036 7590
rect 21092 7588 21116 7590
rect 21172 7588 21196 7590
rect 20956 7568 21252 7588
rect 21284 7546 21312 7783
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 20720 7472 20772 7478
rect 20720 7414 20772 7420
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20536 6928 20588 6934
rect 20536 6870 20588 6876
rect 20548 6458 20576 6870
rect 20536 6452 20588 6458
rect 20536 6394 20588 6400
rect 20536 6316 20588 6322
rect 20536 6258 20588 6264
rect 20548 5914 20576 6258
rect 20824 6186 20852 7142
rect 21456 6928 21508 6934
rect 21456 6870 21508 6876
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 20956 6556 21252 6576
rect 21012 6554 21036 6556
rect 21092 6554 21116 6556
rect 21172 6554 21196 6556
rect 21034 6502 21036 6554
rect 21098 6502 21110 6554
rect 21172 6502 21174 6554
rect 21012 6500 21036 6502
rect 21092 6500 21116 6502
rect 21172 6500 21196 6502
rect 20956 6480 21252 6500
rect 21284 6322 21312 6734
rect 21362 6488 21418 6497
rect 21362 6423 21418 6432
rect 21376 6390 21404 6423
rect 21468 6390 21496 6870
rect 21364 6384 21416 6390
rect 21364 6326 21416 6332
rect 21456 6384 21508 6390
rect 21456 6326 21508 6332
rect 21272 6316 21324 6322
rect 21272 6258 21324 6264
rect 20628 6180 20680 6186
rect 20628 6122 20680 6128
rect 20812 6180 20864 6186
rect 20812 6122 20864 6128
rect 21272 6180 21324 6186
rect 21272 6122 21324 6128
rect 20536 5908 20588 5914
rect 20536 5850 20588 5856
rect 20548 5234 20576 5850
rect 20536 5228 20588 5234
rect 20536 5170 20588 5176
rect 20640 4758 20668 6122
rect 20812 5840 20864 5846
rect 20812 5782 20864 5788
rect 20824 5302 20852 5782
rect 21284 5710 21312 6122
rect 21468 5914 21496 6326
rect 21456 5908 21508 5914
rect 21456 5850 21508 5856
rect 21468 5760 21496 5850
rect 21376 5732 21496 5760
rect 21272 5704 21324 5710
rect 21272 5646 21324 5652
rect 20956 5468 21252 5488
rect 21012 5466 21036 5468
rect 21092 5466 21116 5468
rect 21172 5466 21196 5468
rect 21034 5414 21036 5466
rect 21098 5414 21110 5466
rect 21172 5414 21174 5466
rect 21012 5412 21036 5414
rect 21092 5412 21116 5414
rect 21172 5412 21196 5414
rect 20956 5392 21252 5412
rect 21376 5370 21404 5732
rect 21456 5636 21508 5642
rect 21456 5578 21508 5584
rect 21468 5370 21496 5578
rect 21364 5364 21416 5370
rect 21364 5306 21416 5312
rect 21456 5364 21508 5370
rect 21456 5306 21508 5312
rect 20812 5296 20864 5302
rect 20812 5238 20864 5244
rect 20996 5296 21048 5302
rect 20996 5238 21048 5244
rect 20628 4752 20680 4758
rect 20628 4694 20680 4700
rect 21008 4690 21036 5238
rect 21270 5128 21326 5137
rect 21270 5063 21326 5072
rect 21284 5030 21312 5063
rect 21272 5024 21324 5030
rect 21744 5001 21772 13738
rect 23492 6118 23520 14334
rect 23570 14311 23626 14320
rect 23572 12096 23624 12102
rect 23572 12038 23624 12044
rect 23584 9489 23612 12038
rect 23570 9480 23626 9489
rect 23570 9415 23626 9424
rect 23480 6112 23532 6118
rect 23480 6054 23532 6060
rect 21914 5400 21970 5409
rect 21914 5335 21970 5344
rect 21928 5302 21956 5335
rect 21916 5296 21968 5302
rect 21916 5238 21968 5244
rect 21272 4966 21324 4972
rect 21730 4992 21786 5001
rect 21730 4927 21786 4936
rect 20996 4684 21048 4690
rect 20824 4644 20996 4672
rect 20824 4282 20852 4644
rect 20996 4626 21048 4632
rect 20956 4380 21252 4400
rect 21012 4378 21036 4380
rect 21092 4378 21116 4380
rect 21172 4378 21196 4380
rect 21034 4326 21036 4378
rect 21098 4326 21110 4378
rect 21172 4326 21174 4378
rect 21012 4324 21036 4326
rect 21092 4324 21116 4326
rect 21172 4324 21196 4326
rect 20956 4304 21252 4324
rect 20812 4276 20864 4282
rect 20812 4218 20864 4224
rect 20088 4126 20300 4154
rect 20272 3738 20300 4126
rect 23570 4040 23626 4049
rect 23570 3975 23626 3984
rect 20260 3732 20312 3738
rect 20260 3674 20312 3680
rect 20810 3632 20866 3641
rect 20810 3567 20866 3576
rect 21456 3596 21508 3602
rect 20824 3194 20852 3567
rect 21456 3538 21508 3544
rect 21468 3505 21496 3538
rect 21454 3496 21510 3505
rect 21454 3431 21510 3440
rect 20956 3292 21252 3312
rect 21012 3290 21036 3292
rect 21092 3290 21116 3292
rect 21172 3290 21196 3292
rect 21034 3238 21036 3290
rect 21098 3238 21110 3290
rect 21172 3238 21174 3290
rect 21012 3236 21036 3238
rect 21092 3236 21116 3238
rect 21172 3236 21196 3238
rect 20956 3216 21252 3236
rect 21468 3194 21496 3431
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 21456 3188 21508 3194
rect 21456 3130 21508 3136
rect 22284 2848 22336 2854
rect 22284 2790 22336 2796
rect 19800 2644 19852 2650
rect 19800 2586 19852 2592
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 18878 54 19288 82
rect 19628 82 19656 2382
rect 20444 2372 20496 2378
rect 20444 2314 20496 2320
rect 19798 82 19854 480
rect 19628 54 19854 82
rect 20456 82 20484 2314
rect 20956 2204 21252 2224
rect 21012 2202 21036 2204
rect 21092 2202 21116 2204
rect 21172 2202 21196 2204
rect 21034 2150 21036 2202
rect 21098 2150 21110 2202
rect 21172 2150 21174 2202
rect 21012 2148 21036 2150
rect 21092 2148 21116 2150
rect 21172 2148 21196 2150
rect 20956 2128 21252 2148
rect 21362 1728 21418 1737
rect 21362 1663 21418 1672
rect 20718 82 20774 480
rect 20456 54 20774 82
rect 21376 82 21404 1663
rect 21638 82 21694 480
rect 21376 54 21694 82
rect 22296 82 22324 2790
rect 23204 2304 23256 2310
rect 23204 2246 23256 2252
rect 22558 82 22614 480
rect 22296 54 22614 82
rect 23216 82 23244 2246
rect 23584 1465 23612 3975
rect 23570 1456 23626 1465
rect 23570 1391 23626 1400
rect 23478 82 23534 480
rect 23216 54 23534 82
rect 17958 0 18014 54
rect 18878 0 18934 54
rect 19798 0 19854 54
rect 20718 0 20774 54
rect 21638 0 21694 54
rect 22558 0 22614 54
rect 23478 0 23534 54
<< via2 >>
rect 1306 22480 1362 22536
rect 1582 20712 1638 20768
rect 110 17856 166 17912
rect 110 16224 166 16280
rect 4956 21786 5012 21788
rect 5036 21786 5092 21788
rect 5116 21786 5172 21788
rect 5196 21786 5252 21788
rect 4956 21734 4982 21786
rect 4982 21734 5012 21786
rect 5036 21734 5046 21786
rect 5046 21734 5092 21786
rect 5116 21734 5162 21786
rect 5162 21734 5172 21786
rect 5196 21734 5226 21786
rect 5226 21734 5252 21786
rect 4956 21732 5012 21734
rect 5036 21732 5092 21734
rect 5116 21732 5172 21734
rect 5196 21732 5252 21734
rect 4956 20698 5012 20700
rect 5036 20698 5092 20700
rect 5116 20698 5172 20700
rect 5196 20698 5252 20700
rect 4956 20646 4982 20698
rect 4982 20646 5012 20698
rect 5036 20646 5046 20698
rect 5046 20646 5092 20698
rect 5116 20646 5162 20698
rect 5162 20646 5172 20698
rect 5196 20646 5226 20698
rect 5226 20646 5252 20698
rect 4956 20644 5012 20646
rect 5036 20644 5092 20646
rect 5116 20644 5172 20646
rect 5196 20644 5252 20646
rect 2226 19216 2282 19272
rect 1582 12280 1638 12336
rect 1674 9560 1730 9616
rect 1582 9016 1638 9072
rect 110 8880 166 8936
rect 4956 19610 5012 19612
rect 5036 19610 5092 19612
rect 5116 19610 5172 19612
rect 5196 19610 5252 19612
rect 4956 19558 4982 19610
rect 4982 19558 5012 19610
rect 5036 19558 5046 19610
rect 5046 19558 5092 19610
rect 5116 19558 5162 19610
rect 5162 19558 5172 19610
rect 5196 19558 5226 19610
rect 5226 19558 5252 19610
rect 4956 19556 5012 19558
rect 5036 19556 5092 19558
rect 5116 19556 5172 19558
rect 5196 19556 5252 19558
rect 4956 18522 5012 18524
rect 5036 18522 5092 18524
rect 5116 18522 5172 18524
rect 5196 18522 5252 18524
rect 4956 18470 4982 18522
rect 4982 18470 5012 18522
rect 5036 18470 5046 18522
rect 5046 18470 5092 18522
rect 5116 18470 5162 18522
rect 5162 18470 5172 18522
rect 5196 18470 5226 18522
rect 5226 18470 5252 18522
rect 4956 18468 5012 18470
rect 5036 18468 5092 18470
rect 5116 18468 5172 18470
rect 5196 18468 5252 18470
rect 5814 18264 5870 18320
rect 8956 21242 9012 21244
rect 9036 21242 9092 21244
rect 9116 21242 9172 21244
rect 9196 21242 9252 21244
rect 8956 21190 8982 21242
rect 8982 21190 9012 21242
rect 9036 21190 9046 21242
rect 9046 21190 9092 21242
rect 9116 21190 9162 21242
rect 9162 21190 9172 21242
rect 9196 21190 9226 21242
rect 9226 21190 9252 21242
rect 8956 21188 9012 21190
rect 9036 21188 9092 21190
rect 9116 21188 9172 21190
rect 9196 21188 9252 21190
rect 7102 18128 7158 18184
rect 4956 17434 5012 17436
rect 5036 17434 5092 17436
rect 5116 17434 5172 17436
rect 5196 17434 5252 17436
rect 4956 17382 4982 17434
rect 4982 17382 5012 17434
rect 5036 17382 5046 17434
rect 5046 17382 5092 17434
rect 5116 17382 5162 17434
rect 5162 17382 5172 17434
rect 5196 17382 5226 17434
rect 5226 17382 5252 17434
rect 4956 17380 5012 17382
rect 5036 17380 5092 17382
rect 5116 17380 5172 17382
rect 5196 17380 5252 17382
rect 3514 14728 3570 14784
rect 1582 7112 1638 7168
rect 1582 5344 1638 5400
rect 110 2488 166 2544
rect 1122 1400 1178 1456
rect 3514 9560 3570 9616
rect 2870 6160 2926 6216
rect 2042 1672 2098 1728
rect 4158 9560 4214 9616
rect 4956 16346 5012 16348
rect 5036 16346 5092 16348
rect 5116 16346 5172 16348
rect 5196 16346 5252 16348
rect 4956 16294 4982 16346
rect 4982 16294 5012 16346
rect 5036 16294 5046 16346
rect 5046 16294 5092 16346
rect 5116 16294 5162 16346
rect 5162 16294 5172 16346
rect 5196 16294 5226 16346
rect 5226 16294 5252 16346
rect 4956 16292 5012 16294
rect 5036 16292 5092 16294
rect 5116 16292 5172 16294
rect 5196 16292 5252 16294
rect 4956 15258 5012 15260
rect 5036 15258 5092 15260
rect 5116 15258 5172 15260
rect 5196 15258 5252 15260
rect 4956 15206 4982 15258
rect 4982 15206 5012 15258
rect 5036 15206 5046 15258
rect 5046 15206 5092 15258
rect 5116 15206 5162 15258
rect 5162 15206 5172 15258
rect 5196 15206 5226 15258
rect 5226 15206 5252 15258
rect 4956 15204 5012 15206
rect 5036 15204 5092 15206
rect 5116 15204 5172 15206
rect 5196 15204 5252 15206
rect 4956 14170 5012 14172
rect 5036 14170 5092 14172
rect 5116 14170 5172 14172
rect 5196 14170 5252 14172
rect 4956 14118 4982 14170
rect 4982 14118 5012 14170
rect 5036 14118 5046 14170
rect 5046 14118 5092 14170
rect 5116 14118 5162 14170
rect 5162 14118 5172 14170
rect 5196 14118 5226 14170
rect 5226 14118 5252 14170
rect 4956 14116 5012 14118
rect 5036 14116 5092 14118
rect 5116 14116 5172 14118
rect 5196 14116 5252 14118
rect 5354 13776 5410 13832
rect 5538 13776 5594 13832
rect 4066 8472 4122 8528
rect 4956 13082 5012 13084
rect 5036 13082 5092 13084
rect 5116 13082 5172 13084
rect 5196 13082 5252 13084
rect 4956 13030 4982 13082
rect 4982 13030 5012 13082
rect 5036 13030 5046 13082
rect 5046 13030 5092 13082
rect 5116 13030 5162 13082
rect 5162 13030 5172 13082
rect 5196 13030 5226 13082
rect 5226 13030 5252 13082
rect 4956 13028 5012 13030
rect 5036 13028 5092 13030
rect 5116 13028 5172 13030
rect 5196 13028 5252 13030
rect 4956 11994 5012 11996
rect 5036 11994 5092 11996
rect 5116 11994 5172 11996
rect 5196 11994 5252 11996
rect 4956 11942 4982 11994
rect 4982 11942 5012 11994
rect 5036 11942 5046 11994
rect 5046 11942 5092 11994
rect 5116 11942 5162 11994
rect 5162 11942 5172 11994
rect 5196 11942 5226 11994
rect 5226 11942 5252 11994
rect 4956 11940 5012 11942
rect 5036 11940 5092 11942
rect 5116 11940 5172 11942
rect 5196 11940 5252 11942
rect 4956 10906 5012 10908
rect 5036 10906 5092 10908
rect 5116 10906 5172 10908
rect 5196 10906 5252 10908
rect 4956 10854 4982 10906
rect 4982 10854 5012 10906
rect 5036 10854 5046 10906
rect 5046 10854 5092 10906
rect 5116 10854 5162 10906
rect 5162 10854 5172 10906
rect 5196 10854 5226 10906
rect 5226 10854 5252 10906
rect 4956 10852 5012 10854
rect 5036 10852 5092 10854
rect 5116 10852 5172 10854
rect 5196 10852 5252 10854
rect 4956 9818 5012 9820
rect 5036 9818 5092 9820
rect 5116 9818 5172 9820
rect 5196 9818 5252 9820
rect 4956 9766 4982 9818
rect 4982 9766 5012 9818
rect 5036 9766 5046 9818
rect 5046 9766 5092 9818
rect 5116 9766 5162 9818
rect 5162 9766 5172 9818
rect 5196 9766 5226 9818
rect 5226 9766 5252 9818
rect 4956 9764 5012 9766
rect 5036 9764 5092 9766
rect 5116 9764 5172 9766
rect 5196 9764 5252 9766
rect 5722 9696 5778 9752
rect 4956 8730 5012 8732
rect 5036 8730 5092 8732
rect 5116 8730 5172 8732
rect 5196 8730 5252 8732
rect 4956 8678 4982 8730
rect 4982 8678 5012 8730
rect 5036 8678 5046 8730
rect 5046 8678 5092 8730
rect 5116 8678 5162 8730
rect 5162 8678 5172 8730
rect 5196 8678 5226 8730
rect 5226 8678 5252 8730
rect 4956 8676 5012 8678
rect 5036 8676 5092 8678
rect 5116 8676 5172 8678
rect 5196 8676 5252 8678
rect 4956 7642 5012 7644
rect 5036 7642 5092 7644
rect 5116 7642 5172 7644
rect 5196 7642 5252 7644
rect 4956 7590 4982 7642
rect 4982 7590 5012 7642
rect 5036 7590 5046 7642
rect 5046 7590 5092 7642
rect 5116 7590 5162 7642
rect 5162 7590 5172 7642
rect 5196 7590 5226 7642
rect 5226 7590 5252 7642
rect 4956 7588 5012 7590
rect 5036 7588 5092 7590
rect 5116 7588 5172 7590
rect 5196 7588 5252 7590
rect 4956 6554 5012 6556
rect 5036 6554 5092 6556
rect 5116 6554 5172 6556
rect 5196 6554 5252 6556
rect 4956 6502 4982 6554
rect 4982 6502 5012 6554
rect 5036 6502 5046 6554
rect 5046 6502 5092 6554
rect 5116 6502 5162 6554
rect 5162 6502 5172 6554
rect 5196 6502 5226 6554
rect 5226 6502 5252 6554
rect 4956 6500 5012 6502
rect 5036 6500 5092 6502
rect 5116 6500 5172 6502
rect 5196 6500 5252 6502
rect 4956 5466 5012 5468
rect 5036 5466 5092 5468
rect 5116 5466 5172 5468
rect 5196 5466 5252 5468
rect 4956 5414 4982 5466
rect 4982 5414 5012 5466
rect 5036 5414 5046 5466
rect 5046 5414 5092 5466
rect 5116 5414 5162 5466
rect 5162 5414 5172 5466
rect 5196 5414 5226 5466
rect 5226 5414 5252 5466
rect 4956 5412 5012 5414
rect 5036 5412 5092 5414
rect 5116 5412 5172 5414
rect 5196 5412 5252 5414
rect 4956 4378 5012 4380
rect 5036 4378 5092 4380
rect 5116 4378 5172 4380
rect 5196 4378 5252 4380
rect 4956 4326 4982 4378
rect 4982 4326 5012 4378
rect 5036 4326 5046 4378
rect 5046 4326 5092 4378
rect 5116 4326 5162 4378
rect 5162 4326 5172 4378
rect 5196 4326 5226 4378
rect 5226 4326 5252 4378
rect 4956 4324 5012 4326
rect 5036 4324 5092 4326
rect 5116 4324 5172 4326
rect 5196 4324 5252 4326
rect 6642 17040 6698 17096
rect 7194 16496 7250 16552
rect 8114 15408 8170 15464
rect 5630 5344 5686 5400
rect 4956 3290 5012 3292
rect 5036 3290 5092 3292
rect 5116 3290 5172 3292
rect 5196 3290 5252 3292
rect 4956 3238 4982 3290
rect 4982 3238 5012 3290
rect 5036 3238 5046 3290
rect 5046 3238 5092 3290
rect 5116 3238 5162 3290
rect 5162 3238 5172 3290
rect 5196 3238 5226 3290
rect 5226 3238 5252 3290
rect 4956 3236 5012 3238
rect 5036 3236 5092 3238
rect 5116 3236 5172 3238
rect 5196 3236 5252 3238
rect 4956 2202 5012 2204
rect 5036 2202 5092 2204
rect 5116 2202 5172 2204
rect 5196 2202 5252 2204
rect 4956 2150 4982 2202
rect 4982 2150 5012 2202
rect 5036 2150 5046 2202
rect 5046 2150 5092 2202
rect 5116 2150 5162 2202
rect 5162 2150 5172 2202
rect 5196 2150 5226 2202
rect 5226 2150 5252 2202
rect 4956 2148 5012 2150
rect 5036 2148 5092 2150
rect 5116 2148 5172 2150
rect 5196 2148 5252 2150
rect 6642 5208 6698 5264
rect 8206 14728 8262 14784
rect 7838 13776 7894 13832
rect 7562 7928 7618 7984
rect 7102 1808 7158 1864
rect 7562 40 7618 96
rect 7930 9016 7986 9072
rect 8666 17040 8722 17096
rect 8956 20154 9012 20156
rect 9036 20154 9092 20156
rect 9116 20154 9172 20156
rect 9196 20154 9252 20156
rect 8956 20102 8982 20154
rect 8982 20102 9012 20154
rect 9036 20102 9046 20154
rect 9046 20102 9092 20154
rect 9116 20102 9162 20154
rect 9162 20102 9172 20154
rect 9196 20102 9226 20154
rect 9226 20102 9252 20154
rect 8956 20100 9012 20102
rect 9036 20100 9092 20102
rect 9116 20100 9172 20102
rect 9196 20100 9252 20102
rect 8956 19066 9012 19068
rect 9036 19066 9092 19068
rect 9116 19066 9172 19068
rect 9196 19066 9252 19068
rect 8956 19014 8982 19066
rect 8982 19014 9012 19066
rect 9036 19014 9046 19066
rect 9046 19014 9092 19066
rect 9116 19014 9162 19066
rect 9162 19014 9172 19066
rect 9196 19014 9226 19066
rect 9226 19014 9252 19066
rect 8956 19012 9012 19014
rect 9036 19012 9092 19014
rect 9116 19012 9172 19014
rect 9196 19012 9252 19014
rect 8956 17978 9012 17980
rect 9036 17978 9092 17980
rect 9116 17978 9172 17980
rect 9196 17978 9252 17980
rect 8956 17926 8982 17978
rect 8982 17926 9012 17978
rect 9036 17926 9046 17978
rect 9046 17926 9092 17978
rect 9116 17926 9162 17978
rect 9162 17926 9172 17978
rect 9196 17926 9226 17978
rect 9226 17926 9252 17978
rect 8956 17924 9012 17926
rect 9036 17924 9092 17926
rect 9116 17924 9172 17926
rect 9196 17924 9252 17926
rect 8956 16890 9012 16892
rect 9036 16890 9092 16892
rect 9116 16890 9172 16892
rect 9196 16890 9252 16892
rect 8956 16838 8982 16890
rect 8982 16838 9012 16890
rect 9036 16838 9046 16890
rect 9046 16838 9092 16890
rect 9116 16838 9162 16890
rect 9162 16838 9172 16890
rect 9196 16838 9226 16890
rect 9226 16838 9252 16890
rect 8956 16836 9012 16838
rect 9036 16836 9092 16838
rect 9116 16836 9172 16838
rect 9196 16836 9252 16838
rect 8850 15952 8906 16008
rect 8956 15802 9012 15804
rect 9036 15802 9092 15804
rect 9116 15802 9172 15804
rect 9196 15802 9252 15804
rect 8956 15750 8982 15802
rect 8982 15750 9012 15802
rect 9036 15750 9046 15802
rect 9046 15750 9092 15802
rect 9116 15750 9162 15802
rect 9162 15750 9172 15802
rect 9196 15750 9226 15802
rect 9226 15750 9252 15802
rect 8956 15748 9012 15750
rect 9036 15748 9092 15750
rect 9116 15748 9172 15750
rect 9196 15748 9252 15750
rect 8956 14714 9012 14716
rect 9036 14714 9092 14716
rect 9116 14714 9172 14716
rect 9196 14714 9252 14716
rect 8956 14662 8982 14714
rect 8982 14662 9012 14714
rect 9036 14662 9046 14714
rect 9046 14662 9092 14714
rect 9116 14662 9162 14714
rect 9162 14662 9172 14714
rect 9196 14662 9226 14714
rect 9226 14662 9252 14714
rect 8956 14660 9012 14662
rect 9036 14660 9092 14662
rect 9116 14660 9172 14662
rect 9196 14660 9252 14662
rect 8956 13626 9012 13628
rect 9036 13626 9092 13628
rect 9116 13626 9172 13628
rect 9196 13626 9252 13628
rect 8956 13574 8982 13626
rect 8982 13574 9012 13626
rect 9036 13574 9046 13626
rect 9046 13574 9092 13626
rect 9116 13574 9162 13626
rect 9162 13574 9172 13626
rect 9196 13574 9226 13626
rect 9226 13574 9252 13626
rect 8956 13572 9012 13574
rect 9036 13572 9092 13574
rect 9116 13572 9172 13574
rect 9196 13572 9252 13574
rect 7746 5364 7802 5400
rect 7746 5344 7748 5364
rect 7748 5344 7800 5364
rect 7800 5344 7802 5364
rect 8956 12538 9012 12540
rect 9036 12538 9092 12540
rect 9116 12538 9172 12540
rect 9196 12538 9252 12540
rect 8956 12486 8982 12538
rect 8982 12486 9012 12538
rect 9036 12486 9046 12538
rect 9046 12486 9092 12538
rect 9116 12486 9162 12538
rect 9162 12486 9172 12538
rect 9196 12486 9226 12538
rect 9226 12486 9252 12538
rect 8956 12484 9012 12486
rect 9036 12484 9092 12486
rect 9116 12484 9172 12486
rect 9196 12484 9252 12486
rect 12956 21786 13012 21788
rect 13036 21786 13092 21788
rect 13116 21786 13172 21788
rect 13196 21786 13252 21788
rect 12956 21734 12982 21786
rect 12982 21734 13012 21786
rect 13036 21734 13046 21786
rect 13046 21734 13092 21786
rect 13116 21734 13162 21786
rect 13162 21734 13172 21786
rect 13196 21734 13226 21786
rect 13226 21734 13252 21786
rect 12956 21732 13012 21734
rect 13036 21732 13092 21734
rect 13116 21732 13172 21734
rect 13196 21732 13252 21734
rect 12956 20698 13012 20700
rect 13036 20698 13092 20700
rect 13116 20698 13172 20700
rect 13196 20698 13252 20700
rect 12956 20646 12982 20698
rect 12982 20646 13012 20698
rect 13036 20646 13046 20698
rect 13046 20646 13092 20698
rect 13116 20646 13162 20698
rect 13162 20646 13172 20698
rect 13196 20646 13226 20698
rect 13226 20646 13252 20698
rect 12956 20644 13012 20646
rect 13036 20644 13092 20646
rect 13116 20644 13172 20646
rect 13196 20644 13252 20646
rect 10874 17176 10930 17232
rect 9402 13640 9458 13696
rect 8956 11450 9012 11452
rect 9036 11450 9092 11452
rect 9116 11450 9172 11452
rect 9196 11450 9252 11452
rect 8956 11398 8982 11450
rect 8982 11398 9012 11450
rect 9036 11398 9046 11450
rect 9046 11398 9092 11450
rect 9116 11398 9162 11450
rect 9162 11398 9172 11450
rect 9196 11398 9226 11450
rect 9226 11398 9252 11450
rect 8956 11396 9012 11398
rect 9036 11396 9092 11398
rect 9116 11396 9172 11398
rect 9196 11396 9252 11398
rect 11334 13912 11390 13968
rect 8956 10362 9012 10364
rect 9036 10362 9092 10364
rect 9116 10362 9172 10364
rect 9196 10362 9252 10364
rect 8956 10310 8982 10362
rect 8982 10310 9012 10362
rect 9036 10310 9046 10362
rect 9046 10310 9092 10362
rect 9116 10310 9162 10362
rect 9162 10310 9172 10362
rect 9196 10310 9226 10362
rect 9226 10310 9252 10362
rect 8956 10308 9012 10310
rect 9036 10308 9092 10310
rect 9116 10308 9172 10310
rect 9196 10308 9252 10310
rect 10322 10512 10378 10568
rect 9310 9696 9366 9752
rect 9310 9560 9366 9616
rect 8956 9274 9012 9276
rect 9036 9274 9092 9276
rect 9116 9274 9172 9276
rect 9196 9274 9252 9276
rect 8956 9222 8982 9274
rect 8982 9222 9012 9274
rect 9036 9222 9046 9274
rect 9046 9222 9092 9274
rect 9116 9222 9162 9274
rect 9162 9222 9172 9274
rect 9196 9222 9226 9274
rect 9226 9222 9252 9274
rect 8956 9220 9012 9222
rect 9036 9220 9092 9222
rect 9116 9220 9172 9222
rect 9196 9220 9252 9222
rect 8850 9016 8906 9072
rect 8956 8186 9012 8188
rect 9036 8186 9092 8188
rect 9116 8186 9172 8188
rect 9196 8186 9252 8188
rect 8956 8134 8982 8186
rect 8982 8134 9012 8186
rect 9036 8134 9046 8186
rect 9046 8134 9092 8186
rect 9116 8134 9162 8186
rect 9162 8134 9172 8186
rect 9196 8134 9226 8186
rect 9226 8134 9252 8186
rect 8956 8132 9012 8134
rect 9036 8132 9092 8134
rect 9116 8132 9172 8134
rect 9196 8132 9252 8134
rect 8850 7384 8906 7440
rect 8956 7098 9012 7100
rect 9036 7098 9092 7100
rect 9116 7098 9172 7100
rect 9196 7098 9252 7100
rect 8956 7046 8982 7098
rect 8982 7046 9012 7098
rect 9036 7046 9046 7098
rect 9046 7046 9092 7098
rect 9116 7046 9162 7098
rect 9162 7046 9172 7098
rect 9196 7046 9226 7098
rect 9226 7046 9252 7098
rect 8956 7044 9012 7046
rect 9036 7044 9092 7046
rect 9116 7044 9172 7046
rect 9196 7044 9252 7046
rect 7930 3984 7986 4040
rect 8956 6010 9012 6012
rect 9036 6010 9092 6012
rect 9116 6010 9172 6012
rect 9196 6010 9252 6012
rect 8956 5958 8982 6010
rect 8982 5958 9012 6010
rect 9036 5958 9046 6010
rect 9046 5958 9092 6010
rect 9116 5958 9162 6010
rect 9162 5958 9172 6010
rect 9196 5958 9226 6010
rect 9226 5958 9252 6010
rect 8956 5956 9012 5958
rect 9036 5956 9092 5958
rect 9116 5956 9172 5958
rect 9196 5956 9252 5958
rect 8956 4922 9012 4924
rect 9036 4922 9092 4924
rect 9116 4922 9172 4924
rect 9196 4922 9252 4924
rect 8956 4870 8982 4922
rect 8982 4870 9012 4922
rect 9036 4870 9046 4922
rect 9046 4870 9092 4922
rect 9116 4870 9162 4922
rect 9162 4870 9172 4922
rect 9196 4870 9226 4922
rect 9226 4870 9252 4922
rect 8956 4868 9012 4870
rect 9036 4868 9092 4870
rect 9116 4868 9172 4870
rect 9196 4868 9252 4870
rect 8956 3834 9012 3836
rect 9036 3834 9092 3836
rect 9116 3834 9172 3836
rect 9196 3834 9252 3836
rect 8956 3782 8982 3834
rect 8982 3782 9012 3834
rect 9036 3782 9046 3834
rect 9046 3782 9092 3834
rect 9116 3782 9162 3834
rect 9162 3782 9172 3834
rect 9196 3782 9226 3834
rect 9226 3782 9252 3834
rect 8956 3780 9012 3782
rect 9036 3780 9092 3782
rect 9116 3780 9172 3782
rect 9196 3780 9252 3782
rect 11794 13640 11850 13696
rect 11886 11636 11888 11656
rect 11888 11636 11940 11656
rect 11940 11636 11942 11656
rect 11886 11600 11942 11636
rect 12956 19610 13012 19612
rect 13036 19610 13092 19612
rect 13116 19610 13172 19612
rect 13196 19610 13252 19612
rect 12956 19558 12982 19610
rect 12982 19558 13012 19610
rect 13036 19558 13046 19610
rect 13046 19558 13092 19610
rect 13116 19558 13162 19610
rect 13162 19558 13172 19610
rect 13196 19558 13226 19610
rect 13226 19558 13252 19610
rect 12956 19556 13012 19558
rect 13036 19556 13092 19558
rect 13116 19556 13172 19558
rect 13196 19556 13252 19558
rect 12956 18522 13012 18524
rect 13036 18522 13092 18524
rect 13116 18522 13172 18524
rect 13196 18522 13252 18524
rect 12956 18470 12982 18522
rect 12982 18470 13012 18522
rect 13036 18470 13046 18522
rect 13046 18470 13092 18522
rect 13116 18470 13162 18522
rect 13162 18470 13172 18522
rect 13196 18470 13226 18522
rect 13226 18470 13252 18522
rect 12956 18468 13012 18470
rect 13036 18468 13092 18470
rect 13116 18468 13172 18470
rect 13196 18468 13252 18470
rect 12346 15544 12402 15600
rect 12956 17434 13012 17436
rect 13036 17434 13092 17436
rect 13116 17434 13172 17436
rect 13196 17434 13252 17436
rect 12956 17382 12982 17434
rect 12982 17382 13012 17434
rect 13036 17382 13046 17434
rect 13046 17382 13092 17434
rect 13116 17382 13162 17434
rect 13162 17382 13172 17434
rect 13196 17382 13226 17434
rect 13226 17382 13252 17434
rect 12956 17380 13012 17382
rect 13036 17380 13092 17382
rect 13116 17380 13172 17382
rect 13196 17380 13252 17382
rect 12956 16346 13012 16348
rect 13036 16346 13092 16348
rect 13116 16346 13172 16348
rect 13196 16346 13252 16348
rect 12956 16294 12982 16346
rect 12982 16294 13012 16346
rect 13036 16294 13046 16346
rect 13046 16294 13092 16346
rect 13116 16294 13162 16346
rect 13162 16294 13172 16346
rect 13196 16294 13226 16346
rect 13226 16294 13252 16346
rect 12956 16292 13012 16294
rect 13036 16292 13092 16294
rect 13116 16292 13172 16294
rect 13196 16292 13252 16294
rect 12806 16088 12862 16144
rect 12956 15258 13012 15260
rect 13036 15258 13092 15260
rect 13116 15258 13172 15260
rect 13196 15258 13252 15260
rect 12956 15206 12982 15258
rect 12982 15206 13012 15258
rect 13036 15206 13046 15258
rect 13046 15206 13092 15258
rect 13116 15206 13162 15258
rect 13162 15206 13172 15258
rect 13196 15206 13226 15258
rect 13226 15206 13252 15258
rect 12956 15204 13012 15206
rect 13036 15204 13092 15206
rect 13116 15204 13172 15206
rect 13196 15204 13252 15206
rect 12806 14456 12862 14512
rect 13450 17312 13506 17368
rect 12714 13912 12770 13968
rect 11978 11056 12034 11112
rect 11242 8880 11298 8936
rect 12956 14170 13012 14172
rect 13036 14170 13092 14172
rect 13116 14170 13172 14172
rect 13196 14170 13252 14172
rect 12956 14118 12982 14170
rect 12982 14118 13012 14170
rect 13036 14118 13046 14170
rect 13046 14118 13092 14170
rect 13116 14118 13162 14170
rect 13162 14118 13172 14170
rect 13196 14118 13226 14170
rect 13226 14118 13252 14170
rect 12956 14116 13012 14118
rect 13036 14116 13092 14118
rect 13116 14116 13172 14118
rect 13196 14116 13252 14118
rect 12956 13082 13012 13084
rect 13036 13082 13092 13084
rect 13116 13082 13172 13084
rect 13196 13082 13252 13084
rect 12956 13030 12982 13082
rect 12982 13030 13012 13082
rect 13036 13030 13046 13082
rect 13046 13030 13092 13082
rect 13116 13030 13162 13082
rect 13162 13030 13172 13082
rect 13196 13030 13226 13082
rect 13226 13030 13252 13082
rect 12956 13028 13012 13030
rect 13036 13028 13092 13030
rect 13116 13028 13172 13030
rect 13196 13028 13252 13030
rect 12956 11994 13012 11996
rect 13036 11994 13092 11996
rect 13116 11994 13172 11996
rect 13196 11994 13252 11996
rect 12956 11942 12982 11994
rect 12982 11942 13012 11994
rect 13036 11942 13046 11994
rect 13046 11942 13092 11994
rect 13116 11942 13162 11994
rect 13162 11942 13172 11994
rect 13196 11942 13226 11994
rect 13226 11942 13252 11994
rect 12956 11940 13012 11942
rect 13036 11940 13092 11942
rect 13116 11940 13172 11942
rect 13196 11940 13252 11942
rect 12956 10906 13012 10908
rect 13036 10906 13092 10908
rect 13116 10906 13172 10908
rect 13196 10906 13252 10908
rect 12956 10854 12982 10906
rect 12982 10854 13012 10906
rect 13036 10854 13046 10906
rect 13046 10854 13092 10906
rect 13116 10854 13162 10906
rect 13162 10854 13172 10906
rect 13196 10854 13226 10906
rect 13226 10854 13252 10906
rect 12956 10852 13012 10854
rect 13036 10852 13092 10854
rect 13116 10852 13172 10854
rect 13196 10852 13252 10854
rect 12622 5072 12678 5128
rect 8956 2746 9012 2748
rect 9036 2746 9092 2748
rect 9116 2746 9172 2748
rect 9196 2746 9252 2748
rect 8956 2694 8982 2746
rect 8982 2694 9012 2746
rect 9036 2694 9046 2746
rect 9046 2694 9092 2746
rect 9116 2694 9162 2746
rect 9162 2694 9172 2746
rect 9196 2694 9226 2746
rect 9226 2694 9252 2746
rect 8956 2692 9012 2694
rect 9036 2692 9092 2694
rect 9116 2692 9172 2694
rect 9196 2692 9252 2694
rect 12956 9818 13012 9820
rect 13036 9818 13092 9820
rect 13116 9818 13172 9820
rect 13196 9818 13252 9820
rect 12956 9766 12982 9818
rect 12982 9766 13012 9818
rect 13036 9766 13046 9818
rect 13046 9766 13092 9818
rect 13116 9766 13162 9818
rect 13162 9766 13172 9818
rect 13196 9766 13226 9818
rect 13226 9766 13252 9818
rect 12956 9764 13012 9766
rect 13036 9764 13092 9766
rect 13116 9764 13172 9766
rect 13196 9764 13252 9766
rect 12956 8730 13012 8732
rect 13036 8730 13092 8732
rect 13116 8730 13172 8732
rect 13196 8730 13252 8732
rect 12956 8678 12982 8730
rect 12982 8678 13012 8730
rect 13036 8678 13046 8730
rect 13046 8678 13092 8730
rect 13116 8678 13162 8730
rect 13162 8678 13172 8730
rect 13196 8678 13226 8730
rect 13226 8678 13252 8730
rect 12956 8676 13012 8678
rect 13036 8676 13092 8678
rect 13116 8676 13172 8678
rect 13196 8676 13252 8678
rect 12956 7642 13012 7644
rect 13036 7642 13092 7644
rect 13116 7642 13172 7644
rect 13196 7642 13252 7644
rect 12956 7590 12982 7642
rect 12982 7590 13012 7642
rect 13036 7590 13046 7642
rect 13046 7590 13092 7642
rect 13116 7590 13162 7642
rect 13162 7590 13172 7642
rect 13196 7590 13226 7642
rect 13226 7590 13252 7642
rect 12956 7588 13012 7590
rect 13036 7588 13092 7590
rect 13116 7588 13172 7590
rect 13196 7588 13252 7590
rect 14554 15544 14610 15600
rect 14370 15408 14426 15464
rect 14002 14456 14058 14512
rect 14830 9596 14832 9616
rect 14832 9596 14884 9616
rect 14884 9596 14886 9616
rect 14830 9560 14886 9596
rect 13358 7248 13414 7304
rect 12956 6554 13012 6556
rect 13036 6554 13092 6556
rect 13116 6554 13172 6556
rect 13196 6554 13252 6556
rect 12956 6502 12982 6554
rect 12982 6502 13012 6554
rect 13036 6502 13046 6554
rect 13046 6502 13092 6554
rect 13116 6502 13162 6554
rect 13162 6502 13172 6554
rect 13196 6502 13226 6554
rect 13226 6502 13252 6554
rect 12956 6500 13012 6502
rect 13036 6500 13092 6502
rect 13116 6500 13172 6502
rect 13196 6500 13252 6502
rect 14002 7248 14058 7304
rect 12956 5466 13012 5468
rect 13036 5466 13092 5468
rect 13116 5466 13172 5468
rect 13196 5466 13252 5468
rect 12956 5414 12982 5466
rect 12982 5414 13012 5466
rect 13036 5414 13046 5466
rect 13046 5414 13092 5466
rect 13116 5414 13162 5466
rect 13162 5414 13172 5466
rect 13196 5414 13226 5466
rect 13226 5414 13252 5466
rect 12956 5412 13012 5414
rect 13036 5412 13092 5414
rect 13116 5412 13172 5414
rect 13196 5412 13252 5414
rect 12956 4378 13012 4380
rect 13036 4378 13092 4380
rect 13116 4378 13172 4380
rect 13196 4378 13252 4380
rect 12956 4326 12982 4378
rect 12982 4326 13012 4378
rect 13036 4326 13046 4378
rect 13046 4326 13092 4378
rect 13116 4326 13162 4378
rect 13162 4326 13172 4378
rect 13196 4326 13226 4378
rect 13226 4326 13252 4378
rect 12956 4324 13012 4326
rect 13036 4324 13092 4326
rect 13116 4324 13172 4326
rect 13196 4324 13252 4326
rect 12806 3576 12862 3632
rect 12956 3290 13012 3292
rect 13036 3290 13092 3292
rect 13116 3290 13172 3292
rect 13196 3290 13252 3292
rect 12956 3238 12982 3290
rect 12982 3238 13012 3290
rect 13036 3238 13046 3290
rect 13046 3238 13092 3290
rect 13116 3238 13162 3290
rect 13162 3238 13172 3290
rect 13196 3238 13226 3290
rect 13226 3238 13252 3290
rect 12956 3236 13012 3238
rect 13036 3236 13092 3238
rect 13116 3236 13172 3238
rect 13196 3236 13252 3238
rect 12956 2202 13012 2204
rect 13036 2202 13092 2204
rect 13116 2202 13172 2204
rect 13196 2202 13252 2204
rect 12956 2150 12982 2202
rect 12982 2150 13012 2202
rect 13036 2150 13046 2202
rect 13046 2150 13092 2202
rect 13116 2150 13162 2202
rect 13162 2150 13172 2202
rect 13196 2150 13226 2202
rect 13226 2150 13252 2202
rect 12956 2148 13012 2150
rect 13036 2148 13092 2150
rect 13116 2148 13172 2150
rect 13196 2148 13252 2150
rect 14830 7384 14886 7440
rect 15750 18264 15806 18320
rect 15658 18128 15714 18184
rect 16578 15952 16634 16008
rect 15014 9016 15070 9072
rect 16210 7928 16266 7984
rect 16578 8472 16634 8528
rect 16956 21242 17012 21244
rect 17036 21242 17092 21244
rect 17116 21242 17172 21244
rect 17196 21242 17252 21244
rect 16956 21190 16982 21242
rect 16982 21190 17012 21242
rect 17036 21190 17046 21242
rect 17046 21190 17092 21242
rect 17116 21190 17162 21242
rect 17162 21190 17172 21242
rect 17196 21190 17226 21242
rect 17226 21190 17252 21242
rect 16956 21188 17012 21190
rect 17036 21188 17092 21190
rect 17116 21188 17172 21190
rect 17196 21188 17252 21190
rect 20074 22752 20130 22808
rect 19982 21936 20038 21992
rect 16956 20154 17012 20156
rect 17036 20154 17092 20156
rect 17116 20154 17172 20156
rect 17196 20154 17252 20156
rect 16956 20102 16982 20154
rect 16982 20102 17012 20154
rect 17036 20102 17046 20154
rect 17046 20102 17092 20154
rect 17116 20102 17162 20154
rect 17162 20102 17172 20154
rect 17196 20102 17226 20154
rect 17226 20102 17252 20154
rect 16956 20100 17012 20102
rect 17036 20100 17092 20102
rect 17116 20100 17172 20102
rect 17196 20100 17252 20102
rect 16956 19066 17012 19068
rect 17036 19066 17092 19068
rect 17116 19066 17172 19068
rect 17196 19066 17252 19068
rect 16956 19014 16982 19066
rect 16982 19014 17012 19066
rect 17036 19014 17046 19066
rect 17046 19014 17092 19066
rect 17116 19014 17162 19066
rect 17162 19014 17172 19066
rect 17196 19014 17226 19066
rect 17226 19014 17252 19066
rect 16956 19012 17012 19014
rect 17036 19012 17092 19014
rect 17116 19012 17172 19014
rect 17196 19012 17252 19014
rect 16956 17978 17012 17980
rect 17036 17978 17092 17980
rect 17116 17978 17172 17980
rect 17196 17978 17252 17980
rect 16956 17926 16982 17978
rect 16982 17926 17012 17978
rect 17036 17926 17046 17978
rect 17046 17926 17092 17978
rect 17116 17926 17162 17978
rect 17162 17926 17172 17978
rect 17196 17926 17226 17978
rect 17226 17926 17252 17978
rect 16956 17924 17012 17926
rect 17036 17924 17092 17926
rect 17116 17924 17172 17926
rect 17196 17924 17252 17926
rect 16956 16890 17012 16892
rect 17036 16890 17092 16892
rect 17116 16890 17172 16892
rect 17196 16890 17252 16892
rect 16956 16838 16982 16890
rect 16982 16838 17012 16890
rect 17036 16838 17046 16890
rect 17046 16838 17092 16890
rect 17116 16838 17162 16890
rect 17162 16838 17172 16890
rect 17196 16838 17226 16890
rect 17226 16838 17252 16890
rect 16956 16836 17012 16838
rect 17036 16836 17092 16838
rect 17116 16836 17172 16838
rect 17196 16836 17252 16838
rect 16956 15802 17012 15804
rect 17036 15802 17092 15804
rect 17116 15802 17172 15804
rect 17196 15802 17252 15804
rect 16956 15750 16982 15802
rect 16982 15750 17012 15802
rect 17036 15750 17046 15802
rect 17046 15750 17092 15802
rect 17116 15750 17162 15802
rect 17162 15750 17172 15802
rect 17196 15750 17226 15802
rect 17226 15750 17252 15802
rect 16956 15748 17012 15750
rect 17036 15748 17092 15750
rect 17116 15748 17172 15750
rect 17196 15748 17252 15750
rect 20956 21786 21012 21788
rect 21036 21786 21092 21788
rect 21116 21786 21172 21788
rect 21196 21786 21252 21788
rect 20956 21734 20982 21786
rect 20982 21734 21012 21786
rect 21036 21734 21046 21786
rect 21046 21734 21092 21786
rect 21116 21734 21162 21786
rect 21162 21734 21172 21786
rect 21196 21734 21226 21786
rect 21226 21734 21252 21786
rect 20956 21732 21012 21734
rect 21036 21732 21092 21734
rect 21116 21732 21172 21734
rect 21196 21732 21252 21734
rect 21454 20848 21510 20904
rect 20956 20698 21012 20700
rect 21036 20698 21092 20700
rect 21116 20698 21172 20700
rect 21196 20698 21252 20700
rect 20956 20646 20982 20698
rect 20982 20646 21012 20698
rect 21036 20646 21046 20698
rect 21046 20646 21092 20698
rect 21116 20646 21162 20698
rect 21162 20646 21172 20698
rect 21196 20646 21226 20698
rect 21226 20646 21252 20698
rect 20956 20644 21012 20646
rect 21036 20644 21092 20646
rect 21116 20644 21172 20646
rect 21196 20644 21252 20646
rect 18970 17040 19026 17096
rect 16956 14714 17012 14716
rect 17036 14714 17092 14716
rect 17116 14714 17172 14716
rect 17196 14714 17252 14716
rect 16956 14662 16982 14714
rect 16982 14662 17012 14714
rect 17036 14662 17046 14714
rect 17046 14662 17092 14714
rect 17116 14662 17162 14714
rect 17162 14662 17172 14714
rect 17196 14662 17226 14714
rect 17226 14662 17252 14714
rect 16956 14660 17012 14662
rect 17036 14660 17092 14662
rect 17116 14660 17172 14662
rect 17196 14660 17252 14662
rect 16956 13626 17012 13628
rect 17036 13626 17092 13628
rect 17116 13626 17172 13628
rect 17196 13626 17252 13628
rect 16956 13574 16982 13626
rect 16982 13574 17012 13626
rect 17036 13574 17046 13626
rect 17046 13574 17092 13626
rect 17116 13574 17162 13626
rect 17162 13574 17172 13626
rect 17196 13574 17226 13626
rect 17226 13574 17252 13626
rect 16956 13572 17012 13574
rect 17036 13572 17092 13574
rect 17116 13572 17172 13574
rect 17196 13572 17252 13574
rect 16956 12538 17012 12540
rect 17036 12538 17092 12540
rect 17116 12538 17172 12540
rect 17196 12538 17252 12540
rect 16956 12486 16982 12538
rect 16982 12486 17012 12538
rect 17036 12486 17046 12538
rect 17046 12486 17092 12538
rect 17116 12486 17162 12538
rect 17162 12486 17172 12538
rect 17196 12486 17226 12538
rect 17226 12486 17252 12538
rect 16956 12484 17012 12486
rect 17036 12484 17092 12486
rect 17116 12484 17172 12486
rect 17196 12484 17252 12486
rect 16956 11450 17012 11452
rect 17036 11450 17092 11452
rect 17116 11450 17172 11452
rect 17196 11450 17252 11452
rect 16956 11398 16982 11450
rect 16982 11398 17012 11450
rect 17036 11398 17046 11450
rect 17046 11398 17092 11450
rect 17116 11398 17162 11450
rect 17162 11398 17172 11450
rect 17196 11398 17226 11450
rect 17226 11398 17252 11450
rect 16956 11396 17012 11398
rect 17036 11396 17092 11398
rect 17116 11396 17172 11398
rect 17196 11396 17252 11398
rect 16854 11056 16910 11112
rect 16956 10362 17012 10364
rect 17036 10362 17092 10364
rect 17116 10362 17172 10364
rect 17196 10362 17252 10364
rect 16956 10310 16982 10362
rect 16982 10310 17012 10362
rect 17036 10310 17046 10362
rect 17046 10310 17092 10362
rect 17116 10310 17162 10362
rect 17162 10310 17172 10362
rect 17196 10310 17226 10362
rect 17226 10310 17252 10362
rect 16956 10308 17012 10310
rect 17036 10308 17092 10310
rect 17116 10308 17172 10310
rect 17196 10308 17252 10310
rect 16956 9274 17012 9276
rect 17036 9274 17092 9276
rect 17116 9274 17172 9276
rect 17196 9274 17252 9276
rect 16956 9222 16982 9274
rect 16982 9222 17012 9274
rect 17036 9222 17046 9274
rect 17046 9222 17092 9274
rect 17116 9222 17162 9274
rect 17162 9222 17172 9274
rect 17196 9222 17226 9274
rect 17226 9222 17252 9274
rect 16956 9220 17012 9222
rect 17036 9220 17092 9222
rect 17116 9220 17172 9222
rect 17196 9220 17252 9222
rect 16670 7928 16726 7984
rect 16394 5208 16450 5264
rect 15474 4120 15530 4176
rect 16956 8186 17012 8188
rect 17036 8186 17092 8188
rect 17116 8186 17172 8188
rect 17196 8186 17252 8188
rect 16956 8134 16982 8186
rect 16982 8134 17012 8186
rect 17036 8134 17046 8186
rect 17046 8134 17092 8186
rect 17116 8134 17162 8186
rect 17162 8134 17172 8186
rect 17196 8134 17226 8186
rect 17226 8134 17252 8186
rect 16956 8132 17012 8134
rect 17036 8132 17092 8134
rect 17116 8132 17172 8134
rect 17196 8132 17252 8134
rect 16956 7098 17012 7100
rect 17036 7098 17092 7100
rect 17116 7098 17172 7100
rect 17196 7098 17252 7100
rect 16956 7046 16982 7098
rect 16982 7046 17012 7098
rect 17036 7046 17046 7098
rect 17046 7046 17092 7098
rect 17116 7046 17162 7098
rect 17162 7046 17172 7098
rect 17196 7046 17226 7098
rect 17226 7046 17252 7098
rect 16956 7044 17012 7046
rect 17036 7044 17092 7046
rect 17116 7044 17172 7046
rect 17196 7044 17252 7046
rect 16956 6010 17012 6012
rect 17036 6010 17092 6012
rect 17116 6010 17172 6012
rect 17196 6010 17252 6012
rect 16956 5958 16982 6010
rect 16982 5958 17012 6010
rect 17036 5958 17046 6010
rect 17046 5958 17092 6010
rect 17116 5958 17162 6010
rect 17162 5958 17172 6010
rect 17196 5958 17226 6010
rect 17226 5958 17252 6010
rect 16956 5956 17012 5958
rect 17036 5956 17092 5958
rect 17116 5956 17172 5958
rect 17196 5956 17252 5958
rect 16956 4922 17012 4924
rect 17036 4922 17092 4924
rect 17116 4922 17172 4924
rect 17196 4922 17252 4924
rect 16956 4870 16982 4922
rect 16982 4870 17012 4922
rect 17036 4870 17046 4922
rect 17046 4870 17092 4922
rect 17116 4870 17162 4922
rect 17162 4870 17172 4922
rect 17196 4870 17226 4922
rect 17226 4870 17252 4922
rect 16956 4868 17012 4870
rect 17036 4868 17092 4870
rect 17116 4868 17172 4870
rect 17196 4868 17252 4870
rect 18878 13640 18934 13696
rect 17866 10376 17922 10432
rect 19338 16496 19394 16552
rect 19890 17312 19946 17368
rect 19798 16088 19854 16144
rect 19246 13368 19302 13424
rect 16956 3834 17012 3836
rect 17036 3834 17092 3836
rect 17116 3834 17172 3836
rect 17196 3834 17252 3836
rect 16956 3782 16982 3834
rect 16982 3782 17012 3834
rect 17036 3782 17046 3834
rect 17046 3782 17092 3834
rect 17116 3782 17162 3834
rect 17162 3782 17172 3834
rect 17196 3782 17226 3834
rect 17226 3782 17252 3834
rect 16956 3780 17012 3782
rect 17036 3780 17092 3782
rect 17116 3780 17172 3782
rect 17196 3780 17252 3782
rect 19154 6160 19210 6216
rect 17314 2896 17370 2952
rect 16956 2746 17012 2748
rect 17036 2746 17092 2748
rect 17116 2746 17172 2748
rect 17196 2746 17252 2748
rect 16956 2694 16982 2746
rect 16982 2694 17012 2746
rect 17036 2694 17046 2746
rect 17046 2694 17092 2746
rect 17116 2694 17162 2746
rect 17162 2694 17172 2746
rect 17196 2694 17226 2746
rect 17226 2694 17252 2746
rect 16956 2692 17012 2694
rect 17036 2692 17092 2694
rect 17116 2692 17172 2694
rect 17196 2692 17252 2694
rect 18970 1808 19026 1864
rect 20956 19610 21012 19612
rect 21036 19610 21092 19612
rect 21116 19610 21172 19612
rect 21196 19610 21252 19612
rect 20956 19558 20982 19610
rect 20982 19558 21012 19610
rect 21036 19558 21046 19610
rect 21046 19558 21092 19610
rect 21116 19558 21162 19610
rect 21162 19558 21172 19610
rect 21196 19558 21226 19610
rect 21226 19558 21252 19610
rect 20956 19556 21012 19558
rect 21036 19556 21092 19558
rect 21116 19556 21172 19558
rect 21196 19556 21252 19558
rect 21270 18808 21326 18864
rect 20956 18522 21012 18524
rect 21036 18522 21092 18524
rect 21116 18522 21172 18524
rect 21196 18522 21252 18524
rect 20956 18470 20982 18522
rect 20982 18470 21012 18522
rect 21036 18470 21046 18522
rect 21046 18470 21092 18522
rect 21116 18470 21162 18522
rect 21162 18470 21172 18522
rect 21196 18470 21226 18522
rect 21226 18470 21252 18522
rect 20956 18468 21012 18470
rect 21036 18468 21092 18470
rect 21116 18468 21172 18470
rect 21196 18468 21252 18470
rect 20956 17434 21012 17436
rect 21036 17434 21092 17436
rect 21116 17434 21172 17436
rect 21196 17434 21252 17436
rect 20956 17382 20982 17434
rect 20982 17382 21012 17434
rect 21036 17382 21046 17434
rect 21046 17382 21092 17434
rect 21116 17382 21162 17434
rect 21162 17382 21172 17434
rect 21196 17382 21226 17434
rect 21226 17382 21252 17434
rect 20956 17380 21012 17382
rect 21036 17380 21092 17382
rect 21116 17380 21172 17382
rect 21196 17380 21252 17382
rect 21638 19760 21694 19816
rect 21730 17992 21786 18048
rect 20902 17176 20958 17232
rect 19890 12416 19946 12472
rect 20074 13640 20130 13696
rect 20258 13368 20314 13424
rect 21730 16904 21786 16960
rect 20956 16346 21012 16348
rect 21036 16346 21092 16348
rect 21116 16346 21172 16348
rect 21196 16346 21252 16348
rect 20956 16294 20982 16346
rect 20982 16294 21012 16346
rect 21036 16294 21046 16346
rect 21046 16294 21092 16346
rect 21116 16294 21162 16346
rect 21162 16294 21172 16346
rect 21196 16294 21226 16346
rect 21226 16294 21252 16346
rect 20956 16292 21012 16294
rect 21036 16292 21092 16294
rect 21116 16292 21172 16294
rect 21196 16292 21252 16294
rect 21454 15816 21510 15872
rect 20956 15258 21012 15260
rect 21036 15258 21092 15260
rect 21116 15258 21172 15260
rect 21196 15258 21252 15260
rect 20956 15206 20982 15258
rect 20982 15206 21012 15258
rect 21036 15206 21046 15258
rect 21046 15206 21092 15258
rect 21116 15206 21162 15258
rect 21162 15206 21172 15258
rect 21196 15206 21226 15258
rect 21226 15206 21252 15258
rect 20956 15204 21012 15206
rect 21036 15204 21092 15206
rect 21116 15204 21172 15206
rect 21196 15204 21252 15206
rect 20956 14170 21012 14172
rect 21036 14170 21092 14172
rect 21116 14170 21172 14172
rect 21196 14170 21252 14172
rect 20956 14118 20982 14170
rect 20982 14118 21012 14170
rect 21036 14118 21046 14170
rect 21046 14118 21092 14170
rect 21116 14118 21162 14170
rect 21162 14118 21172 14170
rect 21196 14118 21226 14170
rect 21226 14118 21252 14170
rect 20956 14116 21012 14118
rect 21036 14116 21092 14118
rect 21116 14116 21172 14118
rect 21196 14116 21252 14118
rect 20956 13082 21012 13084
rect 21036 13082 21092 13084
rect 21116 13082 21172 13084
rect 21196 13082 21252 13084
rect 20956 13030 20982 13082
rect 20982 13030 21012 13082
rect 21036 13030 21046 13082
rect 21046 13030 21092 13082
rect 21116 13030 21162 13082
rect 21162 13030 21172 13082
rect 21196 13030 21226 13082
rect 21226 13030 21252 13082
rect 20956 13028 21012 13030
rect 21036 13028 21092 13030
rect 21116 13028 21172 13030
rect 21196 13028 21252 13030
rect 21362 12960 21418 13016
rect 20956 11994 21012 11996
rect 21036 11994 21092 11996
rect 21116 11994 21172 11996
rect 21196 11994 21252 11996
rect 20956 11942 20982 11994
rect 20982 11942 21012 11994
rect 21036 11942 21046 11994
rect 21046 11942 21092 11994
rect 21116 11942 21162 11994
rect 21162 11942 21172 11994
rect 21196 11942 21226 11994
rect 21226 11942 21252 11994
rect 20956 11940 21012 11942
rect 21036 11940 21092 11942
rect 21116 11940 21172 11942
rect 21196 11940 21252 11942
rect 20810 11600 20866 11656
rect 20956 10906 21012 10908
rect 21036 10906 21092 10908
rect 21116 10906 21172 10908
rect 21196 10906 21252 10908
rect 20956 10854 20982 10906
rect 20982 10854 21012 10906
rect 21036 10854 21046 10906
rect 21046 10854 21092 10906
rect 21116 10854 21162 10906
rect 21162 10854 21172 10906
rect 21196 10854 21226 10906
rect 21226 10854 21252 10906
rect 20956 10852 21012 10854
rect 21036 10852 21092 10854
rect 21116 10852 21172 10854
rect 21196 10852 21252 10854
rect 21362 10784 21418 10840
rect 20902 10512 20958 10568
rect 20956 9818 21012 9820
rect 21036 9818 21092 9820
rect 21116 9818 21172 9820
rect 21196 9818 21252 9820
rect 20956 9766 20982 9818
rect 20982 9766 21012 9818
rect 21036 9766 21046 9818
rect 21046 9766 21092 9818
rect 21116 9766 21162 9818
rect 21162 9766 21172 9818
rect 21196 9766 21226 9818
rect 21226 9766 21252 9818
rect 20956 9764 21012 9766
rect 21036 9764 21092 9766
rect 21116 9764 21172 9766
rect 21196 9764 21252 9766
rect 20956 8730 21012 8732
rect 21036 8730 21092 8732
rect 21116 8730 21172 8732
rect 21196 8730 21252 8732
rect 20956 8678 20982 8730
rect 20982 8678 21012 8730
rect 21036 8678 21046 8730
rect 21046 8678 21092 8730
rect 21116 8678 21162 8730
rect 21162 8678 21172 8730
rect 21196 8678 21226 8730
rect 21226 8678 21252 8730
rect 20956 8676 21012 8678
rect 21036 8676 21092 8678
rect 21116 8676 21172 8678
rect 21196 8676 21252 8678
rect 21270 7792 21326 7848
rect 20956 7642 21012 7644
rect 21036 7642 21092 7644
rect 21116 7642 21172 7644
rect 21196 7642 21252 7644
rect 20956 7590 20982 7642
rect 20982 7590 21012 7642
rect 21036 7590 21046 7642
rect 21046 7590 21092 7642
rect 21116 7590 21162 7642
rect 21162 7590 21172 7642
rect 21196 7590 21226 7642
rect 21226 7590 21252 7642
rect 20956 7588 21012 7590
rect 21036 7588 21092 7590
rect 21116 7588 21172 7590
rect 21196 7588 21252 7590
rect 20956 6554 21012 6556
rect 21036 6554 21092 6556
rect 21116 6554 21172 6556
rect 21196 6554 21252 6556
rect 20956 6502 20982 6554
rect 20982 6502 21012 6554
rect 21036 6502 21046 6554
rect 21046 6502 21092 6554
rect 21116 6502 21162 6554
rect 21162 6502 21172 6554
rect 21196 6502 21226 6554
rect 21226 6502 21252 6554
rect 20956 6500 21012 6502
rect 21036 6500 21092 6502
rect 21116 6500 21172 6502
rect 21196 6500 21252 6502
rect 21362 6432 21418 6488
rect 20956 5466 21012 5468
rect 21036 5466 21092 5468
rect 21116 5466 21172 5468
rect 21196 5466 21252 5468
rect 20956 5414 20982 5466
rect 20982 5414 21012 5466
rect 21036 5414 21046 5466
rect 21046 5414 21092 5466
rect 21116 5414 21162 5466
rect 21162 5414 21172 5466
rect 21196 5414 21226 5466
rect 21226 5414 21252 5466
rect 20956 5412 21012 5414
rect 21036 5412 21092 5414
rect 21116 5412 21172 5414
rect 21196 5412 21252 5414
rect 21270 5072 21326 5128
rect 23570 14320 23626 14376
rect 23570 9424 23626 9480
rect 21914 5344 21970 5400
rect 21730 4936 21786 4992
rect 20956 4378 21012 4380
rect 21036 4378 21092 4380
rect 21116 4378 21172 4380
rect 21196 4378 21252 4380
rect 20956 4326 20982 4378
rect 20982 4326 21012 4378
rect 21036 4326 21046 4378
rect 21046 4326 21092 4378
rect 21116 4326 21162 4378
rect 21162 4326 21172 4378
rect 21196 4326 21226 4378
rect 21226 4326 21252 4378
rect 20956 4324 21012 4326
rect 21036 4324 21092 4326
rect 21116 4324 21172 4326
rect 21196 4324 21252 4326
rect 23570 3984 23626 4040
rect 20810 3576 20866 3632
rect 21454 3440 21510 3496
rect 20956 3290 21012 3292
rect 21036 3290 21092 3292
rect 21116 3290 21172 3292
rect 21196 3290 21252 3292
rect 20956 3238 20982 3290
rect 20982 3238 21012 3290
rect 21036 3238 21046 3290
rect 21046 3238 21092 3290
rect 21116 3238 21162 3290
rect 21162 3238 21172 3290
rect 21196 3238 21226 3290
rect 21226 3238 21252 3290
rect 20956 3236 21012 3238
rect 21036 3236 21092 3238
rect 21116 3236 21172 3238
rect 21196 3236 21252 3238
rect 20956 2202 21012 2204
rect 21036 2202 21092 2204
rect 21116 2202 21172 2204
rect 21196 2202 21252 2204
rect 20956 2150 20982 2202
rect 20982 2150 21012 2202
rect 21036 2150 21046 2202
rect 21046 2150 21092 2202
rect 21116 2150 21162 2202
rect 21162 2150 21172 2202
rect 21196 2150 21226 2202
rect 21226 2150 21252 2202
rect 20956 2148 21012 2150
rect 21036 2148 21092 2150
rect 21116 2148 21172 2150
rect 21196 2148 21252 2150
rect 21362 1672 21418 1728
rect 23570 1400 23626 1456
<< metal3 >>
rect 23520 23264 24000 23384
rect 0 22992 480 23112
rect 62 22538 122 22992
rect 20069 22810 20135 22813
rect 23614 22810 23674 23264
rect 20069 22808 23674 22810
rect 20069 22752 20074 22808
rect 20130 22752 23674 22808
rect 20069 22750 23674 22752
rect 20069 22747 20135 22750
rect 1301 22538 1367 22541
rect 62 22536 1367 22538
rect 62 22480 1306 22536
rect 1362 22480 1367 22536
rect 62 22478 1367 22480
rect 1301 22475 1367 22478
rect 23520 22312 24000 22432
rect 19977 21994 20043 21997
rect 23614 21994 23674 22312
rect 19977 21992 23674 21994
rect 19977 21936 19982 21992
rect 20038 21936 23674 21992
rect 19977 21934 23674 21936
rect 19977 21931 20043 21934
rect 4944 21792 5264 21793
rect 4944 21728 4952 21792
rect 5016 21728 5032 21792
rect 5096 21728 5112 21792
rect 5176 21728 5192 21792
rect 5256 21728 5264 21792
rect 4944 21727 5264 21728
rect 12944 21792 13264 21793
rect 12944 21728 12952 21792
rect 13016 21728 13032 21792
rect 13096 21728 13112 21792
rect 13176 21728 13192 21792
rect 13256 21728 13264 21792
rect 12944 21727 13264 21728
rect 20944 21792 21264 21793
rect 20944 21728 20952 21792
rect 21016 21728 21032 21792
rect 21096 21728 21112 21792
rect 21176 21728 21192 21792
rect 21256 21728 21264 21792
rect 20944 21727 21264 21728
rect 23520 21360 24000 21480
rect 0 21224 480 21344
rect 8944 21248 9264 21249
rect 62 20770 122 21224
rect 8944 21184 8952 21248
rect 9016 21184 9032 21248
rect 9096 21184 9112 21248
rect 9176 21184 9192 21248
rect 9256 21184 9264 21248
rect 8944 21183 9264 21184
rect 16944 21248 17264 21249
rect 16944 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17264 21248
rect 16944 21183 17264 21184
rect 21449 20906 21515 20909
rect 23614 20906 23674 21360
rect 21449 20904 23674 20906
rect 21449 20848 21454 20904
rect 21510 20848 23674 20904
rect 21449 20846 23674 20848
rect 21449 20843 21515 20846
rect 1577 20770 1643 20773
rect 62 20768 1643 20770
rect 62 20712 1582 20768
rect 1638 20712 1643 20768
rect 62 20710 1643 20712
rect 1577 20707 1643 20710
rect 4944 20704 5264 20705
rect 4944 20640 4952 20704
rect 5016 20640 5032 20704
rect 5096 20640 5112 20704
rect 5176 20640 5192 20704
rect 5256 20640 5264 20704
rect 4944 20639 5264 20640
rect 12944 20704 13264 20705
rect 12944 20640 12952 20704
rect 13016 20640 13032 20704
rect 13096 20640 13112 20704
rect 13176 20640 13192 20704
rect 13256 20640 13264 20704
rect 12944 20639 13264 20640
rect 20944 20704 21264 20705
rect 20944 20640 20952 20704
rect 21016 20640 21032 20704
rect 21096 20640 21112 20704
rect 21176 20640 21192 20704
rect 21256 20640 21264 20704
rect 20944 20639 21264 20640
rect 23520 20272 24000 20392
rect 8944 20160 9264 20161
rect 8944 20096 8952 20160
rect 9016 20096 9032 20160
rect 9096 20096 9112 20160
rect 9176 20096 9192 20160
rect 9256 20096 9264 20160
rect 8944 20095 9264 20096
rect 16944 20160 17264 20161
rect 16944 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17264 20160
rect 16944 20095 17264 20096
rect 21633 19818 21699 19821
rect 23614 19818 23674 20272
rect 21633 19816 23674 19818
rect 21633 19760 21638 19816
rect 21694 19760 23674 19816
rect 21633 19758 23674 19760
rect 21633 19755 21699 19758
rect 0 19592 480 19712
rect 4944 19616 5264 19617
rect 62 19274 122 19592
rect 4944 19552 4952 19616
rect 5016 19552 5032 19616
rect 5096 19552 5112 19616
rect 5176 19552 5192 19616
rect 5256 19552 5264 19616
rect 4944 19551 5264 19552
rect 12944 19616 13264 19617
rect 12944 19552 12952 19616
rect 13016 19552 13032 19616
rect 13096 19552 13112 19616
rect 13176 19552 13192 19616
rect 13256 19552 13264 19616
rect 12944 19551 13264 19552
rect 20944 19616 21264 19617
rect 20944 19552 20952 19616
rect 21016 19552 21032 19616
rect 21096 19552 21112 19616
rect 21176 19552 21192 19616
rect 21256 19552 21264 19616
rect 20944 19551 21264 19552
rect 23520 19320 24000 19440
rect 2221 19274 2287 19277
rect 62 19272 2287 19274
rect 62 19216 2226 19272
rect 2282 19216 2287 19272
rect 62 19214 2287 19216
rect 2221 19211 2287 19214
rect 8944 19072 9264 19073
rect 8944 19008 8952 19072
rect 9016 19008 9032 19072
rect 9096 19008 9112 19072
rect 9176 19008 9192 19072
rect 9256 19008 9264 19072
rect 8944 19007 9264 19008
rect 16944 19072 17264 19073
rect 16944 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17264 19072
rect 16944 19007 17264 19008
rect 21265 18866 21331 18869
rect 23614 18866 23674 19320
rect 21265 18864 23674 18866
rect 21265 18808 21270 18864
rect 21326 18808 23674 18864
rect 21265 18806 23674 18808
rect 21265 18803 21331 18806
rect 4944 18528 5264 18529
rect 4944 18464 4952 18528
rect 5016 18464 5032 18528
rect 5096 18464 5112 18528
rect 5176 18464 5192 18528
rect 5256 18464 5264 18528
rect 4944 18463 5264 18464
rect 12944 18528 13264 18529
rect 12944 18464 12952 18528
rect 13016 18464 13032 18528
rect 13096 18464 13112 18528
rect 13176 18464 13192 18528
rect 13256 18464 13264 18528
rect 12944 18463 13264 18464
rect 20944 18528 21264 18529
rect 20944 18464 20952 18528
rect 21016 18464 21032 18528
rect 21096 18464 21112 18528
rect 21176 18464 21192 18528
rect 21256 18464 21264 18528
rect 20944 18463 21264 18464
rect 23520 18368 24000 18488
rect 5809 18322 5875 18325
rect 15745 18322 15811 18325
rect 5809 18320 15811 18322
rect 5809 18264 5814 18320
rect 5870 18264 15750 18320
rect 15806 18264 15811 18320
rect 5809 18262 15811 18264
rect 5809 18259 5875 18262
rect 15745 18259 15811 18262
rect 7097 18186 7163 18189
rect 15653 18186 15719 18189
rect 7097 18184 15719 18186
rect 7097 18128 7102 18184
rect 7158 18128 15658 18184
rect 15714 18128 15719 18184
rect 7097 18126 15719 18128
rect 7097 18123 7163 18126
rect 15653 18123 15719 18126
rect 21725 18050 21791 18053
rect 23614 18050 23674 18368
rect 21725 18048 23674 18050
rect 21725 17992 21730 18048
rect 21786 17992 23674 18048
rect 21725 17990 23674 17992
rect 21725 17987 21791 17990
rect 8944 17984 9264 17985
rect 0 17912 480 17944
rect 8944 17920 8952 17984
rect 9016 17920 9032 17984
rect 9096 17920 9112 17984
rect 9176 17920 9192 17984
rect 9256 17920 9264 17984
rect 8944 17919 9264 17920
rect 16944 17984 17264 17985
rect 16944 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17264 17984
rect 16944 17919 17264 17920
rect 0 17856 110 17912
rect 166 17856 480 17912
rect 0 17824 480 17856
rect 4944 17440 5264 17441
rect 4944 17376 4952 17440
rect 5016 17376 5032 17440
rect 5096 17376 5112 17440
rect 5176 17376 5192 17440
rect 5256 17376 5264 17440
rect 4944 17375 5264 17376
rect 12944 17440 13264 17441
rect 12944 17376 12952 17440
rect 13016 17376 13032 17440
rect 13096 17376 13112 17440
rect 13176 17376 13192 17440
rect 13256 17376 13264 17440
rect 12944 17375 13264 17376
rect 20944 17440 21264 17441
rect 20944 17376 20952 17440
rect 21016 17376 21032 17440
rect 21096 17376 21112 17440
rect 21176 17376 21192 17440
rect 21256 17376 21264 17440
rect 20944 17375 21264 17376
rect 13445 17370 13511 17373
rect 19885 17370 19951 17373
rect 13445 17368 19951 17370
rect 13445 17312 13450 17368
rect 13506 17312 19890 17368
rect 19946 17312 19951 17368
rect 13445 17310 19951 17312
rect 13445 17307 13511 17310
rect 19885 17307 19951 17310
rect 23520 17280 24000 17400
rect 10869 17234 10935 17237
rect 20897 17234 20963 17237
rect 10869 17232 20963 17234
rect 10869 17176 10874 17232
rect 10930 17176 20902 17232
rect 20958 17176 20963 17232
rect 10869 17174 20963 17176
rect 10869 17171 10935 17174
rect 20897 17171 20963 17174
rect 6637 17098 6703 17101
rect 8661 17098 8727 17101
rect 18965 17098 19031 17101
rect 6637 17096 19031 17098
rect 6637 17040 6642 17096
rect 6698 17040 8666 17096
rect 8722 17040 18970 17096
rect 19026 17040 19031 17096
rect 6637 17038 19031 17040
rect 6637 17035 6703 17038
rect 8661 17035 8727 17038
rect 18965 17035 19031 17038
rect 21725 16962 21791 16965
rect 23614 16962 23674 17280
rect 21725 16960 23674 16962
rect 21725 16904 21730 16960
rect 21786 16904 23674 16960
rect 21725 16902 23674 16904
rect 21725 16899 21791 16902
rect 8944 16896 9264 16897
rect 8944 16832 8952 16896
rect 9016 16832 9032 16896
rect 9096 16832 9112 16896
rect 9176 16832 9192 16896
rect 9256 16832 9264 16896
rect 8944 16831 9264 16832
rect 16944 16896 17264 16897
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 16944 16831 17264 16832
rect 7189 16554 7255 16557
rect 19333 16554 19399 16557
rect 7189 16552 19399 16554
rect 7189 16496 7194 16552
rect 7250 16496 19338 16552
rect 19394 16496 19399 16552
rect 7189 16494 19399 16496
rect 7189 16491 7255 16494
rect 19333 16491 19399 16494
rect 4944 16352 5264 16353
rect 0 16280 480 16312
rect 4944 16288 4952 16352
rect 5016 16288 5032 16352
rect 5096 16288 5112 16352
rect 5176 16288 5192 16352
rect 5256 16288 5264 16352
rect 4944 16287 5264 16288
rect 12944 16352 13264 16353
rect 12944 16288 12952 16352
rect 13016 16288 13032 16352
rect 13096 16288 13112 16352
rect 13176 16288 13192 16352
rect 13256 16288 13264 16352
rect 12944 16287 13264 16288
rect 20944 16352 21264 16353
rect 20944 16288 20952 16352
rect 21016 16288 21032 16352
rect 21096 16288 21112 16352
rect 21176 16288 21192 16352
rect 21256 16288 21264 16352
rect 23520 16328 24000 16448
rect 20944 16287 21264 16288
rect 0 16224 110 16280
rect 166 16224 480 16280
rect 0 16192 480 16224
rect 12801 16146 12867 16149
rect 19793 16146 19859 16149
rect 12801 16144 19859 16146
rect 12801 16088 12806 16144
rect 12862 16088 19798 16144
rect 19854 16088 19859 16144
rect 12801 16086 19859 16088
rect 12801 16083 12867 16086
rect 19793 16083 19859 16086
rect 8845 16010 8911 16013
rect 16573 16010 16639 16013
rect 8845 16008 16639 16010
rect 8845 15952 8850 16008
rect 8906 15952 16578 16008
rect 16634 15952 16639 16008
rect 8845 15950 16639 15952
rect 8845 15947 8911 15950
rect 16573 15947 16639 15950
rect 21449 15874 21515 15877
rect 23614 15874 23674 16328
rect 21449 15872 23674 15874
rect 21449 15816 21454 15872
rect 21510 15816 23674 15872
rect 21449 15814 23674 15816
rect 21449 15811 21515 15814
rect 8944 15808 9264 15809
rect 8944 15744 8952 15808
rect 9016 15744 9032 15808
rect 9096 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9264 15808
rect 8944 15743 9264 15744
rect 16944 15808 17264 15809
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16944 15743 17264 15744
rect 23606 15738 23612 15740
rect 19290 15678 23612 15738
rect 12341 15602 12407 15605
rect 14549 15602 14615 15605
rect 19290 15602 19350 15678
rect 23606 15676 23612 15678
rect 23676 15676 23682 15740
rect 12341 15600 19350 15602
rect 12341 15544 12346 15600
rect 12402 15544 14554 15600
rect 14610 15544 19350 15600
rect 12341 15542 19350 15544
rect 12341 15539 12407 15542
rect 14549 15539 14615 15542
rect 8109 15466 8175 15469
rect 14365 15466 14431 15469
rect 23520 15468 24000 15496
rect 23520 15466 23612 15468
rect 8109 15464 14431 15466
rect 8109 15408 8114 15464
rect 8170 15408 14370 15464
rect 14426 15408 14431 15464
rect 8109 15406 14431 15408
rect 23484 15406 23612 15466
rect 8109 15403 8175 15406
rect 14365 15403 14431 15406
rect 23520 15404 23612 15406
rect 23676 15404 24000 15468
rect 23520 15376 24000 15404
rect 4944 15264 5264 15265
rect 4944 15200 4952 15264
rect 5016 15200 5032 15264
rect 5096 15200 5112 15264
rect 5176 15200 5192 15264
rect 5256 15200 5264 15264
rect 4944 15199 5264 15200
rect 12944 15264 13264 15265
rect 12944 15200 12952 15264
rect 13016 15200 13032 15264
rect 13096 15200 13112 15264
rect 13176 15200 13192 15264
rect 13256 15200 13264 15264
rect 12944 15199 13264 15200
rect 20944 15264 21264 15265
rect 20944 15200 20952 15264
rect 21016 15200 21032 15264
rect 21096 15200 21112 15264
rect 21176 15200 21192 15264
rect 21256 15200 21264 15264
rect 20944 15199 21264 15200
rect 3509 14786 3575 14789
rect 8201 14786 8267 14789
rect 3509 14784 8267 14786
rect 3509 14728 3514 14784
rect 3570 14728 8206 14784
rect 8262 14728 8267 14784
rect 3509 14726 8267 14728
rect 3509 14723 3575 14726
rect 8201 14723 8267 14726
rect 8944 14720 9264 14721
rect 8944 14656 8952 14720
rect 9016 14656 9032 14720
rect 9096 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9264 14720
rect 8944 14655 9264 14656
rect 16944 14720 17264 14721
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16944 14655 17264 14656
rect 0 14424 480 14544
rect 12801 14514 12867 14517
rect 13997 14514 14063 14517
rect 12801 14512 14063 14514
rect 12801 14456 12806 14512
rect 12862 14456 14002 14512
rect 14058 14456 14063 14512
rect 12801 14454 14063 14456
rect 12801 14451 12867 14454
rect 13997 14451 14063 14454
rect 62 13970 122 14424
rect 23520 14378 24000 14408
rect 23484 14376 24000 14378
rect 23484 14320 23570 14376
rect 23626 14320 24000 14376
rect 23484 14318 24000 14320
rect 23520 14288 24000 14318
rect 4944 14176 5264 14177
rect 4944 14112 4952 14176
rect 5016 14112 5032 14176
rect 5096 14112 5112 14176
rect 5176 14112 5192 14176
rect 5256 14112 5264 14176
rect 4944 14111 5264 14112
rect 12944 14176 13264 14177
rect 12944 14112 12952 14176
rect 13016 14112 13032 14176
rect 13096 14112 13112 14176
rect 13176 14112 13192 14176
rect 13256 14112 13264 14176
rect 12944 14111 13264 14112
rect 20944 14176 21264 14177
rect 20944 14112 20952 14176
rect 21016 14112 21032 14176
rect 21096 14112 21112 14176
rect 21176 14112 21192 14176
rect 21256 14112 21264 14176
rect 20944 14111 21264 14112
rect 11329 13970 11395 13973
rect 12709 13970 12775 13973
rect 62 13968 12775 13970
rect 62 13912 11334 13968
rect 11390 13912 12714 13968
rect 12770 13912 12775 13968
rect 62 13910 12775 13912
rect 11329 13907 11395 13910
rect 12709 13907 12775 13910
rect 5349 13834 5415 13837
rect 5533 13834 5599 13837
rect 7833 13834 7899 13837
rect 5349 13832 7899 13834
rect 5349 13776 5354 13832
rect 5410 13776 5538 13832
rect 5594 13776 7838 13832
rect 7894 13776 7899 13832
rect 5349 13774 7899 13776
rect 5349 13771 5415 13774
rect 5533 13771 5599 13774
rect 7833 13771 7899 13774
rect 9397 13698 9463 13701
rect 11789 13698 11855 13701
rect 9397 13696 11855 13698
rect 9397 13640 9402 13696
rect 9458 13640 11794 13696
rect 11850 13640 11855 13696
rect 9397 13638 11855 13640
rect 9397 13635 9463 13638
rect 11789 13635 11855 13638
rect 18873 13698 18939 13701
rect 20069 13698 20135 13701
rect 18873 13696 20135 13698
rect 18873 13640 18878 13696
rect 18934 13640 20074 13696
rect 20130 13640 20135 13696
rect 18873 13638 20135 13640
rect 18873 13635 18939 13638
rect 20069 13635 20135 13638
rect 8944 13632 9264 13633
rect 8944 13568 8952 13632
rect 9016 13568 9032 13632
rect 9096 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9264 13632
rect 8944 13567 9264 13568
rect 16944 13632 17264 13633
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 13567 17264 13568
rect 19241 13426 19307 13429
rect 20253 13426 20319 13429
rect 19241 13424 20319 13426
rect 19241 13368 19246 13424
rect 19302 13368 20258 13424
rect 20314 13368 20319 13424
rect 19241 13366 20319 13368
rect 19241 13363 19307 13366
rect 20253 13363 20319 13366
rect 23520 13336 24000 13456
rect 4944 13088 5264 13089
rect 4944 13024 4952 13088
rect 5016 13024 5032 13088
rect 5096 13024 5112 13088
rect 5176 13024 5192 13088
rect 5256 13024 5264 13088
rect 4944 13023 5264 13024
rect 12944 13088 13264 13089
rect 12944 13024 12952 13088
rect 13016 13024 13032 13088
rect 13096 13024 13112 13088
rect 13176 13024 13192 13088
rect 13256 13024 13264 13088
rect 12944 13023 13264 13024
rect 20944 13088 21264 13089
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 13023 21264 13024
rect 21357 13018 21423 13021
rect 23614 13018 23674 13336
rect 21357 13016 23674 13018
rect 21357 12960 21362 13016
rect 21418 12960 23674 13016
rect 21357 12958 23674 12960
rect 21357 12955 21423 12958
rect 0 12792 480 12912
rect 62 12338 122 12792
rect 8944 12544 9264 12545
rect 8944 12480 8952 12544
rect 9016 12480 9032 12544
rect 9096 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9264 12544
rect 8944 12479 9264 12480
rect 16944 12544 17264 12545
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16944 12479 17264 12480
rect 19885 12474 19951 12477
rect 23520 12474 24000 12504
rect 19885 12472 24000 12474
rect 19885 12416 19890 12472
rect 19946 12416 24000 12472
rect 19885 12414 24000 12416
rect 19885 12411 19951 12414
rect 23520 12384 24000 12414
rect 1577 12338 1643 12341
rect 62 12336 1643 12338
rect 62 12280 1582 12336
rect 1638 12280 1643 12336
rect 62 12278 1643 12280
rect 1577 12275 1643 12278
rect 4944 12000 5264 12001
rect 4944 11936 4952 12000
rect 5016 11936 5032 12000
rect 5096 11936 5112 12000
rect 5176 11936 5192 12000
rect 5256 11936 5264 12000
rect 4944 11935 5264 11936
rect 12944 12000 13264 12001
rect 12944 11936 12952 12000
rect 13016 11936 13032 12000
rect 13096 11936 13112 12000
rect 13176 11936 13192 12000
rect 13256 11936 13264 12000
rect 12944 11935 13264 11936
rect 20944 12000 21264 12001
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 11935 21264 11936
rect 11881 11658 11947 11661
rect 20805 11658 20871 11661
rect 11881 11656 20871 11658
rect 11881 11600 11886 11656
rect 11942 11600 20810 11656
rect 20866 11600 20871 11656
rect 11881 11598 20871 11600
rect 11881 11595 11947 11598
rect 20805 11595 20871 11598
rect 8944 11456 9264 11457
rect 8944 11392 8952 11456
rect 9016 11392 9032 11456
rect 9096 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9264 11456
rect 8944 11391 9264 11392
rect 16944 11456 17264 11457
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 11391 17264 11392
rect 23520 11296 24000 11416
rect 0 11116 480 11144
rect 0 11052 60 11116
rect 124 11052 480 11116
rect 11973 11114 12039 11117
rect 16849 11114 16915 11117
rect 0 11024 480 11052
rect 1396 11112 16915 11114
rect 1396 11056 11978 11112
rect 12034 11056 16854 11112
rect 16910 11056 16915 11112
rect 1396 11054 16915 11056
rect 54 10780 60 10844
rect 124 10842 130 10844
rect 1396 10842 1456 11054
rect 11973 11051 12039 11054
rect 16849 11051 16915 11054
rect 4944 10912 5264 10913
rect 4944 10848 4952 10912
rect 5016 10848 5032 10912
rect 5096 10848 5112 10912
rect 5176 10848 5192 10912
rect 5256 10848 5264 10912
rect 4944 10847 5264 10848
rect 12944 10912 13264 10913
rect 12944 10848 12952 10912
rect 13016 10848 13032 10912
rect 13096 10848 13112 10912
rect 13176 10848 13192 10912
rect 13256 10848 13264 10912
rect 12944 10847 13264 10848
rect 20944 10912 21264 10913
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 10847 21264 10848
rect 124 10782 1456 10842
rect 21357 10842 21423 10845
rect 23614 10842 23674 11296
rect 21357 10840 23674 10842
rect 21357 10784 21362 10840
rect 21418 10784 23674 10840
rect 21357 10782 23674 10784
rect 124 10780 130 10782
rect 21357 10779 21423 10782
rect 10317 10570 10383 10573
rect 20897 10570 20963 10573
rect 10317 10568 20963 10570
rect 10317 10512 10322 10568
rect 10378 10512 20902 10568
rect 20958 10512 20963 10568
rect 10317 10510 20963 10512
rect 10317 10507 10383 10510
rect 20897 10507 20963 10510
rect 17861 10434 17927 10437
rect 23520 10434 24000 10464
rect 17861 10432 24000 10434
rect 17861 10376 17866 10432
rect 17922 10376 24000 10432
rect 17861 10374 24000 10376
rect 17861 10371 17927 10374
rect 8944 10368 9264 10369
rect 8944 10304 8952 10368
rect 9016 10304 9032 10368
rect 9096 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9264 10368
rect 8944 10303 9264 10304
rect 16944 10368 17264 10369
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 23520 10344 24000 10374
rect 16944 10303 17264 10304
rect 4944 9824 5264 9825
rect 4944 9760 4952 9824
rect 5016 9760 5032 9824
rect 5096 9760 5112 9824
rect 5176 9760 5192 9824
rect 5256 9760 5264 9824
rect 4944 9759 5264 9760
rect 12944 9824 13264 9825
rect 12944 9760 12952 9824
rect 13016 9760 13032 9824
rect 13096 9760 13112 9824
rect 13176 9760 13192 9824
rect 13256 9760 13264 9824
rect 12944 9759 13264 9760
rect 20944 9824 21264 9825
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 9759 21264 9760
rect 5717 9754 5783 9757
rect 9305 9754 9371 9757
rect 5717 9752 9371 9754
rect 5717 9696 5722 9752
rect 5778 9696 9310 9752
rect 9366 9696 9371 9752
rect 5717 9694 9371 9696
rect 5717 9691 5783 9694
rect 9305 9691 9371 9694
rect 1669 9618 1735 9621
rect 3509 9618 3575 9621
rect 4153 9618 4219 9621
rect 1669 9616 4219 9618
rect 1669 9560 1674 9616
rect 1730 9560 3514 9616
rect 3570 9560 4158 9616
rect 4214 9560 4219 9616
rect 1669 9558 4219 9560
rect 1669 9555 1735 9558
rect 3509 9555 3575 9558
rect 4153 9555 4219 9558
rect 9305 9618 9371 9621
rect 14825 9618 14891 9621
rect 9305 9616 14891 9618
rect 9305 9560 9310 9616
rect 9366 9560 14830 9616
rect 14886 9560 14891 9616
rect 9305 9558 14891 9560
rect 9305 9555 9371 9558
rect 14825 9555 14891 9558
rect 23520 9482 24000 9512
rect 23484 9480 24000 9482
rect 23484 9424 23570 9480
rect 23626 9424 24000 9480
rect 23484 9422 24000 9424
rect 23520 9392 24000 9422
rect 0 9348 480 9376
rect 0 9284 60 9348
rect 124 9284 480 9348
rect 0 9256 480 9284
rect 8944 9280 9264 9281
rect 8944 9216 8952 9280
rect 9016 9216 9032 9280
rect 9096 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9264 9280
rect 8944 9215 9264 9216
rect 16944 9280 17264 9281
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 9215 17264 9216
rect 54 9012 60 9076
rect 124 9074 130 9076
rect 1577 9074 1643 9077
rect 124 9072 1643 9074
rect 124 9016 1582 9072
rect 1638 9016 1643 9072
rect 124 9014 1643 9016
rect 124 9012 130 9014
rect 1577 9011 1643 9014
rect 7925 9074 7991 9077
rect 8845 9074 8911 9077
rect 15009 9074 15075 9077
rect 7925 9072 15075 9074
rect 7925 9016 7930 9072
rect 7986 9016 8850 9072
rect 8906 9016 15014 9072
rect 15070 9016 15075 9072
rect 7925 9014 15075 9016
rect 7925 9011 7991 9014
rect 8845 9011 8911 9014
rect 15009 9011 15075 9014
rect 105 8938 171 8941
rect 11237 8938 11303 8941
rect 105 8936 11303 8938
rect 105 8880 110 8936
rect 166 8880 11242 8936
rect 11298 8880 11303 8936
rect 105 8878 11303 8880
rect 105 8875 171 8878
rect 11237 8875 11303 8878
rect 4944 8736 5264 8737
rect 4944 8672 4952 8736
rect 5016 8672 5032 8736
rect 5096 8672 5112 8736
rect 5176 8672 5192 8736
rect 5256 8672 5264 8736
rect 4944 8671 5264 8672
rect 12944 8736 13264 8737
rect 12944 8672 12952 8736
rect 13016 8672 13032 8736
rect 13096 8672 13112 8736
rect 13176 8672 13192 8736
rect 13256 8672 13264 8736
rect 12944 8671 13264 8672
rect 20944 8736 21264 8737
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 8671 21264 8672
rect 4061 8530 4127 8533
rect 16573 8530 16639 8533
rect 4061 8528 16639 8530
rect 4061 8472 4066 8528
rect 4122 8472 16578 8528
rect 16634 8472 16639 8528
rect 4061 8470 16639 8472
rect 4061 8467 4127 8470
rect 16573 8467 16639 8470
rect 23520 8304 24000 8424
rect 8944 8192 9264 8193
rect 8944 8128 8952 8192
rect 9016 8128 9032 8192
rect 9096 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9264 8192
rect 8944 8127 9264 8128
rect 16944 8192 17264 8193
rect 16944 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17264 8192
rect 16944 8127 17264 8128
rect 7557 7986 7623 7989
rect 16205 7986 16271 7989
rect 16665 7986 16731 7989
rect 7557 7984 16731 7986
rect 7557 7928 7562 7984
rect 7618 7928 16210 7984
rect 16266 7928 16670 7984
rect 16726 7928 16731 7984
rect 7557 7926 16731 7928
rect 7557 7923 7623 7926
rect 16205 7923 16271 7926
rect 16665 7923 16731 7926
rect 21265 7850 21331 7853
rect 23614 7850 23674 8304
rect 21265 7848 23674 7850
rect 21265 7792 21270 7848
rect 21326 7792 23674 7848
rect 21265 7790 23674 7792
rect 21265 7787 21331 7790
rect 0 7624 480 7744
rect 4944 7648 5264 7649
rect 62 7170 122 7624
rect 4944 7584 4952 7648
rect 5016 7584 5032 7648
rect 5096 7584 5112 7648
rect 5176 7584 5192 7648
rect 5256 7584 5264 7648
rect 4944 7583 5264 7584
rect 12944 7648 13264 7649
rect 12944 7584 12952 7648
rect 13016 7584 13032 7648
rect 13096 7584 13112 7648
rect 13176 7584 13192 7648
rect 13256 7584 13264 7648
rect 12944 7583 13264 7584
rect 20944 7648 21264 7649
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 7583 21264 7584
rect 8845 7442 8911 7445
rect 14825 7442 14891 7445
rect 23520 7444 24000 7472
rect 23520 7442 23612 7444
rect 8845 7440 14891 7442
rect 8845 7384 8850 7440
rect 8906 7384 14830 7440
rect 14886 7384 14891 7440
rect 8845 7382 14891 7384
rect 23484 7382 23612 7442
rect 8845 7379 8911 7382
rect 14825 7379 14891 7382
rect 23520 7380 23612 7382
rect 23676 7380 24000 7444
rect 23520 7352 24000 7380
rect 13353 7306 13419 7309
rect 13997 7306 14063 7309
rect 13353 7304 19350 7306
rect 13353 7248 13358 7304
rect 13414 7248 14002 7304
rect 14058 7248 19350 7304
rect 13353 7246 19350 7248
rect 13353 7243 13419 7246
rect 13997 7243 14063 7246
rect 1577 7170 1643 7173
rect 62 7168 1643 7170
rect 62 7112 1582 7168
rect 1638 7112 1643 7168
rect 62 7110 1643 7112
rect 19290 7170 19350 7246
rect 23606 7170 23612 7172
rect 19290 7110 23612 7170
rect 1577 7107 1643 7110
rect 23606 7108 23612 7110
rect 23676 7108 23682 7172
rect 8944 7104 9264 7105
rect 8944 7040 8952 7104
rect 9016 7040 9032 7104
rect 9096 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9264 7104
rect 8944 7039 9264 7040
rect 16944 7104 17264 7105
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 7039 17264 7040
rect 4944 6560 5264 6561
rect 4944 6496 4952 6560
rect 5016 6496 5032 6560
rect 5096 6496 5112 6560
rect 5176 6496 5192 6560
rect 5256 6496 5264 6560
rect 4944 6495 5264 6496
rect 12944 6560 13264 6561
rect 12944 6496 12952 6560
rect 13016 6496 13032 6560
rect 13096 6496 13112 6560
rect 13176 6496 13192 6560
rect 13256 6496 13264 6560
rect 12944 6495 13264 6496
rect 20944 6560 21264 6561
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 6495 21264 6496
rect 21357 6490 21423 6493
rect 23520 6490 24000 6520
rect 21357 6488 24000 6490
rect 21357 6432 21362 6488
rect 21418 6432 24000 6488
rect 21357 6430 24000 6432
rect 21357 6427 21423 6430
rect 23520 6400 24000 6430
rect 2865 6218 2931 6221
rect 19149 6218 19215 6221
rect 2865 6216 19215 6218
rect 2865 6160 2870 6216
rect 2926 6160 19154 6216
rect 19210 6160 19215 6216
rect 2865 6158 19215 6160
rect 2865 6155 2931 6158
rect 19149 6155 19215 6158
rect 8944 6016 9264 6017
rect 0 5856 480 5976
rect 8944 5952 8952 6016
rect 9016 5952 9032 6016
rect 9096 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9264 6016
rect 8944 5951 9264 5952
rect 16944 6016 17264 6017
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 5951 17264 5952
rect 62 5402 122 5856
rect 4944 5472 5264 5473
rect 4944 5408 4952 5472
rect 5016 5408 5032 5472
rect 5096 5408 5112 5472
rect 5176 5408 5192 5472
rect 5256 5408 5264 5472
rect 4944 5407 5264 5408
rect 12944 5472 13264 5473
rect 12944 5408 12952 5472
rect 13016 5408 13032 5472
rect 13096 5408 13112 5472
rect 13176 5408 13192 5472
rect 13256 5408 13264 5472
rect 12944 5407 13264 5408
rect 20944 5472 21264 5473
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 5407 21264 5408
rect 1577 5402 1643 5405
rect 62 5400 1643 5402
rect 62 5344 1582 5400
rect 1638 5344 1643 5400
rect 62 5342 1643 5344
rect 1577 5339 1643 5342
rect 5625 5402 5691 5405
rect 7741 5402 7807 5405
rect 5625 5400 7807 5402
rect 5625 5344 5630 5400
rect 5686 5344 7746 5400
rect 7802 5344 7807 5400
rect 5625 5342 7807 5344
rect 5625 5339 5691 5342
rect 7741 5339 7807 5342
rect 21909 5402 21975 5405
rect 23520 5402 24000 5432
rect 21909 5400 24000 5402
rect 21909 5344 21914 5400
rect 21970 5344 24000 5400
rect 21909 5342 24000 5344
rect 21909 5339 21975 5342
rect 23520 5312 24000 5342
rect 6637 5266 6703 5269
rect 16389 5266 16455 5269
rect 6637 5264 16455 5266
rect 6637 5208 6642 5264
rect 6698 5208 16394 5264
rect 16450 5208 16455 5264
rect 6637 5206 16455 5208
rect 6637 5203 6703 5206
rect 16389 5203 16455 5206
rect 12617 5130 12683 5133
rect 21265 5130 21331 5133
rect 12617 5128 21331 5130
rect 12617 5072 12622 5128
rect 12678 5072 21270 5128
rect 21326 5072 21331 5128
rect 12617 5070 21331 5072
rect 12617 5067 12683 5070
rect 21265 5067 21331 5070
rect 21725 4994 21791 4997
rect 21725 4992 23674 4994
rect 21725 4936 21730 4992
rect 21786 4936 23674 4992
rect 21725 4934 23674 4936
rect 21725 4931 21791 4934
rect 8944 4928 9264 4929
rect 8944 4864 8952 4928
rect 9016 4864 9032 4928
rect 9096 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9264 4928
rect 8944 4863 9264 4864
rect 16944 4928 17264 4929
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 4863 17264 4864
rect 23614 4480 23674 4934
rect 4944 4384 5264 4385
rect 0 4316 480 4344
rect 4944 4320 4952 4384
rect 5016 4320 5032 4384
rect 5096 4320 5112 4384
rect 5176 4320 5192 4384
rect 5256 4320 5264 4384
rect 4944 4319 5264 4320
rect 12944 4384 13264 4385
rect 12944 4320 12952 4384
rect 13016 4320 13032 4384
rect 13096 4320 13112 4384
rect 13176 4320 13192 4384
rect 13256 4320 13264 4384
rect 12944 4319 13264 4320
rect 20944 4384 21264 4385
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 23520 4360 24000 4480
rect 20944 4319 21264 4320
rect 0 4252 60 4316
rect 124 4252 480 4316
rect 0 4224 480 4252
rect 15469 4178 15535 4181
rect 614 4176 15535 4178
rect 614 4120 15474 4176
rect 15530 4120 15535 4176
rect 614 4118 15535 4120
rect 54 3980 60 4044
rect 124 4042 130 4044
rect 614 4042 674 4118
rect 15469 4115 15535 4118
rect 124 3982 674 4042
rect 7925 4042 7991 4045
rect 23565 4042 23631 4045
rect 7925 4040 23631 4042
rect 7925 3984 7930 4040
rect 7986 3984 23570 4040
rect 23626 3984 23631 4040
rect 7925 3982 23631 3984
rect 124 3980 130 3982
rect 7925 3979 7991 3982
rect 23565 3979 23631 3982
rect 8944 3840 9264 3841
rect 8944 3776 8952 3840
rect 9016 3776 9032 3840
rect 9096 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9264 3840
rect 8944 3775 9264 3776
rect 16944 3840 17264 3841
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16944 3775 17264 3776
rect 12801 3634 12867 3637
rect 20805 3634 20871 3637
rect 12801 3632 20871 3634
rect 12801 3576 12806 3632
rect 12862 3576 20810 3632
rect 20866 3576 20871 3632
rect 12801 3574 20871 3576
rect 12801 3571 12867 3574
rect 20805 3571 20871 3574
rect 21449 3498 21515 3501
rect 23520 3498 24000 3528
rect 21449 3496 24000 3498
rect 21449 3440 21454 3496
rect 21510 3440 24000 3496
rect 21449 3438 24000 3440
rect 21449 3435 21515 3438
rect 23520 3408 24000 3438
rect 4944 3296 5264 3297
rect 4944 3232 4952 3296
rect 5016 3232 5032 3296
rect 5096 3232 5112 3296
rect 5176 3232 5192 3296
rect 5256 3232 5264 3296
rect 4944 3231 5264 3232
rect 12944 3296 13264 3297
rect 12944 3232 12952 3296
rect 13016 3232 13032 3296
rect 13096 3232 13112 3296
rect 13176 3232 13192 3296
rect 13256 3232 13264 3296
rect 12944 3231 13264 3232
rect 20944 3296 21264 3297
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 3231 21264 3232
rect 17309 2954 17375 2957
rect 17309 2952 23674 2954
rect 17309 2896 17314 2952
rect 17370 2896 23674 2952
rect 17309 2894 23674 2896
rect 17309 2891 17375 2894
rect 8944 2752 9264 2753
rect 8944 2688 8952 2752
rect 9016 2688 9032 2752
rect 9096 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9264 2752
rect 8944 2687 9264 2688
rect 16944 2752 17264 2753
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 16944 2687 17264 2688
rect 0 2544 480 2576
rect 0 2488 110 2544
rect 166 2488 480 2544
rect 0 2456 480 2488
rect 23614 2440 23674 2894
rect 23520 2320 24000 2440
rect 4944 2208 5264 2209
rect 4944 2144 4952 2208
rect 5016 2144 5032 2208
rect 5096 2144 5112 2208
rect 5176 2144 5192 2208
rect 5256 2144 5264 2208
rect 4944 2143 5264 2144
rect 12944 2208 13264 2209
rect 12944 2144 12952 2208
rect 13016 2144 13032 2208
rect 13096 2144 13112 2208
rect 13176 2144 13192 2208
rect 13256 2144 13264 2208
rect 12944 2143 13264 2144
rect 20944 2208 21264 2209
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2143 21264 2144
rect 7097 1866 7163 1869
rect 18965 1866 19031 1869
rect 7097 1864 19031 1866
rect 7097 1808 7102 1864
rect 7158 1808 18970 1864
rect 19026 1808 19031 1864
rect 7097 1806 19031 1808
rect 7097 1803 7163 1806
rect 18965 1803 19031 1806
rect 2037 1730 2103 1733
rect 21357 1730 21423 1733
rect 2037 1728 21423 1730
rect 2037 1672 2042 1728
rect 2098 1672 21362 1728
rect 21418 1672 21423 1728
rect 2037 1670 21423 1672
rect 2037 1667 2103 1670
rect 21357 1667 21423 1670
rect 1117 1458 1183 1461
rect 23520 1458 24000 1488
rect 62 1456 1183 1458
rect 62 1400 1122 1456
rect 1178 1400 1183 1456
rect 62 1398 1183 1400
rect 23484 1456 24000 1458
rect 23484 1400 23570 1456
rect 23626 1400 24000 1456
rect 23484 1398 24000 1400
rect 62 944 122 1398
rect 1117 1395 1183 1398
rect 23520 1368 24000 1398
rect 0 824 480 944
rect 23520 416 24000 536
rect 7557 98 7623 101
rect 23614 98 23674 416
rect 7557 96 23674 98
rect 7557 40 7562 96
rect 7618 40 23674 96
rect 7557 38 23674 40
rect 7557 35 7623 38
<< via3 >>
rect 4952 21788 5016 21792
rect 4952 21732 4956 21788
rect 4956 21732 5012 21788
rect 5012 21732 5016 21788
rect 4952 21728 5016 21732
rect 5032 21788 5096 21792
rect 5032 21732 5036 21788
rect 5036 21732 5092 21788
rect 5092 21732 5096 21788
rect 5032 21728 5096 21732
rect 5112 21788 5176 21792
rect 5112 21732 5116 21788
rect 5116 21732 5172 21788
rect 5172 21732 5176 21788
rect 5112 21728 5176 21732
rect 5192 21788 5256 21792
rect 5192 21732 5196 21788
rect 5196 21732 5252 21788
rect 5252 21732 5256 21788
rect 5192 21728 5256 21732
rect 12952 21788 13016 21792
rect 12952 21732 12956 21788
rect 12956 21732 13012 21788
rect 13012 21732 13016 21788
rect 12952 21728 13016 21732
rect 13032 21788 13096 21792
rect 13032 21732 13036 21788
rect 13036 21732 13092 21788
rect 13092 21732 13096 21788
rect 13032 21728 13096 21732
rect 13112 21788 13176 21792
rect 13112 21732 13116 21788
rect 13116 21732 13172 21788
rect 13172 21732 13176 21788
rect 13112 21728 13176 21732
rect 13192 21788 13256 21792
rect 13192 21732 13196 21788
rect 13196 21732 13252 21788
rect 13252 21732 13256 21788
rect 13192 21728 13256 21732
rect 20952 21788 21016 21792
rect 20952 21732 20956 21788
rect 20956 21732 21012 21788
rect 21012 21732 21016 21788
rect 20952 21728 21016 21732
rect 21032 21788 21096 21792
rect 21032 21732 21036 21788
rect 21036 21732 21092 21788
rect 21092 21732 21096 21788
rect 21032 21728 21096 21732
rect 21112 21788 21176 21792
rect 21112 21732 21116 21788
rect 21116 21732 21172 21788
rect 21172 21732 21176 21788
rect 21112 21728 21176 21732
rect 21192 21788 21256 21792
rect 21192 21732 21196 21788
rect 21196 21732 21252 21788
rect 21252 21732 21256 21788
rect 21192 21728 21256 21732
rect 8952 21244 9016 21248
rect 8952 21188 8956 21244
rect 8956 21188 9012 21244
rect 9012 21188 9016 21244
rect 8952 21184 9016 21188
rect 9032 21244 9096 21248
rect 9032 21188 9036 21244
rect 9036 21188 9092 21244
rect 9092 21188 9096 21244
rect 9032 21184 9096 21188
rect 9112 21244 9176 21248
rect 9112 21188 9116 21244
rect 9116 21188 9172 21244
rect 9172 21188 9176 21244
rect 9112 21184 9176 21188
rect 9192 21244 9256 21248
rect 9192 21188 9196 21244
rect 9196 21188 9252 21244
rect 9252 21188 9256 21244
rect 9192 21184 9256 21188
rect 16952 21244 17016 21248
rect 16952 21188 16956 21244
rect 16956 21188 17012 21244
rect 17012 21188 17016 21244
rect 16952 21184 17016 21188
rect 17032 21244 17096 21248
rect 17032 21188 17036 21244
rect 17036 21188 17092 21244
rect 17092 21188 17096 21244
rect 17032 21184 17096 21188
rect 17112 21244 17176 21248
rect 17112 21188 17116 21244
rect 17116 21188 17172 21244
rect 17172 21188 17176 21244
rect 17112 21184 17176 21188
rect 17192 21244 17256 21248
rect 17192 21188 17196 21244
rect 17196 21188 17252 21244
rect 17252 21188 17256 21244
rect 17192 21184 17256 21188
rect 4952 20700 5016 20704
rect 4952 20644 4956 20700
rect 4956 20644 5012 20700
rect 5012 20644 5016 20700
rect 4952 20640 5016 20644
rect 5032 20700 5096 20704
rect 5032 20644 5036 20700
rect 5036 20644 5092 20700
rect 5092 20644 5096 20700
rect 5032 20640 5096 20644
rect 5112 20700 5176 20704
rect 5112 20644 5116 20700
rect 5116 20644 5172 20700
rect 5172 20644 5176 20700
rect 5112 20640 5176 20644
rect 5192 20700 5256 20704
rect 5192 20644 5196 20700
rect 5196 20644 5252 20700
rect 5252 20644 5256 20700
rect 5192 20640 5256 20644
rect 12952 20700 13016 20704
rect 12952 20644 12956 20700
rect 12956 20644 13012 20700
rect 13012 20644 13016 20700
rect 12952 20640 13016 20644
rect 13032 20700 13096 20704
rect 13032 20644 13036 20700
rect 13036 20644 13092 20700
rect 13092 20644 13096 20700
rect 13032 20640 13096 20644
rect 13112 20700 13176 20704
rect 13112 20644 13116 20700
rect 13116 20644 13172 20700
rect 13172 20644 13176 20700
rect 13112 20640 13176 20644
rect 13192 20700 13256 20704
rect 13192 20644 13196 20700
rect 13196 20644 13252 20700
rect 13252 20644 13256 20700
rect 13192 20640 13256 20644
rect 20952 20700 21016 20704
rect 20952 20644 20956 20700
rect 20956 20644 21012 20700
rect 21012 20644 21016 20700
rect 20952 20640 21016 20644
rect 21032 20700 21096 20704
rect 21032 20644 21036 20700
rect 21036 20644 21092 20700
rect 21092 20644 21096 20700
rect 21032 20640 21096 20644
rect 21112 20700 21176 20704
rect 21112 20644 21116 20700
rect 21116 20644 21172 20700
rect 21172 20644 21176 20700
rect 21112 20640 21176 20644
rect 21192 20700 21256 20704
rect 21192 20644 21196 20700
rect 21196 20644 21252 20700
rect 21252 20644 21256 20700
rect 21192 20640 21256 20644
rect 8952 20156 9016 20160
rect 8952 20100 8956 20156
rect 8956 20100 9012 20156
rect 9012 20100 9016 20156
rect 8952 20096 9016 20100
rect 9032 20156 9096 20160
rect 9032 20100 9036 20156
rect 9036 20100 9092 20156
rect 9092 20100 9096 20156
rect 9032 20096 9096 20100
rect 9112 20156 9176 20160
rect 9112 20100 9116 20156
rect 9116 20100 9172 20156
rect 9172 20100 9176 20156
rect 9112 20096 9176 20100
rect 9192 20156 9256 20160
rect 9192 20100 9196 20156
rect 9196 20100 9252 20156
rect 9252 20100 9256 20156
rect 9192 20096 9256 20100
rect 16952 20156 17016 20160
rect 16952 20100 16956 20156
rect 16956 20100 17012 20156
rect 17012 20100 17016 20156
rect 16952 20096 17016 20100
rect 17032 20156 17096 20160
rect 17032 20100 17036 20156
rect 17036 20100 17092 20156
rect 17092 20100 17096 20156
rect 17032 20096 17096 20100
rect 17112 20156 17176 20160
rect 17112 20100 17116 20156
rect 17116 20100 17172 20156
rect 17172 20100 17176 20156
rect 17112 20096 17176 20100
rect 17192 20156 17256 20160
rect 17192 20100 17196 20156
rect 17196 20100 17252 20156
rect 17252 20100 17256 20156
rect 17192 20096 17256 20100
rect 4952 19612 5016 19616
rect 4952 19556 4956 19612
rect 4956 19556 5012 19612
rect 5012 19556 5016 19612
rect 4952 19552 5016 19556
rect 5032 19612 5096 19616
rect 5032 19556 5036 19612
rect 5036 19556 5092 19612
rect 5092 19556 5096 19612
rect 5032 19552 5096 19556
rect 5112 19612 5176 19616
rect 5112 19556 5116 19612
rect 5116 19556 5172 19612
rect 5172 19556 5176 19612
rect 5112 19552 5176 19556
rect 5192 19612 5256 19616
rect 5192 19556 5196 19612
rect 5196 19556 5252 19612
rect 5252 19556 5256 19612
rect 5192 19552 5256 19556
rect 12952 19612 13016 19616
rect 12952 19556 12956 19612
rect 12956 19556 13012 19612
rect 13012 19556 13016 19612
rect 12952 19552 13016 19556
rect 13032 19612 13096 19616
rect 13032 19556 13036 19612
rect 13036 19556 13092 19612
rect 13092 19556 13096 19612
rect 13032 19552 13096 19556
rect 13112 19612 13176 19616
rect 13112 19556 13116 19612
rect 13116 19556 13172 19612
rect 13172 19556 13176 19612
rect 13112 19552 13176 19556
rect 13192 19612 13256 19616
rect 13192 19556 13196 19612
rect 13196 19556 13252 19612
rect 13252 19556 13256 19612
rect 13192 19552 13256 19556
rect 20952 19612 21016 19616
rect 20952 19556 20956 19612
rect 20956 19556 21012 19612
rect 21012 19556 21016 19612
rect 20952 19552 21016 19556
rect 21032 19612 21096 19616
rect 21032 19556 21036 19612
rect 21036 19556 21092 19612
rect 21092 19556 21096 19612
rect 21032 19552 21096 19556
rect 21112 19612 21176 19616
rect 21112 19556 21116 19612
rect 21116 19556 21172 19612
rect 21172 19556 21176 19612
rect 21112 19552 21176 19556
rect 21192 19612 21256 19616
rect 21192 19556 21196 19612
rect 21196 19556 21252 19612
rect 21252 19556 21256 19612
rect 21192 19552 21256 19556
rect 8952 19068 9016 19072
rect 8952 19012 8956 19068
rect 8956 19012 9012 19068
rect 9012 19012 9016 19068
rect 8952 19008 9016 19012
rect 9032 19068 9096 19072
rect 9032 19012 9036 19068
rect 9036 19012 9092 19068
rect 9092 19012 9096 19068
rect 9032 19008 9096 19012
rect 9112 19068 9176 19072
rect 9112 19012 9116 19068
rect 9116 19012 9172 19068
rect 9172 19012 9176 19068
rect 9112 19008 9176 19012
rect 9192 19068 9256 19072
rect 9192 19012 9196 19068
rect 9196 19012 9252 19068
rect 9252 19012 9256 19068
rect 9192 19008 9256 19012
rect 16952 19068 17016 19072
rect 16952 19012 16956 19068
rect 16956 19012 17012 19068
rect 17012 19012 17016 19068
rect 16952 19008 17016 19012
rect 17032 19068 17096 19072
rect 17032 19012 17036 19068
rect 17036 19012 17092 19068
rect 17092 19012 17096 19068
rect 17032 19008 17096 19012
rect 17112 19068 17176 19072
rect 17112 19012 17116 19068
rect 17116 19012 17172 19068
rect 17172 19012 17176 19068
rect 17112 19008 17176 19012
rect 17192 19068 17256 19072
rect 17192 19012 17196 19068
rect 17196 19012 17252 19068
rect 17252 19012 17256 19068
rect 17192 19008 17256 19012
rect 4952 18524 5016 18528
rect 4952 18468 4956 18524
rect 4956 18468 5012 18524
rect 5012 18468 5016 18524
rect 4952 18464 5016 18468
rect 5032 18524 5096 18528
rect 5032 18468 5036 18524
rect 5036 18468 5092 18524
rect 5092 18468 5096 18524
rect 5032 18464 5096 18468
rect 5112 18524 5176 18528
rect 5112 18468 5116 18524
rect 5116 18468 5172 18524
rect 5172 18468 5176 18524
rect 5112 18464 5176 18468
rect 5192 18524 5256 18528
rect 5192 18468 5196 18524
rect 5196 18468 5252 18524
rect 5252 18468 5256 18524
rect 5192 18464 5256 18468
rect 12952 18524 13016 18528
rect 12952 18468 12956 18524
rect 12956 18468 13012 18524
rect 13012 18468 13016 18524
rect 12952 18464 13016 18468
rect 13032 18524 13096 18528
rect 13032 18468 13036 18524
rect 13036 18468 13092 18524
rect 13092 18468 13096 18524
rect 13032 18464 13096 18468
rect 13112 18524 13176 18528
rect 13112 18468 13116 18524
rect 13116 18468 13172 18524
rect 13172 18468 13176 18524
rect 13112 18464 13176 18468
rect 13192 18524 13256 18528
rect 13192 18468 13196 18524
rect 13196 18468 13252 18524
rect 13252 18468 13256 18524
rect 13192 18464 13256 18468
rect 20952 18524 21016 18528
rect 20952 18468 20956 18524
rect 20956 18468 21012 18524
rect 21012 18468 21016 18524
rect 20952 18464 21016 18468
rect 21032 18524 21096 18528
rect 21032 18468 21036 18524
rect 21036 18468 21092 18524
rect 21092 18468 21096 18524
rect 21032 18464 21096 18468
rect 21112 18524 21176 18528
rect 21112 18468 21116 18524
rect 21116 18468 21172 18524
rect 21172 18468 21176 18524
rect 21112 18464 21176 18468
rect 21192 18524 21256 18528
rect 21192 18468 21196 18524
rect 21196 18468 21252 18524
rect 21252 18468 21256 18524
rect 21192 18464 21256 18468
rect 8952 17980 9016 17984
rect 8952 17924 8956 17980
rect 8956 17924 9012 17980
rect 9012 17924 9016 17980
rect 8952 17920 9016 17924
rect 9032 17980 9096 17984
rect 9032 17924 9036 17980
rect 9036 17924 9092 17980
rect 9092 17924 9096 17980
rect 9032 17920 9096 17924
rect 9112 17980 9176 17984
rect 9112 17924 9116 17980
rect 9116 17924 9172 17980
rect 9172 17924 9176 17980
rect 9112 17920 9176 17924
rect 9192 17980 9256 17984
rect 9192 17924 9196 17980
rect 9196 17924 9252 17980
rect 9252 17924 9256 17980
rect 9192 17920 9256 17924
rect 16952 17980 17016 17984
rect 16952 17924 16956 17980
rect 16956 17924 17012 17980
rect 17012 17924 17016 17980
rect 16952 17920 17016 17924
rect 17032 17980 17096 17984
rect 17032 17924 17036 17980
rect 17036 17924 17092 17980
rect 17092 17924 17096 17980
rect 17032 17920 17096 17924
rect 17112 17980 17176 17984
rect 17112 17924 17116 17980
rect 17116 17924 17172 17980
rect 17172 17924 17176 17980
rect 17112 17920 17176 17924
rect 17192 17980 17256 17984
rect 17192 17924 17196 17980
rect 17196 17924 17252 17980
rect 17252 17924 17256 17980
rect 17192 17920 17256 17924
rect 4952 17436 5016 17440
rect 4952 17380 4956 17436
rect 4956 17380 5012 17436
rect 5012 17380 5016 17436
rect 4952 17376 5016 17380
rect 5032 17436 5096 17440
rect 5032 17380 5036 17436
rect 5036 17380 5092 17436
rect 5092 17380 5096 17436
rect 5032 17376 5096 17380
rect 5112 17436 5176 17440
rect 5112 17380 5116 17436
rect 5116 17380 5172 17436
rect 5172 17380 5176 17436
rect 5112 17376 5176 17380
rect 5192 17436 5256 17440
rect 5192 17380 5196 17436
rect 5196 17380 5252 17436
rect 5252 17380 5256 17436
rect 5192 17376 5256 17380
rect 12952 17436 13016 17440
rect 12952 17380 12956 17436
rect 12956 17380 13012 17436
rect 13012 17380 13016 17436
rect 12952 17376 13016 17380
rect 13032 17436 13096 17440
rect 13032 17380 13036 17436
rect 13036 17380 13092 17436
rect 13092 17380 13096 17436
rect 13032 17376 13096 17380
rect 13112 17436 13176 17440
rect 13112 17380 13116 17436
rect 13116 17380 13172 17436
rect 13172 17380 13176 17436
rect 13112 17376 13176 17380
rect 13192 17436 13256 17440
rect 13192 17380 13196 17436
rect 13196 17380 13252 17436
rect 13252 17380 13256 17436
rect 13192 17376 13256 17380
rect 20952 17436 21016 17440
rect 20952 17380 20956 17436
rect 20956 17380 21012 17436
rect 21012 17380 21016 17436
rect 20952 17376 21016 17380
rect 21032 17436 21096 17440
rect 21032 17380 21036 17436
rect 21036 17380 21092 17436
rect 21092 17380 21096 17436
rect 21032 17376 21096 17380
rect 21112 17436 21176 17440
rect 21112 17380 21116 17436
rect 21116 17380 21172 17436
rect 21172 17380 21176 17436
rect 21112 17376 21176 17380
rect 21192 17436 21256 17440
rect 21192 17380 21196 17436
rect 21196 17380 21252 17436
rect 21252 17380 21256 17436
rect 21192 17376 21256 17380
rect 8952 16892 9016 16896
rect 8952 16836 8956 16892
rect 8956 16836 9012 16892
rect 9012 16836 9016 16892
rect 8952 16832 9016 16836
rect 9032 16892 9096 16896
rect 9032 16836 9036 16892
rect 9036 16836 9092 16892
rect 9092 16836 9096 16892
rect 9032 16832 9096 16836
rect 9112 16892 9176 16896
rect 9112 16836 9116 16892
rect 9116 16836 9172 16892
rect 9172 16836 9176 16892
rect 9112 16832 9176 16836
rect 9192 16892 9256 16896
rect 9192 16836 9196 16892
rect 9196 16836 9252 16892
rect 9252 16836 9256 16892
rect 9192 16832 9256 16836
rect 16952 16892 17016 16896
rect 16952 16836 16956 16892
rect 16956 16836 17012 16892
rect 17012 16836 17016 16892
rect 16952 16832 17016 16836
rect 17032 16892 17096 16896
rect 17032 16836 17036 16892
rect 17036 16836 17092 16892
rect 17092 16836 17096 16892
rect 17032 16832 17096 16836
rect 17112 16892 17176 16896
rect 17112 16836 17116 16892
rect 17116 16836 17172 16892
rect 17172 16836 17176 16892
rect 17112 16832 17176 16836
rect 17192 16892 17256 16896
rect 17192 16836 17196 16892
rect 17196 16836 17252 16892
rect 17252 16836 17256 16892
rect 17192 16832 17256 16836
rect 4952 16348 5016 16352
rect 4952 16292 4956 16348
rect 4956 16292 5012 16348
rect 5012 16292 5016 16348
rect 4952 16288 5016 16292
rect 5032 16348 5096 16352
rect 5032 16292 5036 16348
rect 5036 16292 5092 16348
rect 5092 16292 5096 16348
rect 5032 16288 5096 16292
rect 5112 16348 5176 16352
rect 5112 16292 5116 16348
rect 5116 16292 5172 16348
rect 5172 16292 5176 16348
rect 5112 16288 5176 16292
rect 5192 16348 5256 16352
rect 5192 16292 5196 16348
rect 5196 16292 5252 16348
rect 5252 16292 5256 16348
rect 5192 16288 5256 16292
rect 12952 16348 13016 16352
rect 12952 16292 12956 16348
rect 12956 16292 13012 16348
rect 13012 16292 13016 16348
rect 12952 16288 13016 16292
rect 13032 16348 13096 16352
rect 13032 16292 13036 16348
rect 13036 16292 13092 16348
rect 13092 16292 13096 16348
rect 13032 16288 13096 16292
rect 13112 16348 13176 16352
rect 13112 16292 13116 16348
rect 13116 16292 13172 16348
rect 13172 16292 13176 16348
rect 13112 16288 13176 16292
rect 13192 16348 13256 16352
rect 13192 16292 13196 16348
rect 13196 16292 13252 16348
rect 13252 16292 13256 16348
rect 13192 16288 13256 16292
rect 20952 16348 21016 16352
rect 20952 16292 20956 16348
rect 20956 16292 21012 16348
rect 21012 16292 21016 16348
rect 20952 16288 21016 16292
rect 21032 16348 21096 16352
rect 21032 16292 21036 16348
rect 21036 16292 21092 16348
rect 21092 16292 21096 16348
rect 21032 16288 21096 16292
rect 21112 16348 21176 16352
rect 21112 16292 21116 16348
rect 21116 16292 21172 16348
rect 21172 16292 21176 16348
rect 21112 16288 21176 16292
rect 21192 16348 21256 16352
rect 21192 16292 21196 16348
rect 21196 16292 21252 16348
rect 21252 16292 21256 16348
rect 21192 16288 21256 16292
rect 8952 15804 9016 15808
rect 8952 15748 8956 15804
rect 8956 15748 9012 15804
rect 9012 15748 9016 15804
rect 8952 15744 9016 15748
rect 9032 15804 9096 15808
rect 9032 15748 9036 15804
rect 9036 15748 9092 15804
rect 9092 15748 9096 15804
rect 9032 15744 9096 15748
rect 9112 15804 9176 15808
rect 9112 15748 9116 15804
rect 9116 15748 9172 15804
rect 9172 15748 9176 15804
rect 9112 15744 9176 15748
rect 9192 15804 9256 15808
rect 9192 15748 9196 15804
rect 9196 15748 9252 15804
rect 9252 15748 9256 15804
rect 9192 15744 9256 15748
rect 16952 15804 17016 15808
rect 16952 15748 16956 15804
rect 16956 15748 17012 15804
rect 17012 15748 17016 15804
rect 16952 15744 17016 15748
rect 17032 15804 17096 15808
rect 17032 15748 17036 15804
rect 17036 15748 17092 15804
rect 17092 15748 17096 15804
rect 17032 15744 17096 15748
rect 17112 15804 17176 15808
rect 17112 15748 17116 15804
rect 17116 15748 17172 15804
rect 17172 15748 17176 15804
rect 17112 15744 17176 15748
rect 17192 15804 17256 15808
rect 17192 15748 17196 15804
rect 17196 15748 17252 15804
rect 17252 15748 17256 15804
rect 17192 15744 17256 15748
rect 23612 15676 23676 15740
rect 23612 15404 23676 15468
rect 4952 15260 5016 15264
rect 4952 15204 4956 15260
rect 4956 15204 5012 15260
rect 5012 15204 5016 15260
rect 4952 15200 5016 15204
rect 5032 15260 5096 15264
rect 5032 15204 5036 15260
rect 5036 15204 5092 15260
rect 5092 15204 5096 15260
rect 5032 15200 5096 15204
rect 5112 15260 5176 15264
rect 5112 15204 5116 15260
rect 5116 15204 5172 15260
rect 5172 15204 5176 15260
rect 5112 15200 5176 15204
rect 5192 15260 5256 15264
rect 5192 15204 5196 15260
rect 5196 15204 5252 15260
rect 5252 15204 5256 15260
rect 5192 15200 5256 15204
rect 12952 15260 13016 15264
rect 12952 15204 12956 15260
rect 12956 15204 13012 15260
rect 13012 15204 13016 15260
rect 12952 15200 13016 15204
rect 13032 15260 13096 15264
rect 13032 15204 13036 15260
rect 13036 15204 13092 15260
rect 13092 15204 13096 15260
rect 13032 15200 13096 15204
rect 13112 15260 13176 15264
rect 13112 15204 13116 15260
rect 13116 15204 13172 15260
rect 13172 15204 13176 15260
rect 13112 15200 13176 15204
rect 13192 15260 13256 15264
rect 13192 15204 13196 15260
rect 13196 15204 13252 15260
rect 13252 15204 13256 15260
rect 13192 15200 13256 15204
rect 20952 15260 21016 15264
rect 20952 15204 20956 15260
rect 20956 15204 21012 15260
rect 21012 15204 21016 15260
rect 20952 15200 21016 15204
rect 21032 15260 21096 15264
rect 21032 15204 21036 15260
rect 21036 15204 21092 15260
rect 21092 15204 21096 15260
rect 21032 15200 21096 15204
rect 21112 15260 21176 15264
rect 21112 15204 21116 15260
rect 21116 15204 21172 15260
rect 21172 15204 21176 15260
rect 21112 15200 21176 15204
rect 21192 15260 21256 15264
rect 21192 15204 21196 15260
rect 21196 15204 21252 15260
rect 21252 15204 21256 15260
rect 21192 15200 21256 15204
rect 8952 14716 9016 14720
rect 8952 14660 8956 14716
rect 8956 14660 9012 14716
rect 9012 14660 9016 14716
rect 8952 14656 9016 14660
rect 9032 14716 9096 14720
rect 9032 14660 9036 14716
rect 9036 14660 9092 14716
rect 9092 14660 9096 14716
rect 9032 14656 9096 14660
rect 9112 14716 9176 14720
rect 9112 14660 9116 14716
rect 9116 14660 9172 14716
rect 9172 14660 9176 14716
rect 9112 14656 9176 14660
rect 9192 14716 9256 14720
rect 9192 14660 9196 14716
rect 9196 14660 9252 14716
rect 9252 14660 9256 14716
rect 9192 14656 9256 14660
rect 16952 14716 17016 14720
rect 16952 14660 16956 14716
rect 16956 14660 17012 14716
rect 17012 14660 17016 14716
rect 16952 14656 17016 14660
rect 17032 14716 17096 14720
rect 17032 14660 17036 14716
rect 17036 14660 17092 14716
rect 17092 14660 17096 14716
rect 17032 14656 17096 14660
rect 17112 14716 17176 14720
rect 17112 14660 17116 14716
rect 17116 14660 17172 14716
rect 17172 14660 17176 14716
rect 17112 14656 17176 14660
rect 17192 14716 17256 14720
rect 17192 14660 17196 14716
rect 17196 14660 17252 14716
rect 17252 14660 17256 14716
rect 17192 14656 17256 14660
rect 4952 14172 5016 14176
rect 4952 14116 4956 14172
rect 4956 14116 5012 14172
rect 5012 14116 5016 14172
rect 4952 14112 5016 14116
rect 5032 14172 5096 14176
rect 5032 14116 5036 14172
rect 5036 14116 5092 14172
rect 5092 14116 5096 14172
rect 5032 14112 5096 14116
rect 5112 14172 5176 14176
rect 5112 14116 5116 14172
rect 5116 14116 5172 14172
rect 5172 14116 5176 14172
rect 5112 14112 5176 14116
rect 5192 14172 5256 14176
rect 5192 14116 5196 14172
rect 5196 14116 5252 14172
rect 5252 14116 5256 14172
rect 5192 14112 5256 14116
rect 12952 14172 13016 14176
rect 12952 14116 12956 14172
rect 12956 14116 13012 14172
rect 13012 14116 13016 14172
rect 12952 14112 13016 14116
rect 13032 14172 13096 14176
rect 13032 14116 13036 14172
rect 13036 14116 13092 14172
rect 13092 14116 13096 14172
rect 13032 14112 13096 14116
rect 13112 14172 13176 14176
rect 13112 14116 13116 14172
rect 13116 14116 13172 14172
rect 13172 14116 13176 14172
rect 13112 14112 13176 14116
rect 13192 14172 13256 14176
rect 13192 14116 13196 14172
rect 13196 14116 13252 14172
rect 13252 14116 13256 14172
rect 13192 14112 13256 14116
rect 20952 14172 21016 14176
rect 20952 14116 20956 14172
rect 20956 14116 21012 14172
rect 21012 14116 21016 14172
rect 20952 14112 21016 14116
rect 21032 14172 21096 14176
rect 21032 14116 21036 14172
rect 21036 14116 21092 14172
rect 21092 14116 21096 14172
rect 21032 14112 21096 14116
rect 21112 14172 21176 14176
rect 21112 14116 21116 14172
rect 21116 14116 21172 14172
rect 21172 14116 21176 14172
rect 21112 14112 21176 14116
rect 21192 14172 21256 14176
rect 21192 14116 21196 14172
rect 21196 14116 21252 14172
rect 21252 14116 21256 14172
rect 21192 14112 21256 14116
rect 8952 13628 9016 13632
rect 8952 13572 8956 13628
rect 8956 13572 9012 13628
rect 9012 13572 9016 13628
rect 8952 13568 9016 13572
rect 9032 13628 9096 13632
rect 9032 13572 9036 13628
rect 9036 13572 9092 13628
rect 9092 13572 9096 13628
rect 9032 13568 9096 13572
rect 9112 13628 9176 13632
rect 9112 13572 9116 13628
rect 9116 13572 9172 13628
rect 9172 13572 9176 13628
rect 9112 13568 9176 13572
rect 9192 13628 9256 13632
rect 9192 13572 9196 13628
rect 9196 13572 9252 13628
rect 9252 13572 9256 13628
rect 9192 13568 9256 13572
rect 16952 13628 17016 13632
rect 16952 13572 16956 13628
rect 16956 13572 17012 13628
rect 17012 13572 17016 13628
rect 16952 13568 17016 13572
rect 17032 13628 17096 13632
rect 17032 13572 17036 13628
rect 17036 13572 17092 13628
rect 17092 13572 17096 13628
rect 17032 13568 17096 13572
rect 17112 13628 17176 13632
rect 17112 13572 17116 13628
rect 17116 13572 17172 13628
rect 17172 13572 17176 13628
rect 17112 13568 17176 13572
rect 17192 13628 17256 13632
rect 17192 13572 17196 13628
rect 17196 13572 17252 13628
rect 17252 13572 17256 13628
rect 17192 13568 17256 13572
rect 4952 13084 5016 13088
rect 4952 13028 4956 13084
rect 4956 13028 5012 13084
rect 5012 13028 5016 13084
rect 4952 13024 5016 13028
rect 5032 13084 5096 13088
rect 5032 13028 5036 13084
rect 5036 13028 5092 13084
rect 5092 13028 5096 13084
rect 5032 13024 5096 13028
rect 5112 13084 5176 13088
rect 5112 13028 5116 13084
rect 5116 13028 5172 13084
rect 5172 13028 5176 13084
rect 5112 13024 5176 13028
rect 5192 13084 5256 13088
rect 5192 13028 5196 13084
rect 5196 13028 5252 13084
rect 5252 13028 5256 13084
rect 5192 13024 5256 13028
rect 12952 13084 13016 13088
rect 12952 13028 12956 13084
rect 12956 13028 13012 13084
rect 13012 13028 13016 13084
rect 12952 13024 13016 13028
rect 13032 13084 13096 13088
rect 13032 13028 13036 13084
rect 13036 13028 13092 13084
rect 13092 13028 13096 13084
rect 13032 13024 13096 13028
rect 13112 13084 13176 13088
rect 13112 13028 13116 13084
rect 13116 13028 13172 13084
rect 13172 13028 13176 13084
rect 13112 13024 13176 13028
rect 13192 13084 13256 13088
rect 13192 13028 13196 13084
rect 13196 13028 13252 13084
rect 13252 13028 13256 13084
rect 13192 13024 13256 13028
rect 20952 13084 21016 13088
rect 20952 13028 20956 13084
rect 20956 13028 21012 13084
rect 21012 13028 21016 13084
rect 20952 13024 21016 13028
rect 21032 13084 21096 13088
rect 21032 13028 21036 13084
rect 21036 13028 21092 13084
rect 21092 13028 21096 13084
rect 21032 13024 21096 13028
rect 21112 13084 21176 13088
rect 21112 13028 21116 13084
rect 21116 13028 21172 13084
rect 21172 13028 21176 13084
rect 21112 13024 21176 13028
rect 21192 13084 21256 13088
rect 21192 13028 21196 13084
rect 21196 13028 21252 13084
rect 21252 13028 21256 13084
rect 21192 13024 21256 13028
rect 8952 12540 9016 12544
rect 8952 12484 8956 12540
rect 8956 12484 9012 12540
rect 9012 12484 9016 12540
rect 8952 12480 9016 12484
rect 9032 12540 9096 12544
rect 9032 12484 9036 12540
rect 9036 12484 9092 12540
rect 9092 12484 9096 12540
rect 9032 12480 9096 12484
rect 9112 12540 9176 12544
rect 9112 12484 9116 12540
rect 9116 12484 9172 12540
rect 9172 12484 9176 12540
rect 9112 12480 9176 12484
rect 9192 12540 9256 12544
rect 9192 12484 9196 12540
rect 9196 12484 9252 12540
rect 9252 12484 9256 12540
rect 9192 12480 9256 12484
rect 16952 12540 17016 12544
rect 16952 12484 16956 12540
rect 16956 12484 17012 12540
rect 17012 12484 17016 12540
rect 16952 12480 17016 12484
rect 17032 12540 17096 12544
rect 17032 12484 17036 12540
rect 17036 12484 17092 12540
rect 17092 12484 17096 12540
rect 17032 12480 17096 12484
rect 17112 12540 17176 12544
rect 17112 12484 17116 12540
rect 17116 12484 17172 12540
rect 17172 12484 17176 12540
rect 17112 12480 17176 12484
rect 17192 12540 17256 12544
rect 17192 12484 17196 12540
rect 17196 12484 17252 12540
rect 17252 12484 17256 12540
rect 17192 12480 17256 12484
rect 4952 11996 5016 12000
rect 4952 11940 4956 11996
rect 4956 11940 5012 11996
rect 5012 11940 5016 11996
rect 4952 11936 5016 11940
rect 5032 11996 5096 12000
rect 5032 11940 5036 11996
rect 5036 11940 5092 11996
rect 5092 11940 5096 11996
rect 5032 11936 5096 11940
rect 5112 11996 5176 12000
rect 5112 11940 5116 11996
rect 5116 11940 5172 11996
rect 5172 11940 5176 11996
rect 5112 11936 5176 11940
rect 5192 11996 5256 12000
rect 5192 11940 5196 11996
rect 5196 11940 5252 11996
rect 5252 11940 5256 11996
rect 5192 11936 5256 11940
rect 12952 11996 13016 12000
rect 12952 11940 12956 11996
rect 12956 11940 13012 11996
rect 13012 11940 13016 11996
rect 12952 11936 13016 11940
rect 13032 11996 13096 12000
rect 13032 11940 13036 11996
rect 13036 11940 13092 11996
rect 13092 11940 13096 11996
rect 13032 11936 13096 11940
rect 13112 11996 13176 12000
rect 13112 11940 13116 11996
rect 13116 11940 13172 11996
rect 13172 11940 13176 11996
rect 13112 11936 13176 11940
rect 13192 11996 13256 12000
rect 13192 11940 13196 11996
rect 13196 11940 13252 11996
rect 13252 11940 13256 11996
rect 13192 11936 13256 11940
rect 20952 11996 21016 12000
rect 20952 11940 20956 11996
rect 20956 11940 21012 11996
rect 21012 11940 21016 11996
rect 20952 11936 21016 11940
rect 21032 11996 21096 12000
rect 21032 11940 21036 11996
rect 21036 11940 21092 11996
rect 21092 11940 21096 11996
rect 21032 11936 21096 11940
rect 21112 11996 21176 12000
rect 21112 11940 21116 11996
rect 21116 11940 21172 11996
rect 21172 11940 21176 11996
rect 21112 11936 21176 11940
rect 21192 11996 21256 12000
rect 21192 11940 21196 11996
rect 21196 11940 21252 11996
rect 21252 11940 21256 11996
rect 21192 11936 21256 11940
rect 8952 11452 9016 11456
rect 8952 11396 8956 11452
rect 8956 11396 9012 11452
rect 9012 11396 9016 11452
rect 8952 11392 9016 11396
rect 9032 11452 9096 11456
rect 9032 11396 9036 11452
rect 9036 11396 9092 11452
rect 9092 11396 9096 11452
rect 9032 11392 9096 11396
rect 9112 11452 9176 11456
rect 9112 11396 9116 11452
rect 9116 11396 9172 11452
rect 9172 11396 9176 11452
rect 9112 11392 9176 11396
rect 9192 11452 9256 11456
rect 9192 11396 9196 11452
rect 9196 11396 9252 11452
rect 9252 11396 9256 11452
rect 9192 11392 9256 11396
rect 16952 11452 17016 11456
rect 16952 11396 16956 11452
rect 16956 11396 17012 11452
rect 17012 11396 17016 11452
rect 16952 11392 17016 11396
rect 17032 11452 17096 11456
rect 17032 11396 17036 11452
rect 17036 11396 17092 11452
rect 17092 11396 17096 11452
rect 17032 11392 17096 11396
rect 17112 11452 17176 11456
rect 17112 11396 17116 11452
rect 17116 11396 17172 11452
rect 17172 11396 17176 11452
rect 17112 11392 17176 11396
rect 17192 11452 17256 11456
rect 17192 11396 17196 11452
rect 17196 11396 17252 11452
rect 17252 11396 17256 11452
rect 17192 11392 17256 11396
rect 60 11052 124 11116
rect 60 10780 124 10844
rect 4952 10908 5016 10912
rect 4952 10852 4956 10908
rect 4956 10852 5012 10908
rect 5012 10852 5016 10908
rect 4952 10848 5016 10852
rect 5032 10908 5096 10912
rect 5032 10852 5036 10908
rect 5036 10852 5092 10908
rect 5092 10852 5096 10908
rect 5032 10848 5096 10852
rect 5112 10908 5176 10912
rect 5112 10852 5116 10908
rect 5116 10852 5172 10908
rect 5172 10852 5176 10908
rect 5112 10848 5176 10852
rect 5192 10908 5256 10912
rect 5192 10852 5196 10908
rect 5196 10852 5252 10908
rect 5252 10852 5256 10908
rect 5192 10848 5256 10852
rect 12952 10908 13016 10912
rect 12952 10852 12956 10908
rect 12956 10852 13012 10908
rect 13012 10852 13016 10908
rect 12952 10848 13016 10852
rect 13032 10908 13096 10912
rect 13032 10852 13036 10908
rect 13036 10852 13092 10908
rect 13092 10852 13096 10908
rect 13032 10848 13096 10852
rect 13112 10908 13176 10912
rect 13112 10852 13116 10908
rect 13116 10852 13172 10908
rect 13172 10852 13176 10908
rect 13112 10848 13176 10852
rect 13192 10908 13256 10912
rect 13192 10852 13196 10908
rect 13196 10852 13252 10908
rect 13252 10852 13256 10908
rect 13192 10848 13256 10852
rect 20952 10908 21016 10912
rect 20952 10852 20956 10908
rect 20956 10852 21012 10908
rect 21012 10852 21016 10908
rect 20952 10848 21016 10852
rect 21032 10908 21096 10912
rect 21032 10852 21036 10908
rect 21036 10852 21092 10908
rect 21092 10852 21096 10908
rect 21032 10848 21096 10852
rect 21112 10908 21176 10912
rect 21112 10852 21116 10908
rect 21116 10852 21172 10908
rect 21172 10852 21176 10908
rect 21112 10848 21176 10852
rect 21192 10908 21256 10912
rect 21192 10852 21196 10908
rect 21196 10852 21252 10908
rect 21252 10852 21256 10908
rect 21192 10848 21256 10852
rect 8952 10364 9016 10368
rect 8952 10308 8956 10364
rect 8956 10308 9012 10364
rect 9012 10308 9016 10364
rect 8952 10304 9016 10308
rect 9032 10364 9096 10368
rect 9032 10308 9036 10364
rect 9036 10308 9092 10364
rect 9092 10308 9096 10364
rect 9032 10304 9096 10308
rect 9112 10364 9176 10368
rect 9112 10308 9116 10364
rect 9116 10308 9172 10364
rect 9172 10308 9176 10364
rect 9112 10304 9176 10308
rect 9192 10364 9256 10368
rect 9192 10308 9196 10364
rect 9196 10308 9252 10364
rect 9252 10308 9256 10364
rect 9192 10304 9256 10308
rect 16952 10364 17016 10368
rect 16952 10308 16956 10364
rect 16956 10308 17012 10364
rect 17012 10308 17016 10364
rect 16952 10304 17016 10308
rect 17032 10364 17096 10368
rect 17032 10308 17036 10364
rect 17036 10308 17092 10364
rect 17092 10308 17096 10364
rect 17032 10304 17096 10308
rect 17112 10364 17176 10368
rect 17112 10308 17116 10364
rect 17116 10308 17172 10364
rect 17172 10308 17176 10364
rect 17112 10304 17176 10308
rect 17192 10364 17256 10368
rect 17192 10308 17196 10364
rect 17196 10308 17252 10364
rect 17252 10308 17256 10364
rect 17192 10304 17256 10308
rect 4952 9820 5016 9824
rect 4952 9764 4956 9820
rect 4956 9764 5012 9820
rect 5012 9764 5016 9820
rect 4952 9760 5016 9764
rect 5032 9820 5096 9824
rect 5032 9764 5036 9820
rect 5036 9764 5092 9820
rect 5092 9764 5096 9820
rect 5032 9760 5096 9764
rect 5112 9820 5176 9824
rect 5112 9764 5116 9820
rect 5116 9764 5172 9820
rect 5172 9764 5176 9820
rect 5112 9760 5176 9764
rect 5192 9820 5256 9824
rect 5192 9764 5196 9820
rect 5196 9764 5252 9820
rect 5252 9764 5256 9820
rect 5192 9760 5256 9764
rect 12952 9820 13016 9824
rect 12952 9764 12956 9820
rect 12956 9764 13012 9820
rect 13012 9764 13016 9820
rect 12952 9760 13016 9764
rect 13032 9820 13096 9824
rect 13032 9764 13036 9820
rect 13036 9764 13092 9820
rect 13092 9764 13096 9820
rect 13032 9760 13096 9764
rect 13112 9820 13176 9824
rect 13112 9764 13116 9820
rect 13116 9764 13172 9820
rect 13172 9764 13176 9820
rect 13112 9760 13176 9764
rect 13192 9820 13256 9824
rect 13192 9764 13196 9820
rect 13196 9764 13252 9820
rect 13252 9764 13256 9820
rect 13192 9760 13256 9764
rect 20952 9820 21016 9824
rect 20952 9764 20956 9820
rect 20956 9764 21012 9820
rect 21012 9764 21016 9820
rect 20952 9760 21016 9764
rect 21032 9820 21096 9824
rect 21032 9764 21036 9820
rect 21036 9764 21092 9820
rect 21092 9764 21096 9820
rect 21032 9760 21096 9764
rect 21112 9820 21176 9824
rect 21112 9764 21116 9820
rect 21116 9764 21172 9820
rect 21172 9764 21176 9820
rect 21112 9760 21176 9764
rect 21192 9820 21256 9824
rect 21192 9764 21196 9820
rect 21196 9764 21252 9820
rect 21252 9764 21256 9820
rect 21192 9760 21256 9764
rect 60 9284 124 9348
rect 8952 9276 9016 9280
rect 8952 9220 8956 9276
rect 8956 9220 9012 9276
rect 9012 9220 9016 9276
rect 8952 9216 9016 9220
rect 9032 9276 9096 9280
rect 9032 9220 9036 9276
rect 9036 9220 9092 9276
rect 9092 9220 9096 9276
rect 9032 9216 9096 9220
rect 9112 9276 9176 9280
rect 9112 9220 9116 9276
rect 9116 9220 9172 9276
rect 9172 9220 9176 9276
rect 9112 9216 9176 9220
rect 9192 9276 9256 9280
rect 9192 9220 9196 9276
rect 9196 9220 9252 9276
rect 9252 9220 9256 9276
rect 9192 9216 9256 9220
rect 16952 9276 17016 9280
rect 16952 9220 16956 9276
rect 16956 9220 17012 9276
rect 17012 9220 17016 9276
rect 16952 9216 17016 9220
rect 17032 9276 17096 9280
rect 17032 9220 17036 9276
rect 17036 9220 17092 9276
rect 17092 9220 17096 9276
rect 17032 9216 17096 9220
rect 17112 9276 17176 9280
rect 17112 9220 17116 9276
rect 17116 9220 17172 9276
rect 17172 9220 17176 9276
rect 17112 9216 17176 9220
rect 17192 9276 17256 9280
rect 17192 9220 17196 9276
rect 17196 9220 17252 9276
rect 17252 9220 17256 9276
rect 17192 9216 17256 9220
rect 60 9012 124 9076
rect 4952 8732 5016 8736
rect 4952 8676 4956 8732
rect 4956 8676 5012 8732
rect 5012 8676 5016 8732
rect 4952 8672 5016 8676
rect 5032 8732 5096 8736
rect 5032 8676 5036 8732
rect 5036 8676 5092 8732
rect 5092 8676 5096 8732
rect 5032 8672 5096 8676
rect 5112 8732 5176 8736
rect 5112 8676 5116 8732
rect 5116 8676 5172 8732
rect 5172 8676 5176 8732
rect 5112 8672 5176 8676
rect 5192 8732 5256 8736
rect 5192 8676 5196 8732
rect 5196 8676 5252 8732
rect 5252 8676 5256 8732
rect 5192 8672 5256 8676
rect 12952 8732 13016 8736
rect 12952 8676 12956 8732
rect 12956 8676 13012 8732
rect 13012 8676 13016 8732
rect 12952 8672 13016 8676
rect 13032 8732 13096 8736
rect 13032 8676 13036 8732
rect 13036 8676 13092 8732
rect 13092 8676 13096 8732
rect 13032 8672 13096 8676
rect 13112 8732 13176 8736
rect 13112 8676 13116 8732
rect 13116 8676 13172 8732
rect 13172 8676 13176 8732
rect 13112 8672 13176 8676
rect 13192 8732 13256 8736
rect 13192 8676 13196 8732
rect 13196 8676 13252 8732
rect 13252 8676 13256 8732
rect 13192 8672 13256 8676
rect 20952 8732 21016 8736
rect 20952 8676 20956 8732
rect 20956 8676 21012 8732
rect 21012 8676 21016 8732
rect 20952 8672 21016 8676
rect 21032 8732 21096 8736
rect 21032 8676 21036 8732
rect 21036 8676 21092 8732
rect 21092 8676 21096 8732
rect 21032 8672 21096 8676
rect 21112 8732 21176 8736
rect 21112 8676 21116 8732
rect 21116 8676 21172 8732
rect 21172 8676 21176 8732
rect 21112 8672 21176 8676
rect 21192 8732 21256 8736
rect 21192 8676 21196 8732
rect 21196 8676 21252 8732
rect 21252 8676 21256 8732
rect 21192 8672 21256 8676
rect 8952 8188 9016 8192
rect 8952 8132 8956 8188
rect 8956 8132 9012 8188
rect 9012 8132 9016 8188
rect 8952 8128 9016 8132
rect 9032 8188 9096 8192
rect 9032 8132 9036 8188
rect 9036 8132 9092 8188
rect 9092 8132 9096 8188
rect 9032 8128 9096 8132
rect 9112 8188 9176 8192
rect 9112 8132 9116 8188
rect 9116 8132 9172 8188
rect 9172 8132 9176 8188
rect 9112 8128 9176 8132
rect 9192 8188 9256 8192
rect 9192 8132 9196 8188
rect 9196 8132 9252 8188
rect 9252 8132 9256 8188
rect 9192 8128 9256 8132
rect 16952 8188 17016 8192
rect 16952 8132 16956 8188
rect 16956 8132 17012 8188
rect 17012 8132 17016 8188
rect 16952 8128 17016 8132
rect 17032 8188 17096 8192
rect 17032 8132 17036 8188
rect 17036 8132 17092 8188
rect 17092 8132 17096 8188
rect 17032 8128 17096 8132
rect 17112 8188 17176 8192
rect 17112 8132 17116 8188
rect 17116 8132 17172 8188
rect 17172 8132 17176 8188
rect 17112 8128 17176 8132
rect 17192 8188 17256 8192
rect 17192 8132 17196 8188
rect 17196 8132 17252 8188
rect 17252 8132 17256 8188
rect 17192 8128 17256 8132
rect 4952 7644 5016 7648
rect 4952 7588 4956 7644
rect 4956 7588 5012 7644
rect 5012 7588 5016 7644
rect 4952 7584 5016 7588
rect 5032 7644 5096 7648
rect 5032 7588 5036 7644
rect 5036 7588 5092 7644
rect 5092 7588 5096 7644
rect 5032 7584 5096 7588
rect 5112 7644 5176 7648
rect 5112 7588 5116 7644
rect 5116 7588 5172 7644
rect 5172 7588 5176 7644
rect 5112 7584 5176 7588
rect 5192 7644 5256 7648
rect 5192 7588 5196 7644
rect 5196 7588 5252 7644
rect 5252 7588 5256 7644
rect 5192 7584 5256 7588
rect 12952 7644 13016 7648
rect 12952 7588 12956 7644
rect 12956 7588 13012 7644
rect 13012 7588 13016 7644
rect 12952 7584 13016 7588
rect 13032 7644 13096 7648
rect 13032 7588 13036 7644
rect 13036 7588 13092 7644
rect 13092 7588 13096 7644
rect 13032 7584 13096 7588
rect 13112 7644 13176 7648
rect 13112 7588 13116 7644
rect 13116 7588 13172 7644
rect 13172 7588 13176 7644
rect 13112 7584 13176 7588
rect 13192 7644 13256 7648
rect 13192 7588 13196 7644
rect 13196 7588 13252 7644
rect 13252 7588 13256 7644
rect 13192 7584 13256 7588
rect 20952 7644 21016 7648
rect 20952 7588 20956 7644
rect 20956 7588 21012 7644
rect 21012 7588 21016 7644
rect 20952 7584 21016 7588
rect 21032 7644 21096 7648
rect 21032 7588 21036 7644
rect 21036 7588 21092 7644
rect 21092 7588 21096 7644
rect 21032 7584 21096 7588
rect 21112 7644 21176 7648
rect 21112 7588 21116 7644
rect 21116 7588 21172 7644
rect 21172 7588 21176 7644
rect 21112 7584 21176 7588
rect 21192 7644 21256 7648
rect 21192 7588 21196 7644
rect 21196 7588 21252 7644
rect 21252 7588 21256 7644
rect 21192 7584 21256 7588
rect 23612 7380 23676 7444
rect 23612 7108 23676 7172
rect 8952 7100 9016 7104
rect 8952 7044 8956 7100
rect 8956 7044 9012 7100
rect 9012 7044 9016 7100
rect 8952 7040 9016 7044
rect 9032 7100 9096 7104
rect 9032 7044 9036 7100
rect 9036 7044 9092 7100
rect 9092 7044 9096 7100
rect 9032 7040 9096 7044
rect 9112 7100 9176 7104
rect 9112 7044 9116 7100
rect 9116 7044 9172 7100
rect 9172 7044 9176 7100
rect 9112 7040 9176 7044
rect 9192 7100 9256 7104
rect 9192 7044 9196 7100
rect 9196 7044 9252 7100
rect 9252 7044 9256 7100
rect 9192 7040 9256 7044
rect 16952 7100 17016 7104
rect 16952 7044 16956 7100
rect 16956 7044 17012 7100
rect 17012 7044 17016 7100
rect 16952 7040 17016 7044
rect 17032 7100 17096 7104
rect 17032 7044 17036 7100
rect 17036 7044 17092 7100
rect 17092 7044 17096 7100
rect 17032 7040 17096 7044
rect 17112 7100 17176 7104
rect 17112 7044 17116 7100
rect 17116 7044 17172 7100
rect 17172 7044 17176 7100
rect 17112 7040 17176 7044
rect 17192 7100 17256 7104
rect 17192 7044 17196 7100
rect 17196 7044 17252 7100
rect 17252 7044 17256 7100
rect 17192 7040 17256 7044
rect 4952 6556 5016 6560
rect 4952 6500 4956 6556
rect 4956 6500 5012 6556
rect 5012 6500 5016 6556
rect 4952 6496 5016 6500
rect 5032 6556 5096 6560
rect 5032 6500 5036 6556
rect 5036 6500 5092 6556
rect 5092 6500 5096 6556
rect 5032 6496 5096 6500
rect 5112 6556 5176 6560
rect 5112 6500 5116 6556
rect 5116 6500 5172 6556
rect 5172 6500 5176 6556
rect 5112 6496 5176 6500
rect 5192 6556 5256 6560
rect 5192 6500 5196 6556
rect 5196 6500 5252 6556
rect 5252 6500 5256 6556
rect 5192 6496 5256 6500
rect 12952 6556 13016 6560
rect 12952 6500 12956 6556
rect 12956 6500 13012 6556
rect 13012 6500 13016 6556
rect 12952 6496 13016 6500
rect 13032 6556 13096 6560
rect 13032 6500 13036 6556
rect 13036 6500 13092 6556
rect 13092 6500 13096 6556
rect 13032 6496 13096 6500
rect 13112 6556 13176 6560
rect 13112 6500 13116 6556
rect 13116 6500 13172 6556
rect 13172 6500 13176 6556
rect 13112 6496 13176 6500
rect 13192 6556 13256 6560
rect 13192 6500 13196 6556
rect 13196 6500 13252 6556
rect 13252 6500 13256 6556
rect 13192 6496 13256 6500
rect 20952 6556 21016 6560
rect 20952 6500 20956 6556
rect 20956 6500 21012 6556
rect 21012 6500 21016 6556
rect 20952 6496 21016 6500
rect 21032 6556 21096 6560
rect 21032 6500 21036 6556
rect 21036 6500 21092 6556
rect 21092 6500 21096 6556
rect 21032 6496 21096 6500
rect 21112 6556 21176 6560
rect 21112 6500 21116 6556
rect 21116 6500 21172 6556
rect 21172 6500 21176 6556
rect 21112 6496 21176 6500
rect 21192 6556 21256 6560
rect 21192 6500 21196 6556
rect 21196 6500 21252 6556
rect 21252 6500 21256 6556
rect 21192 6496 21256 6500
rect 8952 6012 9016 6016
rect 8952 5956 8956 6012
rect 8956 5956 9012 6012
rect 9012 5956 9016 6012
rect 8952 5952 9016 5956
rect 9032 6012 9096 6016
rect 9032 5956 9036 6012
rect 9036 5956 9092 6012
rect 9092 5956 9096 6012
rect 9032 5952 9096 5956
rect 9112 6012 9176 6016
rect 9112 5956 9116 6012
rect 9116 5956 9172 6012
rect 9172 5956 9176 6012
rect 9112 5952 9176 5956
rect 9192 6012 9256 6016
rect 9192 5956 9196 6012
rect 9196 5956 9252 6012
rect 9252 5956 9256 6012
rect 9192 5952 9256 5956
rect 16952 6012 17016 6016
rect 16952 5956 16956 6012
rect 16956 5956 17012 6012
rect 17012 5956 17016 6012
rect 16952 5952 17016 5956
rect 17032 6012 17096 6016
rect 17032 5956 17036 6012
rect 17036 5956 17092 6012
rect 17092 5956 17096 6012
rect 17032 5952 17096 5956
rect 17112 6012 17176 6016
rect 17112 5956 17116 6012
rect 17116 5956 17172 6012
rect 17172 5956 17176 6012
rect 17112 5952 17176 5956
rect 17192 6012 17256 6016
rect 17192 5956 17196 6012
rect 17196 5956 17252 6012
rect 17252 5956 17256 6012
rect 17192 5952 17256 5956
rect 4952 5468 5016 5472
rect 4952 5412 4956 5468
rect 4956 5412 5012 5468
rect 5012 5412 5016 5468
rect 4952 5408 5016 5412
rect 5032 5468 5096 5472
rect 5032 5412 5036 5468
rect 5036 5412 5092 5468
rect 5092 5412 5096 5468
rect 5032 5408 5096 5412
rect 5112 5468 5176 5472
rect 5112 5412 5116 5468
rect 5116 5412 5172 5468
rect 5172 5412 5176 5468
rect 5112 5408 5176 5412
rect 5192 5468 5256 5472
rect 5192 5412 5196 5468
rect 5196 5412 5252 5468
rect 5252 5412 5256 5468
rect 5192 5408 5256 5412
rect 12952 5468 13016 5472
rect 12952 5412 12956 5468
rect 12956 5412 13012 5468
rect 13012 5412 13016 5468
rect 12952 5408 13016 5412
rect 13032 5468 13096 5472
rect 13032 5412 13036 5468
rect 13036 5412 13092 5468
rect 13092 5412 13096 5468
rect 13032 5408 13096 5412
rect 13112 5468 13176 5472
rect 13112 5412 13116 5468
rect 13116 5412 13172 5468
rect 13172 5412 13176 5468
rect 13112 5408 13176 5412
rect 13192 5468 13256 5472
rect 13192 5412 13196 5468
rect 13196 5412 13252 5468
rect 13252 5412 13256 5468
rect 13192 5408 13256 5412
rect 20952 5468 21016 5472
rect 20952 5412 20956 5468
rect 20956 5412 21012 5468
rect 21012 5412 21016 5468
rect 20952 5408 21016 5412
rect 21032 5468 21096 5472
rect 21032 5412 21036 5468
rect 21036 5412 21092 5468
rect 21092 5412 21096 5468
rect 21032 5408 21096 5412
rect 21112 5468 21176 5472
rect 21112 5412 21116 5468
rect 21116 5412 21172 5468
rect 21172 5412 21176 5468
rect 21112 5408 21176 5412
rect 21192 5468 21256 5472
rect 21192 5412 21196 5468
rect 21196 5412 21252 5468
rect 21252 5412 21256 5468
rect 21192 5408 21256 5412
rect 8952 4924 9016 4928
rect 8952 4868 8956 4924
rect 8956 4868 9012 4924
rect 9012 4868 9016 4924
rect 8952 4864 9016 4868
rect 9032 4924 9096 4928
rect 9032 4868 9036 4924
rect 9036 4868 9092 4924
rect 9092 4868 9096 4924
rect 9032 4864 9096 4868
rect 9112 4924 9176 4928
rect 9112 4868 9116 4924
rect 9116 4868 9172 4924
rect 9172 4868 9176 4924
rect 9112 4864 9176 4868
rect 9192 4924 9256 4928
rect 9192 4868 9196 4924
rect 9196 4868 9252 4924
rect 9252 4868 9256 4924
rect 9192 4864 9256 4868
rect 16952 4924 17016 4928
rect 16952 4868 16956 4924
rect 16956 4868 17012 4924
rect 17012 4868 17016 4924
rect 16952 4864 17016 4868
rect 17032 4924 17096 4928
rect 17032 4868 17036 4924
rect 17036 4868 17092 4924
rect 17092 4868 17096 4924
rect 17032 4864 17096 4868
rect 17112 4924 17176 4928
rect 17112 4868 17116 4924
rect 17116 4868 17172 4924
rect 17172 4868 17176 4924
rect 17112 4864 17176 4868
rect 17192 4924 17256 4928
rect 17192 4868 17196 4924
rect 17196 4868 17252 4924
rect 17252 4868 17256 4924
rect 17192 4864 17256 4868
rect 4952 4380 5016 4384
rect 4952 4324 4956 4380
rect 4956 4324 5012 4380
rect 5012 4324 5016 4380
rect 4952 4320 5016 4324
rect 5032 4380 5096 4384
rect 5032 4324 5036 4380
rect 5036 4324 5092 4380
rect 5092 4324 5096 4380
rect 5032 4320 5096 4324
rect 5112 4380 5176 4384
rect 5112 4324 5116 4380
rect 5116 4324 5172 4380
rect 5172 4324 5176 4380
rect 5112 4320 5176 4324
rect 5192 4380 5256 4384
rect 5192 4324 5196 4380
rect 5196 4324 5252 4380
rect 5252 4324 5256 4380
rect 5192 4320 5256 4324
rect 12952 4380 13016 4384
rect 12952 4324 12956 4380
rect 12956 4324 13012 4380
rect 13012 4324 13016 4380
rect 12952 4320 13016 4324
rect 13032 4380 13096 4384
rect 13032 4324 13036 4380
rect 13036 4324 13092 4380
rect 13092 4324 13096 4380
rect 13032 4320 13096 4324
rect 13112 4380 13176 4384
rect 13112 4324 13116 4380
rect 13116 4324 13172 4380
rect 13172 4324 13176 4380
rect 13112 4320 13176 4324
rect 13192 4380 13256 4384
rect 13192 4324 13196 4380
rect 13196 4324 13252 4380
rect 13252 4324 13256 4380
rect 13192 4320 13256 4324
rect 20952 4380 21016 4384
rect 20952 4324 20956 4380
rect 20956 4324 21012 4380
rect 21012 4324 21016 4380
rect 20952 4320 21016 4324
rect 21032 4380 21096 4384
rect 21032 4324 21036 4380
rect 21036 4324 21092 4380
rect 21092 4324 21096 4380
rect 21032 4320 21096 4324
rect 21112 4380 21176 4384
rect 21112 4324 21116 4380
rect 21116 4324 21172 4380
rect 21172 4324 21176 4380
rect 21112 4320 21176 4324
rect 21192 4380 21256 4384
rect 21192 4324 21196 4380
rect 21196 4324 21252 4380
rect 21252 4324 21256 4380
rect 21192 4320 21256 4324
rect 60 4252 124 4316
rect 60 3980 124 4044
rect 8952 3836 9016 3840
rect 8952 3780 8956 3836
rect 8956 3780 9012 3836
rect 9012 3780 9016 3836
rect 8952 3776 9016 3780
rect 9032 3836 9096 3840
rect 9032 3780 9036 3836
rect 9036 3780 9092 3836
rect 9092 3780 9096 3836
rect 9032 3776 9096 3780
rect 9112 3836 9176 3840
rect 9112 3780 9116 3836
rect 9116 3780 9172 3836
rect 9172 3780 9176 3836
rect 9112 3776 9176 3780
rect 9192 3836 9256 3840
rect 9192 3780 9196 3836
rect 9196 3780 9252 3836
rect 9252 3780 9256 3836
rect 9192 3776 9256 3780
rect 16952 3836 17016 3840
rect 16952 3780 16956 3836
rect 16956 3780 17012 3836
rect 17012 3780 17016 3836
rect 16952 3776 17016 3780
rect 17032 3836 17096 3840
rect 17032 3780 17036 3836
rect 17036 3780 17092 3836
rect 17092 3780 17096 3836
rect 17032 3776 17096 3780
rect 17112 3836 17176 3840
rect 17112 3780 17116 3836
rect 17116 3780 17172 3836
rect 17172 3780 17176 3836
rect 17112 3776 17176 3780
rect 17192 3836 17256 3840
rect 17192 3780 17196 3836
rect 17196 3780 17252 3836
rect 17252 3780 17256 3836
rect 17192 3776 17256 3780
rect 4952 3292 5016 3296
rect 4952 3236 4956 3292
rect 4956 3236 5012 3292
rect 5012 3236 5016 3292
rect 4952 3232 5016 3236
rect 5032 3292 5096 3296
rect 5032 3236 5036 3292
rect 5036 3236 5092 3292
rect 5092 3236 5096 3292
rect 5032 3232 5096 3236
rect 5112 3292 5176 3296
rect 5112 3236 5116 3292
rect 5116 3236 5172 3292
rect 5172 3236 5176 3292
rect 5112 3232 5176 3236
rect 5192 3292 5256 3296
rect 5192 3236 5196 3292
rect 5196 3236 5252 3292
rect 5252 3236 5256 3292
rect 5192 3232 5256 3236
rect 12952 3292 13016 3296
rect 12952 3236 12956 3292
rect 12956 3236 13012 3292
rect 13012 3236 13016 3292
rect 12952 3232 13016 3236
rect 13032 3292 13096 3296
rect 13032 3236 13036 3292
rect 13036 3236 13092 3292
rect 13092 3236 13096 3292
rect 13032 3232 13096 3236
rect 13112 3292 13176 3296
rect 13112 3236 13116 3292
rect 13116 3236 13172 3292
rect 13172 3236 13176 3292
rect 13112 3232 13176 3236
rect 13192 3292 13256 3296
rect 13192 3236 13196 3292
rect 13196 3236 13252 3292
rect 13252 3236 13256 3292
rect 13192 3232 13256 3236
rect 20952 3292 21016 3296
rect 20952 3236 20956 3292
rect 20956 3236 21012 3292
rect 21012 3236 21016 3292
rect 20952 3232 21016 3236
rect 21032 3292 21096 3296
rect 21032 3236 21036 3292
rect 21036 3236 21092 3292
rect 21092 3236 21096 3292
rect 21032 3232 21096 3236
rect 21112 3292 21176 3296
rect 21112 3236 21116 3292
rect 21116 3236 21172 3292
rect 21172 3236 21176 3292
rect 21112 3232 21176 3236
rect 21192 3292 21256 3296
rect 21192 3236 21196 3292
rect 21196 3236 21252 3292
rect 21252 3236 21256 3292
rect 21192 3232 21256 3236
rect 8952 2748 9016 2752
rect 8952 2692 8956 2748
rect 8956 2692 9012 2748
rect 9012 2692 9016 2748
rect 8952 2688 9016 2692
rect 9032 2748 9096 2752
rect 9032 2692 9036 2748
rect 9036 2692 9092 2748
rect 9092 2692 9096 2748
rect 9032 2688 9096 2692
rect 9112 2748 9176 2752
rect 9112 2692 9116 2748
rect 9116 2692 9172 2748
rect 9172 2692 9176 2748
rect 9112 2688 9176 2692
rect 9192 2748 9256 2752
rect 9192 2692 9196 2748
rect 9196 2692 9252 2748
rect 9252 2692 9256 2748
rect 9192 2688 9256 2692
rect 16952 2748 17016 2752
rect 16952 2692 16956 2748
rect 16956 2692 17012 2748
rect 17012 2692 17016 2748
rect 16952 2688 17016 2692
rect 17032 2748 17096 2752
rect 17032 2692 17036 2748
rect 17036 2692 17092 2748
rect 17092 2692 17096 2748
rect 17032 2688 17096 2692
rect 17112 2748 17176 2752
rect 17112 2692 17116 2748
rect 17116 2692 17172 2748
rect 17172 2692 17176 2748
rect 17112 2688 17176 2692
rect 17192 2748 17256 2752
rect 17192 2692 17196 2748
rect 17196 2692 17252 2748
rect 17252 2692 17256 2748
rect 17192 2688 17256 2692
rect 4952 2204 5016 2208
rect 4952 2148 4956 2204
rect 4956 2148 5012 2204
rect 5012 2148 5016 2204
rect 4952 2144 5016 2148
rect 5032 2204 5096 2208
rect 5032 2148 5036 2204
rect 5036 2148 5092 2204
rect 5092 2148 5096 2204
rect 5032 2144 5096 2148
rect 5112 2204 5176 2208
rect 5112 2148 5116 2204
rect 5116 2148 5172 2204
rect 5172 2148 5176 2204
rect 5112 2144 5176 2148
rect 5192 2204 5256 2208
rect 5192 2148 5196 2204
rect 5196 2148 5252 2204
rect 5252 2148 5256 2204
rect 5192 2144 5256 2148
rect 12952 2204 13016 2208
rect 12952 2148 12956 2204
rect 12956 2148 13012 2204
rect 13012 2148 13016 2204
rect 12952 2144 13016 2148
rect 13032 2204 13096 2208
rect 13032 2148 13036 2204
rect 13036 2148 13092 2204
rect 13092 2148 13096 2204
rect 13032 2144 13096 2148
rect 13112 2204 13176 2208
rect 13112 2148 13116 2204
rect 13116 2148 13172 2204
rect 13172 2148 13176 2204
rect 13112 2144 13176 2148
rect 13192 2204 13256 2208
rect 13192 2148 13196 2204
rect 13196 2148 13252 2204
rect 13252 2148 13256 2204
rect 13192 2144 13256 2148
rect 20952 2204 21016 2208
rect 20952 2148 20956 2204
rect 20956 2148 21012 2204
rect 21012 2148 21016 2204
rect 20952 2144 21016 2148
rect 21032 2204 21096 2208
rect 21032 2148 21036 2204
rect 21036 2148 21092 2204
rect 21092 2148 21096 2204
rect 21032 2144 21096 2148
rect 21112 2204 21176 2208
rect 21112 2148 21116 2204
rect 21116 2148 21172 2204
rect 21172 2148 21176 2204
rect 21112 2144 21176 2148
rect 21192 2204 21256 2208
rect 21192 2148 21196 2204
rect 21196 2148 21252 2204
rect 21252 2148 21256 2204
rect 21192 2144 21256 2148
<< metal4 >>
rect 4944 21792 5264 21808
rect 4944 21728 4952 21792
rect 5016 21728 5032 21792
rect 5096 21728 5112 21792
rect 5176 21728 5192 21792
rect 5256 21728 5264 21792
rect 4944 20704 5264 21728
rect 4944 20640 4952 20704
rect 5016 20640 5032 20704
rect 5096 20640 5112 20704
rect 5176 20640 5192 20704
rect 5256 20640 5264 20704
rect 4944 19616 5264 20640
rect 4944 19552 4952 19616
rect 5016 19552 5032 19616
rect 5096 19552 5112 19616
rect 5176 19552 5192 19616
rect 5256 19552 5264 19616
rect 4944 18528 5264 19552
rect 4944 18464 4952 18528
rect 5016 18464 5032 18528
rect 5096 18464 5112 18528
rect 5176 18464 5192 18528
rect 5256 18464 5264 18528
rect 4944 17440 5264 18464
rect 4944 17376 4952 17440
rect 5016 17376 5032 17440
rect 5096 17376 5112 17440
rect 5176 17376 5192 17440
rect 5256 17376 5264 17440
rect 4944 16352 5264 17376
rect 4944 16288 4952 16352
rect 5016 16288 5032 16352
rect 5096 16288 5112 16352
rect 5176 16288 5192 16352
rect 5256 16288 5264 16352
rect 4944 15264 5264 16288
rect 4944 15200 4952 15264
rect 5016 15200 5032 15264
rect 5096 15200 5112 15264
rect 5176 15200 5192 15264
rect 5256 15200 5264 15264
rect 4944 14176 5264 15200
rect 4944 14112 4952 14176
rect 5016 14112 5032 14176
rect 5096 14112 5112 14176
rect 5176 14112 5192 14176
rect 5256 14112 5264 14176
rect 4944 13088 5264 14112
rect 4944 13024 4952 13088
rect 5016 13024 5032 13088
rect 5096 13024 5112 13088
rect 5176 13024 5192 13088
rect 5256 13024 5264 13088
rect 4944 12000 5264 13024
rect 4944 11936 4952 12000
rect 5016 11936 5032 12000
rect 5096 11936 5112 12000
rect 5176 11936 5192 12000
rect 5256 11936 5264 12000
rect 59 11116 125 11117
rect 59 11052 60 11116
rect 124 11052 125 11116
rect 59 11051 125 11052
rect 62 10845 122 11051
rect 4944 10912 5264 11936
rect 4944 10848 4952 10912
rect 5016 10848 5032 10912
rect 5096 10848 5112 10912
rect 5176 10848 5192 10912
rect 5256 10848 5264 10912
rect 59 10844 125 10845
rect 59 10780 60 10844
rect 124 10780 125 10844
rect 59 10779 125 10780
rect 4944 9824 5264 10848
rect 4944 9760 4952 9824
rect 5016 9760 5032 9824
rect 5096 9760 5112 9824
rect 5176 9760 5192 9824
rect 5256 9760 5264 9824
rect 59 9348 125 9349
rect 59 9284 60 9348
rect 124 9284 125 9348
rect 59 9283 125 9284
rect 62 9077 122 9283
rect 59 9076 125 9077
rect 59 9012 60 9076
rect 124 9012 125 9076
rect 59 9011 125 9012
rect 4944 8736 5264 9760
rect 4944 8672 4952 8736
rect 5016 8672 5032 8736
rect 5096 8672 5112 8736
rect 5176 8672 5192 8736
rect 5256 8672 5264 8736
rect 4944 7648 5264 8672
rect 4944 7584 4952 7648
rect 5016 7584 5032 7648
rect 5096 7584 5112 7648
rect 5176 7584 5192 7648
rect 5256 7584 5264 7648
rect 4944 6560 5264 7584
rect 4944 6496 4952 6560
rect 5016 6496 5032 6560
rect 5096 6496 5112 6560
rect 5176 6496 5192 6560
rect 5256 6496 5264 6560
rect 4944 5472 5264 6496
rect 4944 5408 4952 5472
rect 5016 5408 5032 5472
rect 5096 5408 5112 5472
rect 5176 5408 5192 5472
rect 5256 5408 5264 5472
rect 4944 4384 5264 5408
rect 4944 4320 4952 4384
rect 5016 4320 5032 4384
rect 5096 4320 5112 4384
rect 5176 4320 5192 4384
rect 5256 4320 5264 4384
rect 59 4316 125 4317
rect 59 4252 60 4316
rect 124 4252 125 4316
rect 59 4251 125 4252
rect 62 4045 122 4251
rect 59 4044 125 4045
rect 59 3980 60 4044
rect 124 3980 125 4044
rect 59 3979 125 3980
rect 4944 3296 5264 4320
rect 4944 3232 4952 3296
rect 5016 3232 5032 3296
rect 5096 3232 5112 3296
rect 5176 3232 5192 3296
rect 5256 3232 5264 3296
rect 4944 2208 5264 3232
rect 4944 2144 4952 2208
rect 5016 2144 5032 2208
rect 5096 2144 5112 2208
rect 5176 2144 5192 2208
rect 5256 2144 5264 2208
rect 4944 2128 5264 2144
rect 8944 21248 9264 21808
rect 8944 21184 8952 21248
rect 9016 21184 9032 21248
rect 9096 21184 9112 21248
rect 9176 21184 9192 21248
rect 9256 21184 9264 21248
rect 8944 20160 9264 21184
rect 8944 20096 8952 20160
rect 9016 20096 9032 20160
rect 9096 20096 9112 20160
rect 9176 20096 9192 20160
rect 9256 20096 9264 20160
rect 8944 19072 9264 20096
rect 8944 19008 8952 19072
rect 9016 19008 9032 19072
rect 9096 19008 9112 19072
rect 9176 19008 9192 19072
rect 9256 19008 9264 19072
rect 8944 17984 9264 19008
rect 8944 17920 8952 17984
rect 9016 17920 9032 17984
rect 9096 17920 9112 17984
rect 9176 17920 9192 17984
rect 9256 17920 9264 17984
rect 8944 16896 9264 17920
rect 8944 16832 8952 16896
rect 9016 16832 9032 16896
rect 9096 16832 9112 16896
rect 9176 16832 9192 16896
rect 9256 16832 9264 16896
rect 8944 15808 9264 16832
rect 8944 15744 8952 15808
rect 9016 15744 9032 15808
rect 9096 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9264 15808
rect 8944 14720 9264 15744
rect 8944 14656 8952 14720
rect 9016 14656 9032 14720
rect 9096 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9264 14720
rect 8944 13632 9264 14656
rect 8944 13568 8952 13632
rect 9016 13568 9032 13632
rect 9096 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9264 13632
rect 8944 12544 9264 13568
rect 8944 12480 8952 12544
rect 9016 12480 9032 12544
rect 9096 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9264 12544
rect 8944 11456 9264 12480
rect 8944 11392 8952 11456
rect 9016 11392 9032 11456
rect 9096 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9264 11456
rect 8944 10368 9264 11392
rect 8944 10304 8952 10368
rect 9016 10304 9032 10368
rect 9096 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9264 10368
rect 8944 9280 9264 10304
rect 8944 9216 8952 9280
rect 9016 9216 9032 9280
rect 9096 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9264 9280
rect 8944 8192 9264 9216
rect 8944 8128 8952 8192
rect 9016 8128 9032 8192
rect 9096 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9264 8192
rect 8944 7104 9264 8128
rect 8944 7040 8952 7104
rect 9016 7040 9032 7104
rect 9096 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9264 7104
rect 8944 6016 9264 7040
rect 8944 5952 8952 6016
rect 9016 5952 9032 6016
rect 9096 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9264 6016
rect 8944 4928 9264 5952
rect 8944 4864 8952 4928
rect 9016 4864 9032 4928
rect 9096 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9264 4928
rect 8944 3840 9264 4864
rect 8944 3776 8952 3840
rect 9016 3776 9032 3840
rect 9096 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9264 3840
rect 8944 2752 9264 3776
rect 8944 2688 8952 2752
rect 9016 2688 9032 2752
rect 9096 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9264 2752
rect 8944 2128 9264 2688
rect 12944 21792 13264 21808
rect 12944 21728 12952 21792
rect 13016 21728 13032 21792
rect 13096 21728 13112 21792
rect 13176 21728 13192 21792
rect 13256 21728 13264 21792
rect 12944 20704 13264 21728
rect 12944 20640 12952 20704
rect 13016 20640 13032 20704
rect 13096 20640 13112 20704
rect 13176 20640 13192 20704
rect 13256 20640 13264 20704
rect 12944 19616 13264 20640
rect 12944 19552 12952 19616
rect 13016 19552 13032 19616
rect 13096 19552 13112 19616
rect 13176 19552 13192 19616
rect 13256 19552 13264 19616
rect 12944 18528 13264 19552
rect 12944 18464 12952 18528
rect 13016 18464 13032 18528
rect 13096 18464 13112 18528
rect 13176 18464 13192 18528
rect 13256 18464 13264 18528
rect 12944 17440 13264 18464
rect 12944 17376 12952 17440
rect 13016 17376 13032 17440
rect 13096 17376 13112 17440
rect 13176 17376 13192 17440
rect 13256 17376 13264 17440
rect 12944 16352 13264 17376
rect 12944 16288 12952 16352
rect 13016 16288 13032 16352
rect 13096 16288 13112 16352
rect 13176 16288 13192 16352
rect 13256 16288 13264 16352
rect 12944 15264 13264 16288
rect 12944 15200 12952 15264
rect 13016 15200 13032 15264
rect 13096 15200 13112 15264
rect 13176 15200 13192 15264
rect 13256 15200 13264 15264
rect 12944 14176 13264 15200
rect 12944 14112 12952 14176
rect 13016 14112 13032 14176
rect 13096 14112 13112 14176
rect 13176 14112 13192 14176
rect 13256 14112 13264 14176
rect 12944 13088 13264 14112
rect 12944 13024 12952 13088
rect 13016 13024 13032 13088
rect 13096 13024 13112 13088
rect 13176 13024 13192 13088
rect 13256 13024 13264 13088
rect 12944 12000 13264 13024
rect 12944 11936 12952 12000
rect 13016 11936 13032 12000
rect 13096 11936 13112 12000
rect 13176 11936 13192 12000
rect 13256 11936 13264 12000
rect 12944 10912 13264 11936
rect 12944 10848 12952 10912
rect 13016 10848 13032 10912
rect 13096 10848 13112 10912
rect 13176 10848 13192 10912
rect 13256 10848 13264 10912
rect 12944 9824 13264 10848
rect 12944 9760 12952 9824
rect 13016 9760 13032 9824
rect 13096 9760 13112 9824
rect 13176 9760 13192 9824
rect 13256 9760 13264 9824
rect 12944 8736 13264 9760
rect 12944 8672 12952 8736
rect 13016 8672 13032 8736
rect 13096 8672 13112 8736
rect 13176 8672 13192 8736
rect 13256 8672 13264 8736
rect 12944 7648 13264 8672
rect 12944 7584 12952 7648
rect 13016 7584 13032 7648
rect 13096 7584 13112 7648
rect 13176 7584 13192 7648
rect 13256 7584 13264 7648
rect 12944 6560 13264 7584
rect 12944 6496 12952 6560
rect 13016 6496 13032 6560
rect 13096 6496 13112 6560
rect 13176 6496 13192 6560
rect 13256 6496 13264 6560
rect 12944 5472 13264 6496
rect 12944 5408 12952 5472
rect 13016 5408 13032 5472
rect 13096 5408 13112 5472
rect 13176 5408 13192 5472
rect 13256 5408 13264 5472
rect 12944 4384 13264 5408
rect 12944 4320 12952 4384
rect 13016 4320 13032 4384
rect 13096 4320 13112 4384
rect 13176 4320 13192 4384
rect 13256 4320 13264 4384
rect 12944 3296 13264 4320
rect 12944 3232 12952 3296
rect 13016 3232 13032 3296
rect 13096 3232 13112 3296
rect 13176 3232 13192 3296
rect 13256 3232 13264 3296
rect 12944 2208 13264 3232
rect 12944 2144 12952 2208
rect 13016 2144 13032 2208
rect 13096 2144 13112 2208
rect 13176 2144 13192 2208
rect 13256 2144 13264 2208
rect 12944 2128 13264 2144
rect 16944 21248 17264 21808
rect 16944 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17264 21248
rect 16944 20160 17264 21184
rect 16944 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17264 20160
rect 16944 19072 17264 20096
rect 16944 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17264 19072
rect 16944 17984 17264 19008
rect 16944 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17264 17984
rect 16944 16896 17264 17920
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 16944 15808 17264 16832
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16944 14720 17264 15744
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16944 13632 17264 14656
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 12544 17264 13568
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16944 11456 17264 12480
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 10368 17264 11392
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16944 9280 17264 10304
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 8192 17264 9216
rect 16944 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17264 8192
rect 16944 7104 17264 8128
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 6016 17264 7040
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 4928 17264 5952
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 3840 17264 4864
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16944 2752 17264 3776
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 16944 2128 17264 2688
rect 20944 21792 21264 21808
rect 20944 21728 20952 21792
rect 21016 21728 21032 21792
rect 21096 21728 21112 21792
rect 21176 21728 21192 21792
rect 21256 21728 21264 21792
rect 20944 20704 21264 21728
rect 20944 20640 20952 20704
rect 21016 20640 21032 20704
rect 21096 20640 21112 20704
rect 21176 20640 21192 20704
rect 21256 20640 21264 20704
rect 20944 19616 21264 20640
rect 20944 19552 20952 19616
rect 21016 19552 21032 19616
rect 21096 19552 21112 19616
rect 21176 19552 21192 19616
rect 21256 19552 21264 19616
rect 20944 18528 21264 19552
rect 20944 18464 20952 18528
rect 21016 18464 21032 18528
rect 21096 18464 21112 18528
rect 21176 18464 21192 18528
rect 21256 18464 21264 18528
rect 20944 17440 21264 18464
rect 20944 17376 20952 17440
rect 21016 17376 21032 17440
rect 21096 17376 21112 17440
rect 21176 17376 21192 17440
rect 21256 17376 21264 17440
rect 20944 16352 21264 17376
rect 20944 16288 20952 16352
rect 21016 16288 21032 16352
rect 21096 16288 21112 16352
rect 21176 16288 21192 16352
rect 21256 16288 21264 16352
rect 20944 15264 21264 16288
rect 23611 15740 23677 15741
rect 23611 15676 23612 15740
rect 23676 15676 23677 15740
rect 23611 15675 23677 15676
rect 23614 15469 23674 15675
rect 23611 15468 23677 15469
rect 23611 15404 23612 15468
rect 23676 15404 23677 15468
rect 23611 15403 23677 15404
rect 20944 15200 20952 15264
rect 21016 15200 21032 15264
rect 21096 15200 21112 15264
rect 21176 15200 21192 15264
rect 21256 15200 21264 15264
rect 20944 14176 21264 15200
rect 20944 14112 20952 14176
rect 21016 14112 21032 14176
rect 21096 14112 21112 14176
rect 21176 14112 21192 14176
rect 21256 14112 21264 14176
rect 20944 13088 21264 14112
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 12000 21264 13024
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 10912 21264 11936
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 9824 21264 10848
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 8736 21264 9760
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 7648 21264 8672
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 6560 21264 7584
rect 23611 7444 23677 7445
rect 23611 7380 23612 7444
rect 23676 7380 23677 7444
rect 23611 7379 23677 7380
rect 23614 7173 23674 7379
rect 23611 7172 23677 7173
rect 23611 7108 23612 7172
rect 23676 7108 23677 7172
rect 23611 7107 23677 7108
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 5472 21264 6496
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 4384 21264 5408
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 3296 21264 4320
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 2208 21264 3232
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2128 21264 2144
use scs8hd_fill_2  FILLER_1_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_6
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_buf_2  _160_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_10
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__A
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_11 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_8  _058_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_decap_8  FILLER_0_23 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 3220 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_32
timestamp 1586364061
transform 1 0 4048 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_28
timestamp 1586364061
transform 1 0 3680 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_35
timestamp 1586364061
transform 1 0 4324 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3864 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_72 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_8  _070_
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5704 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_39 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_45
timestamp 1586364061
transform 1 0 5244 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_49 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5612 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_52
timestamp 1586364061
transform 1 0 5888 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 -1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_77
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_73
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_74 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_84
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 314 592
use scs8hd_conb_1  _148_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8556 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_88
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_105
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_101
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_103
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10948 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9568 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use scs8hd_decap_3  FILLER_1_113
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_115
timestamp 1586364061
transform 1 0 11684 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _156_
timestamp 1586364061
transform 1 0 11132 0 1 2720
box -38 -48 406 592
use scs8hd_buf_2  _155_
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_119
timestamp 1586364061
transform 1 0 12052 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11868 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12512 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_133
timestamp 1586364061
transform 1 0 13340 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_137
timestamp 1586364061
transform 1 0 13708 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_138
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13892 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _154_
timestamp 1586364061
transform 1 0 14168 0 -1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 14076 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_146
timestamp 1586364061
transform 1 0 14536 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_156
timestamp 1586364061
transform 1 0 15456 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_152
timestamp 1586364061
transform 1 0 15088 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 1 2720
box -38 -48 866 592
use scs8hd_buf_2  _164_
timestamp 1586364061
transform 1 0 17020 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_165
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_169
timestamp 1586364061
transform 1 0 16652 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_177
timestamp 1586364061
transform 1 0 17388 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_169
timestamp 1586364061
transform 1 0 16652 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_173
timestamp 1586364061
transform 1 0 17020 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_181
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_181
timestamp 1586364061
transform 1 0 17756 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 17572 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_187
timestamp 1586364061
transform 1 0 18308 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_185
timestamp 1586364061
transform 1 0 18124 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _163_
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use scs8hd_conb_1  _142_
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_191
timestamp 1586364061
transform 1 0 18676 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_191
timestamp 1586364061
transform 1 0 18676 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_195
timestamp 1586364061
transform 1 0 19044 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 18860 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 314 592
use scs8hd_buf_2  _170_
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 20056 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_204
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_198
timestamp 1586364061
transform 1 0 19320 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_202
timestamp 1586364061
transform 1 0 19688 0 1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_214
timestamp 1586364061
transform 1 0 20792 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_222
timestamp 1586364061
transform 1 0 21528 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_218
timestamp 1586364061
transform 1 0 21160 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_221
timestamp 1586364061
transform 1 0 21436 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_216
timestamp 1586364061
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_1_226
timestamp 1586364061
transform 1 0 21896 0 1 2720
box -38 -48 590 592
use scs8hd_decap_8  FILLER_0_225
timestamp 1586364061
transform 1 0 21804 0 -1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21712 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 22816 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 22816 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_inv_8  _072_
timestamp 1586364061
transform 1 0 4140 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_42
timestamp 1586364061
transform 1 0 4968 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_46
timestamp 1586364061
transform 1 0 5336 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_6  FILLER_2_53
timestamp 1586364061
transform 1 0 5980 0 -1 3808
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7176 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 6624 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_59
timestamp 1586364061
transform 1 0 6532 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_62
timestamp 1586364061
transform 1 0 6808 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8188 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__C
timestamp 1586364061
transform 1 0 8556 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_75
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_79
timestamp 1586364061
transform 1 0 8372 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_83
timestamp 1586364061
transform 1 0 8740 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_89
timestamp 1586364061
transform 1 0 9292 0 -1 3808
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_104
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11776 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 11592 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_108
timestamp 1586364061
transform 1 0 11040 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_112
timestamp 1586364061
transform 1 0 11408 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_8  _066_
timestamp 1586364061
transform 1 0 13616 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13340 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_127
timestamp 1586364061
transform 1 0 12788 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_131
timestamp 1586364061
transform 1 0 13156 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_135
timestamp 1586364061
transform 1 0 13524 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _165_
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_167
timestamp 1586364061
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_175
timestamp 1586364061
transform 1 0 17204 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17940 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19136 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_186
timestamp 1586364061
transform 1 0 18216 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_2_194
timestamp 1586364061
transform 1 0 18952 0 -1 3808
box -38 -48 222 592
use scs8hd_conb_1  _145_
timestamp 1586364061
transform 1 0 19412 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_198
timestamp 1586364061
transform 1 0 19320 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_218
timestamp 1586364061
transform 1 0 21160 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_2_230
timestamp 1586364061
transform 1 0 22264 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 22816 0 -1 3808
box -38 -48 314 592
use scs8hd_conb_1  _144_
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_6
timestamp 1586364061
transform 1 0 1656 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_10
timestamp 1586364061
transform 1 0 2024 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_14
timestamp 1586364061
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3864 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3680 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3312 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_18
timestamp 1586364061
transform 1 0 2760 0 1 3808
box -38 -48 590 592
use scs8hd_fill_2  FILLER_3_26
timestamp 1586364061
transform 1 0 3496 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5060 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5428 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_41
timestamp 1586364061
transform 1 0 4876 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_45
timestamp 1586364061
transform 1 0 5244 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_52
timestamp 1586364061
transform 1 0 5888 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6072 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7360 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_56
timestamp 1586364061
transform 1 0 6256 0 1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_66
timestamp 1586364061
transform 1 0 7176 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_70
timestamp 1586364061
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _136_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__136__D
timestamp 1586364061
transform 1 0 7728 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _069_
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__C
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_91
timestamp 1586364061
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_95
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__C
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__D
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_108
timestamp 1586364061
transform 1 0 11040 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_112
timestamp 1586364061
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_116
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_120
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _132_
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__132__D
timestamp 1586364061
transform 1 0 13340 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 12972 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_126
timestamp 1586364061
transform 1 0 12696 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_131
timestamp 1586364061
transform 1 0 13156 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__126__D
timestamp 1586364061
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_152
timestamp 1586364061
transform 1 0 15088 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_156
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__C
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_169
timestamp 1586364061
transform 1 0 16652 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_173
timestamp 1586364061
transform 1 0 17020 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_177
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _060_
timestamp 1586364061
transform 1 0 18952 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__060__A
timestamp 1586364061
transform 1 0 18768 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18216 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_181
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_188
timestamp 1586364061
transform 1 0 18400 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19964 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_203
timestamp 1586364061
transform 1 0 19780 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_207
timestamp 1586364061
transform 1 0 20148 0 1 3808
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__059__A
timestamp 1586364061
transform 1 0 20884 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_217
timestamp 1586364061
transform 1 0 21068 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_3_229
timestamp 1586364061
transform 1 0 22172 0 1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 22816 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_16
timestamp 1586364061
transform 1 0 2576 0 -1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4232 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 3680 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__D
timestamp 1586364061
transform 1 0 3312 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_26
timestamp 1586364061
transform 1 0 3496 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_30
timestamp 1586364061
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_43
timestamp 1586364061
transform 1 0 5060 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_4_51
timestamp 1586364061
transform 1 0 5796 0 -1 4896
box -38 -48 314 592
use scs8hd_or3_4  _110_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6624 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 6440 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__C
timestamp 1586364061
transform 1 0 6072 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_69
timestamp 1586364061
transform 1 0 7452 0 -1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8188 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 7912 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 8648 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_73
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_76
timestamp 1586364061
transform 1 0 8096 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 774 592
use scs8hd_nor4_4  _135_
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_nor4_4  _131_
timestamp 1586364061
transform 1 0 11960 0 -1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__131__D
timestamp 1586364061
transform 1 0 11776 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_110
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__132__C
timestamp 1586364061
transform 1 0 13708 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_135
timestamp 1586364061
transform 1 0 13524 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_139
timestamp 1586364061
transform 1 0 13892 0 -1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _126_
timestamp 1586364061
transform 1 0 15548 0 -1 4896
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__125__D
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_143
timestamp 1586364061
transform 1 0 14260 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17388 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_174
timestamp 1586364061
transform 1 0 17112 0 -1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17848 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19136 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18308 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_179
timestamp 1586364061
transform 1 0 17572 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_185
timestamp 1586364061
transform 1 0 18124 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_189
timestamp 1586364061
transform 1 0 18492 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_195
timestamp 1586364061
transform 1 0 19044 0 -1 4896
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_205
timestamp 1586364061
transform 1 0 19964 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_213
timestamp 1586364061
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use scs8hd_inv_8  _059_
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_224
timestamp 1586364061
transform 1 0 21712 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 22816 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_232
timestamp 1586364061
transform 1 0 22448 0 -1 4896
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_12
timestamp 1586364061
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_16
timestamp 1586364061
transform 1 0 2576 0 1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _138_
timestamp 1586364061
transform 1 0 3680 0 1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__138__D
timestamp 1586364061
transform 1 0 3496 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 3128 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 2760 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_20
timestamp 1586364061
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_24
timestamp 1586364061
transform 1 0 3312 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__C
timestamp 1586364061
transform 1 0 5428 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_45
timestamp 1586364061
transform 1 0 5244 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_49
timestamp 1586364061
transform 1 0 5612 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 130 592
use scs8hd_or3_4  _087_
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 6440 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 6072 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_56
timestamp 1586364061
transform 1 0 6256 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_60
timestamp 1586364061
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_71
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _057_
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__057__A
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__056__A
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_75
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_88
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 590 592
use scs8hd_inv_8  _053_
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__053__A
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_94
timestamp 1586364061
transform 1 0 9752 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_97
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_101
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _065_
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 590 592
use scs8hd_inv_8  _054_
timestamp 1586364061
transform 1 0 13984 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__054__A
timestamp 1586364061
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_132
timestamp 1586364061
transform 1 0 13248 0 1 4896
box -38 -48 590 592
use scs8hd_nor4_4  _125_
timestamp 1586364061
transform 1 0 15548 0 1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 15364 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14996 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_149
timestamp 1586364061
transform 1 0 14812 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_153
timestamp 1586364061
transform 1 0 15180 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_174
timestamp 1586364061
transform 1 0 17112 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_178
timestamp 1586364061
transform 1 0 17480 0 1 4896
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_195
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_199
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_212
timestamp 1586364061
transform 1 0 20608 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21804 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21160 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22172 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_216
timestamp 1586364061
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_223
timestamp 1586364061
transform 1 0 21620 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_227
timestamp 1586364061
transform 1 0 21988 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_231
timestamp 1586364061
transform 1 0 22356 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 22816 0 1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_16
timestamp 1586364061
transform 1 0 2576 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_12
timestamp 1586364061
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2668 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 2392 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 1472 0 -1 5984
box -38 -48 1050 592
use scs8hd_inv_8  _071_
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_23
timestamp 1586364061
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_26
timestamp 1586364061
transform 1 0 3496 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_19
timestamp 1586364061
transform 1 0 2852 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 2760 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 3312 0 -1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_32
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_30
timestamp 1586364061
transform 1 0 3864 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__C
timestamp 1586364061
transform 1 0 3680 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_nor4_4  _137_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1602 592
use scs8hd_or3_4  _074_
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_49
timestamp 1586364061
transform 1 0 5612 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_36
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_40
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_55
timestamp 1586364061
transform 1 0 6164 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__095__C
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__C
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_71
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_67
timestamp 1586364061
transform 1 0 7268 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use scs8hd_or3_4  _103_
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use scs8hd_or3_4  _095_
timestamp 1586364061
transform 1 0 6440 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_8  _055_
timestamp 1586364061
transform 1 0 8372 0 1 5984
box -38 -48 866 592
use scs8hd_inv_8  _056_
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__055__A
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_75
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_88
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9384 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_7_92
timestamp 1586364061
transform 1 0 9568 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_106
timestamp 1586364061
transform 1 0 10856 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_122
timestamp 1586364061
transform 1 0 12328 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12512 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_108
timestamp 1586364061
transform 1 0 11040 0 -1 5984
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12512 0 1 5984
box -38 -48 866 592
use scs8hd_or3_4  _111_
timestamp 1586364061
transform 1 0 14076 0 1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 13892 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_126
timestamp 1586364061
transform 1 0 12696 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_6_138
timestamp 1586364061
transform 1 0 13800 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_133
timestamp 1586364061
transform 1 0 13340 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_137
timestamp 1586364061
transform 1 0 13708 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_150
timestamp 1586364061
transform 1 0 14904 0 1 5984
box -38 -48 406 592
use scs8hd_decap_8  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_160
timestamp 1586364061
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_156
timestamp 1586364061
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_159
timestamp 1586364061
transform 1 0 15732 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__133__C
timestamp 1586364061
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 15548 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 15272 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_168
timestamp 1586364061
transform 1 0 16560 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_164
timestamp 1586364061
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_169
timestamp 1586364061
transform 1 0 16652 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_3  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__D
timestamp 1586364061
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__C
timestamp 1586364061
transform 1 0 15916 0 -1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17204 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 5984
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 17388 0 -1 5984
box -38 -48 1050 592
use scs8hd_inv_8  _067_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_188
timestamp 1586364061
transform 1 0 18400 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_194
timestamp 1586364061
transform 1 0 18952 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_193
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_205
timestamp 1586364061
transform 1 0 19964 0 1 5984
box -38 -48 314 592
use scs8hd_decap_6  FILLER_7_197
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19780 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_212
timestamp 1586364061
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_206
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20424 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21436 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21804 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_224
timestamp 1586364061
transform 1 0 21712 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_219
timestamp 1586364061
transform 1 0 21252 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_223
timestamp 1586364061
transform 1 0 21620 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_227
timestamp 1586364061
transform 1 0 21988 0 1 5984
box -38 -48 590 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 22816 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 22816 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_232
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 130 592
use scs8hd_conb_1  _139_
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 314 592
use scs8hd_buf_2  _158_
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1932 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2300 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_7
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_11
timestamp 1586364061
transform 1 0 2116 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4232 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_18
timestamp 1586364061
transform 1 0 2760 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_24
timestamp 1586364061
transform 1 0 3312 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _108_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4416 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__074__C
timestamp 1586364061
transform 1 0 5428 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5980 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_45
timestamp 1586364061
transform 1 0 5244 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_49
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6532 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6348 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_55
timestamp 1586364061
transform 1 0 6164 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_72
timestamp 1586364061
transform 1 0 7728 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_97
timestamp 1586364061
transform 1 0 10028 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_107
timestamp 1586364061
transform 1 0 10948 0 -1 7072
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12144 0 -1 7072
box -38 -48 866 592
use scs8hd_fill_1  FILLER_8_119
timestamp 1586364061
transform 1 0 12052 0 -1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13708 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__111__C
timestamp 1586364061
transform 1 0 14168 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13156 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_133
timestamp 1586364061
transform 1 0 13340 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_140
timestamp 1586364061
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use scs8hd_nor4_4  _133_
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 14536 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_144
timestamp 1586364061
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_148
timestamp 1586364061
transform 1 0 14720 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_152
timestamp 1586364061
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_171
timestamp 1586364061
transform 1 0 16836 0 -1 7072
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 17572 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18768 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_194
timestamp 1586364061
transform 1 0 18952 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_206
timestamp 1586364061
transform 1 0 20056 0 -1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_224
timestamp 1586364061
transform 1 0 21712 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 22816 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_232
timestamp 1586364061
transform 1 0 22448 0 -1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_17
timestamp 1586364061
transform 1 0 2668 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3404 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_21
timestamp 1586364061
transform 1 0 3036 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_34
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_38
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_71
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use scs8hd_or3_4  _118_
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__C
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_75
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_79
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_92
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_97
timestamp 1586364061
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_110
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12604 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_136
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__134__D
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 14904 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_148
timestamp 1586364061
transform 1 0 14720 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_152
timestamp 1586364061
transform 1 0 15088 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_156
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_160
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__C
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_164
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_195
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19872 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20332 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 20700 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_199
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_203
timestamp 1586364061
transform 1 0 19780 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_207
timestamp 1586364061
transform 1 0 20148 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_211
timestamp 1586364061
transform 1 0 20516 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _159_
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__061__A
timestamp 1586364061
transform 1 0 21436 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_219
timestamp 1586364061
transform 1 0 21252 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_223
timestamp 1586364061
transform 1 0 21620 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_231
timestamp 1586364061
transform 1 0 22356 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 22816 0 1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_18
timestamp 1586364061
transform 1 0 2760 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_10_30
timestamp 1586364061
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_6  FILLER_10_52
timestamp 1586364061
transform 1 0 5888 0 -1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6624 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_69
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_73
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_77
timestamp 1586364061
transform 1 0 8188 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_4  FILLER_10_85
timestamp 1586364061
transform 1 0 8924 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_89
timestamp 1586364061
transform 1 0 9292 0 -1 8160
box -38 -48 130 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 866 592
use scs8hd_conb_1  _140_
timestamp 1586364061
transform 1 0 9752 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10396 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_97
timestamp 1586364061
transform 1 0 10028 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_103
timestamp 1586364061
transform 1 0 10580 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12328 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_10_114
timestamp 1586364061
transform 1 0 11592 0 -1 8160
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13524 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_133
timestamp 1586364061
transform 1 0 13340 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_137
timestamp 1586364061
transform 1 0 13708 0 -1 8160
box -38 -48 1142 592
use scs8hd_nor4_4  _134_
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_149
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_171
timestamp 1586364061
transform 1 0 16836 0 -1 8160
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_183
timestamp 1586364061
transform 1 0 17940 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_193
timestamp 1586364061
transform 1 0 18860 0 -1 8160
box -38 -48 222 592
use scs8hd_conb_1  _143_
timestamp 1586364061
transform 1 0 19596 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_197
timestamp 1586364061
transform 1 0 19228 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_8  FILLER_10_204
timestamp 1586364061
transform 1 0 19872 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_212
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_8  _061_
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_224
timestamp 1586364061
transform 1 0 21712 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 22816 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_232
timestamp 1586364061
transform 1 0 22448 0 -1 8160
box -38 -48 130 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 1472 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__079__B
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_13
timestamp 1586364061
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_17
timestamp 1586364061
transform 1 0 2668 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3496 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3956 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 2852 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__C
timestamp 1586364061
transform 1 0 3220 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_21
timestamp 1586364061
transform 1 0 3036 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_25
timestamp 1586364061
transform 1 0 3404 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_29
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_33
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 5612 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_37
timestamp 1586364061
transform 1 0 4508 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_47
timestamp 1586364061
transform 1 0 5428 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_55
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_65
timestamp 1586364061
transform 1 0 7084 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_69
timestamp 1586364061
transform 1 0 7452 0 1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_84
timestamp 1586364061
transform 1 0 8832 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_88
timestamp 1586364061
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9568 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_103
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_107
timestamp 1586364061
transform 1 0 10948 0 1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_111
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 12696 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_128
timestamp 1586364061
transform 1 0 12880 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_139
timestamp 1586364061
transform 1 0 13892 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15824 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15088 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_151
timestamp 1586364061
transform 1 0 14996 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_154
timestamp 1586364061
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_158
timestamp 1586364061
transform 1 0 15640 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16008 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_173
timestamp 1586364061
transform 1 0 17020 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_177
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_194
timestamp 1586364061
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use scs8hd_inv_8  _068_
timestamp 1586364061
transform 1 0 19688 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 19504 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_198
timestamp 1586364061
transform 1 0 19320 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_211
timestamp 1586364061
transform 1 0 20516 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21252 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21712 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22080 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_217
timestamp 1586364061
transform 1 0 21068 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_222
timestamp 1586364061
transform 1 0 21528 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_226
timestamp 1586364061
transform 1 0 21896 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_230
timestamp 1586364061
transform 1 0 22264 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 22816 0 1 8160
box -38 -48 314 592
use scs8hd_or3_4  _079_
timestamp 1586364061
transform 1 0 2024 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_7
timestamp 1586364061
transform 1 0 1748 0 -1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3036 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_19
timestamp 1586364061
transform 1 0 2852 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_35
timestamp 1586364061
transform 1 0 4324 0 -1 9248
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 5336 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 4600 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 4968 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_40
timestamp 1586364061
transform 1 0 4784 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_57
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_61
timestamp 1586364061
transform 1 0 6716 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_64
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 8924 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_74
timestamp 1586364061
transform 1 0 7912 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_12_82
timestamp 1586364061
transform 1 0 8648 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_12_87
timestamp 1586364061
transform 1 0 9108 0 -1 9248
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_91
timestamp 1586364061
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_12_104
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11408 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_115
timestamp 1586364061
transform 1 0 11684 0 -1 9248
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 12696 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__096__C
timestamp 1586364061
transform 1 0 13892 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_125
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_137
timestamp 1586364061
transform 1 0 13708 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 15456 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__C
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 15824 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_149
timestamp 1586364061
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_158
timestamp 1586364061
transform 1 0 15640 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16008 0 -1 9248
box -38 -48 1050 592
use scs8hd_decap_12  FILLER_12_173
timestamp 1586364061
transform 1 0 17020 0 -1 9248
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18400 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18124 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_187
timestamp 1586364061
transform 1 0 18308 0 -1 9248
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20516 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_197
timestamp 1586364061
transform 1 0 19228 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_12_209
timestamp 1586364061
transform 1 0 20332 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_213
timestamp 1586364061
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_224
timestamp 1586364061
transform 1 0 21712 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 22816 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_232
timestamp 1586364061
transform 1 0 22448 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_buf_2  _153_
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_17
timestamp 1586364061
transform 1 0 2668 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_11
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 2300 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_14_25
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_21
timestamp 1586364061
transform 1 0 3036 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_35
timestamp 1586364061
transform 1 0 4324 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_29
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_34
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_31
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4324 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_41
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_44
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 4692 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_45
timestamp 1586364061
transform 1 0 5244 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_49
timestamp 1586364061
transform 1 0 5612 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 5428 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 5428 0 -1 10336
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_14_62
timestamp 1586364061
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_58
timestamp 1586364061
transform 1 0 6440 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6624 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_71
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7176 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_79
timestamp 1586364061
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_75
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_77
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__C
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_87
timestamp 1586364061
transform 1 0 9108 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_83
timestamp 1586364061
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_81
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__D
timestamp 1586364061
transform 1 0 8924 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__C
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_91
timestamp 1586364061
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_94
timestamp 1586364061
transform 1 0 9752 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_104
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_101
timestamp 1586364061
transform 1 0 10396 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_99
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_112
timestamp 1586364061
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_116
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_108
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_119
timestamp 1586364061
transform 1 0 12052 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_128
timestamp 1586364061
transform 1 0 12880 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12696 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_136
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 314 592
use scs8hd_or3_4  _096_
timestamp 1586364061
transform 1 0 13248 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use scs8hd_nor4_4  _127_
timestamp 1586364061
transform 1 0 14996 0 1 9248
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 14812 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__D
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_143
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_147
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_149
timestamp 1586364061
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 16284 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_168
timestamp 1586364061
transform 1 0 16560 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_13_173
timestamp 1586364061
transform 1 0 17020 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_167
timestamp 1586364061
transform 1 0 16468 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_174
timestamp 1586364061
transform 1 0 17112 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_195
timestamp 1586364061
transform 1 0 19044 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_191
timestamp 1586364061
transform 1 0 18676 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18860 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17848 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_205
timestamp 1586364061
transform 1 0 19964 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_201
timestamp 1586364061
transform 1 0 19596 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_204
timestamp 1586364061
transform 1 0 19872 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_201
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_197
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19688 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_213
timestamp 1586364061
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_209
timestamp 1586364061
transform 1 0 20332 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20332 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20516 0 1 9248
box -38 -48 866 592
use scs8hd_buf_2  _169_
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 21528 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_224
timestamp 1586364061
transform 1 0 21712 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_219
timestamp 1586364061
transform 1 0 21252 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_231
timestamp 1586364061
transform 1 0 22356 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 22816 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 22816 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 130 592
use scs8hd_buf_2  _168_
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 2300 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_11
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_25
timestamp 1586364061
transform 1 0 3404 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_30
timestamp 1586364061
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_34
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _104_
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5888 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_47
timestamp 1586364061
transform 1 0 5428 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7084 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 7544 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6256 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_54
timestamp 1586364061
transform 1 0 6072 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_58
timestamp 1586364061
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_68
timestamp 1586364061
transform 1 0 7360 0 1 10336
box -38 -48 222 592
use scs8hd_nor4_4  _129_
timestamp 1586364061
transform 1 0 8096 0 1 10336
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_72
timestamp 1586364061
transform 1 0 7728 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 10488 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_93
timestamp 1586364061
transform 1 0 9660 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_111
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_115
timestamp 1586364061
transform 1 0 11684 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 14168 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_141
timestamp 1586364061
transform 1 0 14076 0 1 10336
box -38 -48 130 592
use scs8hd_nor4_4  _128_
timestamp 1586364061
transform 1 0 15088 0 1 10336
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__128__D
timestamp 1586364061
transform 1 0 14904 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 14536 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_144
timestamp 1586364061
transform 1 0 14352 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_148
timestamp 1586364061
transform 1 0 14720 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_169
timestamp 1586364061
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_173
timestamp 1586364061
transform 1 0 17020 0 1 10336
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_195
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20148 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19964 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_199
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21528 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_216
timestamp 1586364061
transform 1 0 20976 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_224
timestamp 1586364061
transform 1 0 21712 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 22816 0 1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 130 592
use scs8hd_nor2_4  _109_
timestamp 1586364061
transform 1 0 1472 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_13
timestamp 1586364061
transform 1 0 2300 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_17
timestamp 1586364061
transform 1 0 2668 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__073__C
timestamp 1586364061
transform 1 0 4232 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2852 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_21
timestamp 1586364061
transform 1 0 3036 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_29
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _106_
timestamp 1586364061
transform 1 0 4692 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  FILLER_16_36
timestamp 1586364061
transform 1 0 4416 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_48
timestamp 1586364061
transform 1 0 5520 0 -1 11424
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__075__C
timestamp 1586364061
transform 1 0 7636 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_67
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 406 592
use scs8hd_or3_4  _088_
timestamp 1586364061
transform 1 0 8004 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__C
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_73
timestamp 1586364061
transform 1 0 7820 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_88
timestamp 1586364061
transform 1 0 9200 0 -1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10396 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 12144 0 -1 11424
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_16_112
timestamp 1586364061
transform 1 0 11408 0 -1 11424
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 13984 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 13616 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_131
timestamp 1586364061
transform 1 0 13156 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_135
timestamp 1586364061
transform 1 0 13524 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_138
timestamp 1586364061
transform 1 0 13800 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_142
timestamp 1586364061
transform 1 0 14168 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15640 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__128__C
timestamp 1586364061
transform 1 0 15456 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_146
timestamp 1586364061
transform 1 0 14536 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_152
timestamp 1586364061
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_169
timestamp 1586364061
transform 1 0 16652 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_181
timestamp 1586364061
transform 1 0 17756 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_189
timestamp 1586364061
transform 1 0 18492 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_8  _062_
timestamp 1586364061
transform 1 0 19228 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20240 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_210
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_224
timestamp 1586364061
transform 1 0 21712 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 22816 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_232
timestamp 1586364061
transform 1 0 22448 0 -1 11424
box -38 -48 130 592
use scs8hd_inv_8  _051_
timestamp 1586364061
transform 1 0 1564 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__085__C
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_14
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use scs8hd_or3_4  _073_
timestamp 1586364061
transform 1 0 3864 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 3680 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__B
timestamp 1586364061
transform 1 0 3312 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_18
timestamp 1586364061
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_22
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_26
timestamp 1586364061
transform 1 0 3496 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__052__A
timestamp 1586364061
transform 1 0 4876 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 5612 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_43
timestamp 1586364061
transform 1 0 5060 0 1 11424
box -38 -48 590 592
use scs8hd_fill_2  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use scs8hd_or3_4  _077_
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__077__C
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_55
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_71
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use scs8hd_nor4_4  _130_
timestamp 1586364061
transform 1 0 8740 0 1 11424
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__130__D
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__B
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_75
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_79
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10488 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_100
timestamp 1586364061
transform 1 0 10304 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_104
timestamp 1586364061
transform 1 0 10672 0 1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_108
timestamp 1586364061
transform 1 0 11040 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_132
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_138
timestamp 1586364061
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_149
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 590 592
use scs8hd_fill_2  FILLER_17_157
timestamp 1586364061
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_161
timestamp 1586364061
transform 1 0 15916 0 1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 406 592
use scs8hd_conb_1  _146_
timestamp 1586364061
transform 1 0 18952 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18216 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_181
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_188
timestamp 1586364061
transform 1 0 18400 0 1 11424
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19964 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 19688 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_197
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_201
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_204
timestamp 1586364061
transform 1 0 19872 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_214
timestamp 1586364061
transform 1 0 20792 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21528 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21988 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20976 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_218
timestamp 1586364061
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_225
timestamp 1586364061
transform 1 0 21804 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_229
timestamp 1586364061
transform 1 0 22172 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 22816 0 1 11424
box -38 -48 314 592
use scs8hd_or3_4  _085_
timestamp 1586364061
transform 1 0 1748 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__051__A
timestamp 1586364061
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_16
timestamp 1586364061
transform 1 0 2576 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_8  _052_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 2760 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_20
timestamp 1586364061
transform 1 0 2944 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_28
timestamp 1586364061
transform 1 0 3680 0 -1 12512
box -38 -48 130 592
use scs8hd_nor2_4  _082_
timestamp 1586364061
transform 1 0 5612 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_18_41
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 774 592
use scs8hd_or3_4  _075_
timestamp 1586364061
transform 1 0 7636 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__B
timestamp 1586364061
transform 1 0 7176 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_58
timestamp 1586364061
transform 1 0 6440 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_64
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_85
timestamp 1586364061
transform 1 0 8924 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_89
timestamp 1586364061
transform 1 0 9292 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10120 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_97
timestamp 1586364061
transform 1 0 10028 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_101
timestamp 1586364061
transform 1 0 10396 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_6  FILLER_18_107
timestamp 1586364061
transform 1 0 10948 0 -1 12512
box -38 -48 590 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 11592 0 -1 12512
box -38 -48 866 592
use scs8hd_fill_1  FILLER_18_113
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_123
timestamp 1586364061
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _113_
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_127
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_131
timestamp 1586364061
transform 1 0 13156 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_135
timestamp 1586364061
transform 1 0 13524 0 -1 12512
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15364 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16560 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16928 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_170
timestamp 1586364061
transform 1 0 16744 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_174
timestamp 1586364061
transform 1 0 17112 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 17572 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18768 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_194
timestamp 1586364061
transform 1 0 18952 0 -1 12512
box -38 -48 774 592
use scs8hd_buf_2  _167_
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_210
timestamp 1586364061
transform 1 0 20424 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_18_224
timestamp 1586364061
transform 1 0 21712 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 22816 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_232
timestamp 1586364061
transform 1 0 22448 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_17
timestamp 1586364061
transform 1 0 2668 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_13
timestamp 1586364061
transform 1 0 2300 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__B
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__C
timestamp 1586364061
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _086_
timestamp 1586364061
transform 1 0 1472 0 -1 13600
box -38 -48 866 592
use scs8hd_or3_4  _081_
timestamp 1586364061
transform 1 0 1656 0 1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_20_21
timestamp 1586364061
transform 1 0 3036 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_4  FILLER_19_23
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_19
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 2852 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__C
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_or3_4  _083_
timestamp 1586364061
transform 1 0 3772 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _078_
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_8  FILLER_20_41
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_42
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_38
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_49
timestamp 1586364061
transform 1 0 5612 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_52
timestamp 1586364061
transform 1 0 5888 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_46
timestamp 1586364061
transform 1 0 5336 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5704 0 -1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 1 12512
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 5888 0 -1 13600
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_19_60
timestamp 1586364061
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_56
timestamp 1586364061
transform 1 0 6256 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6440 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6072 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_71
timestamp 1586364061
transform 1 0 7636 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_67
timestamp 1586364061
transform 1 0 7268 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_63
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_20_78
timestamp 1586364061
transform 1 0 8280 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_74
timestamp 1586364061
transform 1 0 7912 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_79
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_75
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 8096 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 7728 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_88
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_83
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__094__B
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 13600
box -38 -48 314 592
use scs8hd_nor2_4  _094_
timestamp 1586364061
transform 1 0 8832 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_97
timestamp 1586364061
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_93
timestamp 1586364061
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_104
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_101
timestamp 1586364061
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_20_112
timestamp 1586364061
transform 1 0 11408 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_108
timestamp 1586364061
transform 1 0 11040 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_122
timestamp 1586364061
transform 1 0 12328 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11500 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_3  FILLER_20_130
timestamp 1586364061
transform 1 0 13064 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_130
timestamp 1586364061
transform 1 0 13064 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_126
timestamp 1586364061
transform 1 0 12696 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 13340 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 13340 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_139
timestamp 1586364061
transform 1 0 13892 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_135
timestamp 1586364061
transform 1 0 13524 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_151
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_143
timestamp 1586364061
transform 1 0 14260 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_148
timestamp 1586364061
transform 1 0 14720 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_144
timestamp 1586364061
transform 1 0 14352 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14536 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 14904 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15640 0 -1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 15088 0 1 12512
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_20_168
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_165
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_161
timestamp 1586364061
transform 1 0 15916 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_167
timestamp 1586364061
transform 1 0 16468 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_163
timestamp 1586364061
transform 1 0 16100 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16652 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16284 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_178
timestamp 1586364061
transform 1 0 17480 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_3  FILLER_19_178
timestamp 1586364061
transform 1 0 17480 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_174
timestamp 1586364061
transform 1 0 17112 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17296 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16652 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_193
timestamp 1586364061
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_186
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_202
timestamp 1586364061
transform 1 0 19688 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_198
timestamp 1586364061
transform 1 0 19320 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_197
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19872 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19504 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_19_214
timestamp 1586364061
transform 1 0 20792 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_210
timestamp 1586364061
transform 1 0 20424 0 1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_222
timestamp 1586364061
transform 1 0 21528 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_217
timestamp 1586364061
transform 1 0 21068 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 12512
box -38 -48 222 592
use scs8hd_buf_2  _166_
timestamp 1586364061
transform 1 0 21160 0 1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_224
timestamp 1586364061
transform 1 0 21712 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  FILLER_19_230
timestamp 1586364061
transform 1 0 22264 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_226
timestamp 1586364061
transform 1 0 21896 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 21712 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 22816 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 22816 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_232
timestamp 1586364061
transform 1 0 22448 0 -1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1840 0 1 13600
box -38 -48 1050 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 1656 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3956 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 3772 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 3036 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 3404 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_19
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_23
timestamp 1586364061
transform 1 0 3220 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5520 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5336 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_40
timestamp 1586364061
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_44
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_55
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_65
timestamp 1586364061
transform 1 0 7084 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_69
timestamp 1586364061
transform 1 0 7452 0 1 13600
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9200 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_86
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_90
timestamp 1586364061
transform 1 0 9384 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_94
timestamp 1586364061
transform 1 0 9752 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_97
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 14076 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 13892 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_132
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_136
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_152
timestamp 1586364061
transform 1 0 15088 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_156
timestamp 1586364061
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_160
timestamp 1586364061
transform 1 0 15824 0 1 13600
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18308 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18768 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_190
timestamp 1586364061
transform 1 0 18584 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_194
timestamp 1586364061
transform 1 0 18952 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19320 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20332 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_207
timestamp 1586364061
transform 1 0 20148 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_211
timestamp 1586364061
transform 1 0 20516 0 1 13600
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_218
timestamp 1586364061
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_222
timestamp 1586364061
transform 1 0 21528 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  FILLER_21_230
timestamp 1586364061
transform 1 0 22264 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 22816 0 1 13600
box -38 -48 314 592
use scs8hd_nor2_4  _080_
timestamp 1586364061
transform 1 0 1656 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2668 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_19
timestamp 1586364061
transform 1 0 2852 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_43
timestamp 1586364061
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_47
timestamp 1586364061
transform 1 0 5428 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_51
timestamp 1586364061
transform 1 0 5796 0 -1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6072 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_63
timestamp 1586364061
transform 1 0 6900 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_67
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_71
timestamp 1586364061
transform 1 0 7636 0 -1 14688
box -38 -48 130 592
use scs8hd_nor2_4  _093_
timestamp 1586364061
transform 1 0 7728 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_81
timestamp 1586364061
transform 1 0 8556 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  FILLER_22_89
timestamp 1586364061
transform 1 0 9292 0 -1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 9844 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10212 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_97
timestamp 1586364061
transform 1 0 10028 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_101
timestamp 1586364061
transform 1 0 10396 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_113
timestamp 1586364061
transform 1 0 11500 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_121
timestamp 1586364061
transform 1 0 12236 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _115_
timestamp 1586364061
transform 1 0 13340 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_125
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_142
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 14352 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 14720 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_146
timestamp 1586364061
transform 1 0 14536 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_150
timestamp 1586364061
transform 1 0 14904 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_165
timestamp 1586364061
transform 1 0 16284 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_169
timestamp 1586364061
transform 1 0 16652 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_172
timestamp 1586364061
transform 1 0 16928 0 -1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19136 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_12  FILLER_22_182
timestamp 1586364061
transform 1 0 17848 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_22_194
timestamp 1586364061
transform 1 0 18952 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_205
timestamp 1586364061
transform 1 0 19964 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_213
timestamp 1586364061
transform 1 0 20700 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 590 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 22816 0 -1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 1050 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 1564 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2944 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4324 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3956 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_18
timestamp 1586364061
transform 1 0 2760 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_22
timestamp 1586364061
transform 1 0 3128 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_26
timestamp 1586364061
transform 1 0 3496 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_30
timestamp 1586364061
transform 1 0 3864 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_33
timestamp 1586364061
transform 1 0 4140 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4508 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5520 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_46
timestamp 1586364061
transform 1 0 5336 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_50
timestamp 1586364061
transform 1 0 5704 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_55
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_71
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _091_
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_75
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_88
timestamp 1586364061
transform 1 0 9200 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9936 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 9752 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 9384 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_92
timestamp 1586364061
transform 1 0 9568 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_107
timestamp 1586364061
transform 1 0 10948 0 1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_111
timestamp 1586364061
transform 1 0 11316 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 13984 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_138
timestamp 1586364061
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 14996 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_149
timestamp 1586364061
transform 1 0 14812 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_153
timestamp 1586364061
transform 1 0 15180 0 1 14688
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17296 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_161
timestamp 1586364061
transform 1 0 15916 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_174
timestamp 1586364061
transform 1 0 17112 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_178
timestamp 1586364061
transform 1 0 17480 0 1 14688
box -38 -48 406 592
use scs8hd_conb_1  _141_
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18308 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_182
timestamp 1586364061
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use scs8hd_decap_6  FILLER_23_189
timestamp 1586364061
transform 1 0 18492 0 1 14688
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_198
timestamp 1586364061
transform 1 0 19320 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_202
timestamp 1586364061
transform 1 0 19688 0 1 14688
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_23_214
timestamp 1586364061
transform 1 0 20792 0 1 14688
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_218
timestamp 1586364061
transform 1 0 21160 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_222
timestamp 1586364061
transform 1 0 21528 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  FILLER_23_230
timestamp 1586364061
transform 1 0 22264 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 22816 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1840 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_6
timestamp 1586364061
transform 1 0 1656 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_10
timestamp 1586364061
transform 1 0 2024 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4508 0 -1 15776
box -38 -48 866 592
use scs8hd_fill_1  FILLER_24_36
timestamp 1586364061
transform 1 0 4416 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_46
timestamp 1586364061
transform 1 0 5336 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6348 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  FILLER_24_54
timestamp 1586364061
transform 1 0 6072 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_66
timestamp 1586364061
transform 1 0 7176 0 -1 15776
box -38 -48 774 592
use scs8hd_conb_1  _149_
timestamp 1586364061
transform 1 0 7912 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 8372 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_77
timestamp 1586364061
transform 1 0 8188 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_81
timestamp 1586364061
transform 1 0 8556 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_85
timestamp 1586364061
transform 1 0 8924 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_88
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _090_
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_106
timestamp 1586364061
transform 1 0 10856 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_110
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_121
timestamp 1586364061
transform 1 0 12236 0 -1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _098_
timestamp 1586364061
transform 1 0 13616 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_125
timestamp 1586364061
transform 1 0 12604 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_24_133
timestamp 1586364061
transform 1 0 13340 0 -1 15776
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15732 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_149
timestamp 1586364061
transform 1 0 14812 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_4  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_158
timestamp 1586364061
transform 1 0 15640 0 -1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16744 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16192 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16560 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_162
timestamp 1586364061
transform 1 0 16008 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_166
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18308 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18768 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_179
timestamp 1586364061
transform 1 0 17572 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_183
timestamp 1586364061
transform 1 0 17940 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_190
timestamp 1586364061
transform 1 0 18584 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_194
timestamp 1586364061
transform 1 0 18952 0 -1 15776
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19320 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_201
timestamp 1586364061
transform 1 0 19596 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_205
timestamp 1586364061
transform 1 0 19964 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_6  FILLER_24_208
timestamp 1586364061
transform 1 0 20240 0 -1 15776
box -38 -48 590 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 590 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 22816 0 -1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _076_
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 866 592
use scs8hd_buf_2  _178_
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_7
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_11
timestamp 1586364061
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4048 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 3496 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_24
timestamp 1586364061
transform 1 0 3312 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_28
timestamp 1586364061
transform 1 0 3680 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 5428 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_43
timestamp 1586364061
transform 1 0 5060 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_49
timestamp 1586364061
transform 1 0 5612 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_71
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _089_
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 8832 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_75
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_79
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_83
timestamp 1586364061
transform 1 0 8740 0 1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 10028 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_95
timestamp 1586364061
transform 1 0 9844 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_99
timestamp 1586364061
transform 1 0 10212 0 1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 774 592
use scs8hd_nor2_4  _097_
timestamp 1586364061
transform 1 0 14168 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 13984 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_131
timestamp 1586364061
transform 1 0 13156 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_134
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_138
timestamp 1586364061
transform 1 0 13800 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_151
timestamp 1586364061
transform 1 0 14996 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_156
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_160
timestamp 1586364061
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 16192 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18308 0 1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_179
timestamp 1586364061
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20056 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19872 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19504 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_198
timestamp 1586364061
transform 1 0 19320 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_202
timestamp 1586364061
transform 1 0 19688 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 21068 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_215
timestamp 1586364061
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_219
timestamp 1586364061
transform 1 0 21252 0 1 15776
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_25_231
timestamp 1586364061
transform 1 0 22356 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 22816 0 1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 1 16864
box -38 -48 866 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2024 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_17
timestamp 1586364061
transform 1 0 2668 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_27_9
timestamp 1586364061
transform 1 0 1932 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_25
timestamp 1586364061
transform 1 0 3404 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_21
timestamp 1586364061
transform 1 0 3036 0 1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3496 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_28
timestamp 1586364061
transform 1 0 3680 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_29
timestamp 1586364061
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3864 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_35
timestamp 1586364061
transform 1 0 4324 0 -1 16864
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5428 0 -1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 5060 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 5428 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_41
timestamp 1586364061
transform 1 0 4876 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_45
timestamp 1586364061
transform 1 0 5244 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_49
timestamp 1586364061
transform 1 0 5612 0 1 16864
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_58
timestamp 1586364061
transform 1 0 6440 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_8  FILLER_26_64
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_71
timestamp 1586364061
transform 1 0 7636 0 1 16864
box -38 -48 590 592
use scs8hd_nor2_4  _092_
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_72
timestamp 1586364061
transform 1 0 7728 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_8  FILLER_27_88
timestamp 1586364061
transform 1 0 9200 0 1 16864
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9936 0 -1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 10304 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_26_107
timestamp 1586364061
transform 1 0 10948 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_102
timestamp 1586364061
transform 1 0 10488 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11684 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_124
timestamp 1586364061
transform 1 0 12512 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_113
timestamp 1586364061
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_117
timestamp 1586364061
transform 1 0 11868 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_121
timestamp 1586364061
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use scs8hd_nor2_4  _099_
timestamp 1586364061
transform 1 0 13616 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _100_
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 12880 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 13432 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_132
timestamp 1586364061
transform 1 0 13248 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_126
timestamp 1586364061
transform 1 0 12696 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_130
timestamp 1586364061
transform 1 0 13064 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15272 0 1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15088 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14720 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_4  FILLER_27_143
timestamp 1586364061
transform 1 0 14260 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_147
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_150
timestamp 1586364061
transform 1 0 14904 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 16928 0 -1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16744 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_163
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_26_171
timestamp 1586364061
transform 1 0 16836 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_165
timestamp 1586364061
transform 1 0 16284 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_169
timestamp 1586364061
transform 1 0 16652 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_172
timestamp 1586364061
transform 1 0 16928 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_176
timestamp 1586364061
transform 1 0 17296 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_180
timestamp 1586364061
transform 1 0 17664 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_183
timestamp 1586364061
transform 1 0 17940 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 18308 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_195
timestamp 1586364061
transform 1 0 19044 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_189
timestamp 1586364061
transform 1 0 18492 0 -1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19596 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_200
timestamp 1586364061
transform 1 0 19504 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_26_212
timestamp 1586364061
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_199
timestamp 1586364061
transform 1 0 19412 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_203
timestamp 1586364061
transform 1 0 19780 0 1 16864
box -38 -48 1142 592
use scs8hd_buf_2  _177_
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 21712 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_219
timestamp 1586364061
transform 1 0 21252 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_26_231
timestamp 1586364061
transform 1 0 22356 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_218
timestamp 1586364061
transform 1 0 21160 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_222
timestamp 1586364061
transform 1 0 21528 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_226
timestamp 1586364061
transform 1 0 21896 0 1 16864
box -38 -48 590 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 22816 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 22816 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_232
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 130 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_28_11
timestamp 1586364061
transform 1 0 2116 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_14
timestamp 1586364061
transform 1 0 2392 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_26
timestamp 1586364061
transform 1 0 3496 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_30
timestamp 1586364061
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 774 592
use scs8hd_nor2_4  _084_
timestamp 1586364061
transform 1 0 4876 0 -1 17952
box -38 -48 866 592
use scs8hd_fill_1  FILLER_28_40
timestamp 1586364061
transform 1 0 4784 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_50
timestamp 1586364061
transform 1 0 5704 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6532 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_58
timestamp 1586364061
transform 1 0 6440 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_62
timestamp 1586364061
transform 1 0 6808 0 -1 17952
box -38 -48 1142 592
use scs8hd_conb_1  _151_
timestamp 1586364061
transform 1 0 8556 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__092__B
timestamp 1586364061
transform 1 0 8372 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_74
timestamp 1586364061
transform 1 0 7912 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_78
timestamp 1586364061
transform 1 0 8280 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_84
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 774 592
use scs8hd_buf_2  _175_
timestamp 1586364061
transform 1 0 10304 0 -1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_97
timestamp 1586364061
transform 1 0 10028 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_104
timestamp 1586364061
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11500 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12512 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_108
timestamp 1586364061
transform 1 0 11040 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_112
timestamp 1586364061
transform 1 0 11408 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_122
timestamp 1586364061
transform 1 0 12328 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _102_
timestamp 1586364061
transform 1 0 13616 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 13432 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_126
timestamp 1586364061
transform 1 0 12696 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15732 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_149
timestamp 1586364061
transform 1 0 14812 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_157
timestamp 1586364061
transform 1 0 15548 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16744 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_161
timestamp 1586364061
transform 1 0 15916 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_28_169
timestamp 1586364061
transform 1 0 16652 0 -1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18860 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18216 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_179
timestamp 1586364061
transform 1 0 17572 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_185
timestamp 1586364061
transform 1 0 18124 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_188
timestamp 1586364061
transform 1 0 18400 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_192
timestamp 1586364061
transform 1 0 18768 0 -1 17952
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19872 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_202
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_206
timestamp 1586364061
transform 1 0 20056 0 -1 17952
box -38 -48 774 592
use scs8hd_buf_2  _174_
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_219
timestamp 1586364061
transform 1 0 21252 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_28_231
timestamp 1586364061
transform 1 0 22356 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 22816 0 -1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_6
timestamp 1586364061
transform 1 0 1656 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_10
timestamp 1586364061
transform 1 0 2024 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_14
timestamp 1586364061
transform 1 0 2392 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_26
timestamp 1586364061
transform 1 0 3496 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_38
timestamp 1586364061
transform 1 0 4600 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_50
timestamp 1586364061
transform 1 0 5704 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_58
timestamp 1586364061
transform 1 0 6440 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_29_70
timestamp 1586364061
transform 1 0 7544 0 1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8188 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9200 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_73
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9568 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_90
timestamp 1586364061
transform 1 0 9384 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_103
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_107
timestamp 1586364061
transform 1 0 10948 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14076 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 13708 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_126
timestamp 1586364061
transform 1 0 12696 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_130
timestamp 1586364061
transform 1 0 13064 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_134
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_139
timestamp 1586364061
transform 1 0 13892 0 1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 14260 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15456 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15824 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_154
timestamp 1586364061
transform 1 0 15272 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_158
timestamp 1586364061
transform 1 0 15640 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16468 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16928 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17296 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_162
timestamp 1586364061
transform 1 0 16008 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_166
timestamp 1586364061
transform 1 0 16376 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_170
timestamp 1586364061
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_174
timestamp 1586364061
transform 1 0 17112 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_178
timestamp 1586364061
transform 1 0 17480 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18400 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18216 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17664 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_182
timestamp 1586364061
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_191
timestamp 1586364061
transform 1 0 18676 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_195
timestamp 1586364061
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19412 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 774 592
use scs8hd_buf_2  _171_
timestamp 1586364061
transform 1 0 20976 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 21528 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_224
timestamp 1586364061
transform 1 0 21712 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 22816 0 1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_6
timestamp 1586364061
transform 1 0 1656 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_18
timestamp 1586364061
transform 1 0 2760 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_30_30
timestamp 1586364061
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_82
timestamp 1586364061
transform 1 0 8648 0 -1 19040
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9752 0 -1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_90
timestamp 1586364061
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11500 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_8  FILLER_30_122
timestamp 1586364061
transform 1 0 12328 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13064 0 -1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13524 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_133
timestamp 1586364061
transform 1 0 13340 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_137
timestamp 1586364061
transform 1 0 13708 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_145
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_165
timestamp 1586364061
transform 1 0 16284 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_169
timestamp 1586364061
transform 1 0 16652 0 -1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_8  FILLER_30_182
timestamp 1586364061
transform 1 0 17848 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_200
timestamp 1586364061
transform 1 0 19504 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_204
timestamp 1586364061
transform 1 0 19872 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_212
timestamp 1586364061
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 590 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 22816 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_7
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_19
timestamp 1586364061
transform 1 0 2852 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_31
timestamp 1586364061
transform 1 0 3956 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_43
timestamp 1586364061
transform 1 0 5060 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_55
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 590 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8464 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8280 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_76
timestamp 1586364061
transform 1 0 8096 0 1 19040
box -38 -48 222 592
use scs8hd_inv_8  _064_
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_91
timestamp 1586364061
transform 1 0 9476 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_95
timestamp 1586364061
transform 1 0 9844 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_99
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14076 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_126
timestamp 1586364061
transform 1 0 12696 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_130
timestamp 1586364061
transform 1 0 13064 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_134
timestamp 1586364061
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_139
timestamp 1586364061
transform 1 0 13892 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15364 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15180 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_143
timestamp 1586364061
transform 1 0 14260 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_151
timestamp 1586364061
transform 1 0 14996 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_158
timestamp 1586364061
transform 1 0 15640 0 1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15916 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_163
timestamp 1586364061
transform 1 0 16100 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_175
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use scs8hd_conb_1  _150_
timestamp 1586364061
transform 1 0 18492 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18952 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18308 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_179
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_192
timestamp 1586364061
transform 1 0 18768 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19504 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19320 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20516 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_209
timestamp 1586364061
transform 1 0 20332 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_213
timestamp 1586364061
transform 1 0 20700 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21068 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21528 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_224
timestamp 1586364061
transform 1 0 21712 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 22816 0 1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_6
timestamp 1586364061
transform 1 0 1656 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_18
timestamp 1586364061
transform 1 0 2760 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_32_30
timestamp 1586364061
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 590 592
use scs8hd_inv_8  _063_
timestamp 1586364061
transform 1 0 8004 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9292 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_74
timestamp 1586364061
transform 1 0 7912 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_84
timestamp 1586364061
transform 1 0 8832 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_88
timestamp 1586364061
transform 1 0 9200 0 -1 20128
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_91
timestamp 1586364061
transform 1 0 9476 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_102
timestamp 1586364061
transform 1 0 10488 0 -1 20128
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11500 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12512 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_110
timestamp 1586364061
transform 1 0 11224 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_122
timestamp 1586364061
transform 1 0 12328 0 -1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_4  FILLER_32_126
timestamp 1586364061
transform 1 0 12696 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_139
timestamp 1586364061
transform 1 0 13892 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_151
timestamp 1586364061
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_160
timestamp 1586364061
transform 1 0 15824 0 -1 20128
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15916 0 -1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17112 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_164
timestamp 1586364061
transform 1 0 16192 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_168
timestamp 1586364061
transform 1 0 16560 0 -1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_32_183
timestamp 1586364061
transform 1 0 17940 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_32_195
timestamp 1586364061
transform 1 0 19044 0 -1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_206
timestamp 1586364061
transform 1 0 20056 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_218
timestamp 1586364061
transform 1 0 21160 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_32_230
timestamp 1586364061
transform 1 0 22264 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 22816 0 -1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2116 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2576 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_14
timestamp 1586364061
transform 1 0 2392 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_18
timestamp 1586364061
transform 1 0 2760 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_33_30
timestamp 1586364061
transform 1 0 3864 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_35
timestamp 1586364061
transform 1 0 4324 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4508 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_70
timestamp 1586364061
transform 1 0 7544 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  FILLER_34_76
timestamp 1586364061
transform 1 0 8096 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_6  FILLER_33_80
timestamp 1586364061
transform 1 0 8464 0 1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_76
timestamp 1586364061
transform 1 0 8096 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 8280 0 1 20128
box -38 -48 222 592
use scs8hd_buf_2  _157_
timestamp 1586364061
transform 1 0 7728 0 1 20128
box -38 -48 406 592
use scs8hd_buf_2  _152_
timestamp 1586364061
transform 1 0 8372 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_8  FILLER_34_83
timestamp 1586364061
transform 1 0 8740 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_1  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9292 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_91
timestamp 1586364061
transform 1 0 9476 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_33_114
timestamp 1586364061
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 130 592
use scs8hd_conb_1  _147_
timestamp 1586364061
transform 1 0 11316 0 1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_34_121
timestamp 1586364061
transform 1 0 12236 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_118
timestamp 1586364061
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_buf_2  _162_
timestamp 1586364061
transform 1 0 12328 0 -1 21216
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 866 592
use scs8hd_buf_2  _161_
timestamp 1586364061
transform 1 0 13984 0 1 20128
box -38 -48 406 592
use scs8hd_decap_8  FILLER_33_132
timestamp 1586364061
transform 1 0 13248 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_126
timestamp 1586364061
transform 1 0 12696 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_138
timestamp 1586364061
transform 1 0 13800 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 14536 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_144
timestamp 1586364061
transform 1 0 14352 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_148
timestamp 1586364061
transform 1 0 14720 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_160
timestamp 1586364061
transform 1 0 15824 0 1 20128
box -38 -48 774 592
use scs8hd_decap_3  FILLER_34_150
timestamp 1586364061
transform 1 0 14904 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16652 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17112 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_168
timestamp 1586364061
transform 1 0 16560 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_172
timestamp 1586364061
transform 1 0 16928 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_176
timestamp 1586364061
transform 1 0 17296 0 1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 590 592
use scs8hd_buf_2  _173_
timestamp 1586364061
transform 1 0 18952 0 1 20128
box -38 -48 406 592
use scs8hd_buf_2  _176_
timestamp 1586364061
transform 1 0 18032 0 -1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 18216 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_182
timestamp 1586364061
transform 1 0 17848 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_188
timestamp 1586364061
transform 1 0 18400 0 1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_34_188
timestamp 1586364061
transform 1 0 18400 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_34_200
timestamp 1586364061
transform 1 0 19504 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_202
timestamp 1586364061
transform 1 0 19688 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_198
timestamp 1586364061
transform 1 0 19320 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19872 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 19504 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_34_206
timestamp 1586364061
transform 1 0 20056 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_8  FILLER_33_206
timestamp 1586364061
transform 1 0 20056 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_33_214
timestamp 1586364061
transform 1 0 20792 0 1 20128
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_buf_2  _172_
timestamp 1586364061
transform 1 0 20884 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 21436 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_219
timestamp 1586364061
transform 1 0 21252 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_223
timestamp 1586364061
transform 1 0 21620 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_231
timestamp 1586364061
transform 1 0 22356 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 590 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 22816 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 22816 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_35_32
timestamp 1586364061
transform 1 0 4048 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_44
timestamp 1586364061
transform 1 0 5152 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_56
timestamp 1586364061
transform 1 0 6256 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_63
timestamp 1586364061
transform 1 0 6900 0 1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8464 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8924 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_75
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_79
timestamp 1586364061
transform 1 0 8372 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_83
timestamp 1586364061
transform 1 0 8740 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_87
timestamp 1586364061
transform 1 0 9108 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_94
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_106
timestamp 1586364061
transform 1 0 10856 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_125
timestamp 1586364061
transform 1 0 12604 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_137
timestamp 1586364061
transform 1 0 13708 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_149
timestamp 1586364061
transform 1 0 14812 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_156
timestamp 1586364061
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_168
timestamp 1586364061
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_180
timestamp 1586364061
transform 1 0 17664 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_187
timestamp 1586364061
transform 1 0 18308 0 1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19504 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19964 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_199
timestamp 1586364061
transform 1 0 19412 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_203
timestamp 1586364061
transform 1 0 19780 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_207
timestamp 1586364061
transform 1 0 20148 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_215
timestamp 1586364061
transform 1 0 20884 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_218
timestamp 1586364061
transform 1 0 21160 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_35_230
timestamp 1586364061
transform 1 0 22264 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 22816 0 1 21216
box -38 -48 314 592
<< labels >>
rlabel metal2 s 2318 0 2374 480 6 address[0]
port 0 nsew default input
rlabel metal3 s 23520 416 24000 536 6 address[1]
port 1 nsew default input
rlabel metal2 s 570 23520 626 24000 6 address[2]
port 2 nsew default input
rlabel metal2 s 1766 23520 1822 24000 6 address[3]
port 3 nsew default input
rlabel metal3 s 23520 1368 24000 1488 6 address[4]
port 4 nsew default input
rlabel metal2 s 3238 0 3294 480 6 address[5]
port 5 nsew default input
rlabel metal3 s 23520 2320 24000 2440 6 address[6]
port 6 nsew default input
rlabel metal3 s 23520 6400 24000 6520 6 bottom_left_grid_pin_11_
port 7 nsew default input
rlabel metal2 s 4342 23520 4398 24000 6 bottom_left_grid_pin_13_
port 8 nsew default input
rlabel metal2 s 4158 0 4214 480 6 bottom_left_grid_pin_15_
port 9 nsew default input
rlabel metal3 s 23520 3408 24000 3528 6 bottom_left_grid_pin_1_
port 10 nsew default input
rlabel metal3 s 0 824 480 944 6 bottom_left_grid_pin_3_
port 11 nsew default input
rlabel metal2 s 3054 23520 3110 24000 6 bottom_left_grid_pin_5_
port 12 nsew default input
rlabel metal3 s 23520 4360 24000 4480 6 bottom_left_grid_pin_7_
port 13 nsew default input
rlabel metal3 s 23520 5312 24000 5432 6 bottom_left_grid_pin_9_
port 14 nsew default input
rlabel metal2 s 5078 0 5134 480 6 bottom_right_grid_pin_11_
port 15 nsew default input
rlabel metal2 s 5538 23520 5594 24000 6 chanx_right_in[0]
port 16 nsew default input
rlabel metal2 s 5998 0 6054 480 6 chanx_right_in[1]
port 17 nsew default input
rlabel metal3 s 0 2456 480 2576 6 chanx_right_in[2]
port 18 nsew default input
rlabel metal3 s 0 4224 480 4344 6 chanx_right_in[3]
port 19 nsew default input
rlabel metal2 s 6918 0 6974 480 6 chanx_right_in[4]
port 20 nsew default input
rlabel metal3 s 23520 7352 24000 7472 6 chanx_right_in[5]
port 21 nsew default input
rlabel metal2 s 6826 23520 6882 24000 6 chanx_right_in[6]
port 22 nsew default input
rlabel metal2 s 7838 0 7894 480 6 chanx_right_in[7]
port 23 nsew default input
rlabel metal2 s 8758 0 8814 480 6 chanx_right_in[8]
port 24 nsew default input
rlabel metal3 s 0 5856 480 5976 6 chanx_right_out[0]
port 25 nsew default tristate
rlabel metal3 s 23520 8304 24000 8424 6 chanx_right_out[1]
port 26 nsew default tristate
rlabel metal3 s 0 7624 480 7744 6 chanx_right_out[2]
port 27 nsew default tristate
rlabel metal2 s 8114 23520 8170 24000 6 chanx_right_out[3]
port 28 nsew default tristate
rlabel metal2 s 9678 0 9734 480 6 chanx_right_out[4]
port 29 nsew default tristate
rlabel metal2 s 10598 0 10654 480 6 chanx_right_out[5]
port 30 nsew default tristate
rlabel metal2 s 11518 0 11574 480 6 chanx_right_out[6]
port 31 nsew default tristate
rlabel metal3 s 0 9256 480 9376 6 chanx_right_out[7]
port 32 nsew default tristate
rlabel metal2 s 9402 23520 9458 24000 6 chanx_right_out[8]
port 33 nsew default tristate
rlabel metal2 s 10598 23520 10654 24000 6 chany_bottom_in[0]
port 34 nsew default input
rlabel metal3 s 0 11024 480 11144 6 chany_bottom_in[1]
port 35 nsew default input
rlabel metal2 s 11886 23520 11942 24000 6 chany_bottom_in[2]
port 36 nsew default input
rlabel metal2 s 12438 0 12494 480 6 chany_bottom_in[3]
port 37 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[4]
port 38 nsew default input
rlabel metal3 s 23520 9392 24000 9512 6 chany_bottom_in[5]
port 39 nsew default input
rlabel metal2 s 14278 0 14334 480 6 chany_bottom_in[6]
port 40 nsew default input
rlabel metal3 s 23520 10344 24000 10464 6 chany_bottom_in[7]
port 41 nsew default input
rlabel metal2 s 15198 0 15254 480 6 chany_bottom_in[8]
port 42 nsew default input
rlabel metal3 s 23520 11296 24000 11416 6 chany_bottom_out[0]
port 43 nsew default tristate
rlabel metal3 s 0 12792 480 12912 6 chany_bottom_out[1]
port 44 nsew default tristate
rlabel metal3 s 23520 12384 24000 12504 6 chany_bottom_out[2]
port 45 nsew default tristate
rlabel metal3 s 23520 13336 24000 13456 6 chany_bottom_out[3]
port 46 nsew default tristate
rlabel metal2 s 16118 0 16174 480 6 chany_bottom_out[4]
port 47 nsew default tristate
rlabel metal2 s 17038 0 17094 480 6 chany_bottom_out[5]
port 48 nsew default tristate
rlabel metal2 s 17958 0 18014 480 6 chany_bottom_out[6]
port 49 nsew default tristate
rlabel metal2 s 13174 23520 13230 24000 6 chany_bottom_out[7]
port 50 nsew default tristate
rlabel metal2 s 14462 23520 14518 24000 6 chany_bottom_out[8]
port 51 nsew default tristate
rlabel metal3 s 23520 14288 24000 14408 6 chany_top_in[0]
port 52 nsew default input
rlabel metal2 s 15658 23520 15714 24000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal3 s 0 14424 480 14544 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 18878 0 18934 480 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 16946 23520 17002 24000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 19798 0 19854 480 6 chany_top_in[5]
port 57 nsew default input
rlabel metal3 s 23520 15376 24000 15496 6 chany_top_in[6]
port 58 nsew default input
rlabel metal3 s 23520 16328 24000 16448 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 18234 23520 18290 24000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal3 s 0 16192 480 16312 6 chany_top_out[0]
port 61 nsew default tristate
rlabel metal3 s 23520 17280 24000 17400 6 chany_top_out[1]
port 62 nsew default tristate
rlabel metal2 s 19522 23520 19578 24000 6 chany_top_out[2]
port 63 nsew default tristate
rlabel metal3 s 0 17824 480 17944 6 chany_top_out[3]
port 64 nsew default tristate
rlabel metal3 s 23520 18368 24000 18488 6 chany_top_out[4]
port 65 nsew default tristate
rlabel metal2 s 20718 23520 20774 24000 6 chany_top_out[5]
port 66 nsew default tristate
rlabel metal2 s 22006 23520 22062 24000 6 chany_top_out[6]
port 67 nsew default tristate
rlabel metal3 s 23520 19320 24000 19440 6 chany_top_out[7]
port 68 nsew default tristate
rlabel metal2 s 20718 0 20774 480 6 chany_top_out[8]
port 69 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 data_in
port 70 nsew default input
rlabel metal2 s 478 0 534 480 6 enable
port 71 nsew default input
rlabel metal2 s 23294 23520 23350 24000 6 right_bottom_grid_pin_12_
port 72 nsew default input
rlabel metal2 s 21638 0 21694 480 6 right_top_grid_pin_10_
port 73 nsew default input
rlabel metal3 s 23520 22312 24000 22432 6 top_left_grid_pin_11_
port 74 nsew default input
rlabel metal2 s 23478 0 23534 480 6 top_left_grid_pin_13_
port 75 nsew default input
rlabel metal3 s 0 22992 480 23112 6 top_left_grid_pin_15_
port 76 nsew default input
rlabel metal3 s 0 19592 480 19712 6 top_left_grid_pin_1_
port 77 nsew default input
rlabel metal2 s 22558 0 22614 480 6 top_left_grid_pin_3_
port 78 nsew default input
rlabel metal3 s 23520 20272 24000 20392 6 top_left_grid_pin_5_
port 79 nsew default input
rlabel metal3 s 23520 21360 24000 21480 6 top_left_grid_pin_7_
port 80 nsew default input
rlabel metal3 s 0 21224 480 21344 6 top_left_grid_pin_9_
port 81 nsew default input
rlabel metal3 s 23520 23264 24000 23384 6 top_right_grid_pin_11_
port 82 nsew default input
rlabel metal4 s 4944 2128 5264 21808 6 vpwr
port 83 nsew default input
rlabel metal4 s 8944 2128 9264 21808 6 vgnd
port 84 nsew default input
<< end >>
