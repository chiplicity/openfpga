* NGSPICE file created from sb_0__3_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor3_4 abstract view
.subckt scs8hd_nor3_4 A B C Y vgnd vpwr
.ends

.subckt sb_0__3_ address[0] address[1] address[2] address[3] address[4] address[5]
+ bottom_left_grid_pin_11_ bottom_left_grid_pin_13_ bottom_left_grid_pin_15_ bottom_left_grid_pin_1_
+ bottom_left_grid_pin_3_ bottom_left_grid_pin_5_ bottom_left_grid_pin_7_ bottom_left_grid_pin_9_
+ bottom_right_grid_pin_11_ chanx_right_in[0] chanx_right_in[1] chanx_right_in[2]
+ chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7]
+ chanx_right_in[8] chanx_right_out[0] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8]
+ chany_bottom_in[0] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4]
+ chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_out[0]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ data_in enable right_bottom_grid_pin_12_ right_top_grid_pin_11_ right_top_grid_pin_13_
+ right_top_grid_pin_15_ right_top_grid_pin_1_ right_top_grid_pin_3_ right_top_grid_pin_5_
+ right_top_grid_pin_7_ right_top_grid_pin_9_ vpwr vgnd
Xmem_right_track_12.LATCH_1_.latch data_in _097_/A _143_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_166 vpwr vgnd scs8hd_fill_2
XFILLER_22_177 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 bottom_right_grid_pin_11_ mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_74 vgnd vpwr scs8hd_fill_1
XFILLER_26_41 vgnd vpwr scs8hd_decap_8
XFILLER_9_137 vgnd vpwr scs8hd_decap_8
XFILLER_9_148 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_118 vgnd vpwr scs8hd_decap_6
Xmux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _097_/A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__124__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_200_ _200_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA__209__A _209_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_217 vgnd vpwr scs8hd_decap_12
XFILLER_23_20 vgnd vpwr scs8hd_decap_4
X_131_ _128_/A _131_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_97 vpwr vgnd scs8hd_fill_2
XFILLER_2_143 vgnd vpwr scs8hd_decap_8
XANTENNA__119__A _119_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _209_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ _104_/Y mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_53 vpwr vgnd scs8hd_fill_2
XFILLER_11_220 vgnd vpwr scs8hd_decap_12
X_114_ _114_/A _114_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__121__B address[5] vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _191_/HI _101_/Y mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_227 vgnd vpwr scs8hd_decap_6
XFILLER_6_12 vpwr vgnd scs8hd_fill_2
XFILLER_6_23 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__132__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_19_161 vgnd vpwr scs8hd_decap_3
Xmem_right_track_8.LATCH_1_.latch data_in _093_/A _137_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_32 vgnd vpwr scs8hd_decap_3
XFILLER_25_153 vgnd vpwr scs8hd_fill_1
XFILLER_31_53 vpwr vgnd scs8hd_fill_2
XFILLER_31_42 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ _092_/A mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_0_230 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _118_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_31_134 vgnd vpwr scs8hd_decap_12
XFILLER_31_101 vpwr vgnd scs8hd_fill_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__A address[3] vgnd vpwr scs8hd_diode_2
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _096_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_123 vgnd vpwr scs8hd_decap_3
XFILLER_26_64 vpwr vgnd scs8hd_fill_2
XFILLER_9_116 vpwr vgnd scs8hd_fill_2
XFILLER_13_178 vpwr vgnd scs8hd_fill_2
XFILLER_3_24 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_77 vgnd vpwr scs8hd_decap_12
XFILLER_33_218 vpwr vgnd scs8hd_fill_2
XFILLER_5_196 vgnd vpwr scs8hd_decap_12
XFILLER_5_130 vgnd vpwr scs8hd_decap_4
XANTENNA__124__B _125_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _104_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_15.LATCH_0_.latch_SLEEPB _175_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_229 vgnd vpwr scs8hd_decap_4
X_130_ address[3] _167_/B _123_/C _167_/D _131_/B vgnd vpwr scs8hd_or4_4
XFILLER_0_47 vpwr vgnd scs8hd_fill_2
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
XANTENNA__135__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _120_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_232 vgnd vpwr scs8hd_fill_1
X_113_ _113_/A _113_/Y vgnd vpwr scs8hd_inv_8
XFILLER_15_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _098_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _100_/A mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_29_118 vpwr vgnd scs8hd_fill_2
XFILLER_20_66 vgnd vpwr scs8hd_decap_3
XFILLER_29_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__132__B _131_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_140 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_13.LATCH_1_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_11 vgnd vpwr scs8hd_decap_3
XFILLER_15_55 vpwr vgnd scs8hd_fill_2
XFILLER_15_88 vpwr vgnd scs8hd_fill_2
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_146 vgnd vpwr scs8hd_decap_12
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_16.INVTX1_0_.scs8hd_inv_1 right_bottom_grid_pin_12_ mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _106_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_154 vgnd vpwr scs8hd_decap_3
XFILLER_16_176 vgnd vpwr scs8hd_decap_3
XANTENNA__127__B address[2] vgnd vpwr scs8hd_diode_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_190 vgnd vpwr scs8hd_decap_12
XFILLER_22_146 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _087_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _205_/A vgnd vpwr scs8hd_inv_1
XFILLER_3_58 vgnd vpwr scs8hd_fill_1
XANTENNA__138__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_12_190 vgnd vpwr scs8hd_decap_12
XFILLER_10_127 vgnd vpwr scs8hd_fill_1
XFILLER_12_23 vgnd vpwr scs8hd_decap_8
XFILLER_12_56 vpwr vgnd scs8hd_fill_2
XFILLER_12_89 vgnd vpwr scs8hd_decap_3
XFILLER_5_153 vpwr vgnd scs8hd_fill_2
XANTENNA__140__B _140_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB _146_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_44 vpwr vgnd scs8hd_fill_2
XFILLER_23_55 vpwr vgnd scs8hd_fill_2
XFILLER_23_77 vpwr vgnd scs8hd_fill_2
XFILLER_3_3 vpwr vgnd scs8hd_fill_2
XFILLER_2_167 vgnd vpwr scs8hd_decap_4
XFILLER_9_13 vpwr vgnd scs8hd_fill_2
XFILLER_9_24 vgnd vpwr scs8hd_decap_3
XANTENNA__135__B _135_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_46 vpwr vgnd scs8hd_fill_2
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr
+ scs8hd_diode_2
X_189_ _189_/HI _189_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__151__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XFILLER_18_66 vpwr vgnd scs8hd_fill_2
XFILLER_18_88 vgnd vpwr scs8hd_decap_4
X_112_ _112_/A _112_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__146__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_91 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _089_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _087_/A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_29_98 vpwr vgnd scs8hd_fill_2
XFILLER_28_141 vgnd vpwr scs8hd_decap_12
XFILLER_28_130 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_69 vpwr vgnd scs8hd_fill_2
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
XFILLER_34_111 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1_A bottom_left_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_25_111 vpwr vgnd scs8hd_fill_2
XFILLER_31_22 vgnd vpwr scs8hd_decap_12
XFILLER_31_11 vpwr vgnd scs8hd_fill_2
XFILLER_16_122 vgnd vpwr scs8hd_decap_3
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_158 vgnd vpwr scs8hd_decap_12
XFILLER_31_114 vgnd vpwr scs8hd_decap_6
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_188 vpwr vgnd scs8hd_fill_2
XANTENNA__127__C _123_/C vgnd vpwr scs8hd_diode_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__B _144_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_158 vgnd vpwr scs8hd_decap_8
Xmem_right_track_4.LATCH_1_.latch data_in _089_/A _131_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_107 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
Xmux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _194_/HI _091_/Y mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__138__B _138_/B vgnd vpwr scs8hd_diode_2
XANTENNA__154__A address[0] vgnd vpwr scs8hd_diode_2
Xmux_right_track_14.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_15_ mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_10_106 vgnd vpwr scs8hd_decap_8
XFILLER_5_7 vgnd vpwr scs8hd_fill_1
XFILLER_12_13 vgnd vpwr scs8hd_decap_4
XFILLER_12_35 vpwr vgnd scs8hd_fill_2
XFILLER_5_110 vpwr vgnd scs8hd_fill_2
XANTENNA__149__A address[3] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _119_/A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_23_231 vpwr vgnd scs8hd_fill_2
XFILLER_2_113 vgnd vpwr scs8hd_decap_4
XFILLER_0_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
X_188_ _188_/HI _188_/LO vgnd vpwr scs8hd_conb_1
XFILLER_29_3 vgnd vpwr scs8hd_decap_3
Xmux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _095_/A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__151__B _151_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1_A bottom_left_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_23 vgnd vpwr scs8hd_decap_6
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XFILLER_34_99 vgnd vpwr scs8hd_decap_12
X_111_ _111_/A _111_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__146__B _147_/B vgnd vpwr scs8hd_diode_2
XANTENNA__162__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_70 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_24 vgnd vpwr scs8hd_decap_4
XFILLER_29_44 vpwr vgnd scs8hd_fill_2
XFILLER_29_33 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _195_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_120 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_7.LATCH_0_.latch_SLEEPB _163_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_48 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_13.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_178 vgnd vpwr scs8hd_decap_12
XFILLER_34_123 vgnd vpwr scs8hd_decap_12
XANTENNA__157__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_19_175 vpwr vgnd scs8hd_fill_2
XFILLER_19_197 vpwr vgnd scs8hd_fill_2
Xmux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _190_/HI _099_/Y mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_134 vpwr vgnd scs8hd_fill_2
XFILLER_25_145 vpwr vgnd scs8hd_fill_2
XFILLER_25_156 vgnd vpwr scs8hd_decap_12
XFILLER_31_34 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_126 vpwr vgnd scs8hd_fill_2
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__D _127_/D vgnd vpwr scs8hd_diode_2
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_3 vgnd vpwr scs8hd_fill_1
XFILLER_26_23 vgnd vpwr scs8hd_decap_6
XFILLER_13_126 vpwr vgnd scs8hd_fill_2
XANTENNA__154__B _152_/X vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ _090_/A mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__170__A _167_/A vgnd vpwr scs8hd_diode_2
XANTENNA__080__A address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_5.LATCH_1_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__149__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_32_210 vgnd vpwr scs8hd_decap_4
XANTENNA__165__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_24 vgnd vpwr scs8hd_fill_1
Xmux_right_track_12.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_13_ mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_210 vgnd vpwr scs8hd_decap_4
X_187_ _187_/HI _187_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_191 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _094_/Y mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_20_202 vgnd vpwr scs8hd_decap_12
XFILLER_18_46 vgnd vpwr scs8hd_decap_4
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
X_110_ _110_/A _110_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _117_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _095_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__162__B _162_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_60 vgnd vpwr scs8hd_fill_1
XFILLER_28_154 vgnd vpwr scs8hd_decap_12
XFILLER_6_16 vpwr vgnd scs8hd_fill_2
XFILLER_10_80 vgnd vpwr scs8hd_fill_1
XFILLER_10_91 vgnd vpwr scs8hd_fill_1
XFILLER_13_7 vgnd vpwr scs8hd_decap_3
XFILLER_20_8 vgnd vpwr scs8hd_decap_3
XFILLER_19_121 vgnd vpwr scs8hd_fill_1
XFILLER_34_135 vgnd vpwr scs8hd_decap_12
XANTENNA__157__B _156_/B vgnd vpwr scs8hd_diode_2
XANTENNA__173__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA__083__A enable vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ _098_/A mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_25_168 vgnd vpwr scs8hd_decap_12
XFILLER_31_57 vpwr vgnd scs8hd_fill_2
XFILLER_31_46 vpwr vgnd scs8hd_fill_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_168 vgnd vpwr scs8hd_decap_8
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_190 vgnd vpwr scs8hd_decap_12
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _103_/Y vgnd
+ vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__168__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_68 vgnd vpwr scs8hd_decap_6
XFILLER_21_171 vpwr vgnd scs8hd_fill_2
XFILLER_21_193 vpwr vgnd scs8hd_fill_2
XFILLER_3_39 vpwr vgnd scs8hd_fill_2
XANTENNA__170__B _167_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_230 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _119_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[3] mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_219 vgnd vpwr scs8hd_decap_12
Xmem_right_track_0.LATCH_1_.latch data_in _086_/A _124_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_145 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _097_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ _102_/Y mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__149__C _167_/C vgnd vpwr scs8hd_diode_2
XANTENNA__165__B _165_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_93 vgnd vpwr scs8hd_fill_1
XFILLER_23_211 vgnd vpwr scs8hd_decap_12
XANTENNA__091__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_126 vgnd vpwr scs8hd_decap_8
X_186_ _186_/HI _186_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_91 vpwr vgnd scs8hd_fill_2
XFILLER_1_181 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _090_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__176__A _127_/D vgnd vpwr scs8hd_diode_2
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XANTENNA__086__A _086_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _105_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_10.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_11_ mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_169_ address[0] _168_/B _169_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_7.LATCH_0_.latch data_in _110_/A _163_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_57 vpwr vgnd scs8hd_fill_2
XFILLER_28_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_90 vpwr vgnd scs8hd_fill_2
XFILLER_19_111 vpwr vgnd scs8hd_fill_2
XFILLER_34_147 vgnd vpwr scs8hd_decap_6
XANTENNA__173__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_15_37 vpwr vgnd scs8hd_fill_2
XFILLER_33_191 vgnd vpwr scs8hd_decap_12
XFILLER_15_59 vpwr vgnd scs8hd_fill_2
XFILLER_0_213 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_103 vpwr vgnd scs8hd_fill_2
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _086_/A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_21_80 vgnd vpwr scs8hd_decap_6
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__168__B _168_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_106 vpwr vgnd scs8hd_fill_2
XFILLER_22_128 vgnd vpwr scs8hd_decap_4
XFILLER_13_106 vpwr vgnd scs8hd_fill_2
XANTENNA__094__A _094_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _092_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_154 vgnd vpwr scs8hd_decap_12
XANTENNA__170__C _167_/C vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.tap_buf4_0_.scs8hd_inv_1 mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ _198_/A vgnd vpwr scs8hd_inv_1
XANTENNA__089__A _089_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_168 vgnd vpwr scs8hd_decap_12
XANTENNA__149__D _167_/D vgnd vpwr scs8hd_diode_2
XFILLER_4_50 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _193_/HI _089_/Y mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_59 vpwr vgnd scs8hd_fill_2
XFILLER_23_223 vgnd vpwr scs8hd_decap_8
XFILLER_3_7 vgnd vpwr scs8hd_decap_4
XFILLER_2_105 vgnd vpwr scs8hd_decap_6
XFILLER_9_17 vpwr vgnd scs8hd_fill_2
X_185_ _185_/HI _185_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_81 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[4] mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__176__B _175_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_215 vgnd vpwr scs8hd_decap_12
XFILLER_18_15 vpwr vgnd scs8hd_fill_2
XFILLER_7_208 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _117_/A mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_168_ _128_/A _168_/B _168_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_27_3 vgnd vpwr scs8hd_decap_3
X_099_ _099_/A _099_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_40 vgnd vpwr scs8hd_decap_4
XFILLER_1_62 vgnd vpwr scs8hd_decap_3
XFILLER_28_178 vgnd vpwr scs8hd_decap_12
XANTENNA__097__A _097_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_15.LATCH_0_.latch data_in _118_/A _175_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_93 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_123 vpwr vgnd scs8hd_fill_2
XANTENNA__173__C address[4] vgnd vpwr scs8hd_diode_2
XFILLER_33_181 vpwr vgnd scs8hd_fill_2
XFILLER_15_16 vgnd vpwr scs8hd_decap_3
XFILLER_25_115 vgnd vpwr scs8hd_decap_4
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1 vgnd vpwr scs8hd_decap_3
Xmux_right_track_6.tap_buf4_0_.scs8hd_inv_1 mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ _201_/A vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_17.INVTX1_1_.scs8hd_inv_1 bottom_left_grid_pin_15_ mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_151 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _189_/HI _097_/Y mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_122 vgnd vpwr scs8hd_fill_1
XFILLER_8_166 vgnd vpwr scs8hd_decap_12
XANTENNA__170__D _127_/D vgnd vpwr scs8hd_diode_2
XFILLER_12_39 vpwr vgnd scs8hd_fill_2
XFILLER_5_114 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ _211_/A vgnd vpwr scs8hd_inv_1
XFILLER_17_221 vpwr vgnd scs8hd_fill_2
XFILLER_4_84 vgnd vpwr scs8hd_decap_6
Xmux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _088_/A mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_16 vpwr vgnd scs8hd_fill_2
XFILLER_23_27 vpwr vgnd scs8hd_fill_2
XFILLER_9_29 vpwr vgnd scs8hd_fill_2
X_184_ _184_/HI _184_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_60 vgnd vpwr scs8hd_fill_1
XFILLER_1_161 vpwr vgnd scs8hd_fill_2
XFILLER_1_150 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__176__C _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_227 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_track_15.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_098_ _098_/A _098_/Y vgnd vpwr scs8hd_inv_8
X_167_ _167_/A _167_/B _167_/C _167_/D _168_/B vgnd vpwr scs8hd_or4_4
XFILLER_1_52 vpwr vgnd scs8hd_fill_2
XFILLER_1_74 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[5] mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_15 vpwr vgnd scs8hd_fill_2
XFILLER_20_28 vgnd vpwr scs8hd_fill_1
XFILLER_29_48 vgnd vpwr scs8hd_decap_3
XFILLER_29_37 vgnd vpwr scs8hd_decap_4
XFILLER_28_102 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ _092_/Y mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_10_61 vgnd vpwr scs8hd_fill_1
XFILLER_10_83 vgnd vpwr scs8hd_decap_8
XFILLER_19_157 vpwr vgnd scs8hd_fill_2
XFILLER_19_179 vpwr vgnd scs8hd_fill_2
XANTENNA__173__D _173_/D vgnd vpwr scs8hd_diode_2
XANTENNA__198__A _198_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_138 vpwr vgnd scs8hd_fill_2
XFILLER_25_149 vgnd vpwr scs8hd_decap_4
XFILLER_31_38 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_3.LATCH_0_.latch data_in _106_/A _157_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_204 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_127 vgnd vpwr scs8hd_decap_3
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_2 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ _120_/A mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_15_160 vpwr vgnd scs8hd_fill_2
XFILLER_15_193 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _120_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_7_40 vpwr vgnd scs8hd_fill_2
XFILLER_7_51 vpwr vgnd scs8hd_fill_2
XFILLER_7_62 vpwr vgnd scs8hd_fill_2
XFILLER_7_84 vpwr vgnd scs8hd_fill_2
XFILLER_26_49 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _098_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_82 vpwr vgnd scs8hd_fill_2
XFILLER_16_93 vgnd vpwr scs8hd_fill_1
XFILLER_8_178 vgnd vpwr scs8hd_decap_12
Xmux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ _096_/A mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_35_211 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_126 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_15.INVTX1_1_.scs8hd_inv_1 bottom_left_grid_pin_13_ mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_92 vpwr vgnd scs8hd_fill_2
XFILLER_4_63 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _106_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_0_.scs8hd_inv_1 chanx_right_in[3] mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_183_ _183_/HI _183_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_173 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _100_/Y mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
XFILLER_1_6 vpwr vgnd scs8hd_fill_2
XFILLER_24_93 vpwr vgnd scs8hd_fill_2
X_097_ _097_/A _097_/Y vgnd vpwr scs8hd_inv_8
X_166_ address[0] _165_/B _166_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _100_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_114 vgnd vpwr scs8hd_decap_6
XFILLER_10_51 vgnd vpwr scs8hd_decap_3
XFILLER_19_71 vgnd vpwr scs8hd_decap_4
X_149_ address[3] address[2] _167_/C _167_/D _151_/B vgnd vpwr scs8hd_or4_4
XFILLER_33_150 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ _207_/A vgnd vpwr scs8hd_inv_1
Xmux_right_track_2.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[6] mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_139 vgnd vpwr scs8hd_decap_12
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_bottom_track_11.LATCH_0_.latch data_in _114_/A _169_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_15_172 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _108_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_175 vpwr vgnd scs8hd_fill_2
XFILLER_21_197 vgnd vpwr scs8hd_decap_4
XFILLER_8_102 vgnd vpwr scs8hd_decap_12
XFILLER_12_120 vgnd vpwr scs8hd_decap_12
XFILLER_8_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _089_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_19 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_71 vgnd vpwr scs8hd_decap_8
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB _154_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_171 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_182_ _182_/HI _182_/LO vgnd vpwr scs8hd_conb_1
XFILLER_14_215 vgnd vpwr scs8hd_decap_12
XFILLER_13_62 vpwr vgnd scs8hd_fill_2
XFILLER_13_95 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_13.INVTX1_1_.scs8hd_inv_1 bottom_left_grid_pin_11_ mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__100__A _100_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_230 vgnd vpwr scs8hd_decap_3
Xmux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _192_/HI _087_/Y mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_165_ _128_/A _165_/B _165_/Y vgnd vpwr scs8hd_nor2_4
X_096_ _096_/A _096_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_10 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_7.INVTX1_0_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_87 vpwr vgnd scs8hd_fill_2
XFILLER_10_74 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _091_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_94 vpwr vgnd scs8hd_fill_2
XFILLER_19_115 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _115_/A mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_148_ address[4] _173_/D _167_/C vgnd vpwr scs8hd_nand2_4
XANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_33_173 vgnd vpwr scs8hd_decap_8
XFILLER_31_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_107 vgnd vpwr scs8hd_decap_4
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_62 vgnd vpwr scs8hd_decap_4
XFILLER_30_154 vgnd vpwr scs8hd_decap_12
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_8_114 vgnd vpwr scs8hd_fill_1
XFILLER_8_125 vgnd vpwr scs8hd_fill_1
XFILLER_12_132 vgnd vpwr scs8hd_decap_4
XFILLER_12_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB _176_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_147 vgnd vpwr scs8hd_decap_6
XANTENNA__103__A _103_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[7] mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _182_/HI _119_/Y mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_213 vgnd vpwr scs8hd_fill_1
XFILLER_5_106 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A bottom_right_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_32_227 vgnd vpwr scs8hd_decap_6
Xmux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _188_/HI _095_/Y mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_183 vpwr vgnd scs8hd_fill_2
XFILLER_4_32 vgnd vpwr scs8hd_decap_3
XFILLER_4_10 vpwr vgnd scs8hd_fill_2
XFILLER_14_227 vgnd vpwr scs8hd_decap_6
X_181_ _181_/HI _181_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_52 vpwr vgnd scs8hd_fill_2
XFILLER_13_85 vgnd vpwr scs8hd_decap_4
Xmem_right_track_14.LATCH_0_.latch data_in _100_/A _147_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_18_19 vpwr vgnd scs8hd_fill_2
XFILLER_11_208 vgnd vpwr scs8hd_decap_12
XANTENNA__201__A _201_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ _085_/A mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr
+ scs8hd_diode_2
X_164_ _167_/A address[2] _167_/C _127_/D _165_/B vgnd vpwr scs8hd_or4_4
X_095_ _095_/A _095_/Y vgnd vpwr scs8hd_inv_8
XFILLER_24_84 vpwr vgnd scs8hd_fill_2
XANTENNA__111__A _111_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_44 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A bottom_left_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_12.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_11.INVTX1_1_.scs8hd_inv_1 bottom_left_grid_pin_9_ mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_10_20 vpwr vgnd scs8hd_fill_2
XFILLER_10_64 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_11.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_127 vpwr vgnd scs8hd_fill_2
XFILLER_35_94 vgnd vpwr scs8hd_decap_12
XFILLER_27_182 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__106__A _106_/A vgnd vpwr scs8hd_diode_2
X_147_ address[0] _147_/B _147_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_bottom_track_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _188_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_3 vgnd vpwr scs8hd_decap_3
XFILLER_33_141 vgnd vpwr scs8hd_decap_4
XFILLER_18_182 vgnd vpwr scs8hd_decap_4
XFILLER_25_119 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_5.INVTX1_0_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_218 vgnd vpwr scs8hd_decap_12
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_30_166 vgnd vpwr scs8hd_decap_12
XFILLER_7_21 vgnd vpwr scs8hd_decap_4
Xmux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ _090_/Y mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_26_19 vpwr vgnd scs8hd_fill_2
XFILLER_32_62 vgnd vpwr scs8hd_decap_12
XFILLER_12_166 vgnd vpwr scs8hd_decap_12
XFILLER_16_63 vpwr vgnd scs8hd_fill_2
XFILLER_16_74 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ _118_/A mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_5_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__204__A _204_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_40 vpwr vgnd scs8hd_fill_2
XFILLER_17_225 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB _135_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__114__A _114_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _178_/HI vgnd vpwr
+ scs8hd_diode_2
X_180_ _180_/HI _180_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_42 vgnd vpwr scs8hd_fill_1
XFILLER_1_132 vpwr vgnd scs8hd_fill_2
XFILLER_1_187 vpwr vgnd scs8hd_fill_2
XANTENNA__109__A _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_41 vgnd vpwr scs8hd_decap_3
XFILLER_24_63 vpwr vgnd scs8hd_fill_2
X_094_ _094_/A _094_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_213 vgnd vpwr scs8hd_fill_1
X_163_ address[0] _162_/B _163_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_23 vpwr vgnd scs8hd_fill_2
XFILLER_1_56 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _119_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_19 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _097_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ _098_/Y mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_3_205 vgnd vpwr scs8hd_decap_12
XANTENNA__212__A _212_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_43 vpwr vgnd scs8hd_fill_2
XANTENNA__122__A address[1] vgnd vpwr scs8hd_diode_2
X_146_ _128_/A _147_/B _146_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_131 vgnd vpwr scs8hd_decap_3
XFILLER_33_120 vpwr vgnd scs8hd_fill_2
XFILLER_18_150 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__207__A _207_/A vgnd vpwr scs8hd_diode_2
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_42 vgnd vpwr scs8hd_decap_4
XFILLER_21_53 vpwr vgnd scs8hd_fill_2
XFILLER_21_97 vpwr vgnd scs8hd_fill_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_164 vgnd vpwr scs8hd_decap_8
XFILLER_15_175 vpwr vgnd scs8hd_fill_2
XFILLER_30_178 vgnd vpwr scs8hd_decap_12
XFILLER_7_44 vpwr vgnd scs8hd_fill_2
XFILLER_7_55 vpwr vgnd scs8hd_fill_2
XFILLER_7_66 vgnd vpwr scs8hd_decap_3
XFILLER_7_88 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A _117_/A vgnd vpwr scs8hd_diode_2
X_129_ address[0] _129_/B _129_/Y vgnd vpwr scs8hd_nor2_4
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _111_/A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _105_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_101 vpwr vgnd scs8hd_fill_2
XFILLER_21_123 vgnd vpwr scs8hd_decap_3
XFILLER_21_167 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_7.LATCH_1_.latch data_in _109_/A _162_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_16_86 vgnd vpwr scs8hd_decap_4
XFILLER_32_96 vpwr vgnd scs8hd_fill_2
XFILLER_32_74 vgnd vpwr scs8hd_decap_12
XFILLER_32_52 vgnd vpwr scs8hd_fill_1
XFILLER_32_30 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_3.INVTX1_0_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_145 vgnd vpwr scs8hd_decap_8
XFILLER_12_178 vgnd vpwr scs8hd_decap_12
XFILLER_26_215 vgnd vpwr scs8hd_decap_12
XFILLER_27_96 vpwr vgnd scs8hd_fill_2
XFILLER_4_163 vgnd vpwr scs8hd_decap_8
XFILLER_4_152 vgnd vpwr scs8hd_fill_1
XFILLER_4_67 vpwr vgnd scs8hd_fill_2
XFILLER_4_23 vgnd vpwr scs8hd_decap_8
XANTENNA__130__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _099_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_3 vgnd vpwr scs8hd_decap_3
XFILLER_9_211 vgnd vpwr scs8hd_decap_4
XFILLER_9_222 vgnd vpwr scs8hd_decap_8
XANTENNA__125__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _092_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB _165_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_162_ _128_/A _162_/B _162_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_97 vgnd vpwr scs8hd_decap_3
X_093_ _093_/A _093_/Y vgnd vpwr scs8hd_inv_8
Xmem_right_track_10.LATCH_0_.latch data_in _096_/A _141_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _107_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_217 vgnd vpwr scs8hd_decap_12
XFILLER_19_42 vpwr vgnd scs8hd_fill_2
XFILLER_19_53 vpwr vgnd scs8hd_fill_2
XFILLER_19_107 vpwr vgnd scs8hd_fill_2
XFILLER_35_63 vgnd vpwr scs8hd_decap_12
XFILLER_27_184 vgnd vpwr scs8hd_decap_12
X_145_ _167_/A _167_/B _123_/C _127_/D _147_/B vgnd vpwr scs8hd_or4_4
Xmux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _187_/HI _086_/Y mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_32_7 vgnd vpwr scs8hd_decap_8
XANTENNA__122__B _083_/Y vgnd vpwr scs8hd_diode_2
XFILLER_33_187 vpwr vgnd scs8hd_fill_2
XFILLER_33_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_209 vpwr vgnd scs8hd_fill_2
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_154 vgnd vpwr scs8hd_decap_12
XFILLER_30_135 vgnd vpwr scs8hd_decap_12
XFILLER_30_102 vgnd vpwr scs8hd_decap_3
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_110 vpwr vgnd scs8hd_fill_2
XFILLER_15_198 vgnd vpwr scs8hd_decap_12
XANTENNA__133__A address[3] vgnd vpwr scs8hd_diode_2
X_128_ _128_/A _129_/B _128_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_3 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _113_/A mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_21_135 vpwr vgnd scs8hd_fill_2
XFILLER_21_179 vpwr vgnd scs8hd_fill_2
XFILLER_16_10 vpwr vgnd scs8hd_fill_2
XFILLER_16_32 vgnd vpwr scs8hd_decap_3
XFILLER_32_86 vgnd vpwr scs8hd_decap_6
XFILLER_20_190 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_15.LATCH_1_.latch data_in _117_/A _174_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__128__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_227 vgnd vpwr scs8hd_decap_6
XFILLER_26_205 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _094_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_46 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_0_.scs8hd_inv_1 chanx_right_in[7] mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__130__B _167_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _181_/HI _117_/Y mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_77 vpwr vgnd scs8hd_fill_2
XFILLER_1_112 vgnd vpwr scs8hd_decap_4
Xmem_right_track_6.LATCH_0_.latch data_in _092_/A _135_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__125__B _125_/B vgnd vpwr scs8hd_diode_2
XANTENNA__141__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
XFILLER_10_200 vgnd vpwr scs8hd_decap_12
X_161_ _167_/A address[2] _167_/C _167_/D _162_/B vgnd vpwr scs8hd_or4_4
XFILLER_24_21 vgnd vpwr scs8hd_decap_8
X_092_ _092_/A _092_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_47 vpwr vgnd scs8hd_fill_2
XANTENNA__136__A _167_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_229 vgnd vpwr scs8hd_decap_4
XFILLER_35_75 vgnd vpwr scs8hd_decap_12
XFILLER_27_196 vgnd vpwr scs8hd_decap_12
X_144_ address[0] _144_/B _144_/Y vgnd vpwr scs8hd_nor2_4
X_213_ _213_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_7 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.tap_buf4_0_.scs8hd_inv_1 mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _203_/A vgnd vpwr scs8hd_inv_1
XFILLER_18_141 vgnd vpwr scs8hd_decap_6
XFILLER_18_163 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_166 vgnd vpwr scs8hd_decap_12
XFILLER_21_22 vgnd vpwr scs8hd_fill_1
XFILLER_21_66 vgnd vpwr scs8hd_fill_1
XFILLER_15_100 vgnd vpwr scs8hd_fill_1
XFILLER_30_147 vgnd vpwr scs8hd_decap_6
XFILLER_30_125 vgnd vpwr scs8hd_fill_1
XPHY_8 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_144 vgnd vpwr scs8hd_fill_1
XANTENNA__133__B _167_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_13 vpwr vgnd scs8hd_fill_2
X_127_ address[3] address[2] _123_/C _127_/D _129_/B vgnd vpwr scs8hd_or4_4
Xmux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _213_/A vgnd vpwr scs8hd_inv_1
XFILLER_21_114 vpwr vgnd scs8hd_fill_2
XFILLER_29_214 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_8_118 vgnd vpwr scs8hd_decap_4
XFILLER_16_44 vpwr vgnd scs8hd_fill_2
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XANTENNA__144__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__128__B _129_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_184 vgnd vpwr scs8hd_decap_12
Xmux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _088_/Y mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_27_54 vpwr vgnd scs8hd_fill_2
XFILLER_17_206 vgnd vpwr scs8hd_decap_8
XFILLER_17_217 vpwr vgnd scs8hd_fill_2
XFILLER_4_187 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_3.LATCH_1_.latch data_in _105_/A _156_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__130__C _123_/C vgnd vpwr scs8hd_diode_2
XFILLER_31_220 vgnd vpwr scs8hd_decap_12
XANTENNA__139__A _167_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_12 vpwr vgnd scs8hd_fill_2
XFILLER_13_34 vpwr vgnd scs8hd_fill_2
XFILLER_13_56 vpwr vgnd scs8hd_fill_2
XFILLER_1_168 vgnd vpwr scs8hd_decap_3
XFILLER_1_157 vpwr vgnd scs8hd_fill_2
XFILLER_1_146 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ _116_/A mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_13_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__141__B _140_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_13.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_90 vgnd vpwr scs8hd_fill_1
XFILLER_24_11 vgnd vpwr scs8hd_fill_1
X_091_ _091_/A _091_/Y vgnd vpwr scs8hd_inv_8
X_160_ address[0] _158_/X _160_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_227 vgnd vpwr scs8hd_decap_6
XFILLER_10_212 vpwr vgnd scs8hd_fill_2
XFILLER_24_88 vgnd vpwr scs8hd_decap_4
XANTENNA__136__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__152__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_10_24 vpwr vgnd scs8hd_fill_2
XFILLER_10_57 vgnd vpwr scs8hd_decap_4
XFILLER_19_77 vpwr vgnd scs8hd_fill_2
XFILLER_35_87 vgnd vpwr scs8hd_decap_6
XFILLER_35_32 vgnd vpwr scs8hd_decap_12
X_212_ _212_/A chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
X_143_ _128_/A _144_/B _143_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_145 vgnd vpwr scs8hd_fill_1
XFILLER_33_123 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ _120_/Y mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _189_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__147__A address[0] vgnd vpwr scs8hd_diode_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_145 vpwr vgnd scs8hd_fill_2
XFILLER_24_178 vgnd vpwr scs8hd_decap_12
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_123 vpwr vgnd scs8hd_fill_2
XFILLER_15_134 vpwr vgnd scs8hd_fill_2
Xmux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ _096_/Y mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_156 vpwr vgnd scs8hd_fill_2
XANTENNA__133__C _123_/C vgnd vpwr scs8hd_diode_2
X_126_ address[1] enable _127_/D vgnd vpwr scs8hd_nand2_4
XFILLER_16_23 vgnd vpwr scs8hd_decap_8
XFILLER_32_44 vgnd vpwr scs8hd_decap_8
XFILLER_12_104 vpwr vgnd scs8hd_fill_2
XFILLER_16_67 vpwr vgnd scs8hd_fill_2
XFILLER_16_78 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_13.LATCH_0_.latch_SLEEPB _172_/Y vgnd vpwr scs8hd_diode_2
XFILLER_35_218 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _100_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__144__B _144_/B vgnd vpwr scs8hd_diode_2
X_109_ _109_/A _109_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__160__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_7_196 vgnd vpwr scs8hd_decap_12
XFILLER_8_90 vpwr vgnd scs8hd_fill_2
XFILLER_27_44 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _109_/A mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_4_199 vgnd vpwr scs8hd_decap_12
XFILLER_4_144 vgnd vpwr scs8hd_decap_8
XFILLER_4_133 vgnd vpwr scs8hd_decap_3
XFILLER_4_122 vpwr vgnd scs8hd_fill_2
XANTENNA__130__D _167_/D vgnd vpwr scs8hd_diode_2
XFILLER_31_232 vgnd vpwr scs8hd_fill_1
XANTENNA__155__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA__139__B address[2] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_11.LATCH_1_.latch data_in _113_/A _168_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_136 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _183_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_232 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _108_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_24_67 vgnd vpwr scs8hd_decap_8
X_090_ _090_/A _090_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_27 vpwr vgnd scs8hd_fill_2
XANTENNA__136__C _123_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB _147_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__152__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_11.LATCH_1_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_track_2.LATCH_0_.latch data_in _088_/A _129_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_47 vpwr vgnd scs8hd_fill_2
XFILLER_27_154 vgnd vpwr scs8hd_decap_12
XFILLER_35_44 vgnd vpwr scs8hd_decap_12
X_211_ _211_/A chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
X_142_ _167_/A _167_/B _123_/C _167_/D _144_/B vgnd vpwr scs8hd_or4_4
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _102_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_110 vgnd vpwr scs8hd_decap_4
XFILLER_18_121 vgnd vpwr scs8hd_decap_3
XANTENNA__147__B _147_/B vgnd vpwr scs8hd_diode_2
XANTENNA__163__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_2_81 vpwr vgnd scs8hd_fill_2
XFILLER_24_102 vpwr vgnd scs8hd_fill_2
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_135 vgnd vpwr scs8hd_fill_1
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
XFILLER_7_59 vpwr vgnd scs8hd_fill_2
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
X_125_ address[0] _125_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_30_7 vpwr vgnd scs8hd_fill_2
XANTENNA__133__D _127_/D vgnd vpwr scs8hd_diode_2
XANTENNA__158__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _110_/A vgnd
+ vpwr scs8hd_diode_2
X_108_ _108_/A _108_/Y vgnd vpwr scs8hd_inv_8
XFILLER_7_153 vgnd vpwr scs8hd_decap_12
XFILLER_11_182 vgnd vpwr scs8hd_fill_1
XANTENNA__160__B _158_/X vgnd vpwr scs8hd_diode_2
XFILLER_21_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _091_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _114_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__139__C _123_/C vgnd vpwr scs8hd_diode_2
XANTENNA__155__B _167_/B vgnd vpwr scs8hd_diode_2
XANTENNA__171__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_104 vpwr vgnd scs8hd_fill_2
XANTENNA__081__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _179_/HI vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__166__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_24_46 vgnd vpwr scs8hd_decap_6
XFILLER_6_207 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _180_/HI _115_/Y mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__136__D _167_/D vgnd vpwr scs8hd_diode_2
XANTENNA__152__C _167_/C vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ _112_/A mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_19_46 vpwr vgnd scs8hd_fill_2
XFILLER_35_56 vgnd vpwr scs8hd_decap_6
XFILLER_27_166 vgnd vpwr scs8hd_decap_12
XFILLER_27_100 vgnd vpwr scs8hd_decap_3
XFILLER_19_57 vpwr vgnd scs8hd_fill_2
X_210_ _210_/A chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
X_141_ address[0] _140_/B _141_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_169 vpwr vgnd scs8hd_fill_2
XFILLER_18_188 vpwr vgnd scs8hd_fill_2
XFILLER_18_199 vgnd vpwr scs8hd_decap_12
XANTENNA__163__B _162_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _093_/A vgnd vpwr
+ scs8hd_diode_2
Xmem_right_track_14.LATCH_1_.latch data_in _099_/A _146_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_93 vgnd vpwr scs8hd_decap_3
XFILLER_2_60 vgnd vpwr scs8hd_decap_4
XFILLER_24_125 vpwr vgnd scs8hd_fill_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_14 vpwr vgnd scs8hd_fill_2
XFILLER_21_25 vpwr vgnd scs8hd_fill_2
XFILLER_15_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_27 vpwr vgnd scs8hd_fill_2
X_124_ _128_/A _125_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__158__B _167_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_6 vpwr vgnd scs8hd_fill_2
XANTENNA__174__A _167_/D vgnd vpwr scs8hd_diode_2
XFILLER_21_139 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_217 vgnd vpwr scs8hd_decap_12
XANTENNA__084__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_11_150 vgnd vpwr scs8hd_decap_12
X_107_ _107_/A _107_/Y vgnd vpwr scs8hd_inv_8
XFILLER_7_165 vgnd vpwr scs8hd_decap_12
XFILLER_22_90 vpwr vgnd scs8hd_fill_2
XANTENNA__169__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_27_79 vpwr vgnd scs8hd_fill_2
XFILLER_25_220 vgnd vpwr scs8hd_decap_12
XANTENNA__139__D _127_/D vgnd vpwr scs8hd_diode_2
XFILLER_16_231 vpwr vgnd scs8hd_fill_2
XFILLER_17_90 vpwr vgnd scs8hd_fill_2
XANTENNA__155__C _167_/C vgnd vpwr scs8hd_diode_2
XANTENNA__171__B _170_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_26 vgnd vpwr scs8hd_decap_8
Xmux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ _085_/Y mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1_A bottom_left_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_182 vgnd vpwr scs8hd_decap_4
XFILLER_0_160 vpwr vgnd scs8hd_fill_2
XANTENNA__166__B _165_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_5.LATCH_0_.latch_SLEEPB _160_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__092__A _092_/A vgnd vpwr scs8hd_diode_2
XANTENNA__152__D _127_/D vgnd vpwr scs8hd_diode_2
XANTENNA__177__A _127_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_10.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ _114_/A mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_10_16 vpwr vgnd scs8hd_fill_2
XFILLER_19_25 vpwr vgnd scs8hd_fill_2
XFILLER_27_178 vgnd vpwr scs8hd_decap_4
XANTENNA__087__A _087_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_123 vpwr vgnd scs8hd_fill_2
X_140_ _128_/A _140_/B _140_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_18_167 vgnd vpwr scs8hd_decap_12
XFILLER_33_137 vpwr vgnd scs8hd_fill_2
XFILLER_33_104 vpwr vgnd scs8hd_fill_2
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_24_115 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_107 vgnd vpwr scs8hd_decap_12
XFILLER_7_17 vpwr vgnd scs8hd_fill_2
X_123_ address[3] address[2] _123_/C _167_/D _125_/B vgnd vpwr scs8hd_or4_4
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__158__C _167_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__174__B _175_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
XFILLER_29_229 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ _118_/Y mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_48 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1_A bottom_left_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_3.LATCH_1_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_111 vgnd vpwr scs8hd_decap_4
XFILLER_11_162 vgnd vpwr scs8hd_decap_12
X_106_ _106_/A _106_/Y vgnd vpwr scs8hd_inv_8
XFILLER_7_177 vgnd vpwr scs8hd_decap_6
XFILLER_11_184 vgnd vpwr scs8hd_decap_12
XANTENNA__169__B _168_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_82 vgnd vpwr scs8hd_decap_8
XFILLER_27_58 vgnd vpwr scs8hd_decap_3
XFILLER_27_25 vpwr vgnd scs8hd_fill_2
XFILLER_25_232 vgnd vpwr scs8hd_fill_1
XANTENNA__095__A _095_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_103 vpwr vgnd scs8hd_fill_2
XANTENNA__155__D _167_/D vgnd vpwr scs8hd_diode_2
XFILLER_3_180 vgnd vpwr scs8hd_fill_1
XFILLER_13_16 vgnd vpwr scs8hd_fill_1
XFILLER_13_38 vpwr vgnd scs8hd_fill_2
XFILLER_0_194 vpwr vgnd scs8hd_fill_2
XFILLER_0_172 vgnd vpwr scs8hd_decap_3
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_9_ mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _107_/A mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_10_227 vgnd vpwr scs8hd_decap_6
XFILLER_5_220 vgnd vpwr scs8hd_decap_12
XFILLER_14_70 vgnd vpwr scs8hd_decap_3
XFILLER_30_91 vgnd vpwr scs8hd_fill_1
XFILLER_30_80 vgnd vpwr scs8hd_fill_1
XANTENNA__177__B _175_/B vgnd vpwr scs8hd_diode_2
XFILLER_10_28 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _099_/Y vgnd
+ vpwr scs8hd_diode_2
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_80 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_199_ _199_/A chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _190_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _186_/HI _111_/Y mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_149 vgnd vpwr scs8hd_decap_4
XFILLER_32_182 vgnd vpwr scs8hd_fill_1
XFILLER_21_38 vpwr vgnd scs8hd_fill_2
XFILLER_21_49 vpwr vgnd scs8hd_fill_2
XANTENNA__098__A _098_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_119 vgnd vpwr scs8hd_decap_4
XFILLER_15_138 vgnd vpwr scs8hd_decap_6
X_122_ address[1] _083_/Y _167_/D vgnd vpwr scs8hd_or2_4
XFILLER_11_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__158__D _127_/D vgnd vpwr scs8hd_diode_2
XANTENNA__174__C _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_182 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_208 vgnd vpwr scs8hd_decap_6
XFILLER_12_108 vgnd vpwr scs8hd_decap_12
Xmem_right_track_10.LATCH_1_.latch data_in _095_/A _140_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_130 vpwr vgnd scs8hd_fill_2
XFILLER_20_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _107_/Y vgnd
+ vpwr scs8hd_diode_2
X_105_ _105_/A _105_/Y vgnd vpwr scs8hd_inv_8
XFILLER_7_134 vpwr vgnd scs8hd_fill_2
XFILLER_11_174 vgnd vpwr scs8hd_decap_8
XFILLER_11_196 vgnd vpwr scs8hd_decap_12
XFILLER_27_15 vpwr vgnd scs8hd_fill_2
XFILLER_4_126 vgnd vpwr scs8hd_decap_4
XFILLER_33_91 vgnd vpwr scs8hd_decap_4
XFILLER_3_170 vgnd vpwr scs8hd_decap_4
XANTENNA__196__A _196_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _101_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_218 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _184_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_91 vgnd vpwr scs8hd_fill_1
XFILLER_5_73 vpwr vgnd scs8hd_fill_2
XFILLER_5_51 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _094_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_232 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__177__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_7_ mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_114 vgnd vpwr scs8hd_decap_6
XFILLER_35_180 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _109_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_147 vgnd vpwr scs8hd_fill_1
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_81 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_25_92 vpwr vgnd scs8hd_fill_2
X_198_ _198_/A chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_2_85 vpwr vgnd scs8hd_fill_2
XFILLER_2_30 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _113_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _179_/HI _113_/Y mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_track_6.LATCH_1_.latch data_in _091_/A _134_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ _110_/A mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_121_ address[4] address[5] _123_/C vgnd vpwr scs8hd_or2_4
XFILLER_14_172 vgnd vpwr scs8hd_fill_1
XANTENNA__199__A _199_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _137_/Y vgnd vpwr scs8hd_diode_2
X_104_ _104_/A _104_/Y vgnd vpwr scs8hd_inv_8
XFILLER_22_82 vgnd vpwr scs8hd_decap_8
XFILLER_22_93 vpwr vgnd scs8hd_fill_2
XFILLER_14_6 vpwr vgnd scs8hd_fill_2
XFILLER_4_138 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_17.INVTX1_0_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_71 vgnd vpwr scs8hd_decap_4
XFILLER_33_81 vpwr vgnd scs8hd_fill_2
XFILLER_3_193 vgnd vpwr scs8hd_decap_12
XFILLER_12_3 vgnd vpwr scs8hd_fill_1
XFILLER_22_215 vgnd vpwr scs8hd_decap_12
XFILLER_1_108 vpwr vgnd scs8hd_fill_2
XFILLER_0_141 vpwr vgnd scs8hd_fill_2
XFILLER_28_81 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _180_/HI vgnd
+ vpwr scs8hd_diode_2
XFILLER_35_27 vgnd vpwr scs8hd_decap_4
XFILLER_27_137 vgnd vpwr scs8hd_decap_6
Xmux_right_track_14.tap_buf4_0_.scs8hd_inv_1 mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _197_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _085_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_26_181 vgnd vpwr scs8hd_decap_12
XPHY_82 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_18_126 vpwr vgnd scs8hd_fill_2
XFILLER_18_137 vpwr vgnd scs8hd_fill_2
XFILLER_25_71 vgnd vpwr scs8hd_decap_4
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_197_ _197_/A chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_17_181 vpwr vgnd scs8hd_fill_2
XFILLER_24_129 vgnd vpwr scs8hd_decap_6
XFILLER_21_18 vgnd vpwr scs8hd_decap_4
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
X_120_ _120_/A _120_/Y vgnd vpwr scs8hd_inv_8
XFILLER_23_151 vgnd vpwr scs8hd_decap_12
XFILLER_23_184 vgnd vpwr scs8hd_decap_8
XFILLER_23_195 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_5_ mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_40 vpwr vgnd scs8hd_fill_2
XFILLER_11_62 vpwr vgnd scs8hd_fill_2
XFILLER_11_73 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_154 vpwr vgnd scs8hd_fill_2
XFILLER_11_110 vgnd vpwr scs8hd_decap_12
XFILLER_7_103 vpwr vgnd scs8hd_fill_2
X_103_ _103_/A _103_/Y vgnd vpwr scs8hd_inv_8
XFILLER_34_202 vgnd vpwr scs8hd_decap_12
XFILLER_8_41 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ _116_/Y mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_16_213 vgnd vpwr scs8hd_fill_1
XFILLER_33_60 vgnd vpwr scs8hd_fill_1
XFILLER_17_94 vpwr vgnd scs8hd_fill_2
XFILLER_22_227 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_track_12.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_164 vgnd vpwr scs8hd_decap_8
XFILLER_0_153 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_11.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_86 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_15.INVTX1_0_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_29 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _200_/A vgnd vpwr scs8hd_inv_1
XFILLER_14_62 vpwr vgnd scs8hd_fill_2
XFILLER_14_84 vpwr vgnd scs8hd_fill_2
XANTENNA__101__A _101_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_29 vpwr vgnd scs8hd_fill_2
XFILLER_27_127 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _105_/A mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_6 vpwr vgnd scs8hd_fill_2
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XFILLER_33_108 vgnd vpwr scs8hd_decap_12
XPHY_61 vgnd vpwr scs8hd_decap_3
XFILLER_26_193 vgnd vpwr scs8hd_decap_12
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_83 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_72 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_50 vgnd vpwr scs8hd_decap_3
X_196_ _196_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
Xmux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ _210_/A vgnd vpwr scs8hd_inv_1
XFILLER_17_171 vpwr vgnd scs8hd_fill_2
XFILLER_24_119 vgnd vpwr scs8hd_decap_4
XFILLER_32_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_163 vgnd vpwr scs8hd_decap_12
XFILLER_2_3 vgnd vpwr scs8hd_decap_4
XFILLER_11_85 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_130 vpwr vgnd scs8hd_fill_2
XFILLER_14_141 vgnd vpwr scs8hd_decap_6
X_179_ _179_/HI _179_/LO vgnd vpwr scs8hd_conb_1
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XFILLER_32_18 vgnd vpwr scs8hd_decap_12
XFILLER_20_100 vpwr vgnd scs8hd_fill_2
XFILLER_20_111 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _185_/HI _109_/Y mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_track_2.LATCH_1_.latch data_in _087_/A _128_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_115 vgnd vpwr scs8hd_fill_1
XFILLER_22_51 vgnd vpwr scs8hd_fill_1
X_102_ _102_/A _102_/Y vgnd vpwr scs8hd_inv_8
Xmux_right_track_2.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_3_ mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _102_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_107 vgnd vpwr scs8hd_decap_4
XFILLER_17_40 vpwr vgnd scs8hd_fill_2
XANTENNA__104__A _104_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_206 vgnd vpwr scs8hd_decap_8
XFILLER_0_110 vgnd vpwr scs8hd_decap_6
XFILLER_0_198 vgnd vpwr scs8hd_decap_6
XFILLER_0_187 vgnd vpwr scs8hd_decap_3
XFILLER_5_21 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_9.LATCH_0_.latch data_in _112_/A _166_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_65 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _110_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_84 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _114_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_180 vgnd vpwr scs8hd_decap_3
XFILLER_19_19 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_13.INVTX1_0_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_227 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__202__A _202_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_106 vpwr vgnd scs8hd_fill_2
XFILLER_18_117 vpwr vgnd scs8hd_fill_2
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_84 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_73 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
X_195_ _195_/HI _195_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__112__A _112_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_66 vpwr vgnd scs8hd_fill_2
XFILLER_32_186 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _191_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_175 vgnd vpwr scs8hd_decap_8
XFILLER_11_53 vpwr vgnd scs8hd_fill_2
XFILLER_11_97 vpwr vgnd scs8hd_fill_2
XANTENNA__107__A _107_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_186 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_178_ _178_/HI _178_/LO vgnd vpwr scs8hd_conb_1
XFILLER_28_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_134 vgnd vpwr scs8hd_decap_4
XFILLER_20_167 vgnd vpwr scs8hd_decap_12
XFILLER_7_138 vgnd vpwr scs8hd_decap_4
XFILLER_11_123 vgnd vpwr scs8hd_decap_12
X_101_ _101_/A _101_/Y vgnd vpwr scs8hd_inv_8
XFILLER_22_63 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ _108_/A mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_19_201 vgnd vpwr scs8hd_decap_12
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_6_171 vgnd vpwr scs8hd_decap_12
XFILLER_8_21 vgnd vpwr scs8hd_decap_4
XFILLER_8_65 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _112_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_19 vgnd vpwr scs8hd_decap_4
XANTENNA__210__A _210_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _093_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _116_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_33_95 vgnd vpwr scs8hd_fill_1
XANTENNA__120__A _120_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB _177_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_1_ mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_track_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__205__A _205_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_133 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ _206_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _185_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_55 vpwr vgnd scs8hd_fill_2
XANTENNA__115__A _115_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ _112_/Y mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_10_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _187_/HI vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_track_17.LATCH_0_.latch data_in _120_/A _177_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_41 vgnd vpwr scs8hd_decap_12
XFILLER_30_30 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_74 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr
+ scs8hd_diode_2
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_25_96 vpwr vgnd scs8hd_fill_2
X_194_ _194_/HI _194_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_89 vgnd vpwr scs8hd_decap_3
XFILLER_2_56 vpwr vgnd scs8hd_fill_2
XFILLER_2_23 vgnd vpwr scs8hd_decap_4
XFILLER_32_154 vgnd vpwr scs8hd_decap_12
XFILLER_32_132 vgnd vpwr scs8hd_decap_12
XFILLER_17_184 vpwr vgnd scs8hd_fill_2
XFILLER_17_195 vpwr vgnd scs8hd_fill_2
XFILLER_32_198 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_15.LATCH_1_.latch_SLEEPB _174_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_21 vgnd vpwr scs8hd_decap_3
XANTENNA__213__A _213_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_11.INVTX1_0_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_110 vgnd vpwr scs8hd_decap_8
XFILLER_14_154 vgnd vpwr scs8hd_decap_12
X_177_ _127_/D _175_/B address[0] _177_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_14_198 vgnd vpwr scs8hd_decap_12
XANTENNA__123__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_20_179 vpwr vgnd scs8hd_fill_2
XFILLER_28_202 vgnd vpwr scs8hd_decap_12
X_100_ _100_/A _100_/Y vgnd vpwr scs8hd_inv_8
XFILLER_11_135 vgnd vpwr scs8hd_fill_1
XANTENNA__208__A _208_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_75 vgnd vpwr scs8hd_decap_4
XFILLER_19_213 vgnd vpwr scs8hd_decap_12
XFILLER_34_227 vgnd vpwr scs8hd_decap_6
XANTENNA__118__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_183 vgnd vpwr scs8hd_decap_12
XFILLER_10_190 vgnd vpwr scs8hd_decap_6
XFILLER_16_205 vgnd vpwr scs8hd_decap_8
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_52 vpwr vgnd scs8hd_fill_2
XFILLER_33_30 vpwr vgnd scs8hd_fill_2
XFILLER_31_208 vgnd vpwr scs8hd_decap_12
XFILLER_17_53 vgnd vpwr scs8hd_decap_4
XFILLER_3_153 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_230 vgnd vpwr scs8hd_decap_3
XFILLER_13_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _086_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_178 vpwr vgnd scs8hd_fill_2
XFILLER_0_145 vgnd vpwr scs8hd_decap_8
XFILLER_0_123 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_85 vgnd vpwr scs8hd_decap_4
XFILLER_28_41 vgnd vpwr scs8hd_decap_12
XFILLER_28_30 vgnd vpwr scs8hd_fill_1
XFILLER_5_34 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _181_/HI vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ _114_/Y mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__131__A _128_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[8] mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_10 vpwr vgnd scs8hd_fill_2
XFILLER_14_32 vpwr vgnd scs8hd_fill_2
XFILLER_30_53 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_160 vgnd vpwr scs8hd_decap_12
XANTENNA__126__A address[1] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_5.LATCH_0_.latch data_in _108_/A _160_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_141 vgnd vpwr scs8hd_decap_12
XFILLER_26_130 vpwr vgnd scs8hd_fill_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_25_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A right_bottom_grid_pin_12_ vgnd
+ vpwr scs8hd_diode_2
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_75 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_193_ _193_/HI _193_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mem_bottom_track_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_35 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1_A bottom_left_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_32_166 vgnd vpwr scs8hd_decap_12
XFILLER_32_144 vgnd vpwr scs8hd_decap_8
XFILLER_32_100 vgnd vpwr scs8hd_decap_6
XFILLER_17_152 vpwr vgnd scs8hd_fill_2
XFILLER_23_199 vgnd vpwr scs8hd_decap_12
XFILLER_11_77 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _103_/A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_14_166 vgnd vpwr scs8hd_decap_6
X_176_ _127_/D _175_/B _128_/A _176_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA__123__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_7_107 vpwr vgnd scs8hd_fill_2
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_43 vgnd vpwr scs8hd_decap_8
XFILLER_0_3 vgnd vpwr scs8hd_decap_4
XFILLER_19_225 vgnd vpwr scs8hd_decap_8
XANTENNA__134__A _128_/A vgnd vpwr scs8hd_diode_2
X_159_ _128_/A _158_/X _159_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_195 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr
+ scs8hd_diode_2
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_132 vpwr vgnd scs8hd_fill_2
XFILLER_3_176 vgnd vpwr scs8hd_decap_4
XANTENNA__129__A address[0] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _184_/HI _107_/Y mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_220 vgnd vpwr scs8hd_decap_12
XFILLER_28_20 vgnd vpwr scs8hd_decap_4
XFILLER_28_53 vgnd vpwr scs8hd_decap_3
XFILLER_8_202 vgnd vpwr scs8hd_decap_12
XANTENNA__131__B _131_/B vgnd vpwr scs8hd_diode_2
XFILLER_14_66 vpwr vgnd scs8hd_fill_2
XFILLER_14_88 vpwr vgnd scs8hd_fill_2
XFILLER_29_172 vgnd vpwr scs8hd_decap_8
XANTENNA__126__B enable vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _167_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_208 vgnd vpwr scs8hd_decap_6
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_76 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
X_192_ _192_/HI _192_/LO vgnd vpwr scs8hd_conb_1
Xmux_right_track_14.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[0] mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_bottom_track_13.LATCH_0_.latch data_in _116_/A _172_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB _166_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_131 vpwr vgnd scs8hd_fill_2
XFILLER_32_178 vgnd vpwr scs8hd_decap_4
XFILLER_17_175 vgnd vpwr scs8hd_decap_4
XANTENNA__137__A _128_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _101_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_112 vpwr vgnd scs8hd_fill_2
XFILLER_23_134 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_7 vgnd vpwr scs8hd_fill_1
XFILLER_14_134 vgnd vpwr scs8hd_decap_4
X_175_ _167_/D _175_/B address[0] _175_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA__123__C _123_/C vgnd vpwr scs8hd_diode_2
XFILLER_9_182 vgnd vpwr scs8hd_fill_1
XFILLER_20_115 vgnd vpwr scs8hd_decap_4
XFILLER_28_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_158_ address[3] _167_/B _167_/C _127_/D _158_/X vgnd vpwr scs8hd_or4_4
XANTENNA__134__B _135_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_141 vgnd vpwr scs8hd_decap_3
XFILLER_6_152 vgnd vpwr scs8hd_fill_1
X_089_ _089_/A _089_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _109_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_26_3 vgnd vpwr scs8hd_decap_3
XANTENNA__150__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_11 vgnd vpwr scs8hd_decap_3
XFILLER_17_77 vpwr vgnd scs8hd_fill_2
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_98 vgnd vpwr scs8hd_decap_3
XFILLER_33_87 vpwr vgnd scs8hd_fill_2
XFILLER_33_65 vpwr vgnd scs8hd_fill_2
XFILLER_33_10 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _113_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__129__B _129_/B vgnd vpwr scs8hd_diode_2
XANTENNA__145__A _167_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ _106_/A mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_0_80 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_7.LATCH_1_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_232 vgnd vpwr scs8hd_fill_1
XFILLER_28_65 vpwr vgnd scs8hd_fill_2
XFILLER_5_69 vpwr vgnd scs8hd_fill_2
XFILLER_30_11 vpwr vgnd scs8hd_fill_2
XFILLER_14_23 vpwr vgnd scs8hd_fill_2
XFILLER_14_45 vpwr vgnd scs8hd_fill_2
XFILLER_30_88 vgnd vpwr scs8hd_fill_1
XFILLER_29_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__142__B _167_/B vgnd vpwr scs8hd_diode_2
XFILLER_35_187 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ _110_/Y mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_77 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_25_11 vpwr vgnd scs8hd_fill_2
XFILLER_25_77 vpwr vgnd scs8hd_fill_2
X_191_ _191_/HI _191_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _111_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__137__B _138_/B vgnd vpwr scs8hd_diode_2
XANTENNA__153__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_13 vpwr vgnd scs8hd_fill_2
XFILLER_11_35 vgnd vpwr scs8hd_decap_3
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _115_/A vgnd
+ vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_0_.latch data_in _104_/A _154_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_102 vpwr vgnd scs8hd_fill_2
X_174_ _167_/D _175_/B _128_/A _174_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA__123__D _167_/D vgnd vpwr scs8hd_diode_2
XANTENNA__148__A address[4] vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[1] mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_227 vgnd vpwr scs8hd_decap_6
XFILLER_11_138 vgnd vpwr scs8hd_decap_12
XFILLER_22_23 vgnd vpwr scs8hd_decap_6
X_157_ address[0] _156_/B _157_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_8_69 vpwr vgnd scs8hd_fill_2
X_088_ _088_/A _088_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__150__B _151_/B vgnd vpwr scs8hd_diode_2
XFILLER_25_208 vgnd vpwr scs8hd_decap_12
XFILLER_19_3 vgnd vpwr scs8hd_decap_3
XFILLER_33_230 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _085_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_219 vgnd vpwr scs8hd_decap_12
XFILLER_33_22 vgnd vpwr scs8hd_decap_8
Xmem_right_track_16.LATCH_0_.latch data_in _102_/A _151_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_209_ _209_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA__161__A _167_/A vgnd vpwr scs8hd_diode_2
XANTENNA__145__B _167_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_90 vpwr vgnd scs8hd_fill_2
XFILLER_8_215 vgnd vpwr scs8hd_decap_12
XFILLER_5_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _186_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__156__A _128_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_10.tap_buf4_0_.scs8hd_inv_1 mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ _199_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _192_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__142__C _123_/C vgnd vpwr scs8hd_diode_2
XFILLER_35_199 vgnd vpwr scs8hd_decap_12
XFILLER_6_80 vpwr vgnd scs8hd_fill_2
XPHY_12 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_78 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
X_190_ _190_/HI _190_/LO vgnd vpwr scs8hd_conb_1
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XFILLER_25_34 vpwr vgnd scs8hd_fill_2
XFILLER_2_27 vgnd vpwr scs8hd_fill_1
XFILLER_17_111 vpwr vgnd scs8hd_fill_2
XFILLER_17_199 vgnd vpwr scs8hd_decap_4
XANTENNA__153__B _152_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _088_/A vgnd vpwr
+ scs8hd_diode_2
X_173_ address[3] address[2] address[4] _173_/D _175_/B vgnd vpwr scs8hd_or4_4
XFILLER_28_8 vgnd vpwr scs8hd_decap_3
XANTENNA__148__B _173_/D vgnd vpwr scs8hd_diode_2
XFILLER_9_184 vgnd vpwr scs8hd_decap_12
XANTENNA__164__A _167_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_81 vgnd vpwr scs8hd_decap_4
X_087_ _087_/A _087_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_154 vgnd vpwr scs8hd_decap_3
X_156_ _128_/A _156_/B _156_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_150 vgnd vpwr scs8hd_decap_3
XFILLER_33_6 vpwr vgnd scs8hd_fill_2
XANTENNA__159__A _128_/A vgnd vpwr scs8hd_diode_2
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_10.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[2] mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_33_56 vgnd vpwr scs8hd_decap_4
XFILLER_3_102 vpwr vgnd scs8hd_fill_2
XFILLER_3_157 vpwr vgnd scs8hd_fill_2
XANTENNA__145__C _123_/C vgnd vpwr scs8hd_diode_2
XANTENNA__161__B address[2] vgnd vpwr scs8hd_diode_2
X_139_ _167_/A address[2] _123_/C _127_/D _140_/B vgnd vpwr scs8hd_or4_4
X_208_ _208_/A chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
Xmux_right_track_4.tap_buf4_0_.scs8hd_inv_1 mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ _202_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_116 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_10.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_8_227 vgnd vpwr scs8hd_decap_6
XFILLER_5_38 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _182_/HI vgnd
+ vpwr scs8hd_diode_2
XANTENNA__156__B _156_/B vgnd vpwr scs8hd_diode_2
XANTENNA__172__A address[0] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _183_/HI _105_/Y mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ _212_/A vgnd vpwr scs8hd_inv_1
XFILLER_30_68 vgnd vpwr scs8hd_decap_12
XFILLER_5_208 vgnd vpwr scs8hd_decap_12
XANTENNA__082__A address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__142__D _167_/D vgnd vpwr scs8hd_diode_2
XFILLER_20_90 vpwr vgnd scs8hd_fill_2
XFILLER_35_156 vgnd vpwr scs8hd_decap_12
XANTENNA__167__A _167_/A vgnd vpwr scs8hd_diode_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XPHY_79 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
XFILLER_9_3 vgnd vpwr scs8hd_fill_1
XFILLER_2_39 vgnd vpwr scs8hd_decap_6
XFILLER_32_115 vgnd vpwr scs8hd_decap_8
XFILLER_17_123 vgnd vpwr scs8hd_fill_1
XFILLER_17_167 vpwr vgnd scs8hd_fill_2
XFILLER_31_192 vpwr vgnd scs8hd_fill_2
XFILLER_31_170 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _093_/A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_9.LATCH_1_.latch data_in _111_/A _165_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_track_11.LATCH_0_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
X_172_ address[0] _170_/X _172_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_152 vgnd vpwr scs8hd_decap_12
XANTENNA__164__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_13_170 vgnd vpwr scs8hd_fill_1
XFILLER_9_196 vgnd vpwr scs8hd_fill_1
XANTENNA__090__A _090_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_27 vpwr vgnd scs8hd_fill_2
XFILLER_8_49 vgnd vpwr scs8hd_fill_1
X_155_ address[3] _167_/B _167_/C _167_/D _156_/B vgnd vpwr scs8hd_or4_4
XFILLER_6_133 vgnd vpwr scs8hd_decap_8
X_086_ _086_/A _086_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__159__B _158_/X vgnd vpwr scs8hd_diode_2
XANTENNA__175__A _167_/D vgnd vpwr scs8hd_diode_2
XFILLER_17_25 vpwr vgnd scs8hd_fill_2
XFILLER_17_36 vpwr vgnd scs8hd_fill_2
XFILLER_33_35 vpwr vgnd scs8hd_fill_2
XANTENNA__085__A _085_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_114 vpwr vgnd scs8hd_fill_2
XFILLER_3_136 vgnd vpwr scs8hd_decap_4
XFILLER_15_210 vgnd vpwr scs8hd_decap_4
XFILLER_30_202 vgnd vpwr scs8hd_decap_12
X_207_ _207_/A chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA__145__D _127_/D vgnd vpwr scs8hd_diode_2
X_138_ address[0] _138_/B _138_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__161__C _167_/C vgnd vpwr scs8hd_diode_2
XFILLER_2_180 vpwr vgnd scs8hd_fill_2
XFILLER_24_3 vpwr vgnd scs8hd_fill_2
XFILLER_0_72 vgnd vpwr scs8hd_decap_6
XFILLER_0_94 vgnd vpwr scs8hd_decap_4
XFILLER_12_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_17 vpwr vgnd scs8hd_fill_2
Xmem_right_track_12.LATCH_0_.latch data_in _098_/A _144_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__172__B _170_/X vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ _104_/A mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_29_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _112_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _101_/A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_35_168 vgnd vpwr scs8hd_decap_12
XANTENNA__167__B _167_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _116_/Y vgnd
+ vpwr scs8hd_diode_2
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_157 vgnd vpwr scs8hd_decap_12
XFILLER_26_124 vgnd vpwr scs8hd_decap_4
XFILLER_26_102 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XFILLER_34_190 vgnd vpwr scs8hd_decap_12
XANTENNA__093__A _093_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_135 vpwr vgnd scs8hd_fill_2
XFILLER_23_116 vgnd vpwr scs8hd_decap_4
XFILLER_23_138 vpwr vgnd scs8hd_fill_2
XFILLER_31_182 vgnd vpwr scs8hd_fill_1
XANTENNA__088__A _088_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_149 vgnd vpwr scs8hd_decap_4
X_171_ _128_/A _170_/X _171_/Y vgnd vpwr scs8hd_nor2_4
Xmux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ _108_/Y mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_17.LATCH_1_.latch data_in _119_/A _176_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_120 vpwr vgnd scs8hd_fill_2
XFILLER_9_164 vgnd vpwr scs8hd_decap_12
XANTENNA__164__C _167_/C vgnd vpwr scs8hd_diode_2
XFILLER_13_182 vgnd vpwr scs8hd_fill_1
XFILLER_3_50 vpwr vgnd scs8hd_fill_2
XFILLER_22_15 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_17 vpwr vgnd scs8hd_fill_2
XFILLER_10_130 vgnd vpwr scs8hd_decap_12
X_154_ address[0] _152_/X _154_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_196 vgnd vpwr scs8hd_fill_1
X_085_ _085_/A _085_/Y vgnd vpwr scs8hd_inv_8
XFILLER_33_222 vgnd vpwr scs8hd_decap_8
XANTENNA__175__B _175_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ _208_/A vgnd vpwr scs8hd_inv_1
XFILLER_17_59 vpwr vgnd scs8hd_fill_2
XFILLER_33_69 vgnd vpwr scs8hd_decap_12
XFILLER_33_47 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_0_.latch data_in _094_/A _138_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_206_ _206_/A chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
X_137_ _128_/A _138_/B _137_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__161__D _167_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _118_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_129 vpwr vgnd scs8hd_fill_2
XFILLER_28_69 vgnd vpwr scs8hd_decap_12
XANTENNA__096__A _096_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _096_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_14_27 vpwr vgnd scs8hd_fill_2
XFILLER_14_49 vpwr vgnd scs8hd_fill_2
XFILLER_35_125 vgnd vpwr scs8hd_decap_12
XANTENNA__167__C _167_/C vgnd vpwr scs8hd_diode_2
XFILLER_6_61 vgnd vpwr scs8hd_decap_8
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_26_169 vgnd vpwr scs8hd_decap_12
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XFILLER_25_15 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _104_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_19 vpwr vgnd scs8hd_fill_2
XFILLER_25_180 vgnd vpwr scs8hd_decap_3
XFILLER_15_92 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _086_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_17 vpwr vgnd scs8hd_fill_2
XFILLER_14_106 vpwr vgnd scs8hd_fill_2
X_170_ _167_/A _167_/B _167_/C _127_/D _170_/X vgnd vpwr scs8hd_or4_4
XFILLER_22_194 vgnd vpwr scs8hd_decap_8
XFILLER_9_176 vgnd vpwr scs8hd_decap_6
XANTENNA__164__D _127_/D vgnd vpwr scs8hd_diode_2
XFILLER_3_62 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.INVTX1_1_.scs8hd_inv_1 bottom_left_grid_pin_7_ mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_9 vpwr vgnd scs8hd_fill_2
XANTENNA__099__A _099_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_220 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_5.LATCH_1_.latch data_in _107_/A _159_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_142 vgnd vpwr scs8hd_decap_8
X_153_ _128_/A _152_/X _153_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_146 vgnd vpwr scs8hd_decap_6
XFILLER_12_60 vgnd vpwr scs8hd_decap_6
X_084_ address[0] _128_/A vgnd vpwr scs8hd_inv_8
XANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_18_231 vpwr vgnd scs8hd_fill_2
XANTENNA__175__C address[0] vgnd vpwr scs8hd_diode_2
X_205_ _205_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
X_136_ _167_/A address[2] _123_/C _167_/D _138_/B vgnd vpwr scs8hd_or4_4
XFILLER_23_81 vgnd vpwr scs8hd_decap_12
XFILLER_0_85 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_track_3.LATCH_0_.latch_SLEEPB _157_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_94 vpwr vgnd scs8hd_fill_2
XFILLER_21_204 vpwr vgnd scs8hd_fill_2
XFILLER_28_26 vgnd vpwr scs8hd_decap_4
XFILLER_0_119 vgnd vpwr scs8hd_decap_4
XFILLER_12_215 vgnd vpwr scs8hd_decap_12
XFILLER_18_70 vgnd vpwr scs8hd_decap_3
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _087_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
X_119_ _119_/A _119_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__197__A _197_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _193_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_211 vgnd vpwr scs8hd_decap_3
XFILLER_20_71 vgnd vpwr scs8hd_decap_4
XFILLER_20_93 vgnd vpwr scs8hd_decap_4
XFILLER_35_137 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__167__D _167_/D vgnd vpwr scs8hd_diode_2
XFILLER_6_73 vpwr vgnd scs8hd_fill_2
XFILLER_6_84 vgnd vpwr scs8hd_decap_8
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_25_38 vgnd vpwr scs8hd_decap_4
XFILLER_1_203 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _178_/HI _103_/Y mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_115 vpwr vgnd scs8hd_fill_2
XFILLER_17_148 vpwr vgnd scs8hd_fill_2
XFILLER_15_71 vpwr vgnd scs8hd_fill_2
XFILLER_16_192 vpwr vgnd scs8hd_fill_2
XFILLER_31_184 vgnd vpwr scs8hd_fill_1
XFILLER_14_118 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB _153_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_3 vgnd vpwr scs8hd_fill_1
XFILLER_13_140 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1_A bottom_left_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_199 vgnd vpwr scs8hd_decap_12
XFILLER_13_184 vgnd vpwr scs8hd_decap_12
XFILLER_27_232 vgnd vpwr scs8hd_fill_1
X_083_ enable _083_/Y vgnd vpwr scs8hd_inv_8
X_152_ address[3] address[2] _167_/C _127_/D _152_/X vgnd vpwr scs8hd_or4_4
XFILLER_10_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _091_/A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_5_180 vgnd vpwr scs8hd_decap_3
Xmem_bottom_track_13.LATCH_1_.latch data_in _115_/A _171_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_24_202 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_7.INVTX1_1_.scs8hd_inv_1 bottom_left_grid_pin_5_ mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_106 vgnd vpwr scs8hd_decap_3
X_204_ _204_/A chanx_right_out[0] vgnd vpwr scs8hd_buf_2
X_135_ address[0] _135_/B _135_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_93 vpwr vgnd scs8hd_fill_2
XFILLER_31_7 vpwr vgnd scs8hd_fill_2
XFILLER_9_73 vgnd vpwr scs8hd_decap_6
XFILLER_12_227 vgnd vpwr scs8hd_decap_6
XFILLER_18_93 vpwr vgnd scs8hd_fill_2
XFILLER_7_220 vgnd vpwr scs8hd_decap_12
X_118_ _118_/A _118_/Y vgnd vpwr scs8hd_inv_8
XFILLER_22_3 vgnd vpwr scs8hd_decap_3
Xmem_right_track_4.LATCH_0_.latch data_in _090_/A _132_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_29_102 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A bottom_left_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_35_149 vgnd vpwr scs8hd_decap_6
XFILLER_28_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_15.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_1_215 vgnd vpwr scs8hd_decap_12
XFILLER_17_127 vpwr vgnd scs8hd_fill_2
XFILLER_31_71 vgnd vpwr scs8hd_decap_12
XFILLER_31_130 vpwr vgnd scs8hd_fill_2
XFILLER_31_196 vgnd vpwr scs8hd_decap_12
Xmux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _099_/A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_22_152 vgnd vpwr scs8hd_fill_1
XFILLER_9_123 vgnd vpwr scs8hd_decap_3
XFILLER_13_130 vgnd vpwr scs8hd_decap_8
XFILLER_13_152 vgnd vpwr scs8hd_decap_12
XFILLER_13_174 vpwr vgnd scs8hd_fill_2
XFILLER_13_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_20 vpwr vgnd scs8hd_fill_2
XFILLER_6_159 vgnd vpwr scs8hd_decap_12
XFILLER_10_166 vgnd vpwr scs8hd_decap_12
X_082_ address[2] _167_/B vgnd vpwr scs8hd_inv_8
X_151_ address[0] _151_/B _151_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_203 vgnd vpwr scs8hd_decap_12
XFILLER_18_211 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ _106_/Y mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_17_29 vpwr vgnd scs8hd_fill_2
XFILLER_33_39 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _111_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
XFILLER_15_214 vgnd vpwr scs8hd_fill_1
X_203_ _203_/A chanx_right_out[1] vgnd vpwr scs8hd_buf_2
X_134_ _128_/A _135_/B _134_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_184 vgnd vpwr scs8hd_decap_12
XFILLER_2_151 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_1.LATCH_1_.latch data_in _103_/A _153_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_24_7 vpwr vgnd scs8hd_fill_2
XFILLER_0_32 vpwr vgnd scs8hd_fill_2
XFILLER_0_43 vpwr vgnd scs8hd_fill_2
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XFILLER_0_98 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _115_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _138_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_50 vgnd vpwr scs8hd_fill_1
XFILLER_34_93 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_5.INVTX1_1_.scs8hd_inv_1 bottom_left_grid_pin_3_ mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_7_232 vgnd vpwr scs8hd_fill_1
X_117_ _117_/A _117_/Y vgnd vpwr scs8hd_inv_8
XFILLER_30_18 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _094_/A mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_29_136 vgnd vpwr scs8hd_decap_12
XFILLER_29_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_62 vpwr vgnd scs8hd_fill_2
XFILLER_20_84 vgnd vpwr scs8hd_decap_4
XFILLER_35_106 vgnd vpwr scs8hd_decap_12
XFILLER_29_71 vgnd vpwr scs8hd_decap_12
Xmem_right_track_16.LATCH_1_.latch data_in _101_/A _150_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_25_29 vgnd vpwr scs8hd_decap_3
XFILLER_1_227 vgnd vpwr scs8hd_decap_6
XFILLER_15_51 vpwr vgnd scs8hd_fill_2
XFILLER_31_83 vgnd vpwr scs8hd_fill_1
XANTENNA__102__A _102_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_142 vpwr vgnd scs8hd_fill_2
XFILLER_9_113 vgnd vpwr scs8hd_fill_1
XFILLER_13_164 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _117_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_98 vpwr vgnd scs8hd_fill_2
XFILLER_3_54 vgnd vpwr scs8hd_decap_4
XFILLER_3_43 vpwr vgnd scs8hd_fill_2
XFILLER_8_190 vgnd vpwr scs8hd_decap_12
XFILLER_22_19 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _095_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_10_123 vgnd vpwr scs8hd_decap_4
X_150_ _128_/A _151_/B _150_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_178 vgnd vpwr scs8hd_decap_12
XFILLER_12_52 vpwr vgnd scs8hd_fill_2
X_081_ address[3] _167_/A vgnd vpwr scs8hd_inv_8
XFILLER_24_215 vgnd vpwr scs8hd_decap_12
XANTENNA__200__A _200_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _088_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_218 vgnd vpwr scs8hd_decap_12
X_133_ address[3] _167_/B _123_/C _127_/D _135_/B vgnd vpwr scs8hd_or4_4
X_202_ _202_/A chanx_right_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_23_40 vpwr vgnd scs8hd_fill_2
XFILLER_23_51 vpwr vgnd scs8hd_fill_2
XFILLER_23_62 vgnd vpwr scs8hd_decap_12
XFILLER_2_163 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ _102_/A mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__110__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_196 vgnd vpwr scs8hd_decap_12
XFILLER_0_22 vgnd vpwr scs8hd_decap_3
XFILLER_17_7 vpwr vgnd scs8hd_fill_2
XFILLER_9_42 vpwr vgnd scs8hd_fill_2
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _103_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_84 vpwr vgnd scs8hd_fill_2
XANTENNA__105__A _105_/A vgnd vpwr scs8hd_diode_2
X_116_ _116_/A _116_/Y vgnd vpwr scs8hd_inv_8
XFILLER_29_148 vgnd vpwr scs8hd_decap_12
XFILLER_20_41 vgnd vpwr scs8hd_decap_12
XFILLER_35_118 vgnd vpwr scs8hd_decap_6
XFILLER_29_83 vgnd vpwr scs8hd_decap_4
XFILLER_6_32 vgnd vpwr scs8hd_decap_3
XFILLER_26_107 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_3.INVTX1_1_.scs8hd_inv_1 bottom_left_grid_pin_1_ mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_19 vgnd vpwr scs8hd_decap_3
Xmem_right_track_0.LATCH_0_.latch data_in _085_/A _125_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_107 vpwr vgnd scs8hd_fill_2
XFILLER_25_184 vgnd vpwr scs8hd_decap_12
XFILLER_15_41 vgnd vpwr scs8hd_fill_1
XFILLER_15_96 vpwr vgnd scs8hd_fill_2
XFILLER_31_95 vgnd vpwr scs8hd_decap_4
XFILLER_16_151 vpwr vgnd scs8hd_fill_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_110 vpwr vgnd scs8hd_fill_2
XFILLER_22_132 vgnd vpwr scs8hd_fill_1
XFILLER_22_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _090_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__203__A _203_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_84 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_110 vgnd vpwr scs8hd_decap_12
XANTENNA__113__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_77 vpwr vgnd scs8hd_fill_2
X_080_ address[5] _173_/D vgnd vpwr scs8hd_inv_8
XFILLER_6_106 vgnd vpwr scs8hd_decap_12
XFILLER_5_3 vgnd vpwr scs8hd_decap_4
Xmux_right_track_0.tap_buf4_0_.scs8hd_inv_1 mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _204_/A vgnd vpwr scs8hd_inv_1
XANTENNA__108__A _108_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_227 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_201_ _201_/A chanx_right_out[3] vgnd vpwr scs8hd_buf_2
X_132_ address[0] _131_/B _132_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_74 vgnd vpwr scs8hd_fill_1
Xmux_right_track_16.tap_buf4_0_.scs8hd_inv_1 mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _196_/A vgnd vpwr scs8hd_inv_1
XFILLER_21_208 vgnd vpwr scs8hd_decap_12
Xmux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _089_/A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__211__A _211_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_41 vgnd vpwr scs8hd_decap_3
X_115_ _115_/A _115_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__121__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA__206__A _206_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _194_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_20 vpwr vgnd scs8hd_fill_2
XFILLER_20_97 vgnd vpwr scs8hd_fill_1
XANTENNA__116__A _116_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_44 vpwr vgnd scs8hd_fill_2
XFILLER_20_3 vgnd vpwr scs8hd_decap_3
XFILLER_19_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _195_/HI _093_/Y mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_119 vgnd vpwr scs8hd_decap_3
XFILLER_25_196 vgnd vpwr scs8hd_decap_12
XFILLER_15_75 vpwr vgnd scs8hd_fill_2
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_188 vpwr vgnd scs8hd_fill_2
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

