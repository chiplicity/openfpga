* NGSPICE file created from cby_1__1_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_dfxbp_1 abstract view
.subckt scs8hd_dfxbp_1 CLK D Q QN vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_mux2_1 abstract view
.subckt scs8hd_mux2_1 A0 A1 S X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

.subckt cby_1__1_ ccff_head ccff_tail chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11]
+ chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14] chany_bottom_in[15]
+ chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18] chany_bottom_in[19]
+ chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5]
+ chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_in[9] chany_bottom_out[0]
+ chany_bottom_out[10] chany_bottom_out[11] chany_bottom_out[12] chany_bottom_out[13]
+ chany_bottom_out[14] chany_bottom_out[15] chany_bottom_out[16] chany_bottom_out[17]
+ chany_bottom_out[18] chany_bottom_out[19] chany_bottom_out[1] chany_bottom_out[2]
+ chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6]
+ chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9] chany_top_in[0] chany_top_in[10]
+ chany_top_in[11] chany_top_in[12] chany_top_in[13] chany_top_in[14] chany_top_in[15]
+ chany_top_in[16] chany_top_in[17] chany_top_in[18] chany_top_in[19] chany_top_in[1]
+ chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6]
+ chany_top_in[7] chany_top_in[8] chany_top_in[9] chany_top_out[0] chany_top_out[10]
+ chany_top_out[11] chany_top_out[12] chany_top_out[13] chany_top_out[14] chany_top_out[15]
+ chany_top_out[16] chany_top_out[17] chany_top_out[18] chany_top_out[19] chany_top_out[1]
+ chany_top_out[2] chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6]
+ chany_top_out[7] chany_top_out[8] chany_top_out[9] left_grid_pin_0_ left_grid_pin_10_
+ left_grid_pin_11_ left_grid_pin_12_ left_grid_pin_13_ left_grid_pin_14_ left_grid_pin_15_
+ left_grid_pin_1_ left_grid_pin_2_ left_grid_pin_3_ left_grid_pin_4_ left_grid_pin_5_
+ left_grid_pin_6_ left_grid_pin_7_ left_grid_pin_8_ left_grid_pin_9_ prog_clk right_grid_pin_52_
+ vpwr vgnd
XANTENNA_mux_right_ipin_1.mux_l3_in_0__A1 mux_right_ipin_1.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_85 vgnd vpwr scs8hd_decap_3
XFILLER_42_40 vgnd vpwr scs8hd_decap_4
XFILLER_13_144 vpwr vgnd scs8hd_fill_2
XFILLER_3_45 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.mux_l2_in_1__A1 mux_left_ipin_0.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_63_39 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_ipin_3.mux_l2_in_0__S mux_right_ipin_3.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_125 vpwr vgnd scs8hd_fill_2
XFILLER_12_10 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_4.scs8hd_dfxbp_1_1_ prog_clk mux_right_ipin_4.mux_l1_in_2_/S mux_right_ipin_4.mux_l2_in_3_/S
+ mem_right_ipin_4.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_ipin_8.mux_l4_in_0__A0 mux_right_ipin_8.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_11.mux_l2_in_0_ chany_bottom_in[2] mux_right_ipin_11.mux_l1_in_0_/X
+ mux_right_ipin_11.mux_l2_in_3_/S mux_right_ipin_11.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_37_62 vpwr vgnd scs8hd_fill_2
XFILLER_37_73 vpwr vgnd scs8hd_fill_2
XFILLER_53_50 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_ipin_0.mux_l2_in_0__S mux_left_ipin_0.mux_l2_in_2_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_4.scs8hd_dfxbp_1_2__D mux_right_ipin_4.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_9.mux_l1_in_1__S mux_right_ipin_9.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
X_66_ chany_bottom_in[7] chany_top_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_59_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_2.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_23_53 vpwr vgnd scs8hd_fill_2
XFILLER_23_75 vgnd vpwr scs8hd_decap_4
XFILLER_48_50 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.mux_l3_in_0__A1 mux_left_ipin_0.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_9_22 vgnd vpwr scs8hd_decap_12
XFILLER_9_77 vpwr vgnd scs8hd_fill_2
XFILLER_9_99 vpwr vgnd scs8hd_fill_2
X_49_ chany_top_in[4] chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_ipin_2.mux_l3_in_0__S mux_right_ipin_2.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_62_109 vgnd vpwr scs8hd_decap_12
XFILLER_18_42 vpwr vgnd scs8hd_fill_2
XFILLER_18_64 vgnd vpwr scs8hd_fill_1
XFILLER_18_97 vgnd vpwr scs8hd_fill_1
XFILLER_50_40 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_8.mux_l2_in_1__S mux_right_ipin_8.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_8.mux_l2_in_2__A1 chany_top_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_20_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_11.mux_l1_in_0__S mux_right_ipin_11.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_45_84 vpwr vgnd scs8hd_fill_2
XFILLER_6_23 vpwr vgnd scs8hd_fill_2
XFILLER_6_78 vgnd vpwr scs8hd_fill_1
XFILLER_6_45 vgnd vpwr scs8hd_fill_1
Xmem_right_ipin_14.scs8hd_dfxbp_1_2_ prog_clk mux_right_ipin_14.mux_l2_in_2_/S mux_right_ipin_14.mux_l3_in_0_/S
+ mem_right_ipin_14.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_ipin_3.mux_l2_in_3__S mux_right_ipin_3.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_11.mux_l2_in_0__A1 mux_right_ipin_11.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_1.mux_l4_in_0__S mux_right_ipin_1.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_31_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.mux_l2_in_3__S mux_left_ipin_0.mux_l2_in_2_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_5.mux_l1_in_1__A0 chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_8.mux_l3_in_1__A1 mux_right_ipin_8.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_15.scs8hd_buf_4_0__A mux_right_ipin_15.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_right_ipin_6.scs8hd_dfxbp_1_1__D mux_right_ipin_6.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.mux_l3_in_1__S mux_right_ipin_7.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_112 vpwr vgnd scs8hd_fill_2
XFILLER_26_42 vgnd vpwr scs8hd_decap_3
XFILLER_26_64 vpwr vgnd scs8hd_fill_2
XFILLER_26_75 vgnd vpwr scs8hd_decap_8
XFILLER_26_97 vgnd vpwr scs8hd_decap_3
XFILLER_42_63 vgnd vpwr scs8hd_decap_8
XFILLER_42_30 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_10.mux_l2_in_0__S mux_right_ipin_10.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_57 vpwr vgnd scs8hd_fill_2
XFILLER_3_13 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_5.mux_l2_in_0__A0 mux_right_ipin_5.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_right_ipin_4.scs8hd_dfxbp_1_0_ prog_clk mux_right_ipin_3.mux_l4_in_0_/S mux_right_ipin_4.mux_l1_in_2_/S
+ mem_right_ipin_4.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_ipin_8.mux_l4_in_0__A1 mux_right_ipin_8.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_30 vpwr vgnd scs8hd_fill_2
XFILLER_53_84 vgnd vpwr scs8hd_fill_1
XFILLER_53_62 vgnd vpwr scs8hd_decap_6
X_65_ chany_bottom_in[8] chany_top_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_23_21 vgnd vpwr scs8hd_fill_1
XFILLER_23_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_3.mux_l2_in_2__A0 chany_bottom_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_48_84 vgnd vpwr scs8hd_decap_6
XFILLER_64_94 vgnd vpwr scs8hd_decap_12
XFILLER_0_36 vgnd vpwr scs8hd_decap_4
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
X_48_ chany_top_in[5] chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_60_19 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_11.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_11.mux_l1_in_0_/S
+ mux_right_ipin_11.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_15.mux_l2_in_1__S mux_right_ipin_15.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_32 vgnd vpwr scs8hd_decap_8
XFILLER_34_42 vpwr vgnd scs8hd_fill_2
XFILLER_34_86 vgnd vpwr scs8hd_decap_4
XFILLER_34_97 vgnd vpwr scs8hd_fill_1
XFILLER_50_85 vgnd vpwr scs8hd_decap_6
XFILLER_38_129 vpwr vgnd scs8hd_fill_2
XFILLER_61_143 vgnd vpwr scs8hd_decap_3
XFILLER_61_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_ipin_8.scs8hd_dfxbp_1_0__D mux_right_ipin_7.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_107 vgnd vpwr scs8hd_decap_12
XFILLER_55_19 vgnd vpwr scs8hd_decap_12
XFILLER_52_132 vgnd vpwr scs8hd_decap_12
XFILLER_52_110 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_3.mux_l3_in_1__A0 mux_right_ipin_3.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_140 vgnd vpwr scs8hd_decap_6
XFILLER_20_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_7.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_43_143 vgnd vpwr scs8hd_decap_3
XFILLER_43_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_10.mux_l2_in_3__S mux_right_ipin_10.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_61_40 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_ipin_5.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_14.scs8hd_dfxbp_1_1_ prog_clk mux_right_ipin_14.mux_l1_in_0_/S mux_right_ipin_14.mux_l2_in_2_/S
+ mem_right_ipin_14.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_ipin_14.mux_l3_in_1__S mux_right_ipin_14.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_33 vpwr vgnd scs8hd_fill_2
XFILLER_15_55 vpwr vgnd scs8hd_fill_2
XFILLER_15_66 vgnd vpwr scs8hd_decap_4
XFILLER_25_121 vgnd vpwr scs8hd_fill_1
XFILLER_25_143 vgnd vpwr scs8hd_decap_3
XFILLER_40_102 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_5.mux_l1_in_1__A1 chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_ipin_3.mux_l4_in_0__A0 mux_right_ipin_3.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_135 vgnd vpwr scs8hd_decap_8
XFILLER_22_135 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_ipin_14.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_15.mux_l1_in_0__A0 chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_0__S mux_right_ipin_0.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_32 vgnd vpwr scs8hd_decap_4
XFILLER_26_54 vgnd vpwr scs8hd_decap_4
XFILLER_42_97 vgnd vpwr scs8hd_fill_1
XFILLER_42_75 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_ipin_12.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_2.scs8hd_buf_4_0__A mux_right_ipin_2.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_5.mux_l2_in_0__A1 mux_right_ipin_5.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_23 vgnd vpwr scs8hd_decap_8
XFILLER_12_67 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_13.mux_l1_in_2__A0 chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_37_53 vpwr vgnd scs8hd_fill_2
XFILLER_53_96 vpwr vgnd scs8hd_fill_2
XFILLER_53_74 vpwr vgnd scs8hd_fill_2
XFILLER_5_120 vpwr vgnd scs8hd_fill_2
X_64_ chany_bottom_in[9] chany_top_out[9] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_right_ipin_10.scs8hd_dfxbp_1_1__D mux_right_ipin_10.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_38_6 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_3.mux_l2_in_3_ _31_/HI chany_top_in[16] mux_right_ipin_3.mux_l2_in_3_/S
+ mux_right_ipin_3.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_ipin_8.scs8hd_dfxbp_1_3__D mux_right_ipin_8.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_3 vpwr vgnd scs8hd_fill_2
XFILLER_2_145 vgnd vpwr scs8hd_fill_1
XFILLER_2_101 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_3.mux_l2_in_2__A1 chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_0_15 vpwr vgnd scs8hd_fill_2
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
XFILLER_56_119 vgnd vpwr scs8hd_decap_3
X_47_ chany_top_in[6] chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_ipin_5.mux_l1_in_1__S mux_right_ipin_5.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_13.mux_l2_in_1__A0 chany_bottom_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_18_11 vgnd vpwr scs8hd_fill_1
XFILLER_18_22 vgnd vpwr scs8hd_decap_8
XFILLER_55_130 vgnd vpwr scs8hd_decap_12
XFILLER_34_32 vgnd vpwr scs8hd_decap_8
XFILLER_50_64 vpwr vgnd scs8hd_fill_2
XFILLER_34_65 vpwr vgnd scs8hd_fill_2
XFILLER_59_62 vgnd vpwr scs8hd_decap_4
XFILLER_59_51 vgnd vpwr scs8hd_decap_8
XFILLER_50_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.mux_l1_in_1__A0 chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_3.mux_l3_in_1__A1 mux_right_ipin_3.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_119 vgnd vpwr scs8hd_decap_3
XFILLER_52_144 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_8.scs8hd_buf_4_0_ mux_right_ipin_8.mux_l4_in_0_/X left_grid_pin_8_
+ vgnd vpwr scs8hd_buf_1
XFILLER_20_23 vgnd vpwr scs8hd_decap_8
XFILLER_29_10 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_11.mux_l2_in_3__A0 _25_/HI vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_3.mux_l4_in_0_ mux_right_ipin_3.mux_l3_in_1_/X mux_right_ipin_3.mux_l3_in_0_/X
+ mux_right_ipin_3.mux_l4_in_0_/S mux_right_ipin_3.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_29_54 vgnd vpwr scs8hd_decap_6
XFILLER_45_97 vpwr vgnd scs8hd_fill_2
XFILLER_45_75 vpwr vgnd scs8hd_fill_2
XFILLER_43_111 vpwr vgnd scs8hd_fill_2
XFILLER_20_6 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_13.mux_l3_in_0__A0 mux_right_ipin_13.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_100 vpwr vgnd scs8hd_fill_2
XFILLER_34_122 vgnd vpwr scs8hd_fill_1
XFILLER_34_133 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_14.scs8hd_dfxbp_1_0_ prog_clk mux_right_ipin_13.mux_l4_in_0_/S mux_right_ipin_14.mux_l1_in_0_/S
+ mem_right_ipin_14.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_ipin_4.mux_l2_in_1__S mux_right_ipin_4.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_31_88 vgnd vpwr scs8hd_decap_4
XFILLER_31_99 vgnd vpwr scs8hd_decap_3
XFILLER_56_96 vgnd vpwr scs8hd_decap_4
XFILLER_56_74 vpwr vgnd scs8hd_fill_2
XFILLER_56_30 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_0.mux_l2_in_0__A0 mux_right_ipin_0.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_ipin_3.mux_l4_in_0__A1 mux_right_ipin_3.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_ipin_8.mux_l2_in_3_ _19_/HI chany_top_in[19] mux_right_ipin_8.mux_l2_in_3_/S
+ mux_right_ipin_8.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_ipin_12.scs8hd_dfxbp_1_0__D mux_right_ipin_11.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_right_ipin_3.mux_l3_in_1_ mux_right_ipin_3.mux_l2_in_3_/X mux_right_ipin_3.mux_l2_in_2_/X
+ mux_right_ipin_3.mux_l3_in_1_/S mux_right_ipin_3.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_15.mux_l1_in_0__A1 chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_42_32 vgnd vpwr scs8hd_fill_1
XFILLER_9_107 vpwr vgnd scs8hd_fill_2
XFILLER_13_103 vpwr vgnd scs8hd_fill_2
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
XFILLER_13_136 vpwr vgnd scs8hd_fill_2
XFILLER_3_37 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_14.scs8hd_buf_4_0_ mux_right_ipin_14.mux_l4_in_0_/X left_grid_pin_14_
+ vgnd vpwr scs8hd_buf_1
XANTENNA_mux_right_ipin_3.mux_l3_in_1__S mux_right_ipin_3.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_13.mux_l1_in_2__A1 chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l3_in_1__S mux_left_ipin_0.mux_l3_in_1_/S vgnd vpwr scs8hd_diode_2
XFILLER_45_8 vpwr vgnd scs8hd_fill_2
X_63_ chany_bottom_in[10] chany_top_out[10] vgnd vpwr scs8hd_buf_2
Xmux_right_ipin_3.mux_l2_in_2_ chany_bottom_in[16] chany_top_in[8] mux_right_ipin_3.mux_l2_in_3_/S
+ mux_right_ipin_3.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_9.mux_l2_in_2__S mux_right_ipin_9.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_8.mux_l4_in_0_ mux_right_ipin_8.mux_l3_in_1_/X mux_right_ipin_8.mux_l3_in_0_/X
+ mux_right_ipin_8.mux_l4_in_0_/S mux_right_ipin_8.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_9.mux_l1_in_0__A0 chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_12.mux_l1_in_1__S mux_right_ipin_12.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_48_75 vgnd vpwr scs8hd_decap_3
XFILLER_0_27 vpwr vgnd scs8hd_fill_2
XFILLER_64_63 vgnd vpwr scs8hd_decap_12
XFILLER_9_36 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_7.scs8hd_dfxbp_1_3_ prog_clk mux_right_ipin_7.mux_l3_in_0_/S mux_right_ipin_7.mux_l4_in_0_/S
+ mem_right_ipin_7.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_50_6 vgnd vpwr scs8hd_decap_8
X_46_ chany_top_in[7] chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_ipin_13.mux_l2_in_1__A1 mux_right_ipin_13.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_55_142 vgnd vpwr scs8hd_decap_4
XFILLER_47_109 vpwr vgnd scs8hd_fill_2
XFILLER_18_89 vgnd vpwr scs8hd_decap_3
XFILLER_50_32 vpwr vgnd scs8hd_fill_2
XFILLER_50_21 vpwr vgnd scs8hd_fill_2
XFILLER_61_123 vgnd vpwr scs8hd_decap_12
XFILLER_61_101 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_12.scs8hd_dfxbp_1_3__D mux_right_ipin_12.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_right_ipin_8.mux_l3_in_1_ mux_right_ipin_8.mux_l2_in_3_/X mux_right_ipin_8.mux_l2_in_2_/X
+ mux_right_ipin_8.mux_l3_in_1_/S mux_right_ipin_8.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_0.mux_l1_in_1__A1 chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
X_29_ _29_/HI _29_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_ipin_11.mux_l2_in_3__A1 chany_top_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_20_68 vgnd vpwr scs8hd_fill_1
XFILLER_29_22 vgnd vpwr scs8hd_decap_3
XFILLER_45_43 vgnd vpwr scs8hd_decap_12
XFILLER_43_123 vgnd vpwr scs8hd_decap_12
XFILLER_29_99 vpwr vgnd scs8hd_fill_2
XFILLER_61_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_11.mux_l2_in_1__S mux_right_ipin_11.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_61_97 vpwr vgnd scs8hd_fill_2
XFILLER_6_48 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_13.mux_l3_in_0__A1 mux_right_ipin_13.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_6 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_10.mux_l1_in_0__A0 chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_34_145 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_7.mux_l2_in_1__A0 chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_25_123 vgnd vpwr scs8hd_decap_12
XFILLER_15_46 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.mux_l2_in_0__A1 mux_right_ipin_0.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_145 vgnd vpwr scs8hd_fill_1
XFILLER_31_115 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_8.mux_l2_in_2_ chany_bottom_in[19] chany_top_in[13] mux_right_ipin_8.mux_l2_in_3_/S
+ mux_right_ipin_8.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_3 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_3.mux_l3_in_0_ mux_right_ipin_3.mux_l2_in_1_/X mux_right_ipin_3.mux_l2_in_0_/X
+ mux_right_ipin_3.mux_l3_in_1_/S mux_right_ipin_3.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_5.mux_l2_in_3__A0 _33_/HI vgnd vpwr scs8hd_diode_2
XFILLER_42_22 vgnd vpwr scs8hd_decap_8
XFILLER_9_119 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_10.mux_l3_in_1__S mux_right_ipin_10.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_7.mux_l3_in_0__A0 mux_right_ipin_7.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_10.scs8hd_buf_4_0__A mux_right_ipin_10.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_77 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_62_ chany_bottom_in[11] chany_top_out[11] vgnd vpwr scs8hd_buf_2
Xmux_right_ipin_3.mux_l2_in_1_ chany_bottom_in[8] chany_top_in[2] mux_right_ipin_3.mux_l2_in_3_/S
+ mux_right_ipin_3.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_ipin_14.scs8hd_dfxbp_1_2__D mux_right_ipin_14.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_59_118 vpwr vgnd scs8hd_fill_2
XFILLER_4_81 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_9.mux_l1_in_0__A1 chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_23_24 vpwr vgnd scs8hd_fill_2
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
XFILLER_23_79 vgnd vpwr scs8hd_fill_1
XFILLER_48_32 vgnd vpwr scs8hd_decap_4
XFILLER_48_54 vpwr vgnd scs8hd_fill_2
XFILLER_64_75 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_3.scs8hd_buf_4_0_ mux_right_ipin_3.mux_l4_in_0_/X left_grid_pin_3_
+ vgnd vpwr scs8hd_buf_1
Xmem_right_ipin_7.scs8hd_dfxbp_1_2_ prog_clk mux_right_ipin_7.mux_l2_in_0_/S mux_right_ipin_7.mux_l3_in_0_/S
+ mem_right_ipin_7.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_43_6 vpwr vgnd scs8hd_fill_2
X_45_ chany_top_in[8] chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_18_46 vpwr vgnd scs8hd_fill_2
XFILLER_18_57 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_3.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_34_23 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_12.mux_l2_in_3_ _26_/HI chany_top_in[17] mux_right_ipin_12.mux_l2_in_0_/S
+ mux_right_ipin_12.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_61_135 vgnd vpwr scs8hd_decap_8
XFILLER_61_113 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_ipin_1.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_8.mux_l3_in_0_ mux_right_ipin_8.mux_l2_in_1_/X mux_right_ipin_8.mux_l2_in_0_/X
+ mux_right_ipin_8.mux_l3_in_1_/S mux_right_ipin_8.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
X_28_ _28_/HI _28_/LO vgnd vpwr scs8hd_conb_1
XFILLER_37_132 vpwr vgnd scs8hd_fill_2
XFILLER_52_102 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_ipin_1.scs8hd_dfxbp_1_1__D mux_right_ipin_1.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l1_in_1__S mux_right_ipin_1.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_43_135 vgnd vpwr scs8hd_decap_8
XFILLER_28_143 vgnd vpwr scs8hd_decap_3
XFILLER_61_10 vgnd vpwr scs8hd_decap_8
XFILLER_6_16 vgnd vpwr scs8hd_decap_3
XFILLER_6_27 vpwr vgnd scs8hd_fill_2
XFILLER_19_110 vgnd vpwr scs8hd_decap_4
XFILLER_19_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_10.mux_l1_in_0__A1 chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.mux_l2_in_1__A1 chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_25_113 vgnd vpwr scs8hd_decap_8
XFILLER_25_135 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_ipin_10.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_31_57 vpwr vgnd scs8hd_fill_2
XFILLER_56_32 vpwr vgnd scs8hd_fill_2
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_ipin_8.mux_l2_in_1_ chany_bottom_in[13] mux_right_ipin_8.mux_l1_in_2_/X
+ mux_right_ipin_8.mux_l2_in_3_/S mux_right_ipin_8.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_ipin_12.mux_l4_in_0_ mux_right_ipin_12.mux_l3_in_1_/X mux_right_ipin_12.mux_l3_in_0_/X
+ mux_right_ipin_12.mux_l4_in_0_/S mux_right_ipin_12.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_7_70 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_5.mux_l2_in_3__A1 chany_top_in[16] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l2_in_1__S mux_right_ipin_0.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l1_in_0__A0 chany_top_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.mux_l3_in_0__A1 mux_right_ipin_7.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_15.mux_l2_in_2__A0 chany_bottom_in[12] vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_8.mux_l1_in_2_ chany_top_in[9] chany_bottom_in[9] mux_right_ipin_8.mux_l1_in_2_/S
+ mux_right_ipin_8.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_53_33 vpwr vgnd scs8hd_fill_2
XFILLER_53_11 vgnd vpwr scs8hd_decap_3
XFILLER_5_145 vgnd vpwr scs8hd_fill_1
XFILLER_5_123 vpwr vgnd scs8hd_fill_2
XFILLER_5_112 vpwr vgnd scs8hd_fill_2
X_61_ chany_bottom_in[12] chany_top_out[12] vgnd vpwr scs8hd_buf_2
Xmux_right_ipin_12.mux_l3_in_1_ mux_right_ipin_12.mux_l2_in_3_/X mux_right_ipin_12.mux_l2_in_2_/X
+ mux_right_ipin_12.mux_l3_in_0_/S mux_right_ipin_12.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_ipin_3.mux_l2_in_0_ chany_bottom_in[2] mux_right_ipin_3.mux_l1_in_0_/X
+ mux_right_ipin_3.mux_l2_in_3_/S mux_right_ipin_3.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_93 vgnd vpwr scs8hd_decap_4
XFILLER_23_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_3.scs8hd_dfxbp_1_0__D mux_right_ipin_2.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_137 vgnd vpwr scs8hd_decap_8
XFILLER_2_126 vpwr vgnd scs8hd_fill_2
XFILLER_64_87 vgnd vpwr scs8hd_decap_6
XFILLER_64_32 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_7.scs8hd_dfxbp_1_1_ prog_clk mux_right_ipin_7.mux_l1_in_0_/S mux_right_ipin_7.mux_l2_in_0_/S
+ mem_right_ipin_7.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_ipin_15.mux_l3_in_1__A0 mux_right_ipin_15.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_80 vpwr vgnd scs8hd_fill_2
X_44_ chany_top_in[9] chany_bottom_out[9] vgnd vpwr scs8hd_buf_2
XFILLER_36_6 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_5.mux_l2_in_2__S mux_right_ipin_5.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_14 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_12.mux_l2_in_2_ chany_bottom_in[17] chany_top_in[13] mux_right_ipin_12.mux_l2_in_0_/S
+ mux_right_ipin_12.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_1_3 vgnd vpwr scs8hd_decap_4
XFILLER_59_87 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l2_in_1__A0 chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_46_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_9.mux_l3_in_0__S mux_right_ipin_9.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_3 vpwr vgnd scs8hd_fill_2
X_27_ _27_/HI _27_/LO vgnd vpwr scs8hd_conb_1
XFILLER_37_111 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_15.mux_l4_in_0__A0 mux_right_ipin_15.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_2__D mux_left_ipin_0.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_46 vpwr vgnd scs8hd_fill_2
XFILLER_29_68 vpwr vgnd scs8hd_fill_2
XFILLER_45_12 vpwr vgnd scs8hd_fill_2
XFILLER_61_66 vpwr vgnd scs8hd_fill_2
XANTENNA__34__A chany_top_in[19] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l2_in_3__A0 _22_/HI vgnd vpwr scs8hd_diode_2
XFILLER_34_125 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l3_in_0__A0 mux_right_ipin_2.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_37 vgnd vpwr scs8hd_decap_3
XFILLER_15_59 vpwr vgnd scs8hd_fill_2
XFILLER_56_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_8.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XPHY_120 vgnd vpwr scs8hd_decap_3
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_125 vgnd vpwr scs8hd_decap_12
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_ipin_8.mux_l2_in_0_ mux_right_ipin_8.mux_l1_in_1_/X mux_right_ipin_8.mux_l1_in_0_/X
+ mux_right_ipin_8.mux_l2_in_3_/S mux_right_ipin_8.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_6.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_8.mux_l4_in_0__S mux_right_ipin_8.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_3.scs8hd_dfxbp_1_3__D mux_right_ipin_3.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_13.mux_l1_in_2__S mux_right_ipin_13.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l1_in_0__A1 chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_15.mux_l2_in_2__A1 chany_top_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_15.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_8.mux_l1_in_1_ chany_top_in[3] chany_bottom_in[3] mux_right_ipin_8.mux_l1_in_2_/S
+ mux_right_ipin_8.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_37_13 vpwr vgnd scs8hd_fill_2
XFILLER_37_57 vpwr vgnd scs8hd_fill_2
XFILLER_53_78 vgnd vpwr scs8hd_decap_6
XANTENNA__42__A chany_top_in[11] vgnd vpwr scs8hd_diode_2
X_60_ chany_bottom_in[13] chany_top_out[13] vgnd vpwr scs8hd_buf_2
Xmux_right_ipin_12.mux_l3_in_0_ mux_right_ipin_12.mux_l2_in_1_/X mux_right_ipin_12.mux_l2_in_0_/X
+ mux_right_ipin_12.mux_l3_in_0_/S mux_right_ipin_12.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_ipin_13.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_64_3 vgnd vpwr scs8hd_decap_12
XFILLER_23_15 vgnd vpwr scs8hd_decap_6
XFILLER_48_23 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_12.mux_l2_in_2__S mux_right_ipin_12.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_64_44 vgnd vpwr scs8hd_decap_12
XANTENNA__37__A chany_top_in[16] vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_7.scs8hd_dfxbp_1_0_ prog_clk mux_right_ipin_6.mux_l4_in_0_/S mux_right_ipin_7.mux_l1_in_0_/S
+ mem_right_ipin_7.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_ipin_12.mux_l1_in_1__A0 chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_15.mux_l3_in_1__A1 mux_right_ipin_15.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_64_145 vgnd vpwr scs8hd_fill_1
X_43_ chany_top_in[10] chany_bottom_out[10] vgnd vpwr scs8hd_buf_2
XFILLER_29_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_9.mux_l2_in_2__A0 chany_bottom_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_55_101 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_12.mux_l2_in_1_ chany_bottom_in[13] mux_right_ipin_12.mux_l1_in_2_/X
+ mux_right_ipin_12.mux_l2_in_0_/S mux_right_ipin_12.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_34_69 vpwr vgnd scs8hd_fill_2
XFILLER_59_44 vgnd vpwr scs8hd_decap_4
XFILLER_59_11 vgnd vpwr scs8hd_decap_4
XFILLER_50_68 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l2_in_1__A1 chany_top_in[3] vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_3.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_3.mux_l1_in_0_/S
+ mux_right_ipin_3.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_91 vgnd vpwr scs8hd_fill_1
XFILLER_27_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_0.scs8hd_buf_4_0__A mux_left_ipin_0.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
X_26_ _26_/HI _26_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_62 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_12.mux_l2_in_0__A0 mux_right_ipin_12.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_15.mux_l4_in_0__A1 mux_right_ipin_15.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_45_79 vgnd vpwr scs8hd_decap_3
XFILLER_45_57 vpwr vgnd scs8hd_fill_2
XFILLER_45_35 vpwr vgnd scs8hd_fill_2
XFILLER_43_115 vgnd vpwr scs8hd_decap_6
Xmem_right_ipin_2.scs8hd_dfxbp_1_3_ prog_clk mux_right_ipin_2.mux_l3_in_0_/S mux_right_ipin_2.mux_l4_in_0_/S
+ mem_right_ipin_2.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_right_ipin_5.scs8hd_dfxbp_1_2__D mux_right_ipin_5.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_61_78 vpwr vgnd scs8hd_fill_2
XANTENNA__50__A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_10_71 vpwr vgnd scs8hd_fill_2
XFILLER_10_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_9.mux_l3_in_1__A0 mux_right_ipin_9.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l2_in_3__A1 chany_top_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_19_123 vpwr vgnd scs8hd_fill_2
XFILLER_19_145 vgnd vpwr scs8hd_fill_1
XFILLER_34_104 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_12.mux_l1_in_2_ chany_top_in[7] chany_bottom_in[7] mux_right_ipin_12.mux_l1_in_1_/S
+ mux_right_ipin_12.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_2.mux_l3_in_0__A1 mux_right_ipin_2.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_16 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_15.mux_l4_in_0__S ccff_tail vgnd vpwr scs8hd_diode_2
XFILLER_31_15 vgnd vpwr scs8hd_decap_12
XFILLER_56_78 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_10.mux_l2_in_2__A0 chany_bottom_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_16_137 vgnd vpwr scs8hd_decap_8
XPHY_121 vgnd vpwr scs8hd_decap_3
XPHY_110 vgnd vpwr scs8hd_decap_3
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__45__A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_92 vgnd vpwr scs8hd_decap_3
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_30_140 vgnd vpwr scs8hd_decap_6
XFILLER_26_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_36 vpwr vgnd scs8hd_fill_2
XFILLER_13_107 vpwr vgnd scs8hd_fill_2
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_9.mux_l4_in_0__A0 mux_right_ipin_9.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_70 vgnd vpwr scs8hd_decap_4
XFILLER_8_111 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_7.mux_l1_in_0__S mux_right_ipin_7.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_10.mux_l3_in_1__A0 mux_right_ipin_10.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_8.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_8.mux_l1_in_2_/S
+ mux_right_ipin_8.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_53_46 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_1.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_43_90 vpwr vgnd scs8hd_fill_2
XFILLER_4_51 vpwr vgnd scs8hd_fill_2
XFILLER_23_49 vpwr vgnd scs8hd_fill_2
XFILLER_48_46 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_5.scs8hd_buf_4_0__A mux_right_ipin_5.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_64_56 vgnd vpwr scs8hd_decap_6
XANTENNA__53__A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_7.scs8hd_dfxbp_1_1__D mux_right_ipin_7.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_12.mux_l1_in_1__A1 chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_49_143 vgnd vpwr scs8hd_decap_3
X_42_ chany_top_in[11] chany_bottom_out[11] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_ipin_10.mux_l4_in_0__A0 mux_right_ipin_10.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_9.mux_l2_in_2__A1 chany_top_in[10] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_6.mux_l2_in_0__S mux_right_ipin_6.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_15 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_12.mux_l2_in_0_ mux_right_ipin_12.mux_l1_in_1_/X mux_right_ipin_12.mux_l1_in_0_/X
+ mux_right_ipin_12.mux_l2_in_0_/S mux_right_ipin_12.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_50_36 vgnd vpwr scs8hd_decap_4
XFILLER_50_25 vgnd vpwr scs8hd_decap_6
XFILLER_46_102 vgnd vpwr scs8hd_decap_3
XANTENNA__48__A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_1_30 vpwr vgnd scs8hd_fill_2
X_25_ _25_/HI _25_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_74 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_12.mux_l2_in_0__A1 mux_right_ipin_12.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_right_ipin_2.scs8hd_dfxbp_1_2_ prog_clk mux_right_ipin_2.mux_l2_in_0_/S mux_right_ipin_2.mux_l3_in_0_/S
+ mem_right_ipin_2.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_28_102 vgnd vpwr scs8hd_decap_12
XFILLER_28_135 vgnd vpwr scs8hd_decap_8
XFILLER_61_57 vgnd vpwr scs8hd_decap_4
XFILLER_61_46 vgnd vpwr scs8hd_fill_1
XFILLER_61_24 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l2_in_2__S mux_right_ipin_1.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_9.mux_l3_in_1__A1 mux_right_ipin_9.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_81 vgnd vpwr scs8hd_decap_4
XFILLER_35_91 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_12.mux_l1_in_1_ chany_top_in[3] chany_bottom_in[3] mux_right_ipin_12.mux_l1_in_1_/S
+ mux_right_ipin_12.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_5.mux_l3_in_0__S mux_right_ipin_5.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_31_27 vgnd vpwr scs8hd_decap_12
XFILLER_56_57 vgnd vpwr scs8hd_decap_6
XFILLER_56_46 vpwr vgnd scs8hd_fill_2
XPHY_100 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_10.mux_l2_in_2__A1 chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_16_105 vgnd vpwr scs8hd_decap_12
XPHY_122 vgnd vpwr scs8hd_decap_3
XANTENNA__61__A chany_bottom_in[12] vgnd vpwr scs8hd_diode_2
XPHY_111 vgnd vpwr scs8hd_decap_3
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_119 vgnd vpwr scs8hd_decap_3
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_7 vgnd vpwr scs8hd_decap_3
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_22_108 vpwr vgnd scs8hd_fill_2
XFILLER_7_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_6.mux_l2_in_0__A0 chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_26_38 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_9.mux_l4_in_0__A1 mux_right_ipin_9.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_14.mux_l1_in_0__S mux_right_ipin_14.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA__56__A chany_bottom_in[17] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_9.scs8hd_dfxbp_1_0__D mux_right_ipin_8.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_93 vgnd vpwr scs8hd_decap_12
XFILLER_32_81 vgnd vpwr scs8hd_decap_4
XFILLER_59_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_6.mux_l2_in_3__S mux_right_ipin_6.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l4_in_0__S mux_right_ipin_4.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_10.mux_l3_in_1__A1 mux_right_ipin_10.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_26 vpwr vgnd scs8hd_fill_2
XFILLER_53_58 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_4.mux_l2_in_2__A0 chany_bottom_in[15] vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_12.scs8hd_dfxbp_1_3_ prog_clk mux_right_ipin_12.mux_l3_in_0_/S mux_right_ipin_12.mux_l4_in_0_/S
+ mem_right_ipin_12.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_4_85 vgnd vpwr scs8hd_decap_4
XFILLER_23_28 vpwr vgnd scs8hd_fill_2
XFILLER_3_9 vpwr vgnd scs8hd_fill_2
XFILLER_58_144 vpwr vgnd scs8hd_fill_2
XFILLER_48_36 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_13.mux_l2_in_0__S mux_right_ipin_13.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_10.mux_l4_in_0__A1 mux_right_ipin_10.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
X_41_ chany_top_in[12] chany_bottom_out[12] vgnd vpwr scs8hd_buf_2
XFILLER_64_125 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_4.mux_l3_in_1__A0 mux_right_ipin_4.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_55_114 vpwr vgnd scs8hd_fill_2
XANTENNA__64__A chany_bottom_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_46_136 vgnd vpwr scs8hd_decap_8
XFILLER_41_7 vpwr vgnd scs8hd_fill_2
XFILLER_40_81 vgnd vpwr scs8hd_decap_6
X_24_ _24_/HI _24_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_6.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_37_136 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_2.scs8hd_dfxbp_1_1_ prog_clk mux_right_ipin_2.mux_l1_in_0_/S mux_right_ipin_2.mux_l2_in_0_/S
+ mem_right_ipin_2.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_right_ipin_4.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_28_114 vpwr vgnd scs8hd_fill_2
XFILLER_61_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_11.scs8hd_dfxbp_1_1__D mux_right_ipin_11.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_12.mux_l3_in_0__S mux_right_ipin_12.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_ipin_9.scs8hd_dfxbp_1_3__D mux_right_ipin_9.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA__59__A chany_bottom_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_10_84 vpwr vgnd scs8hd_fill_2
XFILLER_19_71 vgnd vpwr scs8hd_decap_4
XFILLER_19_114 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_4.mux_l4_in_0__A0 mux_right_ipin_4.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_81 vgnd vpwr scs8hd_decap_4
XFILLER_51_80 vpwr vgnd scs8hd_fill_2
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_12.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_12.mux_l1_in_1_/S
+ mux_right_ipin_12.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_31_39 vgnd vpwr scs8hd_decap_12
XFILLER_56_36 vgnd vpwr scs8hd_decap_8
XPHY_123 vgnd vpwr scs8hd_decap_3
XPHY_112 vgnd vpwr scs8hd_decap_3
XPHY_101 vgnd vpwr scs8hd_decap_3
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_117 vgnd vpwr scs8hd_decap_6
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_right_ipin_13.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_7_74 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_11.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_6.mux_l2_in_0__A1 mux_right_ipin_6.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_13.mux_l2_in_3__S mux_right_ipin_13.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_11.mux_l4_in_0__S mux_right_ipin_11.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA__72__A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_32_93 vpwr vgnd scs8hd_fill_2
XFILLER_57_90 vgnd vpwr scs8hd_decap_4
XFILLER_5_127 vgnd vpwr scs8hd_decap_12
XFILLER_5_116 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_4.mux_l2_in_2__A1 chany_top_in[9] vgnd vpwr scs8hd_diode_2
XANTENNA__67__A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_27_71 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_12.scs8hd_dfxbp_1_2_ prog_clk mux_right_ipin_12.mux_l2_in_0_/S mux_right_ipin_12.mux_l3_in_0_/S
+ mem_right_ipin_12.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_4_64 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_14.mux_l2_in_1__A0 chany_bottom_in[11] vgnd vpwr scs8hd_diode_2
XFILLER_48_15 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_ipin_3.mux_l1_in_0__S mux_right_ipin_3.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_ipin_13.scs8hd_dfxbp_1_0__D mux_right_ipin_12.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_62 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_13.scs8hd_buf_4_0__A mux_right_ipin_13.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_49_123 vgnd vpwr scs8hd_decap_12
XFILLER_49_101 vpwr vgnd scs8hd_fill_2
X_40_ chany_top_in[13] chany_bottom_out[13] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_ipin_0.mux_l1_in_0__S mux_left_ipin_0.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_38_70 vgnd vpwr scs8hd_fill_1
XFILLER_64_137 vgnd vpwr scs8hd_decap_8
XFILLER_62_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_1.mux_l1_in_1__A0 chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l3_in_1__A1 mux_right_ipin_4.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_55_126 vpwr vgnd scs8hd_fill_2
XFILLER_18_18 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_9.scs8hd_buf_4_0_ mux_right_ipin_9.mux_l4_in_0_/X left_grid_pin_9_
+ vgnd vpwr scs8hd_buf_1
XFILLER_50_16 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_12.mux_l2_in_3__A0 _26_/HI vgnd vpwr scs8hd_diode_2
XFILLER_1_7 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_4.mux_l2_in_3_ _32_/HI chany_top_in[15] mux_right_ipin_4.mux_l2_in_3_/S
+ mux_right_ipin_4.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_14.mux_l3_in_0__A0 mux_right_ipin_14.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_7 vgnd vpwr scs8hd_decap_8
XFILLER_1_21 vgnd vpwr scs8hd_fill_1
X_23_ _23_/HI _23_/LO vgnd vpwr scs8hd_conb_1
XFILLER_37_115 vgnd vpwr scs8hd_fill_1
XFILLER_43_107 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l2_in_0__S mux_right_ipin_2.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_right_ipin_2.scs8hd_dfxbp_1_0_ prog_clk mux_right_ipin_1.mux_l4_in_0_/S mux_right_ipin_2.mux_l1_in_0_/S
+ mem_right_ipin_2.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_10_30 vgnd vpwr scs8hd_fill_1
XFILLER_10_63 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l2_in_0__A0 mux_right_ipin_1.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l4_in_0__A1 mux_right_ipin_4.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_118 vgnd vpwr scs8hd_decap_4
XFILLER_34_129 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_8.mux_l1_in_1__S mux_right_ipin_8.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_124 vgnd vpwr scs8hd_decap_3
XPHY_113 vgnd vpwr scs8hd_decap_3
XPHY_102 vgnd vpwr scs8hd_decap_3
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_ipin_0.mux_l1_in_1__A0 chany_top_in[2] vgnd vpwr scs8hd_diode_2
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_62 vgnd vpwr scs8hd_decap_4
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_62_91 vgnd vpwr scs8hd_fill_1
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_30_110 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_15.scs8hd_buf_4_0_ mux_right_ipin_15.mux_l4_in_0_/X left_grid_pin_15_
+ vgnd vpwr scs8hd_buf_1
XFILLER_7_53 vpwr vgnd scs8hd_fill_2
XFILLER_21_110 vpwr vgnd scs8hd_fill_2
XFILLER_26_29 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_4.mux_l4_in_0_ mux_right_ipin_4.mux_l3_in_1_/X mux_right_ipin_4.mux_l3_in_0_/X
+ mux_right_ipin_4.mux_l4_in_0_/S mux_right_ipin_4.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_1.mux_l3_in_0__S mux_right_ipin_1.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_ipin_13.scs8hd_dfxbp_1_3__D mux_right_ipin_13.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_9.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_32_72 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_0.mux_l2_in_0__A0 mux_left_ipin_0.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_7.mux_l2_in_1__S mux_right_ipin_7.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_53_16 vpwr vgnd scs8hd_fill_2
XFILLER_5_139 vgnd vpwr scs8hd_decap_6
Xmux_right_ipin_9.mux_l2_in_3_ _20_/HI chany_top_in[14] mux_right_ipin_9.mux_l2_in_1_/S
+ mux_right_ipin_9.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_27_83 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_10.mux_l1_in_0__S mux_right_ipin_10.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_43_71 vgnd vpwr scs8hd_decap_8
XFILLER_57_6 vpwr vgnd scs8hd_fill_2
XFILLER_4_32 vgnd vpwr scs8hd_decap_4
XFILLER_4_10 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_12.scs8hd_dfxbp_1_1_ prog_clk mux_right_ipin_12.mux_l1_in_1_/S mux_right_ipin_12.mux_l2_in_0_/S
+ mem_right_ipin_12.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_right_ipin_4.mux_l3_in_1_ mux_right_ipin_4.mux_l2_in_3_/X mux_right_ipin_4.mux_l2_in_2_/X
+ mux_right_ipin_4.mux_l3_in_1_/S mux_right_ipin_4.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_14.mux_l2_in_1__A1 chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_58_113 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l2_in_3__S mux_right_ipin_2.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_64_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_0.mux_l4_in_0__S mux_right_ipin_0.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_8.mux_l1_in_2__A0 chany_top_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_49_135 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_2__D mux_right_ipin_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_38_82 vgnd vpwr scs8hd_decap_4
XFILLER_55_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l1_in_1__A1 chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_6.mux_l3_in_1__S mux_right_ipin_6.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_59_48 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_12.mux_l2_in_3__A1 chany_top_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_24_62 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_4.mux_l2_in_2_ chany_bottom_in[15] chany_top_in[9] mux_right_ipin_4.mux_l2_in_3_/S
+ mux_right_ipin_4.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_40_61 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_14.mux_l3_in_0__A1 mux_right_ipin_14.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_49_70 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_11.mux_l1_in_0__A0 chany_top_in[0] vgnd vpwr scs8hd_diode_2
X_22_ _22_/HI _22_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_ipin_8.mux_l2_in_1__A0 chany_bottom_in[13] vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_9.mux_l4_in_0_ mux_right_ipin_9.mux_l3_in_1_/X mux_right_ipin_9.mux_l3_in_0_/X
+ mux_right_ipin_9.mux_l4_in_0_/S mux_right_ipin_9.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_0.scs8hd_buf_4_0__A mux_right_ipin_0.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_45_39 vpwr vgnd scs8hd_fill_2
XFILLER_10_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_15.scs8hd_dfxbp_1_2__D mux_right_ipin_15.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_1.mux_l2_in_0__A1 mux_right_ipin_1.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_127 vgnd vpwr scs8hd_decap_12
XFILLER_51_71 vgnd vpwr scs8hd_decap_3
XFILLER_18_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_6.mux_l2_in_3__A0 _17_/HI vgnd vpwr scs8hd_diode_2
XPHY_125 vgnd vpwr scs8hd_decap_3
XPHY_114 vgnd vpwr scs8hd_decap_3
XPHY_103 vgnd vpwr scs8hd_decap_3
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_ipin_0.mux_l1_in_1__A1 chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_130 vgnd vpwr scs8hd_decap_12
XPHY_5 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_8.mux_l3_in_0__A0 mux_right_ipin_8.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_9.mux_l3_in_1_ mux_right_ipin_9.mux_l2_in_3_/X mux_right_ipin_9.mux_l2_in_2_/X
+ mux_right_ipin_9.mux_l3_in_0_/S mux_right_ipin_9.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_7_87 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_14.mux_l2_in_1__S mux_right_ipin_14.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_30 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_ipin_2.scs8hd_dfxbp_1_1__D mux_right_ipin_2.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_left_ipin_0.scs8hd_buf_4_0_ mux_left_ipin_0.mux_l4_in_0_/X right_grid_pin_52_
+ vgnd vpwr scs8hd_buf_1
XANTENNA_mux_left_ipin_0.mux_l2_in_0__A1 mux_left_ipin_0.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_9.mux_l2_in_2_ chany_bottom_in[14] chany_top_in[10] mux_right_ipin_9.mux_l2_in_1_/S
+ mux_right_ipin_9.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_43_50 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_4.scs8hd_buf_4_0_ mux_right_ipin_4.mux_l4_in_0_/X left_grid_pin_4_
+ vgnd vpwr scs8hd_buf_1
XFILLER_27_51 vpwr vgnd scs8hd_fill_2
XFILLER_43_94 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_12.scs8hd_dfxbp_1_0_ prog_clk mux_right_ipin_11.mux_l4_in_0_/S mux_right_ipin_12.mux_l1_in_1_/S
+ mem_right_ipin_12.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_4_99 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_4.mux_l3_in_0_ mux_right_ipin_4.mux_l2_in_1_/X mux_right_ipin_4.mux_l2_in_0_/X
+ mux_right_ipin_4.mux_l3_in_1_/S mux_right_ipin_4.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_58_136 vgnd vpwr scs8hd_decap_8
XFILLER_64_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_8.mux_l1_in_2__A1 chany_bottom_in[9] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_13.mux_l3_in_1__S mux_right_ipin_13.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_53 vpwr vgnd scs8hd_fill_2
XFILLER_49_114 vpwr vgnd scs8hd_fill_2
XFILLER_1_132 vpwr vgnd scs8hd_fill_2
XFILLER_64_106 vgnd vpwr scs8hd_decap_12
XFILLER_54_93 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_2.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_48_3 vgnd vpwr scs8hd_decap_12
XFILLER_34_19 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_24_41 vpwr vgnd scs8hd_fill_2
XFILLER_24_85 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_ipin_11.mux_l1_in_0__A1 chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_4.mux_l2_in_1_ chany_bottom_in[9] mux_right_ipin_4.mux_l1_in_2_/X
+ mux_right_ipin_4.mux_l2_in_3_/S mux_right_ipin_4.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_96 vgnd vpwr scs8hd_decap_6
XFILLER_49_60 vgnd vpwr scs8hd_fill_1
X_21_ _21_/HI _21_/LO vgnd vpwr scs8hd_conb_1
XFILLER_60_120 vgnd vpwr scs8hd_decap_3
XFILLER_1_78 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_8.mux_l2_in_1__A1 mux_right_ipin_8.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_61_28 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_10.scs8hd_buf_4_0_ mux_right_ipin_10.mux_l4_in_0_/X left_grid_pin_10_
+ vgnd vpwr scs8hd_buf_1
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
XFILLER_19_106 vpwr vgnd scs8hd_fill_2
XFILLER_19_117 vpwr vgnd scs8hd_fill_2
XFILLER_19_139 vgnd vpwr scs8hd_decap_6
XFILLER_35_40 vpwr vgnd scs8hd_fill_2
XFILLER_35_95 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_4.scs8hd_dfxbp_1_0__D mux_right_ipin_3.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_25_109 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_13.mux_l2_in_3_ _27_/HI chany_top_in[18] mux_right_ipin_13.mux_l2_in_3_/S
+ mux_right_ipin_13.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_ipin_4.mux_l1_in_2_ chany_top_in[5] chany_bottom_in[5] mux_right_ipin_4.mux_l1_in_2_/S
+ mux_right_ipin_4.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_6.mux_l2_in_3__A1 chany_top_in[19] vgnd vpwr scs8hd_diode_2
XPHY_126 vgnd vpwr scs8hd_decap_3
XPHY_115 vgnd vpwr scs8hd_decap_3
XPHY_104 vgnd vpwr scs8hd_decap_3
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_142 vgnd vpwr scs8hd_decap_4
XFILLER_21_53 vpwr vgnd scs8hd_fill_2
XFILLER_21_97 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_5.scs8hd_dfxbp_1_3_ prog_clk mux_right_ipin_5.mux_l3_in_0_/S mux_right_ipin_5.mux_l4_in_0_/S
+ mem_right_ipin_5.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_ipin_5.mux_l1_in_0__A0 chany_top_in[0] vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_8.mux_l3_in_0__A1 mux_right_ipin_8.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_9.mux_l3_in_0_ mux_right_ipin_9.mux_l2_in_1_/X mux_right_ipin_9.mux_l2_in_0_/X
+ mux_right_ipin_9.mux_l3_in_0_/S mux_right_ipin_9.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_7_33 vgnd vpwr scs8hd_fill_1
XFILLER_30_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_4.mux_l1_in_1__S mux_right_ipin_4.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_53 vpwr vgnd scs8hd_fill_2
XFILLER_8_138 vgnd vpwr scs8hd_decap_8
XFILLER_12_134 vpwr vgnd scs8hd_fill_2
XFILLER_32_85 vgnd vpwr scs8hd_fill_1
XFILLER_53_29 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_9.mux_l2_in_1_ chany_bottom_in[10] mux_right_ipin_9.mux_l1_in_2_/X
+ mux_right_ipin_9.mux_l2_in_1_/S mux_right_ipin_9.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_ipin_13.mux_l4_in_0_ mux_right_ipin_13.mux_l3_in_1_/X mux_right_ipin_13.mux_l3_in_0_/X
+ mux_right_ipin_13.mux_l4_in_0_/S mux_right_ipin_13.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_89 vgnd vpwr scs8hd_fill_1
XFILLER_4_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_3.mux_l2_in_1__S mux_right_ipin_3.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_3.mux_l2_in_1__A0 chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_13_32 vpwr vgnd scs8hd_fill_2
XFILLER_13_76 vpwr vgnd scs8hd_fill_2
XFILLER_1_144 vpwr vgnd scs8hd_fill_2
XFILLER_64_118 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_ipin_0.mux_l2_in_1__S mux_left_ipin_0.mux_l2_in_2_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_4.scs8hd_dfxbp_1_3__D mux_right_ipin_4.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_9.mux_l1_in_2__S mux_right_ipin_9.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_55_118 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_9.mux_l1_in_2_ chany_top_in[4] chany_bottom_in[4] mux_right_ipin_9.mux_l1_in_2_/S
+ mux_right_ipin_9.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_59_17 vgnd vpwr scs8hd_decap_6
XFILLER_46_107 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_13.mux_l3_in_1_ mux_right_ipin_13.mux_l2_in_3_/X mux_right_ipin_13.mux_l2_in_2_/X
+ mux_right_ipin_13.mux_l3_in_1_/S mux_right_ipin_13.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_75 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_4.mux_l2_in_0_ mux_right_ipin_4.mux_l1_in_1_/X mux_right_ipin_4.mux_l1_in_0_/X
+ mux_right_ipin_4.mux_l2_in_3_/S mux_right_ipin_4.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_40_41 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_1.mux_l2_in_3__A0 _23_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_8.scs8hd_buf_4_0__A mux_right_ipin_8.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
X_20_ _20_/HI _20_/LO vgnd vpwr scs8hd_conb_1
XFILLER_37_107 vpwr vgnd scs8hd_fill_2
XFILLER_37_118 vpwr vgnd scs8hd_fill_2
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_3.mux_l3_in_0__A0 mux_right_ipin_3.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_61_18 vpwr vgnd scs8hd_fill_2
XFILLER_51_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_2.mux_l3_in_1__S mux_right_ipin_2.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_11 vgnd vpwr scs8hd_decap_3
XFILLER_10_88 vpwr vgnd scs8hd_fill_2
XFILLER_19_31 vpwr vgnd scs8hd_fill_2
XFILLER_19_53 vpwr vgnd scs8hd_fill_2
XFILLER_51_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_7.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_25_6 vpwr vgnd scs8hd_fill_2
XFILLER_33_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_8.mux_l2_in_2__S mux_right_ipin_8.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_56_18 vgnd vpwr scs8hd_decap_12
XPHY_116 vgnd vpwr scs8hd_decap_3
XPHY_105 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_13.mux_l2_in_2_ chany_bottom_in[18] chany_top_in[14] mux_right_ipin_13.mux_l2_in_3_/S
+ mux_right_ipin_13.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_ipin_4.mux_l1_in_1_ chany_top_in[3] chany_bottom_in[3] mux_right_ipin_4.mux_l1_in_2_/S
+ mux_right_ipin_4.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_ipin_5.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XPHY_127 vgnd vpwr scs8hd_decap_3
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_right_ipin_5.scs8hd_dfxbp_1_2_ prog_clk mux_right_ipin_5.mux_l2_in_0_/S mux_right_ipin_5.mux_l3_in_0_/S
+ mem_right_ipin_5.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_21_43 vpwr vgnd scs8hd_fill_2
XFILLER_46_51 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_5.mux_l1_in_0__A1 chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_132 vgnd vpwr scs8hd_decap_12
XFILLER_30_102 vpwr vgnd scs8hd_fill_2
XFILLER_23_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_0.mux_l2_in_3__A0 _21_/HI vgnd vpwr scs8hd_diode_2
XFILLER_16_32 vgnd vpwr scs8hd_decap_8
XFILLER_32_64 vgnd vpwr scs8hd_decap_8
XFILLER_32_75 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_14.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_6.scs8hd_dfxbp_1_2__D mux_right_ipin_6.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_12.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_9.mux_l2_in_0_ mux_right_ipin_9.mux_l1_in_1_/X mux_right_ipin_9.mux_l1_in_0_/X
+ mux_right_ipin_9.mux_l2_in_1_/S mux_right_ipin_9.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_27_75 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_13.mux_l1_in_1__A0 chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_43_30 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_10.mux_l2_in_1__S mux_right_ipin_10.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_131 vgnd vpwr scs8hd_decap_12
XFILLER_4_68 vpwr vgnd scs8hd_fill_2
XFILLER_13_11 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_3.mux_l2_in_1__A1 chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_1_101 vpwr vgnd scs8hd_fill_2
XFILLER_38_41 vgnd vpwr scs8hd_decap_6
XFILLER_38_63 vgnd vpwr scs8hd_fill_1
XFILLER_54_51 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_9.mux_l1_in_1_ chany_top_in[2] chany_bottom_in[2] mux_right_ipin_9.mux_l1_in_2_/S
+ mux_right_ipin_9.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmem_right_ipin_15.scs8hd_dfxbp_1_3_ prog_clk mux_right_ipin_15.mux_l3_in_0_/S ccff_tail
+ mem_right_ipin_15.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_ipin_13.mux_l2_in_0__A0 mux_right_ipin_13.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_13.mux_l3_in_0_ mux_right_ipin_13.mux_l2_in_1_/X mux_right_ipin_13.mux_l2_in_0_/X
+ mux_right_ipin_13.mux_l3_in_1_/S mux_right_ipin_13.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_40_53 vgnd vpwr scs8hd_decap_8
XFILLER_40_64 vpwr vgnd scs8hd_fill_2
XFILLER_49_62 vgnd vpwr scs8hd_decap_6
XFILLER_1_14 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_1.mux_l2_in_3__A1 chany_top_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_53_3 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_0.mux_l1_in_0__A0 chany_top_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_3.mux_l3_in_0__A1 mux_right_ipin_3.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_130 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_15.mux_l2_in_2__S mux_right_ipin_15.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_67 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_11.mux_l2_in_2__A0 chany_bottom_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_19_43 vgnd vpwr scs8hd_fill_1
XFILLER_42_144 vpwr vgnd scs8hd_fill_2
XFILLER_42_100 vgnd vpwr scs8hd_decap_12
XFILLER_35_53 vpwr vgnd scs8hd_fill_2
XFILLER_33_111 vpwr vgnd scs8hd_fill_2
XFILLER_33_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_8.scs8hd_dfxbp_1_1__D mux_right_ipin_8.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_right_ipin_13.mux_l2_in_1_ chany_bottom_in[14] mux_right_ipin_13.mux_l1_in_2_/X
+ mux_right_ipin_13.mux_l2_in_3_/S mux_right_ipin_13.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_ipin_4.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_4.mux_l1_in_2_/S
+ mux_right_ipin_4.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XPHY_128 vgnd vpwr scs8hd_decap_3
XPHY_117 vgnd vpwr scs8hd_decap_3
XPHY_106 vgnd vpwr scs8hd_decap_3
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_66 vgnd vpwr scs8hd_fill_1
Xmem_right_ipin_5.scs8hd_dfxbp_1_1_ prog_clk mux_right_ipin_5.mux_l1_in_0_/S mux_right_ipin_5.mux_l2_in_0_/S
+ mem_right_ipin_5.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_46_85 vgnd vpwr scs8hd_fill_1
XFILLER_62_51 vgnd vpwr scs8hd_decap_12
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_144 vpwr vgnd scs8hd_fill_2
XFILLER_7_57 vpwr vgnd scs8hd_fill_2
XFILLER_16_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_11.mux_l3_in_1__A0 mux_right_ipin_11.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_3__A1 chany_top_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_21_114 vpwr vgnd scs8hd_fill_2
XFILLER_16_66 vpwr vgnd scs8hd_fill_2
XFILLER_16_77 vgnd vpwr scs8hd_decap_12
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XFILLER_57_62 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_13.mux_l1_in_2_ chany_top_in[8] chany_bottom_in[8] mux_right_ipin_13.mux_l1_in_1_/S
+ mux_right_ipin_13.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_1__S mux_right_ipin_0.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_13.mux_l1_in_1__A1 chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_43_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_11.mux_l4_in_0__A0 mux_right_ipin_11.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_143 vgnd vpwr scs8hd_decap_3
XFILLER_4_110 vpwr vgnd scs8hd_fill_2
XFILLER_4_47 vpwr vgnd scs8hd_fill_2
XFILLER_13_45 vpwr vgnd scs8hd_fill_2
XFILLER_1_113 vgnd vpwr scs8hd_decap_3
XFILLER_38_86 vgnd vpwr scs8hd_fill_1
XFILLER_54_85 vpwr vgnd scs8hd_fill_2
XFILLER_54_63 vpwr vgnd scs8hd_fill_2
XFILLER_54_30 vgnd vpwr scs8hd_fill_1
XFILLER_55_7 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_10.scs8hd_dfxbp_1_2__D mux_right_ipin_10.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_right_ipin_9.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_9.mux_l1_in_2_/S
+ mux_right_ipin_9.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_13.mux_l2_in_0__A1 mux_right_ipin_13.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_right_ipin_15.scs8hd_dfxbp_1_2_ prog_clk mux_right_ipin_15.mux_l2_in_0_/S mux_right_ipin_15.mux_l3_in_0_/S
+ mem_right_ipin_15.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_49_52 vpwr vgnd scs8hd_fill_2
XFILLER_49_74 vpwr vgnd scs8hd_fill_2
XFILLER_1_26 vpwr vgnd scs8hd_fill_2
XFILLER_60_145 vgnd vpwr scs8hd_fill_1
XFILLER_60_112 vgnd vpwr scs8hd_decap_8
XFILLER_46_3 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_0.mux_l1_in_0__A1 chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_51_123 vgnd vpwr scs8hd_decap_12
XFILLER_51_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_5.mux_l1_in_2__S mux_right_ipin_5.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_142 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_11.mux_l2_in_2__A1 chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_19_77 vpwr vgnd scs8hd_fill_2
XFILLER_42_112 vgnd vpwr scs8hd_decap_12
XFILLER_35_87 vpwr vgnd scs8hd_fill_2
XFILLER_51_53 vpwr vgnd scs8hd_fill_2
XFILLER_18_7 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_9.mux_l2_in_0__S mux_right_ipin_9.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_13.mux_l2_in_0_ mux_right_ipin_13.mux_l1_in_1_/X mux_right_ipin_13.mux_l1_in_0_/X
+ mux_right_ipin_13.mux_l2_in_3_/S mux_right_ipin_13.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_7.mux_l2_in_0__A0 chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XPHY_129 vgnd vpwr scs8hd_decap_3
XPHY_118 vgnd vpwr scs8hd_decap_3
XPHY_107 vgnd vpwr scs8hd_decap_3
Xmem_right_ipin_5.scs8hd_dfxbp_1_0_ prog_clk mux_right_ipin_4.mux_l4_in_0_/S mux_right_ipin_5.mux_l1_in_0_/S
+ mem_right_ipin_5.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_46_64 vgnd vpwr scs8hd_decap_6
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_62_63 vgnd vpwr scs8hd_decap_12
XFILLER_7_36 vpwr vgnd scs8hd_fill_2
XFILLER_7_25 vgnd vpwr scs8hd_decap_8
XFILLER_21_126 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_11.mux_l3_in_1__A1 mux_right_ipin_11.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l2_in_2__S mux_right_ipin_4.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_23 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_5.mux_l2_in_2__A0 chany_bottom_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_16_89 vgnd vpwr scs8hd_decap_3
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XFILLER_32_88 vgnd vpwr scs8hd_decap_4
XFILLER_57_96 vpwr vgnd scs8hd_fill_2
XFILLER_57_30 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_13.mux_l1_in_1_ chany_top_in[2] chany_bottom_in[2] mux_right_ipin_13.mux_l1_in_1_/S
+ mux_right_ipin_13.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_ipin_12.scs8hd_dfxbp_1_1__D mux_right_ipin_12.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_8.mux_l3_in_0__S mux_right_ipin_8.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_right_ipin_0.scs8hd_dfxbp_1_3_ prog_clk mux_right_ipin_0.mux_l3_in_1_/S mux_right_ipin_0.mux_l4_in_0_/S
+ mem_right_ipin_0.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_43_10 vgnd vpwr scs8hd_decap_12
XFILLER_27_55 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_11.mux_l4_in_0__A1 mux_right_ipin_11.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_5.mux_l3_in_1__A0 mux_right_ipin_5.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XFILLER_8_6 vpwr vgnd scs8hd_fill_2
XFILLER_1_136 vgnd vpwr scs8hd_decap_8
XFILLER_57_140 vpwr vgnd scs8hd_fill_2
XFILLER_49_118 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_9.mux_l2_in_3__S mux_right_ipin_9.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_63_143 vgnd vpwr scs8hd_decap_3
XFILLER_63_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_7.mux_l4_in_0__S mux_right_ipin_7.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_right_ipin_15.scs8hd_dfxbp_1_1_ prog_clk mux_right_ipin_15.mux_l1_in_0_/S mux_right_ipin_15.mux_l2_in_0_/S
+ mem_right_ipin_15.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_54_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_ipin_5.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_24_23 vgnd vpwr scs8hd_decap_3
XFILLER_24_45 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_12.mux_l1_in_2__S mux_right_ipin_12.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_40_11 vpwr vgnd scs8hd_fill_2
XFILLER_40_77 vpwr vgnd scs8hd_fill_2
XFILLER_49_97 vpwr vgnd scs8hd_fill_2
XFILLER_45_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_5.mux_l4_in_0__A0 mux_right_ipin_5.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_ipin_3.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_39_3 vgnd vpwr scs8hd_decap_12
XFILLER_51_135 vgnd vpwr scs8hd_decap_8
XFILLER_27_143 vgnd vpwr scs8hd_decap_3
XFILLER_42_124 vgnd vpwr scs8hd_decap_12
XFILLER_51_76 vpwr vgnd scs8hd_fill_2
XFILLER_18_121 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_14.scs8hd_dfxbp_1_0__D mux_right_ipin_13.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_12.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.mux_l2_in_0__A1 mux_right_ipin_7.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_119 vgnd vpwr scs8hd_decap_3
XPHY_108 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_3.scs8hd_buf_4_0__A mux_right_ipin_3.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_11.mux_l2_in_2__S mux_right_ipin_11.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_ipin_10.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_62_97 vgnd vpwr scs8hd_decap_12
XFILLER_62_75 vgnd vpwr scs8hd_decap_12
XFILLER_30_116 vgnd vpwr scs8hd_decap_12
XFILLER_21_138 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_15.mux_l3_in_0__S mux_right_ipin_15.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_5.mux_l2_in_2__A1 chany_top_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_12_138 vgnd vpwr scs8hd_decap_8
XFILLER_32_56 vgnd vpwr scs8hd_decap_6
XFILLER_57_53 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_13.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_13.mux_l1_in_1_/S
+ mux_right_ipin_13.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_21_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_15.mux_l2_in_1__A0 chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_8_80 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_0.scs8hd_dfxbp_1_2_ prog_clk mux_right_ipin_0.mux_l2_in_0_/S mux_right_ipin_0.mux_l3_in_1_/S
+ mem_right_ipin_0.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_27_23 vpwr vgnd scs8hd_fill_2
XFILLER_43_33 vpwr vgnd scs8hd_fill_2
XFILLER_43_22 vgnd vpwr scs8hd_decap_8
XFILLER_4_27 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_0.mux_l2_in_3_ _22_/HI chany_top_in[17] mux_right_ipin_0.mux_l2_in_0_/S
+ mux_right_ipin_0.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_5.mux_l3_in_1__A1 mux_right_ipin_5.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_13.mux_l2_in_3__A0 _27_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_14.mux_l4_in_0__S mux_right_ipin_14.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_66 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_15.mux_l3_in_0__A0 mux_right_ipin_15.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_ipin_14.scs8hd_dfxbp_1_3__D mux_right_ipin_14.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_right_ipin_15.scs8hd_dfxbp_1_0_ prog_clk mux_right_ipin_14.mux_l4_in_0_/S mux_right_ipin_15.mux_l1_in_0_/S
+ mem_right_ipin_15.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_5_70 vgnd vpwr scs8hd_decap_4
XFILLER_54_144 vpwr vgnd scs8hd_fill_2
XFILLER_54_111 vpwr vgnd scs8hd_fill_2
XFILLER_24_57 vgnd vpwr scs8hd_decap_3
XFILLER_40_89 vgnd vpwr scs8hd_decap_3
XFILLER_49_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l2_in_0__A0 chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_60_125 vgnd vpwr scs8hd_decap_12
XFILLER_45_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_5.mux_l4_in_0__A1 mux_right_ipin_5.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_60_7 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_6.mux_l1_in_0__S mux_right_ipin_6.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_26 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_0.mux_l4_in_0_ mux_right_ipin_0.mux_l3_in_1_/X mux_right_ipin_0.mux_l3_in_0_/X
+ mux_right_ipin_0.mux_l4_in_0_/S mux_right_ipin_0.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_19_35 vpwr vgnd scs8hd_fill_2
XFILLER_42_136 vgnd vpwr scs8hd_decap_8
XFILLER_19_57 vpwr vgnd scs8hd_fill_2
XFILLER_27_111 vgnd vpwr scs8hd_decap_4
XFILLER_35_12 vpwr vgnd scs8hd_fill_2
XFILLER_51_88 vpwr vgnd scs8hd_fill_2
XFILLER_18_100 vpwr vgnd scs8hd_fill_2
XFILLER_18_133 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_0.mux_l2_in_2__A0 chany_bottom_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_33_136 vgnd vpwr scs8hd_decap_8
Xmem_right_ipin_10.scs8hd_dfxbp_1_3_ prog_clk mux_right_ipin_10.mux_l3_in_1_/S mux_right_ipin_10.mux_l4_in_0_/S
+ mem_right_ipin_10.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_51_3 vgnd vpwr scs8hd_decap_6
X_59_ chany_bottom_in[14] chany_top_out[14] vgnd vpwr scs8hd_buf_2
XFILLER_2_71 vpwr vgnd scs8hd_fill_2
XFILLER_24_114 vgnd vpwr scs8hd_fill_1
XPHY_109 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_1.scs8hd_dfxbp_1_2__D mux_right_ipin_1.mux_l2_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_47 vgnd vpwr scs8hd_decap_4
XFILLER_21_69 vpwr vgnd scs8hd_fill_2
XFILLER_46_11 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_1.mux_l1_in_2__S mux_right_ipin_1.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_5.mux_l2_in_3_ _33_/HI chany_top_in[16] mux_right_ipin_5.mux_l2_in_0_/S
+ mux_right_ipin_5.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_62_32 vgnd vpwr scs8hd_decap_12
XFILLER_46_88 vpwr vgnd scs8hd_fill_2
XFILLER_30_106 vpwr vgnd scs8hd_fill_2
XFILLER_30_128 vgnd vpwr scs8hd_decap_12
XFILLER_62_87 vgnd vpwr scs8hd_decap_4
XFILLER_7_49 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_8.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l3_in_1_ mux_right_ipin_0.mux_l2_in_3_/X mux_right_ipin_0.mux_l2_in_2_/X
+ mux_right_ipin_0.mux_l3_in_1_/S mux_right_ipin_0.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_5.mux_l2_in_0__S mux_right_ipin_5.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l3_in_1__A0 mux_right_ipin_0.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_57_10 vpwr vgnd scs8hd_fill_2
XFILLER_57_21 vgnd vpwr scs8hd_decap_6
XFILLER_7_121 vgnd vpwr scs8hd_fill_1
Xmem_right_ipin_8.scs8hd_dfxbp_1_3_ prog_clk mux_right_ipin_8.mux_l3_in_1_/S mux_right_ipin_8.mux_l4_in_0_/S
+ mem_right_ipin_8.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_14_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_15.mux_l2_in_1__A1 chany_top_in[2] vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_0.scs8hd_dfxbp_1_1_ prog_clk mux_right_ipin_0.mux_l1_in_2_/S mux_right_ipin_0.mux_l2_in_0_/S
+ mem_right_ipin_0.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_0__D ccff_head vgnd vpwr scs8hd_diode_2
XFILLER_27_46 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_9.mux_l1_in_2__A0 chany_top_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l2_in_2__S mux_right_ipin_0.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_ipin_15.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l2_in_2_ chany_bottom_in[17] chany_top_in[11] mux_right_ipin_0.mux_l2_in_0_/S
+ mux_right_ipin_0.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_58_109 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.mux_l4_in_0__A0 mux_right_ipin_0.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_5.mux_l4_in_0_ mux_right_ipin_5.mux_l3_in_1_/X mux_right_ipin_5.mux_l3_in_0_/X
+ mux_right_ipin_5.mux_l4_in_0_/S mux_right_ipin_5.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_13_15 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_4.mux_l3_in_0__S mux_right_ipin_4.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_13.mux_l2_in_3__A1 chany_top_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_1_105 vpwr vgnd scs8hd_fill_2
XFILLER_54_55 vpwr vgnd scs8hd_fill_2
XFILLER_54_22 vgnd vpwr scs8hd_decap_8
XFILLER_38_89 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_12.mux_l1_in_0__A0 chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_54_77 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_15.mux_l3_in_0__A1 mux_right_ipin_15.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_63_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_9.mux_l2_in_1__A0 chany_bottom_in[10] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_3.scs8hd_dfxbp_1_1__D mux_right_ipin_3.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_13.mux_l1_in_0__S mux_right_ipin_13.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_45_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l2_in_0__A1 mux_right_ipin_2.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_18 vgnd vpwr scs8hd_fill_1
XFILLER_60_137 vgnd vpwr scs8hd_decap_8
XFILLER_14_80 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_5.mux_l3_in_1_ mux_right_ipin_5.mux_l2_in_3_/X mux_right_ipin_5.mux_l2_in_2_/X
+ mux_right_ipin_5.mux_l3_in_0_/S mux_right_ipin_5.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_30_90 vpwr vgnd scs8hd_fill_2
XFILLER_51_115 vpwr vgnd scs8hd_fill_2
XFILLER_10_16 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_5.mux_l2_in_3__S mux_right_ipin_5.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_3.mux_l4_in_0__S mux_right_ipin_3.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_7.mux_l2_in_3__A0 _18_/HI vgnd vpwr scs8hd_diode_2
XFILLER_27_123 vgnd vpwr scs8hd_decap_12
XFILLER_35_57 vpwr vgnd scs8hd_fill_2
XFILLER_51_34 vpwr vgnd scs8hd_fill_2
XFILLER_51_12 vpwr vgnd scs8hd_fill_2
XANTENNA__40__A chany_top_in[13] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l4_in_0__S mux_left_ipin_0.mux_l4_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_18_145 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_9.mux_l3_in_0__A0 mux_right_ipin_9.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_90 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_0.mux_l2_in_2__A1 chany_top_in[11] vgnd vpwr scs8hd_diode_2
XFILLER_33_115 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_9.mux_l3_in_1__S mux_right_ipin_9.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_right_ipin_10.scs8hd_dfxbp_1_2_ prog_clk mux_right_ipin_10.mux_l2_in_2_/S mux_right_ipin_10.mux_l3_in_1_/S
+ mem_right_ipin_10.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_44_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_50 vpwr vgnd scs8hd_fill_2
X_58_ chany_bottom_in[15] chany_top_out[15] vgnd vpwr scs8hd_buf_2
XFILLER_24_104 vpwr vgnd scs8hd_fill_2
XFILLER_24_126 vpwr vgnd scs8hd_fill_2
XFILLER_21_15 vgnd vpwr scs8hd_decap_3
XFILLER_46_23 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_3__D mux_left_ipin_0.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_5.mux_l2_in_2_ chany_bottom_in[16] chany_top_in[10] mux_right_ipin_5.mux_l2_in_0_/S
+ mux_right_ipin_5.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_62_44 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_12.mux_l2_in_0__S mux_right_ipin_12.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA__35__A chany_top_in[18] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_10.mux_l2_in_1__A0 chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_11.scs8hd_buf_4_0__A mux_right_ipin_11.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l3_in_0_ mux_right_ipin_0.mux_l2_in_1_/X mux_right_ipin_0.mux_l2_in_0_/X
+ mux_right_ipin_0.mux_l3_in_1_/S mux_right_ipin_0.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
XFILLER_12_107 vgnd vpwr scs8hd_decap_8
XFILLER_16_15 vgnd vpwr scs8hd_decap_8
XFILLER_16_26 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_0.mux_l3_in_1__A1 mux_right_ipin_0.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_57_66 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_5.scs8hd_buf_4_0_ mux_right_ipin_5.mux_l4_in_0_/X left_grid_pin_5_
+ vgnd vpwr scs8hd_buf_1
Xmem_right_ipin_8.scs8hd_dfxbp_1_2_ prog_clk mux_right_ipin_8.mux_l2_in_3_/S mux_right_ipin_8.mux_l3_in_1_/S
+ mem_right_ipin_8.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_8_93 vgnd vpwr scs8hd_decap_4
Xmem_right_ipin_0.scs8hd_dfxbp_1_0_ prog_clk mux_left_ipin_0.mux_l4_in_0_/S mux_right_ipin_0.mux_l1_in_2_/S
+ mem_right_ipin_0.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_ipin_10.mux_l3_in_0__A0 mux_right_ipin_10.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_9.mux_l1_in_2__A1 chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_43_57 vpwr vgnd scs8hd_fill_2
XFILLER_43_46 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_5.scs8hd_dfxbp_1_0__D mux_right_ipin_4.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_11.mux_l3_in_0__S mux_right_ipin_11.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_114 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_0.mux_l2_in_1_ chany_bottom_in[11] mux_right_ipin_0.mux_l1_in_2_/X
+ mux_right_ipin_0.mux_l2_in_0_/S mux_right_ipin_0.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_ipin_0.mux_l4_in_0__A1 mux_right_ipin_0.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_ipin_1.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_13_49 vpwr vgnd scs8hd_fill_2
XFILLER_57_132 vpwr vgnd scs8hd_fill_2
XFILLER_54_89 vgnd vpwr scs8hd_decap_3
XFILLER_54_67 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_12.mux_l1_in_0__A1 chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__43__A chany_top_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_63_135 vgnd vpwr scs8hd_decap_8
XFILLER_28_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_9.mux_l2_in_1__A1 mux_right_ipin_9.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_39_143 vgnd vpwr scs8hd_decap_3
XFILLER_39_110 vpwr vgnd scs8hd_fill_2
XFILLER_54_124 vgnd vpwr scs8hd_decap_12
XFILLER_24_15 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_11.scs8hd_buf_4_0_ mux_right_ipin_11.mux_l4_in_0_/X left_grid_pin_11_
+ vgnd vpwr scs8hd_buf_1
Xmux_right_ipin_0.mux_l1_in_2_ chany_top_in[5] chany_bottom_in[5] mux_right_ipin_0.mux_l1_in_2_/S
+ mux_right_ipin_0.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_49_56 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_12.mux_l2_in_3__S mux_right_ipin_12.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA__38__A chany_top_in[15] vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_5.mux_l3_in_0_ mux_right_ipin_5.mux_l2_in_1_/X mux_right_ipin_5.mux_l2_in_0_/X
+ mux_right_ipin_5.mux_l3_in_0_/S mux_right_ipin_5.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_10.mux_l4_in_0__S mux_right_ipin_10.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_51_105 vpwr vgnd scs8hd_fill_2
XFILLER_36_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_7.mux_l2_in_3__A1 chany_top_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_27_135 vgnd vpwr scs8hd_decap_8
XFILLER_35_36 vpwr vgnd scs8hd_fill_2
XFILLER_51_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_6.mux_l1_in_0__A0 chany_top_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_9.mux_l3_in_0__A1 mux_right_ipin_9.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_105 vgnd vpwr scs8hd_decap_4
XPHY_91 vgnd vpwr scs8hd_decap_3
Xmem_right_ipin_10.scs8hd_dfxbp_1_1_ prog_clk mux_right_ipin_10.mux_l1_in_0_/S mux_right_ipin_10.mux_l2_in_2_/S
+ mem_right_ipin_10.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XPHY_80 vgnd vpwr scs8hd_decap_3
XFILLER_2_84 vpwr vgnd scs8hd_fill_2
XFILLER_37_3 vpwr vgnd scs8hd_fill_2
X_57_ chany_bottom_in[16] chany_top_out[16] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_ipin_2.mux_l1_in_0__S mux_right_ipin_2.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_46_79 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_ipin_5.scs8hd_dfxbp_1_3__D mux_right_ipin_5.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_right_ipin_5.mux_l2_in_1_ chany_bottom_in[10] mux_right_ipin_5.mux_l1_in_2_/X
+ mux_right_ipin_5.mux_l2_in_0_/S mux_right_ipin_5.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_10.mux_l2_in_1__A1 chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__51__A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l1_in_2__A0 chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_16_49 vpwr vgnd scs8hd_fill_2
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
XANTENNA__46__A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_7_145 vgnd vpwr scs8hd_fill_1
XFILLER_7_123 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_8.scs8hd_dfxbp_1_1_ prog_clk mux_right_ipin_8.mux_l1_in_2_/S mux_right_ipin_8.mux_l2_in_3_/S
+ mem_right_ipin_8.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_right_ipin_14.mux_l2_in_3_ _28_/HI chany_top_in[19] mux_right_ipin_14.mux_l2_in_2_/S
+ mux_right_ipin_14.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_ipin_5.mux_l1_in_2_ chany_top_in[6] chany_bottom_in[6] mux_right_ipin_5.mux_l1_in_0_/S
+ mux_right_ipin_5.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_10.mux_l3_in_0__A1 mux_right_ipin_10.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_15 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_1.mux_l2_in_0__S mux_right_ipin_1.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l2_in_1__A0 chany_bottom_in[9] vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l2_in_0_ mux_right_ipin_0.mux_l1_in_1_/X mux_right_ipin_0.mux_l1_in_0_/X
+ mux_right_ipin_0.mux_l2_in_0_/S mux_right_ipin_0.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_81 vgnd vpwr scs8hd_decap_12
XFILLER_13_28 vpwr vgnd scs8hd_fill_2
XFILLER_1_118 vpwr vgnd scs8hd_fill_2
XFILLER_57_144 vpwr vgnd scs8hd_fill_2
XFILLER_57_100 vpwr vgnd scs8hd_fill_2
XFILLER_38_14 vgnd vpwr scs8hd_decap_3
XFILLER_38_47 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_2.mux_l2_in_3__A0 _30_/HI vgnd vpwr scs8hd_diode_2
XFILLER_44_90 vpwr vgnd scs8hd_fill_2
XFILLER_5_95 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_4.mux_l3_in_0__A0 mux_right_ipin_4.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_54_136 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_0.mux_l1_in_1_ chany_top_in[3] chany_bottom_in[3] mux_right_ipin_0.mux_l1_in_2_/S
+ mux_right_ipin_0.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_40_15 vpwr vgnd scs8hd_fill_2
XFILLER_49_35 vpwr vgnd scs8hd_fill_2
XFILLER_6_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.mux_l3_in_0__S mux_right_ipin_0.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_45_136 vgnd vpwr scs8hd_decap_8
XFILLER_45_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_7.scs8hd_dfxbp_1_2__D mux_right_ipin_7.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA__54__A chany_bottom_in[19] vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_14.mux_l4_in_0_ mux_right_ipin_14.mux_l3_in_1_/X mux_right_ipin_14.mux_l3_in_0_/X
+ mux_right_ipin_14.mux_l4_in_0_/S mux_right_ipin_14.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_14_93 vgnd vpwr scs8hd_decap_8
X_73_ chany_bottom_in[0] chany_top_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_36_125 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_6.mux_l2_in_1__S mux_right_ipin_6.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_ipin_6.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA__49__A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_6.mux_l1_in_0__A1 chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_4.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XPHY_92 vgnd vpwr scs8hd_decap_3
XPHY_81 vgnd vpwr scs8hd_decap_3
XFILLER_25_92 vpwr vgnd scs8hd_fill_2
XPHY_70 vgnd vpwr scs8hd_decap_3
Xmem_right_ipin_10.scs8hd_dfxbp_1_0_ prog_clk mux_right_ipin_9.mux_l4_in_0_/S mux_right_ipin_10.mux_l1_in_0_/S
+ mem_right_ipin_10.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
X_56_ chany_bottom_in[17] chany_top_out[17] vgnd vpwr scs8hd_buf_2
Xmux_right_ipin_0.scs8hd_buf_4_0_ mux_right_ipin_0.mux_l4_in_0_/X left_grid_pin_0_
+ vgnd vpwr scs8hd_buf_1
XFILLER_21_39 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_14.mux_l3_in_1_ mux_right_ipin_14.mux_l2_in_3_/X mux_right_ipin_14.mux_l2_in_2_/X
+ mux_right_ipin_14.mux_l3_in_0_/S mux_right_ipin_14.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_ipin_5.mux_l2_in_0_ mux_right_ipin_5.mux_l1_in_1_/X mux_right_ipin_5.mux_l1_in_0_/X
+ mux_right_ipin_5.mux_l2_in_0_/S mux_right_ipin_5.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_1.mux_l2_in_3__S mux_right_ipin_1.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_117 vgnd vpwr scs8hd_decap_3
XFILLER_16_9 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_4.mux_l1_in_2__A1 chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_36_80 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_ipin_13.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_39_ chany_top_in[14] chany_bottom_out[14] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_ipin_5.mux_l3_in_1__S mux_right_ipin_5.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_11.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA__62__A chany_bottom_in[11] vgnd vpwr scs8hd_diode_2
XFILLER_22_93 vgnd vpwr scs8hd_decap_4
Xmem_right_ipin_8.scs8hd_dfxbp_1_0_ prog_clk mux_right_ipin_7.mux_l4_in_0_/S mux_right_ipin_8.mux_l1_in_2_/S
+ mem_right_ipin_8.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_right_ipin_14.mux_l2_in_2_ chany_bottom_in[19] chany_top_in[11] mux_right_ipin_14.mux_l2_in_2_/S
+ mux_right_ipin_14.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_ipin_5.mux_l1_in_1_ chany_top_in[2] chany_bottom_in[2] mux_right_ipin_5.mux_l1_in_0_/S
+ mux_right_ipin_5.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_8_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_4.mux_l2_in_1__A1 mux_right_ipin_4.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_127 vpwr vgnd scs8hd_fill_2
XANTENNA__57__A chany_bottom_in[16] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_9.scs8hd_dfxbp_1_1__D mux_right_ipin_9.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_93 vgnd vpwr scs8hd_decap_8
XFILLER_12_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_14.mux_l2_in_0__A0 chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_38_59 vgnd vpwr scs8hd_decap_4
Xmem_right_ipin_3.scs8hd_dfxbp_1_3_ prog_clk mux_right_ipin_3.mux_l3_in_1_/S mux_right_ipin_3.mux_l4_in_0_/S
+ mem_right_ipin_3.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_48_101 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_2.mux_l2_in_3__A1 chany_top_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_44_80 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_1.mux_l1_in_0__A0 chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_54_115 vgnd vpwr scs8hd_decap_6
XFILLER_39_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_4.mux_l3_in_0__A1 mux_right_ipin_4.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_0.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_0.mux_l1_in_2_/S
+ mux_right_ipin_0.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_28 vgnd vpwr scs8hd_decap_3
XFILLER_49_14 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_12.mux_l2_in_2__A0 chany_bottom_in[17] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_13.mux_l2_in_1__S mux_right_ipin_13.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA__70__A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_30_71 vpwr vgnd scs8hd_fill_2
XFILLER_30_82 vgnd vpwr scs8hd_decap_8
X_72_ chany_bottom_in[1] chany_top_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_19_39 vpwr vgnd scs8hd_fill_2
XFILLER_27_115 vgnd vpwr scs8hd_fill_1
XFILLER_35_16 vgnd vpwr scs8hd_fill_1
XANTENNA__65__A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_93 vgnd vpwr scs8hd_decap_3
XFILLER_41_92 vgnd vpwr scs8hd_decap_12
XFILLER_41_70 vgnd vpwr scs8hd_fill_1
X_55_ chany_bottom_in[18] chany_top_out[18] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_ipin_12.mux_l3_in_1__A0 mux_right_ipin_12.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_97 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_14.mux_l3_in_0_ mux_right_ipin_14.mux_l2_in_1_/X mux_right_ipin_14.mux_l2_in_0_/X
+ mux_right_ipin_14.mux_l3_in_0_/S mux_right_ipin_14.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_46_59 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_ipin_0.mux_l1_in_0__A0 chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_11.scs8hd_dfxbp_1_2__D mux_right_ipin_11.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_12.mux_l3_in_1__S mux_right_ipin_12.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_62 vgnd vpwr scs8hd_decap_3
XFILLER_11_84 vpwr vgnd scs8hd_fill_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_8
X_38_ chany_top_in[15] chany_bottom_out[15] vgnd vpwr scs8hd_buf_2
XFILLER_57_58 vgnd vpwr scs8hd_decap_3
XFILLER_57_14 vgnd vpwr scs8hd_decap_4
XFILLER_11_132 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_6.scs8hd_buf_4_0__A mux_right_ipin_6.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_12.mux_l4_in_0__A0 mux_right_ipin_12.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_72 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_9.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_14.mux_l2_in_1_ chany_bottom_in[11] chany_top_in[3] mux_right_ipin_14.mux_l2_in_2_/S
+ mux_right_ipin_14.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_8_74 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_5.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_5.mux_l1_in_0_/S
+ mux_right_ipin_5.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__73__A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_60 vgnd vpwr scs8hd_fill_1
XFILLER_33_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_14.mux_l2_in_0__A1 mux_right_ipin_14.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_57_113 vgnd vpwr scs8hd_decap_4
XFILLER_54_15 vgnd vpwr scs8hd_decap_4
XFILLER_54_59 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_3.scs8hd_dfxbp_1_2_ prog_clk mux_right_ipin_3.mux_l2_in_3_/S mux_right_ipin_3.mux_l3_in_1_/S
+ mem_right_ipin_3.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_ipin_8.mux_l1_in_1__A0 chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__68__A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_0_142 vpwr vgnd scs8hd_fill_2
XFILLER_28_82 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_ipin_1.mux_l1_in_0__A1 chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XFILLER_5_42 vgnd vpwr scs8hd_decap_4
XFILLER_39_135 vgnd vpwr scs8hd_decap_8
XFILLER_49_26 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_ipin_12.mux_l2_in_2__A1 chany_top_in[13] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_13.scs8hd_dfxbp_1_1__D mux_right_ipin_13.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l1_in_1__S mux_left_ipin_0.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
X_71_ chany_bottom_in[2] chany_top_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_51_119 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_8.mux_l2_in_0__A0 mux_right_ipin_8.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_51_38 vgnd vpwr scs8hd_decap_4
XFILLER_51_16 vgnd vpwr scs8hd_decap_3
XFILLER_50_130 vgnd vpwr scs8hd_decap_12
XFILLER_4_6 vpwr vgnd scs8hd_fill_2
XPHY_94 vgnd vpwr scs8hd_decap_3
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XFILLER_33_119 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XFILLER_2_32 vpwr vgnd scs8hd_fill_2
X_54_ chany_bottom_in[19] chany_top_out[19] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_ipin_12.mux_l3_in_1__A1 mux_right_ipin_12.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_54 vpwr vgnd scs8hd_fill_2
XFILLER_24_108 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_ipin_6.mux_l2_in_2__A0 chany_bottom_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_62_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_2.mux_l2_in_1__S mux_right_ipin_2.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l1_in_0__A1 chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_2_3 vpwr vgnd scs8hd_fill_2
XFILLER_11_52 vgnd vpwr scs8hd_decap_3
XFILLER_52_70 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_0__D mux_left_ipin_0.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_8.mux_l1_in_2__S mux_right_ipin_8.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_3 vgnd vpwr scs8hd_decap_3
Xmem_right_ipin_13.scs8hd_dfxbp_1_3_ prog_clk mux_right_ipin_13.mux_l3_in_1_/S mux_right_ipin_13.mux_l4_in_0_/S
+ mem_right_ipin_13.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
X_37_ chany_top_in[16] chany_bottom_out[16] vgnd vpwr scs8hd_buf_2
XFILLER_20_111 vgnd vpwr scs8hd_decap_4
XFILLER_20_144 vpwr vgnd scs8hd_fill_2
XFILLER_11_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_12.mux_l4_in_0__A1 mux_right_ipin_12.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_84 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_14.mux_l2_in_0_ chany_bottom_in[3] mux_right_ipin_14.mux_l1_in_0_/X
+ mux_right_ipin_14.mux_l2_in_2_/S mux_right_ipin_14.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_8_42 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_6.mux_l3_in_1__A0 mux_right_ipin_6.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_1.mux_l3_in_1__S mux_right_ipin_1.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_ipin_15.scs8hd_dfxbp_1_0__D mux_right_ipin_14.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_83 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_7.mux_l2_in_2__S mux_right_ipin_7.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_57_136 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_3.scs8hd_dfxbp_1_1_ prog_clk mux_right_ipin_3.mux_l1_in_0_/S mux_right_ipin_3.mux_l2_in_3_/S
+ mem_right_ipin_3.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_ipin_8.mux_l1_in_1__A1 chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_0_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_6.mux_l4_in_0__A0 mux_right_ipin_6.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_72 vgnd vpwr scs8hd_decap_4
XFILLER_44_93 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_4.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_39_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_2.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_70_ chany_bottom_in[3] chany_top_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_51_109 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_3__D mux_right_ipin_0.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_106 vpwr vgnd scs8hd_fill_2
XFILLER_39_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_8.mux_l2_in_0__A1 mux_right_ipin_8.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_50_142 vgnd vpwr scs8hd_decap_4
XFILLER_51_28 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_11.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XPHY_95 vgnd vpwr scs8hd_decap_3
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_40 vgnd vpwr scs8hd_decap_3
XFILLER_25_51 vpwr vgnd scs8hd_fill_2
XFILLER_25_62 vpwr vgnd scs8hd_fill_2
XPHY_51 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XFILLER_51_9 vgnd vpwr scs8hd_fill_1
X_53_ chany_top_in[0] chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_2_11 vpwr vgnd scs8hd_fill_2
XFILLER_37_7 vgnd vpwr scs8hd_decap_4
XFILLER_2_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_6.mux_l2_in_2__A1 chany_top_in[11] vgnd vpwr scs8hd_diode_2
XFILLER_62_27 vgnd vpwr scs8hd_decap_4
XFILLER_15_109 vgnd vpwr scs8hd_decap_8
XFILLER_11_20 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_15.scs8hd_dfxbp_1_3__D mux_right_ipin_15.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_14_120 vgnd vpwr scs8hd_decap_3
XFILLER_36_83 vpwr vgnd scs8hd_fill_2
X_36_ chany_top_in[17] chany_bottom_out[17] vgnd vpwr scs8hd_buf_2
XFILLER_28_3 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_13.scs8hd_dfxbp_1_2_ prog_clk mux_right_ipin_13.mux_l2_in_3_/S mux_right_ipin_13.mux_l3_in_1_/S
+ mem_right_ipin_13.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_57_27 vgnd vpwr scs8hd_fill_1
XFILLER_7_127 vgnd vpwr scs8hd_decap_12
XFILLER_11_101 vpwr vgnd scs8hd_fill_2
XFILLER_22_30 vgnd vpwr scs8hd_fill_1
XFILLER_47_82 vpwr vgnd scs8hd_fill_2
XFILLER_14_9 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_14.scs8hd_buf_4_0__A mux_right_ipin_14.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_32 vgnd vpwr scs8hd_decap_8
XFILLER_8_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_6.mux_l3_in_1__A1 mux_right_ipin_6.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
X_19_ _19_/HI _19_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_ipin_14.mux_l2_in_3__A0 _28_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_14.mux_l2_in_2__S mux_right_ipin_14.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_2.scs8hd_dfxbp_1_2__D mux_right_ipin_2.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_right_ipin_3.scs8hd_dfxbp_1_0_ prog_clk mux_right_ipin_2.mux_l4_in_0_/S mux_right_ipin_3.mux_l1_in_0_/S
+ mem_right_ipin_3.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_ipin_3.mux_l2_in_0__A0 chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_6.mux_l4_in_0__A1 mux_right_ipin_6.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_14.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_14.mux_l1_in_0_/S
+ mux_right_ipin_14.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_48_126 vgnd vpwr scs8hd_decap_12
XFILLER_44_83 vgnd vpwr scs8hd_decap_4
XFILLER_44_72 vpwr vgnd scs8hd_fill_2
XFILLER_44_61 vpwr vgnd scs8hd_fill_2
XFILLER_5_11 vpwr vgnd scs8hd_fill_2
XFILLER_5_99 vpwr vgnd scs8hd_fill_2
XFILLER_5_66 vpwr vgnd scs8hd_fill_2
XFILLER_10_3 vgnd vpwr scs8hd_decap_8
XFILLER_54_107 vpwr vgnd scs8hd_fill_2
XFILLER_40_19 vgnd vpwr scs8hd_decap_12
XFILLER_49_39 vpwr vgnd scs8hd_fill_2
XFILLER_45_118 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_1.mux_l2_in_3_ _23_/HI chany_top_in[18] mux_right_ipin_1.mux_l2_in_2_/S
+ mux_right_ipin_1.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_14_64 vgnd vpwr scs8hd_decap_3
XFILLER_14_86 vgnd vpwr scs8hd_decap_6
XFILLER_30_63 vgnd vpwr scs8hd_decap_8
XFILLER_39_83 vpwr vgnd scs8hd_fill_2
XFILLER_55_82 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l2_in_2__A0 chany_bottom_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_58_3 vpwr vgnd scs8hd_fill_2
XFILLER_27_107 vpwr vgnd scs8hd_fill_2
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_143 vgnd vpwr scs8hd_decap_3
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_25_96 vpwr vgnd scs8hd_fill_2
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_74 vgnd vpwr scs8hd_decap_3
XFILLER_41_62 vgnd vpwr scs8hd_decap_8
XFILLER_41_51 vpwr vgnd scs8hd_fill_2
X_52_ chany_top_in[1] chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_2_67 vpwr vgnd scs8hd_fill_2
XFILLER_2_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_9.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_7.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_1.mux_l3_in_1__A0 mux_right_ipin_1.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_132 vpwr vgnd scs8hd_fill_2
XFILLER_52_83 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_4.scs8hd_dfxbp_1_1__D mux_right_ipin_4.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_9.mux_l1_in_0__S mux_right_ipin_9.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_right_ipin_13.scs8hd_dfxbp_1_1_ prog_clk mux_right_ipin_13.mux_l1_in_1_/S mux_right_ipin_13.mux_l2_in_3_/S
+ mem_right_ipin_13.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
X_35_ chany_top_in[18] chany_bottom_out[18] vgnd vpwr scs8hd_buf_2
Xmux_right_ipin_1.mux_l4_in_0_ mux_right_ipin_1.mux_l3_in_1_/X mux_right_ipin_1.mux_l3_in_0_/X
+ mux_right_ipin_1.mux_l4_in_0_/S mux_right_ipin_1.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_20_124 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_0.mux_l2_in_2__A0 chany_bottom_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_7_139 vgnd vpwr scs8hd_decap_6
XFILLER_7_106 vgnd vpwr scs8hd_decap_12
XFILLER_11_113 vpwr vgnd scs8hd_fill_2
XFILLER_22_64 vpwr vgnd scs8hd_fill_2
XFILLER_8_88 vpwr vgnd scs8hd_fill_2
XFILLER_8_99 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_14.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_1.mux_l4_in_0__A0 mux_right_ipin_1.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_40_3 vgnd vpwr scs8hd_decap_8
X_18_ _18_/HI _18_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_ipin_14.mux_l2_in_3__A1 chany_top_in[19] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l1_in_2__S mux_right_ipin_4.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_6.mux_l2_in_3_ _17_/HI chany_top_in[19] mux_right_ipin_6.mux_l2_in_3_/S
+ mux_right_ipin_6.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_ipin_13.mux_l1_in_0__A0 chany_top_in[0] vgnd vpwr scs8hd_diode_2
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_53 vpwr vgnd scs8hd_fill_2
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_52 vgnd vpwr scs8hd_decap_8
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_120 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_1.mux_l3_in_1_ mux_right_ipin_1.mux_l2_in_3_/X mux_right_ipin_1.mux_l2_in_2_/X
+ mux_right_ipin_1.mux_l3_in_1_/S mux_right_ipin_1.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_ipin_0.mux_l3_in_1__A0 mux_left_ipin_0.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_58_93 vpwr vgnd scs8hd_fill_2
XFILLER_12_7 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_8.mux_l2_in_0__S mux_right_ipin_8.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_19 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_1.scs8hd_buf_4_0__A mux_right_ipin_1.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_134 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_3.mux_l2_in_0__A1 mux_right_ipin_3.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_48_138 vgnd vpwr scs8hd_decap_8
XFILLER_60_72 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_8.mux_l2_in_3__A0 _19_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_3.mux_l2_in_2__S mux_right_ipin_3.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_32 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_1.mux_l2_in_2_ chany_bottom_in[18] chany_top_in[12] mux_right_ipin_1.mux_l2_in_2_/S
+ mux_right_ipin_1.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_ipin_0.mux_l4_in_0__A0 mux_left_ipin_0.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_1.mux_l2_in_2__A1 chany_top_in[12] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_2__S mux_left_ipin_0.mux_l2_in_2_/S vgnd vpwr scs8hd_diode_2
XFILLER_44_130 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_6.mux_l4_in_0_ mux_right_ipin_6.mux_l3_in_1_/X mux_right_ipin_6.mux_l3_in_0_/X
+ mux_right_ipin_6.mux_l4_in_0_/S mux_right_ipin_6.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_36_119 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_6.scs8hd_dfxbp_1_0__D mux_right_ipin_5.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.mux_l3_in_0__S mux_right_ipin_7.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_11.mux_l2_in_1__A0 chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XPHY_20 vgnd vpwr scs8hd_decap_3
Xmem_left_ipin_0.scs8hd_dfxbp_1_3_ prog_clk mux_left_ipin_0.mux_l3_in_1_/S mux_left_ipin_0.mux_l4_in_0_/S
+ mem_left_ipin_0.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_97 vgnd vpwr scs8hd_decap_3
XPHY_86 vgnd vpwr scs8hd_decap_3
XFILLER_41_30 vpwr vgnd scs8hd_fill_2
XFILLER_25_75 vpwr vgnd scs8hd_fill_2
XPHY_75 vgnd vpwr scs8hd_decap_3
X_51_ chany_top_in[2] chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_32_133 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_1.mux_l3_in_1__A1 mux_right_ipin_1.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_144 vpwr vgnd scs8hd_fill_2
XFILLER_11_33 vpwr vgnd scs8hd_fill_2
XFILLER_11_44 vgnd vpwr scs8hd_decap_8
XFILLER_11_88 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_6.mux_l3_in_1_ mux_right_ipin_6.mux_l2_in_3_/X mux_right_ipin_6.mux_l2_in_2_/X
+ mux_right_ipin_6.mux_l3_in_1_/S mux_right_ipin_6.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_ipin_6.scs8hd_buf_4_0_ mux_right_ipin_6.mux_l4_in_0_/X left_grid_pin_6_
+ vgnd vpwr scs8hd_buf_1
XFILLER_36_63 vgnd vpwr scs8hd_fill_1
Xmem_right_ipin_13.scs8hd_dfxbp_1_0_ prog_clk mux_right_ipin_12.mux_l4_in_0_/S mux_right_ipin_13.mux_l1_in_1_/S
+ mem_right_ipin_13.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
X_34_ chany_top_in[19] chany_bottom_out[19] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_ipin_8.mux_l2_in_3__S mux_right_ipin_8.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_11.mux_l3_in_0__A0 mux_right_ipin_11.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_2__A1 chany_top_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_20_136 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_6.mux_l4_in_0__S mux_right_ipin_6.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_57_18 vgnd vpwr scs8hd_fill_1
XFILLER_7_118 vgnd vpwr scs8hd_fill_1
XFILLER_22_32 vpwr vgnd scs8hd_fill_2
XFILLER_22_43 vgnd vpwr scs8hd_decap_12
XFILLER_0_3 vgnd vpwr scs8hd_decap_4
XFILLER_47_62 vgnd vpwr scs8hd_decap_4
XFILLER_47_51 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_1.mux_l4_in_0__A1 mux_right_ipin_1.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_3 vgnd vpwr scs8hd_decap_12
X_17_ _17_/HI _17_/LO vgnd vpwr scs8hd_conb_1
Xmux_right_ipin_6.mux_l2_in_2_ chany_bottom_in[19] chany_top_in[11] mux_right_ipin_6.mux_l2_in_3_/S
+ mux_right_ipin_6.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_15.mux_l2_in_0__S mux_right_ipin_15.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_32 vpwr vgnd scs8hd_fill_2
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_ipin_13.mux_l1_in_0__A1 chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_33_75 vpwr vgnd scs8hd_fill_2
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_ipin_1.mux_l3_in_0_ mux_right_ipin_1.mux_l2_in_1_/X mux_right_ipin_1.mux_l2_in_0_/X
+ mux_right_ipin_1.mux_l3_in_1_/S mux_right_ipin_1.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_3_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.mux_l3_in_1__A1 mux_left_ipin_0.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_ipin_6.scs8hd_dfxbp_1_3__D mux_right_ipin_6.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_54_19 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_12.scs8hd_buf_4_0_ mux_right_ipin_12.mux_l4_in_0_/X left_grid_pin_12_
+ vgnd vpwr scs8hd_buf_1
XFILLER_0_113 vpwr vgnd scs8hd_fill_2
XFILLER_44_30 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_10.mux_l2_in_2__S mux_right_ipin_10.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_60_84 vgnd vpwr scs8hd_decap_6
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XFILLER_5_46 vgnd vpwr scs8hd_fill_1
XFILLER_39_106 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_8.mux_l2_in_3__A1 chany_top_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_53_142 vgnd vpwr scs8hd_decap_4
XFILLER_53_120 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_1.mux_l2_in_1_ chany_bottom_in[12] mux_right_ipin_1.mux_l1_in_2_/X
+ mux_right_ipin_1.mux_l2_in_2_/S mux_right_ipin_1.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_14.mux_l3_in_0__S mux_right_ipin_14.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l4_in_0__A1 mux_left_ipin_0.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_7.mux_l1_in_0__A0 chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_6.scs8hd_dfxbp_1_3_ prog_clk mux_right_ipin_6.mux_l3_in_1_/S mux_right_ipin_6.mux_l4_in_0_/S
+ mem_right_ipin_6.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_39_52 vgnd vpwr scs8hd_decap_3
XFILLER_55_95 vgnd vpwr scs8hd_decap_4
XFILLER_55_62 vgnd vpwr scs8hd_decap_3
XFILLER_55_40 vpwr vgnd scs8hd_fill_2
XFILLER_44_142 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_11.mux_l2_in_1__A1 chany_top_in[2] vgnd vpwr scs8hd_diode_2
XPHY_98 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_decap_3
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
Xmem_left_ipin_0.scs8hd_dfxbp_1_2_ prog_clk mux_left_ipin_0.mux_l2_in_2_/S mux_left_ipin_0.mux_l3_in_1_/S
+ mem_left_ipin_0.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XFILLER_25_10 vpwr vgnd scs8hd_fill_2
XFILLER_25_43 vpwr vgnd scs8hd_fill_2
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_76 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_5.mux_l1_in_2__A0 chany_top_in[6] vgnd vpwr scs8hd_diode_2
X_50_ chany_top_in[3] chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_2_36 vgnd vpwr scs8hd_decap_3
XFILLER_17_120 vpwr vgnd scs8hd_fill_2
XFILLER_32_145 vgnd vpwr scs8hd_fill_1
XFILLER_63_3 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_10.mux_l2_in_3_ _24_/HI chany_top_in[15] mux_right_ipin_10.mux_l2_in_2_/S
+ mux_right_ipin_10.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_ipin_1.mux_l1_in_2_ chany_top_in[6] chany_bottom_in[6] mux_right_ipin_1.mux_l1_in_0_/S
+ mux_right_ipin_1.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_15.mux_l2_in_3__S mux_right_ipin_15.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_12 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_13.mux_l4_in_0__S mux_right_ipin_13.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_6.mux_l3_in_0_ mux_right_ipin_6.mux_l2_in_1_/X mux_right_ipin_6.mux_l2_in_0_/X
+ mux_right_ipin_6.mux_l3_in_1_/S mux_right_ipin_6.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_52_41 vpwr vgnd scs8hd_fill_2
XFILLER_14_145 vgnd vpwr scs8hd_fill_1
X_33_ _33_/HI _33_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mem_right_ipin_10.scs8hd_dfxbp_1_0__D mux_right_ipin_9.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_11.mux_l3_in_0__A1 mux_right_ipin_11.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_ipin_8.scs8hd_dfxbp_1_2__D mux_right_ipin_8.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_5.mux_l2_in_1__A0 chany_bottom_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_22_22 vgnd vpwr scs8hd_decap_8
XFILLER_22_88 vgnd vpwr scs8hd_decap_4
XFILLER_47_30 vgnd vpwr scs8hd_decap_6
XFILLER_63_62 vgnd vpwr scs8hd_decap_12
XFILLER_8_68 vgnd vpwr scs8hd_decap_4
XFILLER_8_46 vgnd vpwr scs8hd_decap_3
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_6.mux_l2_in_1_ chany_bottom_in[11] chany_top_in[3] mux_right_ipin_6.mux_l2_in_3_/S
+ mux_right_ipin_6.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_5.mux_l1_in_0__S mux_right_ipin_5.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_ipin_10.mux_l4_in_0_ mux_right_ipin_10.mux_l3_in_1_/X mux_right_ipin_10.mux_l3_in_0_/X
+ mux_right_ipin_10.mux_l4_in_0_/S mux_right_ipin_10.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_3_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_3.mux_l2_in_3__A0 _31_/HI vgnd vpwr scs8hd_diode_2
XFILLER_58_40 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_9.scs8hd_buf_4_0__A mux_right_ipin_9.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_5.mux_l3_in_0__A0 mux_right_ipin_5.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_2__S mux_right_ipin_0.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_32 vpwr vgnd scs8hd_fill_2
XFILLER_60_41 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_15.mux_l2_in_3_ _29_/HI chany_top_in[12] mux_right_ipin_15.mux_l2_in_0_/S
+ mux_right_ipin_15.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_62_121 vgnd vpwr scs8hd_decap_12
XFILLER_39_118 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_4.mux_l2_in_0__S mux_right_ipin_4.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_1.mux_l2_in_0_ mux_right_ipin_1.mux_l1_in_1_/X mux_right_ipin_1.mux_l1_in_0_/X
+ mux_right_ipin_1.mux_l2_in_2_/S mux_right_ipin_1.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_ipin_10.mux_l3_in_1_ mux_right_ipin_10.mux_l2_in_3_/X mux_right_ipin_10.mux_l2_in_2_/X
+ mux_right_ipin_10.mux_l3_in_1_/S mux_right_ipin_10.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_14_23 vgnd vpwr scs8hd_decap_8
XFILLER_14_56 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_7.mux_l1_in_0__A1 chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_39_31 vgnd vpwr scs8hd_fill_1
XFILLER_39_42 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_ipin_5.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_6.scs8hd_dfxbp_1_2_ prog_clk mux_right_ipin_6.mux_l2_in_3_/S mux_right_ipin_6.mux_l3_in_1_/S
+ mem_right_ipin_6.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_39_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_10.scs8hd_dfxbp_1_3__D mux_right_ipin_10.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_right_ipin_1.scs8hd_buf_4_0_ mux_right_ipin_1.mux_l4_in_0_/X left_grid_pin_1_
+ vgnd vpwr scs8hd_buf_1
XFILLER_35_132 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_3.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_0.scs8hd_dfxbp_1_1_ prog_clk mux_left_ipin_0.mux_l1_in_0_/S mux_left_ipin_0.mux_l2_in_2_/S
+ mem_left_ipin_0.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_26_121 vgnd vpwr scs8hd_decap_12
XPHY_99 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_decap_3
XFILLER_41_135 vgnd vpwr scs8hd_decap_8
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_25_22 vpwr vgnd scs8hd_fill_2
XFILLER_25_55 vgnd vpwr scs8hd_decap_4
XPHY_55 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_77 vgnd vpwr scs8hd_decap_3
XFILLER_2_15 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_5.mux_l1_in_2__A1 chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_17_143 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_10.mux_l2_in_2_ chany_bottom_in[15] chany_top_in[7] mux_right_ipin_10.mux_l2_in_2_/S
+ mux_right_ipin_10.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_ipin_1.mux_l1_in_1_ chany_top_in[2] chany_bottom_in[2] mux_right_ipin_1.mux_l1_in_0_/S
+ mux_right_ipin_1.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_3.mux_l3_in_0__S mux_right_ipin_3.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_15.mux_l4_in_0_ mux_right_ipin_15.mux_l3_in_1_/X mux_right_ipin_15.mux_l3_in_0_/X
+ ccff_tail mux_right_ipin_15.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_ipin_12.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_36_32 vpwr vgnd scs8hd_fill_2
XFILLER_36_76 vgnd vpwr scs8hd_decap_4
XFILLER_36_87 vgnd vpwr scs8hd_decap_3
XFILLER_52_53 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_0.mux_l3_in_0__S mux_left_ipin_0.mux_l3_in_1_/S vgnd vpwr scs8hd_diode_2
X_32_ _32_/HI _32_/LO vgnd vpwr scs8hd_conb_1
XFILLER_35_8 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_10.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_9.mux_l2_in_1__S mux_right_ipin_9.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_105 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_5.mux_l2_in_1__A1 mux_right_ipin_5.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_12.mux_l1_in_0__S mux_right_ipin_12.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_63_74 vgnd vpwr scs8hd_decap_12
XFILLER_47_86 vpwr vgnd scs8hd_fill_2
XFILLER_19_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_15.mux_l2_in_0__A0 chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_15.mux_l3_in_1_ mux_right_ipin_15.mux_l2_in_3_/X mux_right_ipin_15.mux_l2_in_2_/X
+ mux_right_ipin_15.mux_l3_in_0_/S mux_right_ipin_15.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_ipin_6.mux_l2_in_0_ chany_bottom_in[3] mux_right_ipin_6.mux_l1_in_0_/X
+ mux_right_ipin_6.mux_l2_in_3_/S mux_right_ipin_6.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_4.mux_l2_in_3__S mux_right_ipin_4.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_2.mux_l4_in_0__S mux_right_ipin_2.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_ipin_3.mux_l2_in_3__A1 chany_top_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_3_112 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l1_in_0__A0 chany_top_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_5.mux_l3_in_0__A1 mux_right_ipin_5.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_8.mux_l3_in_1__S mux_right_ipin_8.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_57_119 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_12.scs8hd_dfxbp_1_2__D mux_right_ipin_12.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_13.mux_l2_in_2__A0 chany_bottom_in[18] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_11.mux_l2_in_0__S mux_right_ipin_11.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_44_87 vgnd vpwr scs8hd_fill_1
XFILLER_44_76 vgnd vpwr scs8hd_decap_4
XFILLER_44_65 vgnd vpwr scs8hd_decap_4
XFILLER_44_32 vgnd vpwr scs8hd_decap_4
XFILLER_60_53 vgnd vpwr scs8hd_decap_12
XFILLER_5_15 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_15.mux_l2_in_2_ chany_bottom_in[12] chany_top_in[4] mux_right_ipin_15.mux_l2_in_0_/S
+ mux_right_ipin_15.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_62_133 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_0.mux_l1_in_2__A0 chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_53_100 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_10.mux_l3_in_0_ mux_right_ipin_10.mux_l2_in_1_/X mux_right_ipin_10.mux_l2_in_0_/X
+ mux_right_ipin_10.mux_l3_in_1_/S mux_right_ipin_10.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_55_53 vpwr vgnd scs8hd_fill_2
XFILLER_55_31 vgnd vpwr scs8hd_decap_3
Xmem_right_ipin_6.scs8hd_dfxbp_1_1_ prog_clk mux_right_ipin_6.mux_l1_in_0_/S mux_right_ipin_6.mux_l2_in_3_/S
+ mem_right_ipin_6.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_ipin_13.mux_l3_in_1__A0 mux_right_ipin_13.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_144 vpwr vgnd scs8hd_fill_2
XFILLER_6_91 vgnd vpwr scs8hd_fill_1
Xmem_left_ipin_0.scs8hd_dfxbp_1_0_ prog_clk ccff_head mux_left_ipin_0.mux_l1_in_0_/S
+ mem_left_ipin_0.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_26_133 vgnd vpwr scs8hd_decap_12
XPHY_89 vgnd vpwr scs8hd_decap_3
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_78 vgnd vpwr scs8hd_decap_3
XFILLER_41_55 vgnd vpwr scs8hd_decap_6
XFILLER_2_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_10.mux_l3_in_0__S mux_right_ipin_10.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l2_in_1__A0 chany_bottom_in[11] vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_1.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_1.mux_l1_in_0_/S
+ mux_right_ipin_1.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_ipin_10.mux_l2_in_1_ chany_bottom_in[7] chany_top_in[3] mux_right_ipin_10.mux_l2_in_2_/S
+ mux_right_ipin_10.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_114 vpwr vgnd scs8hd_fill_2
XFILLER_23_136 vgnd vpwr scs8hd_decap_8
XFILLER_14_125 vgnd vpwr scs8hd_decap_3
XFILLER_36_66 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_13.mux_l4_in_0__A0 mux_right_ipin_13.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
X_31_ _31_/HI _31_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mem_right_ipin_14.scs8hd_dfxbp_1_1__D mux_right_ipin_14.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_92 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_8.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_11_117 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_0.mux_l3_in_0__A0 mux_right_ipin_0.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_68 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_11.mux_l2_in_3__S mux_right_ipin_11.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_47_54 vpwr vgnd scs8hd_fill_2
XFILLER_47_43 vpwr vgnd scs8hd_fill_2
XFILLER_63_86 vgnd vpwr scs8hd_decap_12
XFILLER_63_53 vgnd vpwr scs8hd_decap_8
XFILLER_6_110 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_15.mux_l2_in_0__A1 mux_right_ipin_15.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_15.mux_l3_in_0_ mux_right_ipin_15.mux_l2_in_1_/X mux_right_ipin_15.mux_l2_in_0_/X
+ mux_right_ipin_15.mux_l3_in_0_/S mux_right_ipin_15.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_15.mux_l3_in_1__S mux_right_ipin_15.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_ipin_9.mux_l1_in_1__A0 chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_33_45 vgnd vpwr scs8hd_fill_1
XFILLER_58_97 vgnd vpwr scs8hd_decap_3
XFILLER_58_75 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_2.mux_l1_in_0__A1 chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_15.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
XFILLER_0_71 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_13.mux_l2_in_2__A1 chany_top_in[14] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_1.scs8hd_dfxbp_1_0__D mux_right_ipin_0.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_138 vpwr vgnd scs8hd_fill_2
XFILLER_56_131 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_1.mux_l1_in_0__S mux_right_ipin_1.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_45 vgnd vpwr scs8hd_decap_8
XFILLER_28_78 vpwr vgnd scs8hd_fill_2
XFILLER_44_99 vpwr vgnd scs8hd_fill_2
XFILLER_44_22 vgnd vpwr scs8hd_decap_8
XFILLER_60_76 vgnd vpwr scs8hd_decap_4
XFILLER_60_65 vgnd vpwr scs8hd_decap_3
XFILLER_60_32 vgnd vpwr scs8hd_decap_4
XFILLER_5_38 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_15.mux_l2_in_1_ chany_bottom_in[4] chany_top_in[2] mux_right_ipin_15.mux_l2_in_0_/S
+ mux_right_ipin_15.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_ipin_6.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_6.mux_l1_in_0_/S
+ mux_right_ipin_6.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_62_145 vgnd vpwr scs8hd_fill_1
Xmux_left_ipin_0.mux_l2_in_3_ _21_/HI chany_top_in[16] mux_left_ipin_0.mux_l2_in_2_/S
+ mux_left_ipin_0.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_9.mux_l2_in_0__A0 mux_right_ipin_9.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_2__A1 chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_53_123 vgnd vpwr scs8hd_decap_12
XFILLER_14_69 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_6.scs8hd_dfxbp_1_0_ prog_clk mux_right_ipin_5.mux_l4_in_0_/S mux_right_ipin_6.mux_l1_in_0_/S
+ mem_right_ipin_6.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_ipin_13.mux_l3_in_1__A1 mux_right_ipin_13.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_112 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_7.mux_l2_in_2__A0 chany_bottom_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_41_104 vgnd vpwr scs8hd_decap_12
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XFILLER_25_35 vgnd vpwr scs8hd_decap_6
XFILLER_26_145 vgnd vpwr scs8hd_fill_1
XFILLER_41_34 vpwr vgnd scs8hd_fill_2
XPHY_79 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_0.mux_l2_in_0__S mux_right_ipin_0.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_79 vpwr vgnd scs8hd_fill_2
XPHY_57 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XFILLER_17_101 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_0.mux_l2_in_1__A1 mux_right_ipin_0.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_123 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_10.mux_l2_in_0_ chany_bottom_in[3] mux_right_ipin_10.mux_l1_in_0_/X
+ mux_right_ipin_10.mux_l2_in_2_/S mux_right_ipin_10.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_11_37 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_1.scs8hd_dfxbp_1_3_ prog_clk mux_right_ipin_1.mux_l3_in_1_/S mux_right_ipin_1.mux_l4_in_0_/S
+ mem_right_ipin_1.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_52_11 vgnd vpwr scs8hd_decap_3
XFILLER_14_137 vgnd vpwr scs8hd_decap_8
XFILLER_36_23 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_ipin_10.mux_l2_in_0__A0 chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_13.mux_l4_in_0__A1 mux_right_ipin_13.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_52_66 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_0.mux_l4_in_0_ mux_left_ipin_0.mux_l3_in_1_/X mux_left_ipin_0.mux_l3_in_0_/X
+ mux_left_ipin_0.mux_l4_in_0_/S mux_left_ipin_0.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
X_30_ _30_/HI _30_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_ipin_7.mux_l3_in_1__A0 mux_right_ipin_7.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_107 vpwr vgnd scs8hd_fill_2
XFILLER_3_71 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_1.scs8hd_dfxbp_1_3__D mux_right_ipin_1.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l3_in_0__A1 mux_right_ipin_0.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_47_99 vgnd vpwr scs8hd_decap_8
XFILLER_47_66 vgnd vpwr scs8hd_fill_1
XFILLER_63_98 vgnd vpwr scs8hd_decap_12
XFILLER_6_133 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_5.mux_l2_in_1__S mux_right_ipin_5.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_left_ipin_0.mux_l3_in_1_ mux_left_ipin_0.mux_l2_in_3_/X mux_left_ipin_0.mux_l2_in_2_/X
+ mux_left_ipin_0.mux_l3_in_1_/S mux_left_ipin_0.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_17_36 vpwr vgnd scs8hd_fill_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_ipin_9.mux_l1_in_1__A1 chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.mux_l4_in_0__A0 mux_right_ipin_7.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_79 vgnd vpwr scs8hd_decap_4
XFILLER_58_87 vgnd vpwr scs8hd_decap_3
XFILLER_3_136 vgnd vpwr scs8hd_decap_8
XFILLER_24_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_3.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_9_81 vpwr vgnd scs8hd_fill_2
XFILLER_0_117 vgnd vpwr scs8hd_decap_4
XFILLER_56_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_1__D mux_left_ipin_0.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_44_45 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_ipin_1.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l2_in_3__S mux_right_ipin_0.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_15.mux_l2_in_0_ chany_bottom_in[2] mux_right_ipin_15.mux_l1_in_0_/X
+ mux_right_ipin_15.mux_l2_in_0_/S mux_right_ipin_15.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_47_143 vgnd vpwr scs8hd_decap_3
XFILLER_47_121 vgnd vpwr scs8hd_fill_1
Xmux_left_ipin_0.mux_l2_in_2_ chany_bottom_in[16] chany_top_in[10] mux_left_ipin_0.mux_l2_in_2_/S
+ mux_left_ipin_0.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_9.mux_l2_in_0__A1 mux_right_ipin_9.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l3_in_1__S mux_right_ipin_4.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_4.scs8hd_buf_4_0__A mux_right_ipin_4.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_143 vgnd vpwr scs8hd_decap_3
XFILLER_39_34 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_10.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_6_93 vpwr vgnd scs8hd_fill_2
XFILLER_6_71 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_7.mux_l2_in_2__A1 chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_41_116 vgnd vpwr scs8hd_decap_6
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XFILLER_25_47 vgnd vpwr scs8hd_fill_1
XPHY_58 vgnd vpwr scs8hd_decap_3
XPHY_69 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_3.scs8hd_dfxbp_1_2__D mux_right_ipin_3.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_13.mux_l1_in_1__S mux_right_ipin_13.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_135 vgnd vpwr scs8hd_decap_8
XFILLER_56_6 vgnd vpwr scs8hd_decap_12
XFILLER_11_16 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_1.scs8hd_dfxbp_1_2_ prog_clk mux_right_ipin_1.mux_l2_in_2_/S mux_right_ipin_1.mux_l3_in_1_/S
+ mem_right_ipin_1.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_52_45 vpwr vgnd scs8hd_fill_2
XFILLER_52_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_10.mux_l2_in_0__A1 mux_right_ipin_10.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_52_89 vgnd vpwr scs8hd_decap_3
XANTENNA__41__A chany_top_in[12] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l1_in_1__A0 chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.mux_l3_in_1__A1 mux_right_ipin_7.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_90 vpwr vgnd scs8hd_fill_2
XFILLER_54_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_15.mux_l2_in_3__A0 _29_/HI vgnd vpwr scs8hd_diode_2
XFILLER_22_15 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_12.mux_l2_in_1__S mux_right_ipin_12.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA__36__A chany_top_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_8_17 vgnd vpwr scs8hd_decap_12
XFILLER_10_141 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_10.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_10.mux_l1_in_0_/S
+ mux_right_ipin_10.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_6_145 vgnd vpwr scs8hd_fill_1
Xmux_left_ipin_0.mux_l3_in_0_ mux_left_ipin_0.mux_l2_in_1_/X mux_left_ipin_0.mux_l2_in_0_/X
+ mux_left_ipin_0.mux_l3_in_1_/S mux_left_ipin_0.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_ipin_4.mux_l2_in_0__A0 mux_right_ipin_4.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_7.mux_l4_in_0__A1 mux_right_ipin_7.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_58_11 vgnd vpwr scs8hd_decap_8
XFILLER_0_40 vgnd vpwr scs8hd_fill_1
XFILLER_17_3 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_ipin_5.scs8hd_dfxbp_1_1__D mux_right_ipin_5.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_11.mux_l3_in_1__S mux_right_ipin_11.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_2.mux_l2_in_2__A0 chany_bottom_in[15] vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.mux_l2_in_1_ chany_bottom_in[10] mux_left_ipin_0.mux_l1_in_2_/X mux_left_ipin_0.mux_l2_in_2_/S
+ mux_left_ipin_0.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmem_right_ipin_11.scs8hd_dfxbp_1_3_ prog_clk mux_right_ipin_11.mux_l3_in_0_/S mux_right_ipin_11.mux_l4_in_0_/S
+ mem_right_ipin_11.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_38_133 vgnd vpwr scs8hd_decap_12
XFILLER_30_15 vgnd vpwr scs8hd_decap_12
XFILLER_44_103 vpwr vgnd scs8hd_fill_2
XFILLER_39_57 vpwr vgnd scs8hd_fill_2
XFILLER_39_79 vpwr vgnd scs8hd_fill_2
XFILLER_55_78 vpwr vgnd scs8hd_fill_2
XFILLER_55_67 vpwr vgnd scs8hd_fill_2
XANTENNA__44__A chany_top_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_6_83 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_8.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_15.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_15.mux_l1_in_0_/S
+ mux_right_ipin_15.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_2.mux_l3_in_1__A0 mux_right_ipin_2.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_41_47 vpwr vgnd scs8hd_fill_2
XANTENNA__39__A chany_top_in[14] vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.mux_l1_in_2_ chany_top_in[4] chany_bottom_in[4] mux_left_ipin_0.mux_l1_in_0_/S
+ mux_left_ipin_0.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_ipin_6.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_15_70 vgnd vpwr scs8hd_fill_1
XFILLER_32_106 vgnd vpwr scs8hd_decap_8
XFILLER_49_6 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_9.scs8hd_dfxbp_1_3_ prog_clk mux_right_ipin_9.mux_l3_in_0_/S mux_right_ipin_9.mux_l4_in_0_/S
+ mem_right_ipin_9.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
Xmem_right_ipin_1.scs8hd_dfxbp_1_1_ prog_clk mux_right_ipin_1.mux_l1_in_0_/S mux_right_ipin_1.mux_l2_in_2_/S
+ mem_right_ipin_1.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_right_ipin_2.mux_l2_in_3_ _30_/HI chany_top_in[15] mux_right_ipin_2.mux_l2_in_0_/S
+ mux_right_ipin_2.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_36_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_4.mux_l1_in_1__A1 chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_9_143 vgnd vpwr scs8hd_decap_3
XFILLER_47_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_15.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_2.mux_l4_in_0__A0 mux_right_ipin_2.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_15.mux_l2_in_3__A1 chany_top_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_11_109 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_13.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_14.mux_l1_in_0__A0 chany_top_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_7.scs8hd_dfxbp_1_0__D mux_right_ipin_6.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_29 vpwr vgnd scs8hd_fill_2
XANTENNA__52__A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_12_93 vgnd vpwr scs8hd_decap_4
XFILLER_37_90 vpwr vgnd scs8hd_fill_2
XFILLER_17_49 vpwr vgnd scs8hd_fill_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_ipin_4.mux_l2_in_0__A1 mux_right_ipin_4.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_15 vgnd vpwr scs8hd_decap_12
XFILLER_33_48 vpwr vgnd scs8hd_fill_2
XFILLER_3_116 vpwr vgnd scs8hd_fill_2
XFILLER_58_23 vpwr vgnd scs8hd_fill_2
XANTENNA__47__A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_12.mux_l1_in_2__A0 chany_top_in[7] vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_2.mux_l4_in_0_ mux_right_ipin_2.mux_l3_in_1_/X mux_right_ipin_2.mux_l3_in_0_/X
+ mux_right_ipin_2.mux_l4_in_0_/S mux_right_ipin_2.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_9.mux_l2_in_3__A0 _20_/HI vgnd vpwr scs8hd_diode_2
XFILLER_28_15 vgnd vpwr scs8hd_decap_12
XFILLER_44_36 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_1.mux_l2_in_1__S mux_right_ipin_1.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_2.mux_l2_in_2__A1 chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_47_123 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_11.scs8hd_dfxbp_1_2_ prog_clk mux_right_ipin_11.mux_l2_in_3_/S mux_right_ipin_11.mux_l3_in_0_/S
+ mem_right_ipin_11.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_left_ipin_0.mux_l2_in_0_ mux_left_ipin_0.mux_l1_in_1_/X mux_left_ipin_0.mux_l1_in_0_/X
+ mux_left_ipin_0.mux_l2_in_2_/S mux_left_ipin_0.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_ipin_7.mux_l2_in_3_ _18_/HI chany_top_in[12] mux_right_ipin_7.mux_l2_in_0_/S
+ mux_right_ipin_7.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_38_112 vgnd vpwr scs8hd_decap_8
XFILLER_38_145 vgnd vpwr scs8hd_fill_1
XFILLER_53_104 vpwr vgnd scs8hd_fill_2
XFILLER_30_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_12.mux_l2_in_1__A0 chany_bottom_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_55_57 vpwr vgnd scs8hd_fill_2
XFILLER_44_126 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_2.mux_l3_in_1_ mux_right_ipin_2.mux_l2_in_3_/X mux_right_ipin_2.mux_l2_in_2_/X
+ mux_right_ipin_2.mux_l3_in_0_/S mux_right_ipin_2.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_29_123 vgnd vpwr scs8hd_decap_12
XANTENNA__60__A chany_bottom_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_20_60 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_12.scs8hd_buf_4_0__A mux_right_ipin_12.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_71 vpwr vgnd scs8hd_fill_2
XFILLER_20_93 vgnd vpwr scs8hd_decap_3
XFILLER_50_118 vgnd vpwr scs8hd_decap_12
XPHY_16 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_2.mux_l3_in_1__A1 mux_right_ipin_2.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_7.scs8hd_buf_4_0_ mux_right_ipin_7.mux_l4_in_0_/X left_grid_pin_7_
+ vgnd vpwr scs8hd_buf_1
XANTENNA_mux_right_ipin_0.mux_l3_in_1__S mux_right_ipin_0.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_7.scs8hd_dfxbp_1_3__D mux_right_ipin_7.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA__55__A chany_bottom_in[18] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_10.mux_l2_in_3__A0 _24_/HI vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.mux_l1_in_1_ chany_top_in[2] chany_bottom_in[2] mux_left_ipin_0.mux_l1_in_0_/S
+ mux_left_ipin_0.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_17_104 vpwr vgnd scs8hd_fill_2
XFILLER_31_92 vgnd vpwr scs8hd_fill_1
Xmem_right_ipin_9.scs8hd_dfxbp_1_2_ prog_clk mux_right_ipin_9.mux_l2_in_1_/S mux_right_ipin_9.mux_l3_in_0_/S
+ mem_right_ipin_9.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_ipin_12.mux_l3_in_0__A0 mux_right_ipin_12.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_6.mux_l2_in_2__S mux_right_ipin_6.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_2.mux_l2_in_2_ chany_bottom_in[15] chany_top_in[7] mux_right_ipin_2.mux_l2_in_0_/S
+ mux_right_ipin_2.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
Xmem_right_ipin_1.scs8hd_dfxbp_1_0_ prog_clk mux_right_ipin_0.mux_l4_in_0_/S mux_right_ipin_1.mux_l1_in_0_/S
+ mem_right_ipin_1.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_36_59 vgnd vpwr scs8hd_decap_4
XFILLER_7_3 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_7.mux_l4_in_0_ mux_right_ipin_7.mux_l3_in_1_/X mux_right_ipin_7.mux_l3_in_0_/X
+ mux_right_ipin_7.mux_l4_in_0_/S mux_right_ipin_7.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_13_140 vpwr vgnd scs8hd_fill_2
XFILLER_61_6 vpwr vgnd scs8hd_fill_2
XFILLER_42_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_2.mux_l4_in_0__A1 mux_right_ipin_2.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_111 vgnd vpwr scs8hd_decap_8
XFILLER_3_41 vpwr vgnd scs8hd_fill_2
XFILLER_3_96 vgnd vpwr scs8hd_fill_1
XFILLER_47_69 vpwr vgnd scs8hd_fill_2
XFILLER_47_58 vgnd vpwr scs8hd_decap_3
XFILLER_47_47 vgnd vpwr scs8hd_decap_4
XFILLER_47_36 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_14.mux_l1_in_0__A1 chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_10_110 vgnd vpwr scs8hd_decap_12
XFILLER_19_8 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_13.scs8hd_buf_4_0_ mux_right_ipin_13.mux_l4_in_0_/X left_grid_pin_13_
+ vgnd vpwr scs8hd_buf_1
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_ipin_7.mux_l3_in_1_ mux_right_ipin_7.mux_l2_in_3_/X mux_right_ipin_7.mux_l2_in_2_/X
+ mux_right_ipin_7.mux_l3_in_0_/S mux_right_ipin_7.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_27 vgnd vpwr scs8hd_decap_12
XFILLER_59_132 vgnd vpwr scs8hd_decap_12
XANTENNA__63__A chany_bottom_in[10] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_12.mux_l1_in_2__A1 chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_23_71 vpwr vgnd scs8hd_fill_2
XFILLER_23_82 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_9.mux_l4_in_0__S mux_right_ipin_9.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_40 vpwr vgnd scs8hd_fill_2
XFILLER_9_62 vpwr vgnd scs8hd_fill_2
XFILLER_9_73 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_9.mux_l2_in_3__A1 chany_top_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_56_102 vgnd vpwr scs8hd_decap_3
XFILLER_44_48 vpwr vgnd scs8hd_fill_2
XFILLER_44_15 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_8.mux_l1_in_0__A0 chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_60_36 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_ipin_11.scs8hd_dfxbp_1_0__D mux_right_ipin_10.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA__58__A chany_bottom_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_47_113 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_ipin_9.scs8hd_dfxbp_1_2__D mux_right_ipin_9.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_47_135 vgnd vpwr scs8hd_decap_8
XFILLER_18_93 vgnd vpwr scs8hd_decap_4
XFILLER_50_91 vgnd vpwr scs8hd_fill_1
Xmem_right_ipin_11.scs8hd_dfxbp_1_1_ prog_clk mux_right_ipin_11.mux_l1_in_0_/S mux_right_ipin_11.mux_l2_in_3_/S
+ mem_right_ipin_11.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_right_ipin_7.mux_l2_in_2_ chany_bottom_in[12] chany_top_in[4] mux_right_ipin_7.mux_l2_in_0_/S
+ mux_right_ipin_7.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_22_3 vgnd vpwr scs8hd_decap_12
XFILLER_53_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_12.mux_l2_in_1__A1 mux_right_ipin_12.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_39_15 vgnd vpwr scs8hd_decap_12
XFILLER_55_36 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_2.mux_l3_in_0_ mux_right_ipin_2.mux_l2_in_1_/X mux_right_ipin_2.mux_l2_in_0_/X
+ mux_right_ipin_2.mux_l3_in_0_/S mux_right_ipin_2.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_29_135 vgnd vpwr scs8hd_decap_8
XFILLER_61_90 vgnd vpwr scs8hd_fill_1
XFILLER_6_41 vgnd vpwr scs8hd_decap_4
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_25_17 vgnd vpwr scs8hd_decap_3
XPHY_39 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_13.mux_l2_in_2__S mux_right_ipin_13.mux_l2_in_3_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_left_ipin_0.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_left_ipin_0.mux_l1_in_0_/S
+ mux_left_ipin_0.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_10.mux_l2_in_3__A1 chany_top_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_15_50 vgnd vpwr scs8hd_decap_3
XANTENNA__71__A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_40_130 vgnd vpwr scs8hd_decap_12
XFILLER_31_71 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_9.scs8hd_dfxbp_1_1_ prog_clk mux_right_ipin_9.mux_l1_in_2_/S mux_right_ipin_9.mux_l2_in_1_/S
+ mem_right_ipin_9.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_ipin_12.mux_l3_in_0__A1 mux_right_ipin_12.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_2.mux_l2_in_1_ chany_bottom_in[7] chany_top_in[3] mux_right_ipin_2.mux_l2_in_0_/S
+ mux_right_ipin_2.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_6.mux_l2_in_1__A0 chany_bottom_in[11] vgnd vpwr scs8hd_diode_2
XANTENNA__66__A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_9_123 vgnd vpwr scs8hd_decap_12
XFILLER_26_60 vpwr vgnd scs8hd_fill_2
XFILLER_26_93 vpwr vgnd scs8hd_fill_2
XFILLER_3_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_11.scs8hd_dfxbp_1_3__D mux_right_ipin_11.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l2_in_3__A0 _32_/HI vgnd vpwr scs8hd_diode_2
XFILLER_10_122 vgnd vpwr scs8hd_fill_1
XFILLER_12_51 vgnd vpwr scs8hd_decap_12
XFILLER_12_73 vpwr vgnd scs8hd_fill_2
XFILLER_12_84 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_11.mux_l2_in_3_ _25_/HI chany_top_in[16] mux_right_ipin_11.mux_l2_in_3_/S
+ mux_right_ipin_11.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_6.mux_l3_in_0__A0 mux_right_ipin_6.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_52_3 vgnd vpwr scs8hd_decap_8
X_69_ chany_bottom_in[4] chany_top_out[4] vgnd vpwr scs8hd_buf_2
Xmux_right_ipin_7.mux_l3_in_0_ mux_right_ipin_7.mux_l2_in_1_/X mux_right_ipin_7.mux_l2_in_0_/X
+ mux_right_ipin_7.mux_l3_in_0_/S mux_right_ipin_7.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_33_39 vgnd vpwr scs8hd_decap_6
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_59_144 vpwr vgnd scs8hd_fill_2
XFILLER_58_36 vpwr vgnd scs8hd_fill_2
XFILLER_48_80 vpwr vgnd scs8hd_fill_2
XFILLER_0_43 vpwr vgnd scs8hd_fill_2
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XFILLER_9_85 vgnd vpwr scs8hd_decap_3
XFILLER_56_114 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_8.mux_l1_in_0__A1 chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_18_61 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_2.scs8hd_buf_4_0_ mux_right_ipin_2.mux_l4_in_0_/X left_grid_pin_2_
+ vgnd vpwr scs8hd_buf_1
XFILLER_34_82 vpwr vgnd scs8hd_fill_2
XFILLER_34_93 vgnd vpwr scs8hd_decap_4
XFILLER_50_81 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_11.scs8hd_dfxbp_1_0_ prog_clk mux_right_ipin_10.mux_l4_in_0_/S mux_right_ipin_11.mux_l1_in_0_/S
+ mem_right_ipin_11.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_right_ipin_7.mux_l2_in_1_ chany_bottom_in[4] chany_top_in[2] mux_right_ipin_7.mux_l2_in_0_/S
+ mux_right_ipin_7.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_15_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_4.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_8.mux_l1_in_0__S mux_right_ipin_8.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_103 vpwr vgnd scs8hd_fill_2
XFILLER_39_27 vgnd vpwr scs8hd_decap_4
XFILLER_39_38 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_11.mux_l4_in_0_ mux_right_ipin_11.mux_l3_in_1_/X mux_right_ipin_11.mux_l3_in_0_/X
+ mux_right_ipin_11.mux_l4_in_0_/S mux_right_ipin_11.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_ipin_2.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA__69__A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_20_40 vgnd vpwr scs8hd_fill_1
XFILLER_20_84 vpwr vgnd scs8hd_fill_2
XFILLER_29_60 vgnd vpwr scs8hd_fill_1
XFILLER_6_75 vgnd vpwr scs8hd_fill_1
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_13.scs8hd_dfxbp_1_2__D mux_right_ipin_13.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_142 vgnd vpwr scs8hd_decap_4
XFILLER_15_62 vpwr vgnd scs8hd_fill_2
XFILLER_15_73 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_0.mux_l1_in_2__S mux_left_ipin_0.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_9.scs8hd_dfxbp_1_0_ prog_clk mux_right_ipin_8.mux_l4_in_0_/S mux_right_ipin_9.mux_l1_in_2_/S
+ mem_right_ipin_9.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_right_ipin_11.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.mux_l2_in_0__S mux_right_ipin_7.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_11.mux_l3_in_1_ mux_right_ipin_11.mux_l2_in_3_/X mux_right_ipin_11.mux_l2_in_2_/X
+ mux_right_ipin_11.mux_l3_in_0_/S mux_right_ipin_11.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_ipin_2.mux_l2_in_0_ chany_bottom_in[3] mux_right_ipin_2.mux_l1_in_0_/X
+ mux_right_ipin_2.mux_l2_in_0_/S mux_right_ipin_2.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_52_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_6.mux_l2_in_1__A1 chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_52_49 vpwr vgnd scs8hd_fill_2
XFILLER_42_71 vpwr vgnd scs8hd_fill_2
XFILLER_9_135 vgnd vpwr scs8hd_decap_8
XFILLER_42_93 vgnd vpwr scs8hd_decap_4
XFILLER_22_19 vgnd vpwr scs8hd_fill_1
XFILLER_63_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_2.mux_l2_in_2__S mux_right_ipin_2.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l2_in_3__A1 chany_top_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_10_145 vgnd vpwr scs8hd_fill_1
XFILLER_12_63 vgnd vpwr scs8hd_fill_1
Xmem_right_ipin_4.scs8hd_dfxbp_1_3_ prog_clk mux_right_ipin_4.mux_l3_in_1_/S mux_right_ipin_4.mux_l4_in_0_/S
+ mem_right_ipin_4.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_right_ipin_11.mux_l2_in_2_ chany_bottom_in[16] chany_top_in[8] mux_right_ipin_11.mux_l2_in_3_/S
+ mux_right_ipin_11.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_1__D mux_right_ipin_0.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_53_70 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_3.mux_l1_in_0__A0 chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_6.mux_l3_in_0__A1 mux_right_ipin_6.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_45_3 vgnd vpwr scs8hd_decap_3
X_68_ chany_bottom_in[5] chany_top_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_ipin_6.mux_l3_in_0__S mux_right_ipin_6.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_14.mux_l2_in_2__A0 chany_bottom_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_3_108 vpwr vgnd scs8hd_fill_2
XFILLER_58_48 vgnd vpwr scs8hd_decap_8
XFILLER_23_95 vgnd vpwr scs8hd_decap_4
XFILLER_2_130 vpwr vgnd scs8hd_fill_2
XFILLER_0_11 vpwr vgnd scs8hd_fill_2
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l1_in_2__A0 chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_28_29 vpwr vgnd scs8hd_fill_2
XFILLER_44_39 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_ipin_15.mux_l1_in_0__S mux_right_ipin_15.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_ipin_15.scs8hd_dfxbp_1_1__D mux_right_ipin_15.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_84 vgnd vpwr scs8hd_decap_3
XFILLER_50_93 vpwr vgnd scs8hd_fill_2
XFILLER_50_60 vpwr vgnd scs8hd_fill_2
XFILLER_59_91 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_14.mux_l3_in_1__A0 mux_right_ipin_14.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_7.mux_l2_in_0_ chany_bottom_in[2] mux_right_ipin_7.mux_l1_in_0_/X
+ mux_right_ipin_7.mux_l2_in_0_/S mux_right_ipin_7.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_7.mux_l2_in_3__S mux_right_ipin_7.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_5.mux_l4_in_0__S mux_right_ipin_5.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_1.mux_l2_in_1__A0 chany_bottom_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_29_50 vpwr vgnd scs8hd_fill_2
XFILLER_29_72 vpwr vgnd scs8hd_fill_2
XFILLER_35_107 vgnd vpwr scs8hd_decap_3
XFILLER_35_118 vpwr vgnd scs8hd_fill_2
XFILLER_61_70 vgnd vpwr scs8hd_decap_4
XFILLER_45_71 vpwr vgnd scs8hd_fill_2
XFILLER_6_87 vpwr vgnd scs8hd_fill_2
XPHY_19 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_14.mux_l2_in_0__S mux_right_ipin_14.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l1_in_2__A0 chany_top_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_14.mux_l4_in_0__A0 mux_right_ipin_14.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_85 vgnd vpwr scs8hd_decap_12
XFILLER_40_110 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_7.scs8hd_buf_4_0__A mux_right_ipin_7.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_31_51 vgnd vpwr scs8hd_decap_4
XFILLER_31_95 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_2.scs8hd_dfxbp_1_0__D mux_right_ipin_1.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_143 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_11.mux_l3_in_0_ mux_right_ipin_11.mux_l2_in_1_/X mux_right_ipin_11.mux_l2_in_0_/X
+ mux_right_ipin_11.mux_l3_in_0_/S mux_right_ipin_11.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_ipin_9.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_22_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_1.mux_l3_in_0__A0 mux_right_ipin_1.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_ipin_7.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_42_83 vgnd vpwr scs8hd_decap_8
XFILLER_9_103 vpwr vgnd scs8hd_fill_2
XFILLER_13_132 vpwr vgnd scs8hd_fill_2
XFILLER_3_88 vpwr vgnd scs8hd_fill_2
XFILLER_3_77 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.mux_l2_in_1__A0 chany_bottom_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_47_17 vpwr vgnd scs8hd_fill_2
XFILLER_63_49 vpwr vgnd scs8hd_fill_2
XFILLER_63_27 vgnd vpwr scs8hd_decap_12
XFILLER_47_39 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_13.mux_l3_in_0__S mux_right_ipin_13.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_106 vpwr vgnd scs8hd_fill_2
XFILLER_12_97 vgnd vpwr scs8hd_fill_1
Xmem_right_ipin_4.scs8hd_dfxbp_1_2_ prog_clk mux_right_ipin_4.mux_l2_in_3_/S mux_right_ipin_4.mux_l3_in_1_/S
+ mem_right_ipin_4.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_right_ipin_11.mux_l2_in_1_ chany_bottom_in[8] chany_top_in[2] mux_right_ipin_11.mux_l2_in_3_/S
+ mux_right_ipin_11.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_ipin_2.mux_l1_in_0_ chany_top_in[1] chany_bottom_in[1] mux_right_ipin_2.mux_l1_in_0_/S
+ mux_right_ipin_2.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_3.mux_l1_in_0__A1 chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_37_94 vpwr vgnd scs8hd_fill_2
X_67_ chany_bottom_in[6] chany_top_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_ipin_14.mux_l2_in_2__A1 chany_top_in[11] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_14.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_58_27 vgnd vpwr scs8hd_decap_4
XFILLER_48_93 vgnd vpwr scs8hd_decap_6
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XFILLER_0_67 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.mux_l3_in_0__A0 mux_left_ipin_0.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_89 vpwr vgnd scs8hd_fill_2
XFILLER_9_10 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_1.mux_l1_in_2__A1 chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_44_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_14.mux_l2_in_3__S mux_right_ipin_14.mux_l2_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_12.mux_l4_in_0__S mux_right_ipin_12.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_30 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_14.mux_l3_in_1__A1 mux_right_ipin_14.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_ipin_2.scs8hd_dfxbp_1_3__D mux_right_ipin_2.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_53_108 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_8.mux_l2_in_2__A0 chany_bottom_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_20_64 vgnd vpwr scs8hd_decap_4
XFILLER_29_62 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_1.mux_l2_in_1__A1 mux_right_ipin_1.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_95 vpwr vgnd scs8hd_fill_2
XFILLER_61_82 vgnd vpwr scs8hd_decap_8
XFILLER_6_11 vgnd vpwr scs8hd_decap_3
Xmem_right_ipin_14.scs8hd_dfxbp_1_3_ prog_clk mux_right_ipin_14.mux_l3_in_0_/S mux_right_ipin_14.mux_l4_in_0_/S
+ mem_right_ipin_14.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_ipin_4.mux_l1_in_0__S mux_right_ipin_4.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_14.mux_l4_in_0__A1 mux_right_ipin_14.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_11.mux_l2_in_0__A0 chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l1_in_2__A1 chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_17_108 vgnd vpwr scs8hd_decap_12
XFILLER_15_20 vpwr vgnd scs8hd_fill_2
XFILLER_15_42 vpwr vgnd scs8hd_fill_2
XFILLER_15_97 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_7.mux_l1_in_0_ chany_top_in[0] chany_bottom_in[0] mux_right_ipin_7.mux_l1_in_0_/S
+ mux_right_ipin_7.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_ipin_8.mux_l3_in_1__A0 mux_right_ipin_8.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_31_111 vpwr vgnd scs8hd_fill_2
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

