* NGSPICE file created from grid_clb.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_mux2_1 abstract view
.subckt scs8hd_mux2_1 A0 A1 S X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_dfxbp_1 abstract view
.subckt scs8hd_dfxbp_1 CLK D Q QN vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_sdfxbp_1 abstract view
.subckt scs8hd_sdfxbp_1 CLK D Q QN SCD SCE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_1 abstract view
.subckt scs8hd_or2_1 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_clkbuf_16 abstract view
.subckt scs8hd_clkbuf_16 A X vgnd vpwr
.ends

.subckt grid_clb Test_en bottom_width_0_height_0__pin_16_ bottom_width_0_height_0__pin_17_
+ bottom_width_0_height_0__pin_18_ bottom_width_0_height_0__pin_19_ bottom_width_0_height_0__pin_20_
+ bottom_width_0_height_0__pin_21_ bottom_width_0_height_0__pin_22_ bottom_width_0_height_0__pin_23_
+ bottom_width_0_height_0__pin_24_ bottom_width_0_height_0__pin_25_ bottom_width_0_height_0__pin_26_
+ bottom_width_0_height_0__pin_27_ bottom_width_0_height_0__pin_28_ bottom_width_0_height_0__pin_29_
+ bottom_width_0_height_0__pin_30_ bottom_width_0_height_0__pin_31_ bottom_width_0_height_0__pin_42_lower
+ bottom_width_0_height_0__pin_42_upper bottom_width_0_height_0__pin_43_lower bottom_width_0_height_0__pin_43_upper
+ bottom_width_0_height_0__pin_44_lower bottom_width_0_height_0__pin_44_upper bottom_width_0_height_0__pin_45_lower
+ bottom_width_0_height_0__pin_45_upper bottom_width_0_height_0__pin_46_lower bottom_width_0_height_0__pin_46_upper
+ bottom_width_0_height_0__pin_47_lower bottom_width_0_height_0__pin_47_upper bottom_width_0_height_0__pin_48_lower
+ bottom_width_0_height_0__pin_48_upper bottom_width_0_height_0__pin_49_lower bottom_width_0_height_0__pin_49_upper
+ bottom_width_0_height_0__pin_50_ bottom_width_0_height_0__pin_51_ ccff_head ccff_tail
+ clk left_width_0_height_0__pin_52_ prog_clk right_width_0_height_0__pin_0_ right_width_0_height_0__pin_10_
+ right_width_0_height_0__pin_11_ right_width_0_height_0__pin_12_ right_width_0_height_0__pin_13_
+ right_width_0_height_0__pin_14_ right_width_0_height_0__pin_15_ right_width_0_height_0__pin_1_
+ right_width_0_height_0__pin_2_ right_width_0_height_0__pin_34_lower right_width_0_height_0__pin_34_upper
+ right_width_0_height_0__pin_35_lower right_width_0_height_0__pin_35_upper right_width_0_height_0__pin_36_lower
+ right_width_0_height_0__pin_36_upper right_width_0_height_0__pin_37_lower right_width_0_height_0__pin_37_upper
+ right_width_0_height_0__pin_38_lower right_width_0_height_0__pin_38_upper right_width_0_height_0__pin_39_lower
+ right_width_0_height_0__pin_39_upper right_width_0_height_0__pin_3_ right_width_0_height_0__pin_40_lower
+ right_width_0_height_0__pin_40_upper right_width_0_height_0__pin_41_lower right_width_0_height_0__pin_41_upper
+ right_width_0_height_0__pin_4_ right_width_0_height_0__pin_5_ right_width_0_height_0__pin_6_
+ right_width_0_height_0__pin_7_ right_width_0_height_0__pin_8_ right_width_0_height_0__pin_9_
+ top_width_0_height_0__pin_32_ top_width_0_height_0__pin_33_ vpwr vgnd
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_266 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_10_328 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_ _62_/HI
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_406 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_ _36_/HI
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ bottom_width_0_height_0__pin_43_lower vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_239 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_310 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_13_144 vpwr vgnd scs8hd_fill_2
XFILLER_13_188 vgnd vpwr scs8hd_decap_3
XFILLER_3_56 vgnd vpwr scs8hd_decap_3
XFILLER_3_34 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_1__f_clk/X vgnd vpwr scs8hd_diode_2
XFILLER_59_306 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_39 vgnd vpwr scs8hd_decap_12
XFILLER_27_236 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_6_129 vpwr vgnd scs8hd_fill_2
XFILLER_10_125 vgnd vpwr scs8hd_fill_1
XFILLER_12_32 vgnd vpwr scs8hd_decap_12
XFILLER_2_368 vpwr vgnd scs8hd_fill_2
XFILLER_58_361 vpwr vgnd scs8hd_fill_2
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XFILLER_37_51 vgnd vpwr scs8hd_decap_8
XFILLER_18_203 vpwr vgnd scs8hd_fill_2
XFILLER_33_217 vpwr vgnd scs8hd_fill_2
XFILLER_26_280 vpwr vgnd scs8hd_fill_2
XFILLER_18_269 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_294 vpwr vgnd scs8hd_fill_2
XFILLER_5_184 vpwr vgnd scs8hd_fill_2
XFILLER_64_397 vgnd vpwr scs8hd_decap_6
XFILLER_64_342 vgnd vpwr scs8hd_decap_12
X_66_ bottom_width_0_height_0__pin_44_lower bottom_width_0_height_0__pin_44_upper
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
+ clkbuf_1_1__f_clk/X ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en vgnd vpwr scs8hd_sdfxbp_1
XFILLER_59_147 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_386 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
+ right_width_0_height_0__pin_4_ vgnd vpwr scs8hd_diode_2
XFILLER_23_250 vpwr vgnd scs8hd_fill_2
XFILLER_15_206 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_53 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
+ bottom_width_0_height_0__pin_29_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_2_154 vpwr vgnd scs8hd_fill_2
XFILLER_46_386 vgnd vpwr scs8hd_decap_8
XFILLER_46_375 vpwr vgnd scs8hd_fill_2
XFILLER_0_13 vgnd vpwr scs8hd_fill_1
XFILLER_61_367 vgnd vpwr scs8hd_decap_6
XFILLER_9_11 vgnd vpwr scs8hd_decap_3
XFILLER_9_44 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_56_117 vgnd vpwr scs8hd_decap_12
XFILLER_37_331 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
X_49_ _49_/HI _49_/LO vgnd vpwr scs8hd_conb_1
XFILLER_20_286 vgnd vpwr scs8hd_decap_3
XFILLER_20_242 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_43_301 vpwr vgnd scs8hd_fill_2
XPHY_554 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_543 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_532 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_521 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_510 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_242 vpwr vgnd scs8hd_fill_2
XFILLER_7_279 vpwr vgnd scs8hd_fill_2
XFILLER_11_297 vgnd vpwr scs8hd_decap_8
XFILLER_38_117 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_40_337 vgnd vpwr scs8hd_decap_6
XFILLER_25_367 vgnd vpwr scs8hd_decap_4
XFILLER_20_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_238 vpwr vgnd scs8hd_fill_2
XFILLER_29_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_62 vgnd vpwr scs8hd_decap_12
XFILLER_45_51 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_mux2_1
XPHY_395 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_384 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_373 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_362 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_351 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_340 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_293 vpwr vgnd scs8hd_fill_2
XFILLER_6_45 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_13_3 vgnd vpwr scs8hd_decap_12
XFILLER_22_337 vgnd vpwr scs8hd_decap_3
XFILLER_57_245 vgnd vpwr scs8hd_decap_12
XFILLER_25_142 vgnd vpwr scs8hd_decap_12
XFILLER_13_304 vgnd vpwr scs8hd_fill_1
XFILLER_40_178 vgnd vpwr scs8hd_decap_12
XFILLER_15_98 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _35_/HI vgnd vpwr scs8hd_diode_2
XFILLER_31_86 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_0_241 vgnd vpwr scs8hd_decap_4
XFILLER_31_123 vgnd vpwr scs8hd_decap_12
XFILLER_16_186 vpwr vgnd scs8hd_fill_2
XFILLER_16_175 vgnd vpwr scs8hd_decap_8
XFILLER_16_131 vgnd vpwr scs8hd_decap_4
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_396 vgnd vpwr scs8hd_fill_1
XFILLER_54_215 vgnd vpwr scs8hd_decap_12
XFILLER_39_278 vgnd vpwr scs8hd_decap_3
XFILLER_39_245 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_22_101 vpwr vgnd scs8hd_fill_2
XFILLER_10_318 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_281 vgnd vpwr scs8hd_decap_12
XFILLER_26_64 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_101 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XFILLER_5_322 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_8_193 vgnd vpwr scs8hd_decap_4
XFILLER_27_204 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_50_251 vgnd vpwr scs8hd_decap_12
XFILLER_35_292 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_6_108 vgnd vpwr scs8hd_decap_6
XFILLER_12_44 vgnd vpwr scs8hd_decap_12
XFILLER_12_99 vgnd vpwr scs8hd_decap_6
XFILLER_58_384 vgnd vpwr scs8hd_decap_12
XFILLER_37_74 vgnd vpwr scs8hd_decap_12
XFILLER_18_215 vpwr vgnd scs8hd_fill_2
XFILLER_53_62 vgnd vpwr scs8hd_decap_12
XFILLER_53_51 vgnd vpwr scs8hd_decap_8
XFILLER_41_273 vpwr vgnd scs8hd_fill_2
XFILLER_5_163 vgnd vpwr scs8hd_decap_3
XFILLER_49_362 vpwr vgnd scs8hd_fill_2
XFILLER_49_351 vgnd vpwr scs8hd_fill_1
XFILLER_1_380 vgnd vpwr scs8hd_decap_12
XFILLER_64_354 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_229 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
X_65_ bottom_width_0_height_0__pin_43_lower bottom_width_0_height_0__pin_43_upper
+ vgnd vpwr scs8hd_buf_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XFILLER_32_284 vgnd vpwr scs8hd_decap_12
XFILLER_32_251 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_159 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_55_398 vpwr vgnd scs8hd_fill_2
XFILLER_23_273 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_23_87 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
+ bottom_width_0_height_0__pin_28_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_2_100 vpwr vgnd scs8hd_fill_2
XFILLER_2_144 vpwr vgnd scs8hd_fill_2
XFILLER_64_94 vgnd vpwr scs8hd_decap_12
XFILLER_61_335 vgnd vpwr scs8hd_decap_12
XFILLER_46_398 vgnd vpwr scs8hd_decap_8
XFILLER_46_354 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_14_273 vpwr vgnd scs8hd_fill_2
XFILLER_43_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_56_129 vgnd vpwr scs8hd_decap_12
X_48_ _48_/HI _48_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_298 vpwr vgnd scs8hd_fill_2
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XPHY_500 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_55_184 vgnd vpwr scs8hd_decap_12
XFILLER_43_346 vgnd vpwr scs8hd_fill_1
XFILLER_28_398 vgnd vpwr scs8hd_decap_8
XFILLER_28_354 vpwr vgnd scs8hd_fill_2
XFILLER_28_332 vgnd vpwr scs8hd_fill_1
XFILLER_18_32 vgnd vpwr scs8hd_decap_12
XPHY_555 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_544 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_533 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_522 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_511 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_203 vpwr vgnd scs8hd_fill_2
XFILLER_7_236 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_258 vpwr vgnd scs8hd_fill_2
XFILLER_38_129 vgnd vpwr scs8hd_decap_12
XFILLER_19_332 vgnd vpwr scs8hd_decap_4
XFILLER_61_110 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_184 vgnd vpwr scs8hd_decap_12
XFILLER_25_346 vpwr vgnd scs8hd_fill_2
XFILLER_25_335 vpwr vgnd scs8hd_fill_2
XFILLER_25_324 vpwr vgnd scs8hd_fill_2
XFILLER_25_302 vgnd vpwr scs8hd_decap_3
XFILLER_52_154 vgnd vpwr scs8hd_decap_12
XFILLER_40_349 vpwr vgnd scs8hd_fill_2
XFILLER_40_316 vpwr vgnd scs8hd_fill_2
XFILLER_20_99 vgnd vpwr scs8hd_decap_4
XFILLER_0_401 vpwr vgnd scs8hd_fill_2
XFILLER_4_206 vpwr vgnd scs8hd_fill_2
XFILLER_29_86 vgnd vpwr scs8hd_decap_12
XFILLER_45_74 vgnd vpwr scs8hd_decap_12
XFILLER_43_110 vgnd vpwr scs8hd_decap_12
XPHY_352 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_338 vgnd vpwr scs8hd_decap_3
XPHY_341 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_330 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_28_195 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_16_335 vgnd vpwr scs8hd_fill_1
XFILLER_16_302 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XFILLER_61_62 vgnd vpwr scs8hd_decap_12
XFILLER_61_51 vgnd vpwr scs8hd_decap_8
XPHY_396 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_385 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_374 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_363 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_68 vpwr vgnd scs8hd_fill_2
XFILLER_19_184 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_57_257 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_154 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_88 vgnd vpwr scs8hd_decap_8
XFILLER_9_309 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_98 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
+ bottom_width_0_height_0__pin_18_ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_202 vgnd vpwr scs8hd_decap_12
XFILLER_0_275 vpwr vgnd scs8hd_fill_2
XFILLER_31_135 vgnd vpwr scs8hd_decap_12
XFILLER_16_154 vpwr vgnd scs8hd_fill_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_227 vgnd vpwr scs8hd_decap_12
XFILLER_22_113 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_190 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_9 vpwr vgnd scs8hd_fill_2
XFILLER_45_249 vgnd vpwr scs8hd_fill_1
XFILLER_45_238 vgnd vpwr scs8hd_fill_1
XFILLER_45_216 vgnd vpwr scs8hd_decap_3
XFILLER_38_290 vgnd vpwr scs8hd_fill_1
XFILLER_26_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_293 vgnd vpwr scs8hd_fill_1
XFILLER_9_117 vgnd vpwr scs8hd_decap_3
XFILLER_5_345 vgnd vpwr scs8hd_decap_4
XFILLER_5_367 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_208 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_8_172 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_50_263 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
+ right_width_0_height_0__pin_1_ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_10_138 vpwr vgnd scs8hd_fill_2
XFILLER_12_56 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_396 vgnd vpwr scs8hd_fill_1
XFILLER_37_86 vgnd vpwr scs8hd_decap_12
XFILLER_33_208 vgnd vpwr scs8hd_decap_6
XFILLER_26_260 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_74 vgnd vpwr scs8hd_decap_12
XFILLER_41_230 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_5_175 vpwr vgnd scs8hd_fill_2
XFILLER_64_311 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
X_64_ bottom_width_0_height_0__pin_42_lower bottom_width_0_height_0__pin_42_upper
+ vgnd vpwr scs8hd_buf_2
XFILLER_1_392 vgnd vpwr scs8hd_decap_12
XFILLER_64_366 vgnd vpwr scs8hd_decap_6
XFILLER_32_274 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_333 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _61_/HI vgnd vpwr scs8hd_diode_2
XFILLER_23_285 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
+ top_width_0_height_0__pin_33_ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_2_123 vpwr vgnd scs8hd_fill_2
XFILLER_46_311 vpwr vgnd scs8hd_fill_2
XFILLER_61_347 vgnd vpwr scs8hd_decap_12
XFILLER_0_59 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XFILLER_49_171 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
X_47_ _47_/HI _47_/LO vgnd vpwr scs8hd_conb_1
XFILLER_52_347 vpwr vgnd scs8hd_fill_2
XFILLER_20_266 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XPHY_534 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_523 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_512 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_501 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_55_196 vgnd vpwr scs8hd_decap_12
XFILLER_43_358 vpwr vgnd scs8hd_fill_2
XFILLER_43_314 vpwr vgnd scs8hd_fill_2
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_556 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_545 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_215 vpwr vgnd scs8hd_fill_2
XFILLER_11_222 vgnd vpwr scs8hd_decap_12
XFILLER_59_62 vgnd vpwr scs8hd_decap_12
XFILLER_59_51 vgnd vpwr scs8hd_decap_8
XFILLER_46_141 vgnd vpwr scs8hd_decap_12
XFILLER_34_369 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_57_406 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_166 vgnd vpwr scs8hd_decap_12
XFILLER_37_196 vgnd vpwr scs8hd_decap_8
XFILLER_25_358 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
+ clkbuf_1_0__f_clk/X ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 Test_en
+ vgnd vpwr scs8hd_sdfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_33_380 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_89 vgnd vpwr scs8hd_decap_3
XFILLER_48_406 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_29_98 vgnd vpwr scs8hd_decap_12
XFILLER_28_152 vgnd vpwr scs8hd_fill_1
XFILLER_28_130 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_45_86 vgnd vpwr scs8hd_decap_12
XPHY_386 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_375 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_364 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_353 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_306 vgnd vpwr scs8hd_decap_3
XPHY_342 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_331 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_320 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_74 vgnd vpwr scs8hd_decap_12
XPHY_397 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_406 vgnd vpwr scs8hd_fill_1
XFILLER_3_240 vpwr vgnd scs8hd_fill_2
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
XFILLER_30_383 vgnd vpwr scs8hd_decap_12
XFILLER_57_269 vgnd vpwr scs8hd_decap_12
XFILLER_25_166 vgnd vpwr scs8hd_decap_12
XFILLER_13_306 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
+ bottom_width_0_height_0__pin_17_ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_100 vpwr vgnd scs8hd_fill_2
XFILLER_31_147 vgnd vpwr scs8hd_decap_12
XFILLER_16_199 vpwr vgnd scs8hd_fill_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_354 vgnd vpwr scs8hd_decap_8
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_372 vpwr vgnd scs8hd_fill_2
XFILLER_12_383 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_398 vgnd vpwr scs8hd_decap_8
XFILLER_39_214 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_ _48_/HI
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ bottom_width_0_height_0__pin_49_lower vgnd vpwr scs8hd_mux2_1
XFILLER_54_239 vgnd vpwr scs8hd_decap_12
XFILLER_22_158 vgnd vpwr scs8hd_decap_6
XFILLER_22_125 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_90 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
+ bottom_width_0_height_0__pin_29_ vgnd vpwr scs8hd_diode_2
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
XFILLER_13_136 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_5_302 vgnd vpwr scs8hd_decap_3
XFILLER_5_379 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
X_80_ right_width_0_height_0__pin_41_lower right_width_0_height_0__pin_41_upper vgnd
+ vpwr scs8hd_buf_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
+ clkbuf_1_1__f_clk/X ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en vgnd vpwr scs8hd_sdfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_26 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_10_128 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_305 vgnd vpwr scs8hd_fill_1
XFILLER_5_7 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_98 vgnd vpwr scs8hd_decap_12
XFILLER_26_272 vgnd vpwr scs8hd_decap_3
XFILLER_26_250 vgnd vpwr scs8hd_fill_1
XFILLER_53_86 vgnd vpwr scs8hd_decap_12
XFILLER_41_286 vpwr vgnd scs8hd_fill_2
XFILLER_41_253 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_64_323 vgnd vpwr scs8hd_decap_12
XFILLER_49_386 vgnd vpwr scs8hd_decap_12
XFILLER_49_331 vgnd vpwr scs8hd_decap_6
X_63_ _63_/HI _63_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_231 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_301 vpwr vgnd scs8hd_fill_2
XFILLER_55_345 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_231 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_23_297 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XFILLER_11_404 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_0_27 vpwr vgnd scs8hd_fill_2
XFILLER_64_63 vgnd vpwr scs8hd_decap_12
XFILLER_61_359 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_29_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XFILLER_1_190 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_359 vgnd vpwr scs8hd_fill_1
XFILLER_52_337 vgnd vpwr scs8hd_fill_1
XFILLER_37_367 vgnd vpwr scs8hd_decap_3
XFILLER_37_334 vpwr vgnd scs8hd_fill_2
XFILLER_37_301 vpwr vgnd scs8hd_fill_2
X_46_ _46_/HI _46_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XFILLER_20_234 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _47_/HI ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_mux2_1
XFILLER_28_323 vgnd vpwr scs8hd_fill_1
XFILLER_18_56 vgnd vpwr scs8hd_decap_4
XPHY_557 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_546 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_535 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_524 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_513 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_502 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_337 vgnd vpwr scs8hd_decap_3
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_32 vgnd vpwr scs8hd_decap_12
XFILLER_11_234 vgnd vpwr scs8hd_decap_8
XFILLER_11_245 vgnd vpwr scs8hd_decap_4
XFILLER_59_74 vgnd vpwr scs8hd_decap_12
XFILLER_61_123 vgnd vpwr scs8hd_decap_12
XFILLER_34_337 vpwr vgnd scs8hd_fill_2
XFILLER_34_326 vgnd vpwr scs8hd_decap_8
XFILLER_34_315 vpwr vgnd scs8hd_fill_2
XFILLER_19_367 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_52_178 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _56_/HI vgnd vpwr scs8hd_diode_2
XFILLER_20_46 vgnd vpwr scs8hd_decap_4
XFILLER_43_123 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_61_86 vgnd vpwr scs8hd_decap_12
XFILLER_45_98 vgnd vpwr scs8hd_decap_12
XPHY_398 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_387 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_376 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_365 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_354 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_343 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_332 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_321 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_310 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
+ bottom_width_0_height_0__pin_23_ vgnd vpwr scs8hd_diode_2
XFILLER_6_26 vpwr vgnd scs8hd_fill_2
XFILLER_19_131 vgnd vpwr scs8hd_decap_6
XFILLER_19_120 vpwr vgnd scs8hd_fill_2
XFILLER_3_285 vgnd vpwr scs8hd_fill_1
XFILLER_10_90 vpwr vgnd scs8hd_fill_2
XFILLER_34_178 vgnd vpwr scs8hd_decap_12
XFILLER_19_175 vpwr vgnd scs8hd_fill_2
XFILLER_30_395 vpwr vgnd scs8hd_fill_2
XFILLER_30_362 vgnd vpwr scs8hd_decap_4
XFILLER_15_392 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_178 vgnd vpwr scs8hd_decap_4
XFILLER_21_362 vgnd vpwr scs8hd_fill_1
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
+ bottom_width_0_height_0__pin_16_ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_48_215 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_31_159 vgnd vpwr scs8hd_decap_12
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_388 vgnd vpwr scs8hd_decap_8
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_395 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_281 vgnd vpwr scs8hd_decap_8
XFILLER_39_237 vpwr vgnd scs8hd_fill_2
XFILLER_11_3 vgnd vpwr scs8hd_decap_12
XFILLER_62_251 vgnd vpwr scs8hd_decap_12
XFILLER_22_137 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_56 vgnd vpwr scs8hd_decap_8
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_148 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _63_/HI ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_mux2_1
XFILLER_3_38 vpwr vgnd scs8hd_fill_2
XFILLER_5_314 vpwr vgnd scs8hd_fill_2
XFILLER_44_295 vgnd vpwr scs8hd_decap_3
XFILLER_44_240 vgnd vpwr scs8hd_decap_6
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_59_3 vgnd vpwr scs8hd_decap_12
XFILLER_8_152 vgnd vpwr scs8hd_fill_1
XFILLER_12_170 vpwr vgnd scs8hd_fill_2
XFILLER_12_181 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_240 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_50_276 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_328 vpwr vgnd scs8hd_fill_2
XFILLER_58_398 vgnd vpwr scs8hd_decap_8
XFILLER_18_207 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_284 vpwr vgnd scs8hd_fill_2
XFILLER_53_98 vgnd vpwr scs8hd_decap_12
XFILLER_41_298 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_5_111 vgnd vpwr scs8hd_decap_4
XFILLER_5_155 vpwr vgnd scs8hd_fill_2
XFILLER_49_310 vpwr vgnd scs8hd_fill_2
XFILLER_1_350 vpwr vgnd scs8hd_fill_2
XFILLER_64_335 vgnd vpwr scs8hd_decap_6
XFILLER_49_398 vgnd vpwr scs8hd_decap_8
X_62_ _62_/HI _62_/LO vgnd vpwr scs8hd_conb_1
XFILLER_17_240 vpwr vgnd scs8hd_fill_2
XFILLER_32_298 vgnd vpwr scs8hd_decap_8
XFILLER_32_276 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_0__f_clk/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
XFILLER_48_32 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
+ right_width_0_height_0__pin_6_ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_2_169 vpwr vgnd scs8hd_fill_2
XFILLER_2_158 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ccff_tail vgnd vpwr scs8hd_diode_2
XFILLER_46_379 vgnd vpwr scs8hd_decap_4
XFILLER_46_346 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_ _57_/HI
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ right_width_0_height_0__pin_36_lower vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_75 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_48 vgnd vpwr scs8hd_fill_1
XFILLER_14_265 vgnd vpwr scs8hd_decap_8
XFILLER_14_276 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_49_184 vgnd vpwr scs8hd_decap_12
XFILLER_64_187 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_357 vgnd vpwr scs8hd_decap_3
X_45_ _45_/HI _45_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_371 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_55_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_28_335 vgnd vpwr scs8hd_fill_1
XFILLER_28_313 vpwr vgnd scs8hd_fill_2
XFILLER_18_79 vgnd vpwr scs8hd_decap_12
XPHY_558 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_547 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_536 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_525 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_514 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_503 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
XFILLER_50_44 vgnd vpwr scs8hd_decap_12
XFILLER_59_86 vgnd vpwr scs8hd_decap_12
XFILLER_19_302 vgnd vpwr scs8hd_decap_3
XFILLER_61_135 vgnd vpwr scs8hd_decap_12
XFILLER_46_154 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_19_357 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _55_/HI vgnd vpwr scs8hd_diode_2
XFILLER_6_272 vgnd vpwr scs8hd_decap_3
XFILLER_37_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_82 vpwr vgnd scs8hd_fill_2
XFILLER_60_190 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_69 vpwr vgnd scs8hd_fill_2
XFILLER_0_404 vgnd vpwr scs8hd_decap_3
XFILLER_43_135 vgnd vpwr scs8hd_decap_12
XFILLER_28_154 vgnd vpwr scs8hd_decap_12
XPHY_300 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_61_98 vgnd vpwr scs8hd_decap_12
XPHY_399 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_388 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_377 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_366 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_355 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_344 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_333 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_322 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_311 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_264 vpwr vgnd scs8hd_fill_2
XFILLER_6_49 vgnd vpwr scs8hd_decap_4
XFILLER_3_297 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_190 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_clkbuf_0_clk_A clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_25_113 vpwr vgnd scs8hd_fill_2
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_21_330 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
+ bottom_width_0_height_0__pin_26_ vgnd vpwr scs8hd_diode_2
XFILLER_63_208 vgnd vpwr scs8hd_decap_12
XFILLER_56_32 vgnd vpwr scs8hd_decap_12
XFILLER_48_227 vgnd vpwr scs8hd_decap_12
XFILLER_0_245 vgnd vpwr scs8hd_fill_1
XFILLER_24_190 vgnd vpwr scs8hd_decap_6
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_334 vpwr vgnd scs8hd_fill_2
XFILLER_8_367 vpwr vgnd scs8hd_fill_2
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_39_249 vpwr vgnd scs8hd_fill_2
XFILLER_39_227 vpwr vgnd scs8hd_fill_2
XFILLER_62_263 vgnd vpwr scs8hd_decap_12
XFILLER_22_149 vgnd vpwr scs8hd_decap_4
XFILLER_22_105 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_208 vgnd vpwr scs8hd_decap_8
XFILLER_53_296 vpwr vgnd scs8hd_fill_2
XFILLER_38_282 vgnd vpwr scs8hd_decap_6
XFILLER_26_68 vgnd vpwr scs8hd_decap_3
XFILLER_42_56 vgnd vpwr scs8hd_decap_12
XFILLER_5_326 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_8_120 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_35_296 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_12_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_219 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_5_123 vpwr vgnd scs8hd_fill_2
X_61_ _61_/HI _61_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_362 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_255 vgnd vpwr scs8hd_decap_12
XFILLER_20_406 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_55_358 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_71 vpwr vgnd scs8hd_fill_2
XFILLER_63_391 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_141 vgnd vpwr scs8hd_decap_12
XFILLER_48_44 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
+ right_width_0_height_0__pin_5_ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_2_148 vpwr vgnd scs8hd_fill_2
XFILLER_64_87 vgnd vpwr scs8hd_decap_6
XFILLER_64_32 vgnd vpwr scs8hd_decap_12
XFILLER_61_306 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_14_200 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
+ clkbuf_1_1__f_clk/X ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 Test_en
+ vgnd vpwr scs8hd_sdfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_16 vpwr vgnd scs8hd_fill_2
XFILLER_14_288 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_13_80 vpwr vgnd scs8hd_fill_2
XFILLER_49_196 vgnd vpwr scs8hd_decap_12
XFILLER_37_325 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_diode_2
X_44_ _44_/HI _44_/LO vgnd vpwr scs8hd_conb_1
XFILLER_64_199 vgnd vpwr scs8hd_decap_12
XFILLER_60_383 vgnd vpwr scs8hd_decap_12
XFILLER_52_328 vgnd vpwr scs8hd_decap_3
XFILLER_52_306 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_270 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_28_358 vpwr vgnd scs8hd_fill_2
XPHY_559 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_548 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_537 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_526 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_515 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_504 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XFILLER_7_207 vgnd vpwr scs8hd_decap_8
XFILLER_11_214 vpwr vgnd scs8hd_fill_2
XFILLER_50_56 vgnd vpwr scs8hd_decap_12
XFILLER_1_3 vpwr vgnd scs8hd_fill_2
XFILLER_59_98 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _45_/HI vgnd vpwr scs8hd_diode_2
XFILLER_61_147 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_46_166 vgnd vpwr scs8hd_decap_12
XFILLER_27_380 vgnd vpwr scs8hd_decap_4
XFILLER_42_394 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_251 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XFILLER_25_339 vgnd vpwr scs8hd_decap_3
XFILLER_25_328 vgnd vpwr scs8hd_decap_4
XFILLER_25_306 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_380 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_20_15 vgnd vpwr scs8hd_decap_12
XFILLER_43_147 vgnd vpwr scs8hd_decap_12
XPHY_334 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_323 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_28_166 vgnd vpwr scs8hd_decap_12
XPHY_312 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_301 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_350 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_389 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_378 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_367 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_356 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_345 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_24_383 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_320 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_117 vgnd vpwr scs8hd_decap_12
XFILLER_15_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
+ clkbuf_1_1__f_clk/X ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en vgnd vpwr scs8hd_sdfxbp_1
XFILLER_0_213 vpwr vgnd scs8hd_fill_2
XFILLER_56_44 vgnd vpwr scs8hd_decap_12
XFILLER_48_239 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_120 vgnd vpwr scs8hd_decap_3
XFILLER_56_294 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_80 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_206 vpwr vgnd scs8hd_fill_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
+ bottom_width_0_height_0__pin_20_ vgnd vpwr scs8hd_diode_2
XFILLER_7_71 vpwr vgnd scs8hd_fill_2
XFILLER_53_220 vgnd vpwr scs8hd_decap_12
XFILLER_41_404 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_68 vgnd vpwr scs8hd_decap_12
XFILLER_21_194 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_16_91 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ bottom_width_0_height_0__pin_31_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/A
+ vgnd vpwr scs8hd_or2_1
XFILLER_8_176 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_209 vpwr vgnd scs8hd_fill_2
XFILLER_23_404 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_27 vgnd vpwr scs8hd_decap_4
XFILLER_58_301 vgnd vpwr scs8hd_decap_8
XFILLER_2_308 vgnd vpwr scs8hd_fill_1
XFILLER_58_356 vgnd vpwr scs8hd_decap_3
XFILLER_26_264 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_5_179 vpwr vgnd scs8hd_fill_2
XFILLER_64_304 vgnd vpwr scs8hd_decap_6
XFILLER_49_323 vpwr vgnd scs8hd_fill_2
XFILLER_49_301 vpwr vgnd scs8hd_fill_2
X_60_ _60_/HI _60_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XFILLER_17_297 vpwr vgnd scs8hd_fill_2
XFILLER_17_286 vpwr vgnd scs8hd_fill_2
XFILLER_64_3 vgnd vpwr scs8hd_decap_12
XFILLER_32_267 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_289 vpwr vgnd scs8hd_fill_2
XFILLER_23_278 vgnd vpwr scs8hd_decap_3
XFILLER_23_245 vgnd vpwr scs8hd_decap_3
XFILLER_23_234 vpwr vgnd scs8hd_fill_2
XFILLER_23_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
+ right_width_0_height_0__pin_4_ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_2_127 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_48_56 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_44 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_54_381 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_39 vgnd vpwr scs8hd_decap_3
XFILLER_13_92 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_64_156 vgnd vpwr scs8hd_decap_12
X_43_ _43_/HI _43_/LO vgnd vpwr scs8hd_conb_1
XFILLER_60_395 vpwr vgnd scs8hd_fill_2
XFILLER_60_351 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XFILLER_18_15 vgnd vpwr scs8hd_decap_12
XPHY_516 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_505 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_55_123 vgnd vpwr scs8hd_decap_12
XFILLER_28_337 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XPHY_549 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_538 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_527 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_219 vpwr vgnd scs8hd_fill_2
XFILLER_50_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_403 vgnd vpwr scs8hd_decap_4
XFILLER_19_315 vpwr vgnd scs8hd_fill_2
XFILLER_61_159 vgnd vpwr scs8hd_decap_12
XFILLER_46_178 vgnd vpwr scs8hd_decap_12
XFILLER_27_392 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_80 vpwr vgnd scs8hd_fill_2
XFILLER_6_285 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_123 vgnd vpwr scs8hd_decap_12
XFILLER_1_62 vgnd vpwr scs8hd_fill_1
XFILLER_33_384 vpwr vgnd scs8hd_fill_2
XFILLER_33_362 vpwr vgnd scs8hd_fill_2
XFILLER_33_351 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/A
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
XFILLER_28_134 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_43_159 vgnd vpwr scs8hd_decap_12
XPHY_368 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_357 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_346 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_335 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_324 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_28_178 vgnd vpwr scs8hd_decap_12
XPHY_313 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_302 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_395 vpwr vgnd scs8hd_fill_2
XFILLER_24_362 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_379 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_288 vgnd vpwr scs8hd_fill_1
XFILLER_10_82 vgnd vpwr scs8hd_decap_8
XFILLER_10_93 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_281 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_19_112 vpwr vgnd scs8hd_fill_2
XFILLER_30_398 vgnd vpwr scs8hd_decap_8
XFILLER_15_351 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_53_402 vgnd vpwr scs8hd_decap_4
XFILLER_40_129 vgnd vpwr scs8hd_decap_12
XFILLER_15_27 vgnd vpwr scs8hd_decap_12
XFILLER_31_59 vpwr vgnd scs8hd_fill_2
XFILLER_31_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_365 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_56_251 vgnd vpwr scs8hd_decap_12
XFILLER_56_56 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_16_104 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
XPHY_121 vgnd vpwr scs8hd_decap_3
XPHY_110 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _40_/HI vgnd vpwr scs8hd_diode_2
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_314 vgnd vpwr scs8hd_decap_12
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_12_398 vgnd vpwr scs8hd_decap_8
XFILLER_62_276 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_15_192 vpwr vgnd scs8hd_fill_2
XFILLER_7_83 vgnd vpwr scs8hd_decap_4
XFILLER_7_94 vpwr vgnd scs8hd_fill_2
XFILLER_7_380 vgnd vpwr scs8hd_decap_12
XFILLER_53_232 vgnd vpwr scs8hd_decap_12
XFILLER_38_295 vpwr vgnd scs8hd_fill_2
XFILLER_38_251 vpwr vgnd scs8hd_fill_2
XFILLER_26_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_184 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_295 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_32_80 vgnd vpwr scs8hd_decap_12
XFILLER_8_133 vpwr vgnd scs8hd_fill_2
XFILLER_8_144 vgnd vpwr scs8hd_decap_8
XFILLER_12_195 vpwr vgnd scs8hd_fill_2
XFILLER_4_350 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_ _38_/HI
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XFILLER_50_202 vgnd vpwr scs8hd_decap_12
XFILLER_35_265 vpwr vgnd scs8hd_fill_2
XFILLER_35_254 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_243 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_257 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_0__f_clk/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_202 vgnd vpwr scs8hd_decap_12
XFILLER_57_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_84 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_0__f_clk/X vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_ _37_/HI
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ bottom_width_0_height_0__pin_42_lower vgnd vpwr scs8hd_mux2_1
XFILLER_23_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_154 vgnd vpwr scs8hd_decap_12
XFILLER_48_68 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_64_56 vgnd vpwr scs8hd_decap_6
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_54_393 vgnd vpwr scs8hd_decap_4
XFILLER_14_235 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_49_110 vgnd vpwr scs8hd_decap_12
XFILLER_1_194 vpwr vgnd scs8hd_fill_2
XFILLER_64_168 vgnd vpwr scs8hd_decap_12
X_42_ _42_/HI _42_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_27 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XPHY_539 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_528 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_517 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_506 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_55_135 vgnd vpwr scs8hd_decap_12
XFILLER_51_341 vpwr vgnd scs8hd_fill_2
XFILLER_51_330 vgnd vpwr scs8hd_fill_1
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_34_319 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_190 vgnd vpwr scs8hd_decap_12
XFILLER_42_352 vpwr vgnd scs8hd_fill_2
XFILLER_42_330 vgnd vpwr scs8hd_decap_4
XFILLER_40_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_30 vpwr vgnd scs8hd_fill_2
XFILLER_52_105 vgnd vpwr scs8hd_decap_12
XFILLER_37_135 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_29_15 vgnd vpwr scs8hd_decap_12
XFILLER_29_59 vpwr vgnd scs8hd_fill_2
XFILLER_28_146 vgnd vpwr scs8hd_decap_6
XFILLER_16_319 vgnd vpwr scs8hd_decap_12
XFILLER_16_308 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_51_171 vgnd vpwr scs8hd_decap_12
XFILLER_36_190 vgnd vpwr scs8hd_decap_12
XPHY_369 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_358 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_347 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_336 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_325 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_314 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_303 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_61 vpwr vgnd scs8hd_fill_2
XFILLER_59_293 vgnd vpwr scs8hd_decap_8
XFILLER_34_105 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_19_179 vpwr vgnd scs8hd_fill_2
XFILLER_19_81 vpwr vgnd scs8hd_fill_2
XFILLER_15_363 vgnd vpwr scs8hd_decap_3
XFILLER_30_366 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
+ bottom_width_0_height_0__pin_17_ vgnd vpwr scs8hd_diode_2
XFILLER_57_208 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_33_171 vgnd vpwr scs8hd_decap_12
XFILLER_21_322 vgnd vpwr scs8hd_decap_8
XFILLER_15_39 vgnd vpwr scs8hd_decap_12
XFILLER_31_27 vgnd vpwr scs8hd_decap_12
XFILLER_0_237 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_56_263 vgnd vpwr scs8hd_decap_12
XFILLER_56_68 vgnd vpwr scs8hd_decap_12
XPHY_100 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_16_127 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XPHY_122 vgnd vpwr scs8hd_decap_3
XPHY_111 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_326 vgnd vpwr scs8hd_decap_8
XFILLER_8_337 vgnd vpwr scs8hd_decap_6
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_366 vgnd vpwr scs8hd_decap_4
XFILLER_21_93 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_62_288 vgnd vpwr scs8hd_decap_12
XFILLER_50_406 vgnd vpwr scs8hd_fill_1
Xclkbuf_0_clk clk clkbuf_0_clk/X vgnd vpwr scs8hd_clkbuf_16
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_30_141 vgnd vpwr scs8hd_decap_12
XFILLER_7_40 vpwr vgnd scs8hd_fill_2
XFILLER_7_392 vgnd vpwr scs8hd_decap_12
XFILLER_38_263 vgnd vpwr scs8hd_decap_12
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_32_406 vgnd vpwr scs8hd_fill_1
XFILLER_16_93 vgnd vpwr scs8hd_decap_3
XFILLER_8_189 vpwr vgnd scs8hd_fill_2
XFILLER_12_174 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
+ clkbuf_1_1__f_clk/X ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 Test_en
+ vgnd vpwr scs8hd_sdfxbp_1
XFILLER_37_15 vgnd vpwr scs8hd_decap_12
XFILLER_37_59 vpwr vgnd scs8hd_fill_2
XFILLER_26_288 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_14_406 vgnd vpwr scs8hd_fill_1
XFILLER_41_269 vpwr vgnd scs8hd_fill_2
XFILLER_5_115 vgnd vpwr scs8hd_fill_1
XFILLER_1_376 vpwr vgnd scs8hd_fill_2
XFILLER_1_354 vpwr vgnd scs8hd_fill_2
XFILLER_5_159 vpwr vgnd scs8hd_fill_2
XFILLER_49_358 vpwr vgnd scs8hd_fill_2
XFILLER_27_70 vpwr vgnd scs8hd_fill_2
XFILLER_17_222 vgnd vpwr scs8hd_decap_12
XFILLER_17_200 vgnd vpwr scs8hd_decap_3
XFILLER_40_280 vgnd vpwr scs8hd_decap_4
XFILLER_55_306 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_39 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_58_166 vgnd vpwr scs8hd_decap_12
XFILLER_39_380 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XFILLER_14_247 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_22_291 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
X_41_ _41_/HI _41_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_184 vpwr vgnd scs8hd_fill_2
XFILLER_64_125 vgnd vpwr scs8hd_decap_12
XFILLER_38_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_60_375 vgnd vpwr scs8hd_decap_4
XFILLER_20_206 vgnd vpwr scs8hd_decap_8
XFILLER_9_240 vpwr vgnd scs8hd_fill_2
XFILLER_55_147 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
+ right_width_0_height_0__pin_11_ vgnd vpwr scs8hd_diode_2
XFILLER_28_328 vgnd vpwr scs8hd_decap_4
XFILLER_28_317 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_buf_2
XPHY_529 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_518 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_507 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_386 vgnd vpwr scs8hd_decap_12
XFILLER_51_364 vpwr vgnd scs8hd_fill_2
XFILLER_36_350 vgnd vpwr scs8hd_fill_1
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
XFILLER_50_15 vgnd vpwr scs8hd_decap_12
XFILLER_19_328 vpwr vgnd scs8hd_fill_2
XANTENNA__64__A bottom_width_0_height_0__pin_42_lower vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_386 vgnd vpwr scs8hd_decap_8
XFILLER_42_342 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ bottom_width_0_height_0__pin_19_ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/A
+ vgnd vpwr scs8hd_or2_1
XFILLER_10_261 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_10_294 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_147 vgnd vpwr scs8hd_decap_12
XFILLER_1_53 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
+ clkbuf_1_0__f_clk/X ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en vgnd vpwr scs8hd_sdfxbp_1
XFILLER_52_117 vgnd vpwr scs8hd_decap_12
XFILLER_33_320 vgnd vpwr scs8hd_decap_8
XFILLER_18_361 vgnd vpwr scs8hd_decap_8
XFILLER_1_86 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_27 vgnd vpwr scs8hd_decap_12
XFILLER_45_59 vpwr vgnd scs8hd_fill_2
XFILLER_45_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_359 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_348 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_337 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_326 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_315 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_304 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_224 vpwr vgnd scs8hd_fill_2
XFILLER_3_268 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_117 vgnd vpwr scs8hd_decap_12
XFILLER_27_180 vgnd vpwr scs8hd_decap_3
XFILLER_19_93 vpwr vgnd scs8hd_fill_2
XFILLER_15_331 vgnd vpwr scs8hd_decap_6
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_30_334 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
XFILLER_25_117 vgnd vpwr scs8hd_decap_3
XFILLER_21_367 vgnd vpwr scs8hd_decap_3
XFILLER_18_191 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_0_249 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XPHY_123 vgnd vpwr scs8hd_decap_3
XPHY_112 vgnd vpwr scs8hd_decap_3
XPHY_101 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_16_139 vgnd vpwr scs8hd_decap_12
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_312 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_72 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_297 vpwr vgnd scs8hd_fill_2
XFILLER_47_220 vgnd vpwr scs8hd_decap_12
XFILLER_46_80 vgnd vpwr scs8hd_decap_12
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_53_245 vgnd vpwr scs8hd_decap_12
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_21_175 vpwr vgnd scs8hd_fill_2
XFILLER_21_153 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_44_267 vgnd vpwr scs8hd_decap_8
XANTENNA__72__A bottom_width_0_height_0__pin_50_ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_32_93 vgnd vpwr scs8hd_decap_12
XFILLER_8_157 vgnd vpwr scs8hd_decap_12
XFILLER_4_396 vgnd vpwr scs8hd_fill_1
XFILLER_50_215 vgnd vpwr scs8hd_decap_12
XFILLER_35_212 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ bottom_width_0_height_0__pin_50_ vgnd vpwr scs8hd_diode_2
XFILLER_37_27 vgnd vpwr scs8hd_decap_12
XFILLER_53_59 vpwr vgnd scs8hd_fill_2
XFILLER_53_15 vgnd vpwr scs8hd_decap_12
XFILLER_41_204 vgnd vpwr scs8hd_fill_1
XFILLER_26_223 vgnd vpwr scs8hd_fill_1
XFILLER_5_127 vpwr vgnd scs8hd_fill_2
XANTENNA__67__A bottom_width_0_height_0__pin_45_lower vgnd vpwr scs8hd_diode_2
XFILLER_1_322 vpwr vgnd scs8hd_fill_2
XFILLER_1_300 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_93 vgnd vpwr scs8hd_decap_8
XFILLER_17_245 vgnd vpwr scs8hd_decap_3
XFILLER_17_234 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XFILLER_55_329 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_381 vgnd vpwr scs8hd_decap_4
XFILLER_23_215 vgnd vpwr scs8hd_decap_12
XFILLER_31_281 vgnd vpwr scs8hd_decap_12
XFILLER_48_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_58_178 vgnd vpwr scs8hd_decap_12
XFILLER_54_373 vgnd vpwr scs8hd_decap_4
XFILLER_46_318 vgnd vpwr scs8hd_decap_12
XFILLER_46_307 vpwr vgnd scs8hd_fill_2
XFILLER_14_204 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_22_270 vgnd vpwr scs8hd_decap_3
XFILLER_13_51 vgnd vpwr scs8hd_decap_8
XFILLER_14_215 vgnd vpwr scs8hd_fill_1
XFILLER_14_259 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_13_62 vgnd vpwr scs8hd_decap_4
XFILLER_13_84 vgnd vpwr scs8hd_decap_8
XFILLER_49_123 vgnd vpwr scs8hd_decap_12
XFILLER_1_163 vpwr vgnd scs8hd_fill_2
X_40_ _40_/HI _40_/LO vgnd vpwr scs8hd_conb_1
XFILLER_64_137 vgnd vpwr scs8hd_decap_12
XFILLER_54_80 vgnd vpwr scs8hd_decap_12
XFILLER_45_362 vpwr vgnd scs8hd_fill_2
XANTENNA_clkbuf_1_1__f_clk_A clkbuf_0_clk/X vgnd vpwr scs8hd_diode_2
XFILLER_62_3 vgnd vpwr scs8hd_decap_12
XFILLER_60_398 vgnd vpwr scs8hd_decap_8
XFILLER_9_274 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_55_159 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XPHY_519 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_508 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_398 vgnd vpwr scs8hd_decap_8
XFILLER_11_218 vpwr vgnd scs8hd_fill_2
XFILLER_50_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_27_351 vgnd vpwr scs8hd_fill_1
XANTENNA__80__A right_width_0_height_0__pin_41_lower vgnd vpwr scs8hd_diode_2
XFILLER_42_398 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
+ right_width_0_height_0__pin_14_ vgnd vpwr scs8hd_diode_2
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_255 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_37_159 vgnd vpwr scs8hd_decap_12
XFILLER_52_129 vgnd vpwr scs8hd_decap_12
XFILLER_33_376 vpwr vgnd scs8hd_fill_2
XFILLER_18_384 vgnd vpwr scs8hd_decap_12
XFILLER_29_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_45_27 vgnd vpwr scs8hd_decap_12
XPHY_316 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_305 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_354 vpwr vgnd scs8hd_fill_2
XFILLER_24_332 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_61_59 vpwr vgnd scs8hd_fill_2
XFILLER_61_15 vgnd vpwr scs8hd_decap_12
XFILLER_51_184 vgnd vpwr scs8hd_decap_12
XPHY_349 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_338 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_327 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_398 vgnd vpwr scs8hd_decap_8
XFILLER_3_236 vpwr vgnd scs8hd_fill_2
XFILLER_10_30 vgnd vpwr scs8hd_fill_1
XANTENNA__75__A right_width_0_height_0__pin_36_lower vgnd vpwr scs8hd_diode_2
XFILLER_19_148 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_129 vgnd vpwr scs8hd_decap_12
XFILLER_15_343 vpwr vgnd scs8hd_fill_2
XFILLER_30_379 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
XFILLER_33_184 vgnd vpwr scs8hd_decap_12
XFILLER_21_335 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_56_15 vgnd vpwr scs8hd_decap_12
XFILLER_29_402 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_124 vgnd vpwr scs8hd_decap_3
XPHY_113 vgnd vpwr scs8hd_decap_3
XFILLER_56_276 vgnd vpwr scs8hd_decap_12
XPHY_102 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_62 vgnd vpwr scs8hd_fill_1
XFILLER_21_40 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_84 vgnd vpwr scs8hd_decap_3
XFILLER_62_202 vgnd vpwr scs8hd_decap_12
XFILLER_47_232 vgnd vpwr scs8hd_decap_12
XFILLER_35_405 vpwr vgnd scs8hd_fill_2
XFILLER_62_80 vgnd vpwr scs8hd_decap_12
XFILLER_30_154 vgnd vpwr scs8hd_decap_12
XPHY_4 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_53 vpwr vgnd scs8hd_fill_2
XFILLER_7_75 vpwr vgnd scs8hd_fill_2
XFILLER_38_210 vpwr vgnd scs8hd_fill_2
XFILLER_53_257 vgnd vpwr scs8hd_decap_12
XFILLER_38_276 vgnd vpwr scs8hd_decap_4
XFILLER_21_110 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_21_198 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_ _60_/HI
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ right_width_0_height_0__pin_39_lower vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_202 vgnd vpwr scs8hd_decap_12
XFILLER_29_287 vgnd vpwr scs8hd_decap_6
XFILLER_29_265 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_405 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_16_84 vgnd vpwr scs8hd_decap_4
XFILLER_12_154 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_50_227 vgnd vpwr scs8hd_decap_12
XFILLER_35_235 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_37_39 vgnd vpwr scs8hd_decap_12
XFILLER_26_202 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_249 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_327 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_227 vgnd vpwr scs8hd_decap_4
XFILLER_40_293 vgnd vpwr scs8hd_decap_4
XFILLER_25_290 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_ _49_/HI
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ bottom_width_0_height_0__pin_48_lower vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_32 vpwr vgnd scs8hd_fill_2
XFILLER_4_43 vpwr vgnd scs8hd_fill_2
XFILLER_4_172 vpwr vgnd scs8hd_fill_2
XFILLER_63_330 vgnd vpwr scs8hd_decap_12
XFILLER_23_238 vgnd vpwr scs8hd_decap_4
XFILLER_23_227 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_293 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_48_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _43_/HI vgnd vpwr scs8hd_diode_2
XFILLER_64_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_54_341 vgnd vpwr scs8hd_decap_4
XANTENNA__78__A right_width_0_height_0__pin_39_lower vgnd vpwr scs8hd_diode_2
XFILLER_1_131 vpwr vgnd scs8hd_fill_2
XFILLER_64_149 vgnd vpwr scs8hd_decap_6
XFILLER_49_135 vgnd vpwr scs8hd_decap_12
XFILLER_38_93 vgnd vpwr scs8hd_decap_12
XFILLER_1_175 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_60_300 vgnd vpwr scs8hd_decap_12
XFILLER_45_352 vgnd vpwr scs8hd_decap_4
XFILLER_55_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_264 vgnd vpwr scs8hd_decap_4
XFILLER_9_297 vpwr vgnd scs8hd_fill_2
XFILLER_13_282 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_63_171 vgnd vpwr scs8hd_decap_12
XFILLER_48_190 vgnd vpwr scs8hd_decap_12
XFILLER_36_385 vpwr vgnd scs8hd_fill_2
XPHY_509 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_333 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_59_59 vpwr vgnd scs8hd_fill_2
XFILLER_59_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _57_/HI vgnd vpwr scs8hd_diode_2
XFILLER_46_105 vgnd vpwr scs8hd_decap_12
XFILLER_19_319 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_42_300 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XFILLER_24_84 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_234 vpwr vgnd scs8hd_fill_2
XFILLER_6_267 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_289 vpwr vgnd scs8hd_fill_2
XFILLER_45_171 vgnd vpwr scs8hd_decap_12
XFILLER_18_341 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_141 vgnd vpwr scs8hd_decap_12
XFILLER_33_388 vgnd vpwr scs8hd_decap_12
XFILLER_33_355 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_396 vgnd vpwr scs8hd_fill_1
XFILLER_45_39 vgnd vpwr scs8hd_decap_12
XPHY_339 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_328 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_317 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_306 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_366 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_61_27 vgnd vpwr scs8hd_decap_12
XFILLER_51_196 vgnd vpwr scs8hd_decap_12
XFILLER_10_97 vgnd vpwr scs8hd_decap_3
XFILLER_62_406 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
+ right_width_0_height_0__pin_8_ vgnd vpwr scs8hd_diode_2
XFILLER_27_160 vgnd vpwr scs8hd_decap_12
XFILLER_19_127 vpwr vgnd scs8hd_fill_2
XFILLER_19_116 vpwr vgnd scs8hd_fill_2
XFILLER_42_141 vgnd vpwr scs8hd_decap_12
XFILLER_30_369 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_18_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_281 vpwr vgnd scs8hd_fill_2
XFILLER_53_406 vgnd vpwr scs8hd_fill_1
XFILLER_21_303 vpwr vgnd scs8hd_fill_2
XFILLER_33_196 vgnd vpwr scs8hd_decap_12
XFILLER_21_358 vgnd vpwr scs8hd_decap_4
XFILLER_21_314 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_56_288 vgnd vpwr scs8hd_decap_4
XFILLER_56_27 vgnd vpwr scs8hd_decap_4
XFILLER_44_406 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_125 vgnd vpwr scs8hd_decap_3
XPHY_114 vgnd vpwr scs8hd_decap_3
XPHY_103 vgnd vpwr scs8hd_decap_3
XFILLER_24_152 vgnd vpwr scs8hd_fill_1
XFILLER_24_130 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_93 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
+ clkbuf_1_1__f_clk/X ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 Test_en
+ vgnd vpwr scs8hd_sdfxbp_1
XFILLER_15_152 vpwr vgnd scs8hd_fill_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_166 vgnd vpwr scs8hd_decap_12
XFILLER_15_196 vgnd vpwr scs8hd_fill_1
XFILLER_7_32 vpwr vgnd scs8hd_fill_2
XFILLER_7_351 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_7_87 vgnd vpwr scs8hd_fill_1
XFILLER_38_255 vpwr vgnd scs8hd_fill_2
XFILLER_26_406 vgnd vpwr scs8hd_fill_1
XFILLER_53_269 vgnd vpwr scs8hd_decap_12
XFILLER_38_299 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_29_299 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ right_width_0_height_0__pin_7_ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ vgnd vpwr scs8hd_or2_1
XFILLER_8_137 vpwr vgnd scs8hd_fill_2
XFILLER_12_111 vpwr vgnd scs8hd_fill_2
XFILLER_12_199 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_4_354 vgnd vpwr scs8hd_decap_3
XFILLER_4_376 vgnd vpwr scs8hd_decap_12
XFILLER_4_398 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_50_239 vgnd vpwr scs8hd_decap_12
XFILLER_35_269 vpwr vgnd scs8hd_fill_2
XFILLER_35_258 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_58_328 vgnd vpwr scs8hd_decap_6
XFILLER_26_247 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_5_107 vpwr vgnd scs8hd_fill_2
XFILLER_5_118 vpwr vgnd scs8hd_fill_2
XFILLER_57_350 vpwr vgnd scs8hd_fill_2
XFILLER_49_339 vgnd vpwr scs8hd_decap_12
XFILLER_49_306 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_27_62 vgnd vpwr scs8hd_decap_8
XFILLER_27_51 vgnd vpwr scs8hd_decap_8
XFILLER_40_261 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_22 vpwr vgnd scs8hd_fill_2
XFILLER_4_55 vpwr vgnd scs8hd_fill_2
XFILLER_4_88 vpwr vgnd scs8hd_fill_2
XFILLER_4_195 vgnd vpwr scs8hd_decap_4
XFILLER_63_342 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_280 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_39_350 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_27 vgnd vpwr scs8hd_decap_4
XFILLER_54_353 vgnd vpwr scs8hd_decap_4
XFILLER_13_97 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_106 vgnd vpwr scs8hd_decap_12
XFILLER_49_147 vgnd vpwr scs8hd_decap_12
XFILLER_54_93 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_1__f_clk/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_294 vgnd vpwr scs8hd_decap_8
XFILLER_48_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_51_345 vpwr vgnd scs8hd_fill_2
XFILLER_51_301 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_353 vpwr vgnd scs8hd_fill_2
XFILLER_36_320 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_117 vgnd vpwr scs8hd_decap_12
XFILLER_27_342 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ bottom_width_0_height_0__pin_50_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_0__f_clk/X vgnd vpwr scs8hd_diode_2
XFILLER_42_356 vgnd vpwr scs8hd_decap_4
XFILLER_27_364 vpwr vgnd scs8hd_fill_2
XFILLER_6_202 vpwr vgnd scs8hd_fill_2
XFILLER_10_231 vgnd vpwr scs8hd_decap_8
XFILLER_10_286 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_334 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_61_39 vgnd vpwr scs8hd_decap_12
XPHY_329 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_318 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_307 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_301 vgnd vpwr scs8hd_decap_4
XFILLER_59_220 vgnd vpwr scs8hd_decap_12
XFILLER_10_32 vpwr vgnd scs8hd_fill_2
XFILLER_10_65 vpwr vgnd scs8hd_fill_2
XFILLER_35_51 vgnd vpwr scs8hd_decap_8
XFILLER_27_172 vgnd vpwr scs8hd_decap_8
XFILLER_19_85 vpwr vgnd scs8hd_fill_2
XFILLER_19_52 vpwr vgnd scs8hd_fill_2
XFILLER_15_301 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
XFILLER_30_337 vgnd vpwr scs8hd_decap_6
XFILLER_30_326 vgnd vpwr scs8hd_decap_8
XFILLER_15_367 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_260 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _52_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XPHY_126 vgnd vpwr scs8hd_decap_3
XPHY_115 vgnd vpwr scs8hd_decap_3
XPHY_104 vgnd vpwr scs8hd_decap_3
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_337 vgnd vpwr scs8hd_decap_3
XFILLER_21_53 vpwr vgnd scs8hd_fill_2
XFILLER_47_245 vgnd vpwr scs8hd_decap_12
XFILLER_62_215 vgnd vpwr scs8hd_decap_12
XFILLER_47_289 vgnd vpwr scs8hd_decap_3
XFILLER_15_175 vgnd vpwr scs8hd_decap_8
XPHY_6 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_93 vgnd vpwr scs8hd_decap_12
XFILLER_30_178 vgnd vpwr scs8hd_decap_12
XFILLER_7_44 vgnd vpwr scs8hd_fill_1
XFILLER_7_363 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_11_392 vgnd vpwr scs8hd_decap_12
XFILLER_30_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_234 vpwr vgnd scs8hd_fill_2
XFILLER_61_281 vgnd vpwr scs8hd_decap_12
XFILLER_21_123 vgnd vpwr scs8hd_decap_12
XFILLER_29_245 vgnd vpwr scs8hd_decap_12
XFILLER_29_212 vgnd vpwr scs8hd_decap_12
XFILLER_44_215 vpwr vgnd scs8hd_fill_2
XFILLER_16_64 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_8_116 vpwr vgnd scs8hd_fill_2
XFILLER_12_134 vpwr vgnd scs8hd_fill_2
XFILLER_12_145 vgnd vpwr scs8hd_decap_8
XFILLER_12_178 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_4_388 vgnd vpwr scs8hd_decap_8
XFILLER_35_204 vpwr vgnd scs8hd_fill_2
XPHY_490 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_207 vpwr vgnd scs8hd_fill_2
XFILLER_26_215 vgnd vpwr scs8hd_decap_6
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
+ bottom_width_0_height_0__pin_26_ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_buf_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_358 vpwr vgnd scs8hd_fill_2
XFILLER_57_362 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_43_62 vgnd vpwr scs8hd_decap_12
XFILLER_43_51 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_284 vgnd vpwr scs8hd_fill_1
XFILLER_40_273 vpwr vgnd scs8hd_fill_2
XFILLER_4_141 vpwr vgnd scs8hd_fill_2
XFILLER_4_67 vpwr vgnd scs8hd_fill_2
XFILLER_4_163 vgnd vpwr scs8hd_decap_3
XFILLER_63_354 vgnd vpwr scs8hd_decap_12
XFILLER_48_362 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_39_384 vpwr vgnd scs8hd_fill_2
XFILLER_39_362 vpwr vgnd scs8hd_fill_2
XFILLER_54_398 vgnd vpwr scs8hd_decap_8
XFILLER_22_295 vpwr vgnd scs8hd_fill_2
XFILLER_6_406 vgnd vpwr scs8hd_fill_1
XFILLER_13_76 vpwr vgnd scs8hd_fill_2
XFILLER_8_3 vgnd vpwr scs8hd_decap_4
XFILLER_64_118 vgnd vpwr scs8hd_decap_6
XFILLER_49_159 vgnd vpwr scs8hd_decap_12
XFILLER_45_387 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_63_184 vgnd vpwr scs8hd_decap_12
XFILLER_36_398 vgnd vpwr scs8hd_decap_8
XFILLER_36_332 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_402 vgnd vpwr scs8hd_decap_4
XFILLER_59_39 vgnd vpwr scs8hd_decap_12
XFILLER_46_129 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
+ right_width_0_height_0__pin_5_ vgnd vpwr scs8hd_diode_2
XFILLER_27_376 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_10_265 vpwr vgnd scs8hd_fill_2
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
XFILLER_60_154 vgnd vpwr scs8hd_decap_12
XFILLER_45_184 vgnd vpwr scs8hd_decap_12
XFILLER_33_302 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_398 vgnd vpwr scs8hd_decap_8
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
XFILLER_60_3 vgnd vpwr scs8hd_decap_12
XFILLER_28_107 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_51_110 vgnd vpwr scs8hd_decap_12
XPHY_319 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_308 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_379 vpwr vgnd scs8hd_fill_2
XFILLER_24_324 vgnd vpwr scs8hd_decap_8
XFILLER_3_228 vpwr vgnd scs8hd_fill_2
XFILLER_10_22 vgnd vpwr scs8hd_decap_8
XFILLER_59_232 vgnd vpwr scs8hd_decap_12
XFILLER_42_154 vgnd vpwr scs8hd_decap_12
XFILLER_35_74 vgnd vpwr scs8hd_decap_12
XFILLER_27_184 vgnd vpwr scs8hd_decap_12
XFILLER_19_97 vgnd vpwr scs8hd_decap_4
XFILLER_51_62 vgnd vpwr scs8hd_decap_12
XFILLER_51_51 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_33_110 vgnd vpwr scs8hd_decap_12
XFILLER_18_195 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_202 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_209 vpwr vgnd scs8hd_fill_2
XPHY_116 vgnd vpwr scs8hd_decap_3
XPHY_105 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_127 vgnd vpwr scs8hd_decap_3
XFILLER_24_198 vgnd vpwr scs8hd_decap_12
XFILLER_24_154 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_316 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_21_76 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _35_/HI ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_47_257 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_227 vgnd vpwr scs8hd_decap_12
XFILLER_15_132 vgnd vpwr scs8hd_decap_3
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_7_342 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_38_202 vgnd vpwr scs8hd_decap_8
XFILLER_23_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_ _40_/HI
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ bottom_width_0_height_0__pin_45_lower vgnd vpwr scs8hd_mux2_1
XFILLER_61_293 vgnd vpwr scs8hd_decap_12
XFILLER_21_179 vpwr vgnd scs8hd_fill_2
XFILLER_21_135 vgnd vpwr scs8hd_decap_12
XFILLER_29_257 vgnd vpwr scs8hd_decap_8
XFILLER_29_224 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_32 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_4_334 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_290 vgnd vpwr scs8hd_decap_4
XPHY_491 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_480 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_271 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_271 vpwr vgnd scs8hd_fill_2
XFILLER_19_290 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
+ bottom_width_0_height_0__pin_25_ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_17_205 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_74 vgnd vpwr scs8hd_decap_12
XFILLER_58_105 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_333 vgnd vpwr scs8hd_decap_3
XFILLER_54_311 vgnd vpwr scs8hd_decap_3
XFILLER_54_300 vpwr vgnd scs8hd_fill_2
XFILLER_14_208 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_13_66 vgnd vpwr scs8hd_fill_1
XFILLER_1_167 vpwr vgnd scs8hd_fill_2
XFILLER_60_314 vpwr vgnd scs8hd_fill_2
XFILLER_57_171 vgnd vpwr scs8hd_decap_12
XFILLER_45_399 vgnd vpwr scs8hd_decap_8
XFILLER_9_223 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _51_/HI ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_196 vgnd vpwr scs8hd_decap_12
XFILLER_51_358 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_141 vgnd vpwr scs8hd_decap_12
XFILLER_39_171 vgnd vpwr scs8hd_decap_12
XFILLER_27_388 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_76 vpwr vgnd scs8hd_fill_2
XFILLER_24_54 vgnd vpwr scs8hd_fill_1
XFILLER_24_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XFILLER_6_259 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_49_62 vgnd vpwr scs8hd_decap_12
XFILLER_49_51 vgnd vpwr scs8hd_decap_8
XFILLER_18_322 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_60_166 vgnd vpwr scs8hd_decap_12
XFILLER_45_196 vgnd vpwr scs8hd_decap_12
XFILLER_53_3 vgnd vpwr scs8hd_decap_12
XFILLER_41_380 vpwr vgnd scs8hd_fill_2
XFILLER_5_281 vpwr vgnd scs8hd_fill_2
X_79_ right_width_0_height_0__pin_40_lower right_width_0_height_0__pin_40_upper vgnd
+ vpwr scs8hd_buf_2
XFILLER_56_406 vgnd vpwr scs8hd_fill_1
XFILLER_36_141 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_buf_2
XPHY_309 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_369 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
+ clkbuf_1_1__f_clk/X ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_/QN
+ top_width_0_height_0__pin_33_ Test_en vgnd vpwr scs8hd_sdfxbp_1
XFILLER_10_78 vpwr vgnd scs8hd_fill_2
XFILLER_42_166 vgnd vpwr scs8hd_decap_12
XFILLER_35_86 vgnd vpwr scs8hd_decap_12
XFILLER_27_196 vgnd vpwr scs8hd_decap_8
XFILLER_15_347 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _41_/HI vgnd vpwr scs8hd_diode_2
XFILLER_51_74 vgnd vpwr scs8hd_decap_12
XFILLER_23_380 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_38_406 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_18_174 vgnd vpwr scs8hd_decap_8
XFILLER_18_141 vgnd vpwr scs8hd_decap_12
XFILLER_21_306 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_29_406 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_280 vgnd vpwr scs8hd_decap_12
XPHY_128 vgnd vpwr scs8hd_decap_3
XPHY_117 vgnd vpwr scs8hd_decap_3
XPHY_106 vgnd vpwr scs8hd_decap_3
XFILLER_24_166 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_328 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_239 vgnd vpwr scs8hd_decap_12
XFILLER_47_269 vgnd vpwr scs8hd_decap_12
XFILLER_15_188 vpwr vgnd scs8hd_fill_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_7_57 vpwr vgnd scs8hd_fill_2
XFILLER_7_310 vpwr vgnd scs8hd_fill_2
XFILLER_7_376 vpwr vgnd scs8hd_fill_2
XFILLER_16_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_147 vgnd vpwr scs8hd_decap_6
XFILLER_21_114 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_29_236 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_88 vgnd vpwr scs8hd_fill_1
XFILLER_16_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_158 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XFILLER_4_346 vpwr vgnd scs8hd_fill_2
XFILLER_57_62 vgnd vpwr scs8hd_decap_12
XFILLER_57_51 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _63_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XPHY_492 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_481 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_470 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_294 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
+ bottom_width_0_height_0__pin_27_ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_261 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
+ bottom_width_0_height_0__pin_24_ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_buf_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_ _46_/HI
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_386 vgnd vpwr scs8hd_decap_12
XFILLER_25_250 vpwr vgnd scs8hd_fill_2
XFILLER_43_86 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_9_405 vpwr vgnd scs8hd_fill_2
XFILLER_4_47 vpwr vgnd scs8hd_fill_2
XFILLER_4_110 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_393 vgnd vpwr scs8hd_decap_8
XFILLER_0_382 vpwr vgnd scs8hd_fill_2
XFILLER_63_367 vgnd vpwr scs8hd_decap_12
XFILLER_31_220 vgnd vpwr scs8hd_decap_12
XFILLER_16_250 vgnd vpwr scs8hd_decap_3
XFILLER_58_117 vgnd vpwr scs8hd_decap_12
XFILLER_54_323 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
+ right_width_0_height_0__pin_2_ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_1_113 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_301 vpwr vgnd scs8hd_fill_2
XFILLER_1_135 vpwr vgnd scs8hd_fill_2
XFILLER_1_179 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_359 vgnd vpwr scs8hd_fill_1
XFILLER_60_337 vgnd vpwr scs8hd_decap_12
XFILLER_45_367 vgnd vpwr scs8hd_fill_1
XFILLER_13_242 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_1__f_clk/X vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_ _58_/HI
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_326 vgnd vpwr scs8hd_decap_4
XFILLER_36_389 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_27_301 vpwr vgnd scs8hd_fill_2
XFILLER_42_337 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_1__f_clk/X vgnd vpwr scs8hd_diode_2
XFILLER_50_381 vgnd vpwr scs8hd_decap_12
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
XFILLER_24_88 vpwr vgnd scs8hd_fill_2
XFILLER_6_238 vpwr vgnd scs8hd_fill_2
XFILLER_49_74 vgnd vpwr scs8hd_decap_12
XFILLER_18_345 vpwr vgnd scs8hd_fill_2
XFILLER_18_334 vpwr vgnd scs8hd_fill_2
XFILLER_1_26 vpwr vgnd scs8hd_fill_2
XFILLER_60_178 vgnd vpwr scs8hd_decap_12
XFILLER_33_359 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_271 vgnd vpwr scs8hd_decap_4
XFILLER_46_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
X_78_ right_width_0_height_0__pin_39_lower right_width_0_height_0__pin_39_upper vgnd
+ vpwr scs8hd_buf_2
XFILLER_51_123 vgnd vpwr scs8hd_decap_12
XFILLER_24_337 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
+ right_width_0_height_0__pin_14_ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_245 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_178 vgnd vpwr scs8hd_decap_12
XFILLER_35_98 vgnd vpwr scs8hd_decap_12
XFILLER_23_392 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_86 vgnd vpwr scs8hd_decap_12
XFILLER_2_285 vgnd vpwr scs8hd_decap_4
XFILLER_2_274 vgnd vpwr scs8hd_fill_1
XFILLER_33_123 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_318 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_215 vgnd vpwr scs8hd_decap_12
XPHY_129 vgnd vpwr scs8hd_decap_3
XFILLER_64_292 vgnd vpwr scs8hd_decap_12
XPHY_118 vgnd vpwr scs8hd_decap_3
XPHY_107 vgnd vpwr scs8hd_decap_3
XFILLER_24_178 vgnd vpwr scs8hd_decap_12
XFILLER_24_134 vgnd vpwr scs8hd_decap_12
XFILLER_12_307 vgnd vpwr scs8hd_decap_3
XFILLER_21_89 vpwr vgnd scs8hd_fill_2
XFILLER_20_362 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_55_281 vgnd vpwr scs8hd_decap_12
XFILLER_15_112 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_36 vpwr vgnd scs8hd_fill_2
XFILLER_7_300 vpwr vgnd scs8hd_fill_2
XFILLER_7_322 vgnd vpwr scs8hd_decap_12
XFILLER_11_362 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_7_355 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_270 vgnd vpwr scs8hd_decap_4
XFILLER_52_251 vgnd vpwr scs8hd_decap_12
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XFILLER_16_56 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_20_192 vpwr vgnd scs8hd_fill_2
XFILLER_4_303 vgnd vpwr scs8hd_decap_3
XFILLER_4_325 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _36_/HI vgnd vpwr scs8hd_diode_2
XFILLER_57_74 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_493 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_482 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_471 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_460 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_192 vgnd vpwr scs8hd_fill_1
XFILLER_3_391 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_295 vgnd vpwr scs8hd_fill_1
XFILLER_1_306 vgnd vpwr scs8hd_decap_3
XFILLER_8_90 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_398 vgnd vpwr scs8hd_decap_8
XFILLER_40_210 vgnd vpwr scs8hd_fill_1
XFILLER_25_273 vpwr vgnd scs8hd_fill_2
XFILLER_25_240 vpwr vgnd scs8hd_fill_2
XFILLER_17_218 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
+ bottom_width_0_height_0__pin_30_ vgnd vpwr scs8hd_diode_2
XFILLER_43_98 vgnd vpwr scs8hd_decap_12
XFILLER_40_276 vpwr vgnd scs8hd_fill_2
XFILLER_40_265 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_4_26 vgnd vpwr scs8hd_decap_3
XFILLER_4_59 vpwr vgnd scs8hd_fill_2
XFILLER_4_199 vgnd vpwr scs8hd_fill_1
XFILLER_48_398 vgnd vpwr scs8hd_decap_8
XFILLER_48_343 vgnd vpwr scs8hd_decap_12
XFILLER_63_379 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_262 vgnd vpwr scs8hd_decap_4
XPHY_290 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_129 vgnd vpwr scs8hd_decap_12
XFILLER_54_357 vgnd vpwr scs8hd_fill_1
XFILLER_39_376 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_287 vpwr vgnd scs8hd_fill_2
XFILLER_22_276 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_57_184 vgnd vpwr scs8hd_decap_12
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_53_390 vgnd vpwr scs8hd_decap_12
XFILLER_9_203 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_236 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_357 vpwr vgnd scs8hd_fill_2
XFILLER_36_346 vgnd vpwr scs8hd_decap_4
XFILLER_36_324 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_280 vpwr vgnd scs8hd_fill_2
XFILLER_39_184 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_54_154 vgnd vpwr scs8hd_decap_12
XFILLER_35_390 vgnd vpwr scs8hd_decap_4
XFILLER_50_393 vgnd vpwr scs8hd_decap_4
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_206 vgnd vpwr scs8hd_decap_8
XFILLER_10_213 vgnd vpwr scs8hd_fill_1
XFILLER_49_86 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_45_110 vgnd vpwr scs8hd_decap_12
XFILLER_33_316 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_33_338 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_294 vpwr vgnd scs8hd_fill_2
XFILLER_39_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
+ ccff_head vgnd vpwr scs8hd_diode_2
X_77_ right_width_0_height_0__pin_38_lower right_width_0_height_0__pin_38_upper vgnd
+ vpwr scs8hd_buf_2
XFILLER_51_135 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
+ right_width_0_height_0__pin_13_ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_36_154 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_36 vgnd vpwr scs8hd_decap_6
XFILLER_59_257 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XFILLER_27_132 vpwr vgnd scs8hd_fill_2
XFILLER_19_56 vgnd vpwr scs8hd_decap_3
XFILLER_50_190 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_98 vgnd vpwr scs8hd_decap_12
XFILLER_2_264 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_33_135 vgnd vpwr scs8hd_decap_12
XFILLER_18_154 vgnd vpwr scs8hd_fill_1
XFILLER_18_110 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_227 vgnd vpwr scs8hd_decap_12
XFILLER_24_102 vgnd vpwr scs8hd_decap_6
XPHY_119 vgnd vpwr scs8hd_decap_3
XPHY_108 vgnd vpwr scs8hd_decap_3
XFILLER_32_190 vgnd vpwr scs8hd_decap_12
XFILLER_24_146 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_20_341 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
XFILLER_21_35 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_55_293 vgnd vpwr scs8hd_decap_6
XFILLER_46_32 vgnd vpwr scs8hd_decap_12
XFILLER_30_105 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_7_334 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_7_367 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_53_208 vgnd vpwr scs8hd_decap_12
XFILLER_38_238 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_219 vpwr vgnd scs8hd_fill_2
XFILLER_37_293 vpwr vgnd scs8hd_fill_2
XFILLER_52_263 vgnd vpwr scs8hd_decap_12
XFILLER_32_56 vgnd vpwr scs8hd_decap_12
XFILLER_12_138 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_86 vgnd vpwr scs8hd_decap_12
XFILLER_35_208 vpwr vgnd scs8hd_fill_2
XPHY_461 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_450 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_494 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_483 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_472 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_175 vpwr vgnd scs8hd_fill_2
XFILLER_21_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_285 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_1_318 vpwr vgnd scs8hd_fill_2
XFILLER_57_333 vpwr vgnd scs8hd_fill_2
XFILLER_40_244 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_48_311 vgnd vpwr scs8hd_decap_3
XFILLER_4_145 vpwr vgnd scs8hd_fill_2
XFILLER_48_377 vpwr vgnd scs8hd_fill_2
XFILLER_48_366 vgnd vpwr scs8hd_fill_1
XFILLER_48_355 vgnd vpwr scs8hd_decap_4
XPHY_291 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_54_369 vpwr vgnd scs8hd_fill_2
XFILLER_39_388 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_299 vgnd vpwr scs8hd_decap_12
XFILLER_22_244 vgnd vpwr scs8hd_fill_1
XFILLER_10_406 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
+ bottom_width_0_height_0__pin_24_ vgnd vpwr scs8hd_diode_2
XFILLER_13_69 vgnd vpwr scs8hd_decap_3
XFILLER_8_7 vgnd vpwr scs8hd_fill_1
XFILLER_57_196 vgnd vpwr scs8hd_decap_12
XFILLER_54_32 vgnd vpwr scs8hd_decap_12
XFILLER_45_358 vpwr vgnd scs8hd_fill_2
XFILLER_45_325 vpwr vgnd scs8hd_fill_2
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XFILLER_60_328 vgnd vpwr scs8hd_decap_8
XFILLER_9_215 vpwr vgnd scs8hd_fill_2
XFILLER_48_141 vgnd vpwr scs8hd_decap_12
XFILLER_51_306 vgnd vpwr scs8hd_fill_1
XFILLER_36_303 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_59_406 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_39_196 vgnd vpwr scs8hd_decap_8
XFILLER_27_358 vgnd vpwr scs8hd_decap_4
XFILLER_27_347 vgnd vpwr scs8hd_decap_4
XFILLER_27_325 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_166 vgnd vpwr scs8hd_decap_12
XFILLER_24_46 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_269 vgnd vpwr scs8hd_decap_4
XFILLER_49_98 vgnd vpwr scs8hd_decap_12
XFILLER_33_328 vgnd vpwr scs8hd_decap_3
XFILLER_33_306 vgnd vpwr scs8hd_fill_1
XFILLER_18_369 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_240 vpwr vgnd scs8hd_fill_2
X_76_ right_width_0_height_0__pin_37_lower right_width_0_height_0__pin_37_upper vgnd
+ vpwr scs8hd_buf_2
XFILLER_51_147 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
+ right_width_0_height_0__pin_12_ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_36_166 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_15 vgnd vpwr scs8hd_decap_4
XFILLER_59_269 vgnd vpwr scs8hd_decap_12
XFILLER_15_306 vgnd vpwr scs8hd_decap_4
XFILLER_2_232 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_33_147 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_199 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XFILLER_51_3 vgnd vpwr scs8hd_decap_12
XFILLER_64_261 vgnd vpwr scs8hd_decap_12
XFILLER_56_239 vgnd vpwr scs8hd_decap_12
X_59_ _59_/HI _59_/LO vgnd vpwr scs8hd_conb_1
XPHY_109 vgnd vpwr scs8hd_decap_3
XFILLER_62_32 vgnd vpwr scs8hd_decap_12
XFILLER_46_44 vgnd vpwr scs8hd_decap_12
XFILLER_30_117 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_7_49 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_61_220 vgnd vpwr scs8hd_decap_12
XFILLER_46_294 vpwr vgnd scs8hd_fill_2
XFILLER_46_261 vgnd vpwr scs8hd_decap_12
XFILLER_21_106 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_98 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XPHY_495 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_484 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_473 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_462 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_451 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_440 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_150 vgnd vpwr scs8hd_decap_6
XFILLER_7_132 vpwr vgnd scs8hd_fill_2
XFILLER_14_3 vgnd vpwr scs8hd_decap_12
XFILLER_19_294 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
+ right_width_0_height_0__pin_2_ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_301 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_289 vpwr vgnd scs8hd_fill_2
XFILLER_4_102 vgnd vpwr scs8hd_decap_8
XFILLER_48_323 vgnd vpwr scs8hd_decap_12
XFILLER_0_363 vgnd vpwr scs8hd_decap_3
XFILLER_4_168 vpwr vgnd scs8hd_fill_2
XFILLER_48_389 vgnd vpwr scs8hd_decap_8
XFILLER_16_242 vpwr vgnd scs8hd_fill_2
XFILLER_31_245 vgnd vpwr scs8hd_decap_12
XFILLER_31_234 vpwr vgnd scs8hd_fill_2
XPHY_292 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XFILLER_54_337 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_ _61_/HI
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ right_width_0_height_0__pin_38_lower vgnd vpwr scs8hd_mux2_1
XFILLER_39_301 vpwr vgnd scs8hd_fill_2
XFILLER_13_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_127 vpwr vgnd scs8hd_fill_2
XFILLER_60_318 vgnd vpwr scs8hd_fill_1
XFILLER_54_44 vgnd vpwr scs8hd_decap_12
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
XFILLER_13_234 vgnd vpwr scs8hd_decap_8
XFILLER_13_245 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_123 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_271 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_5_71 vgnd vpwr scs8hd_decap_4
XFILLER_54_178 vgnd vpwr scs8hd_decap_12
XFILLER_42_318 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_50_373 vpwr vgnd scs8hd_fill_2
XFILLER_50_351 vpwr vgnd scs8hd_fill_2
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_123 vgnd vpwr scs8hd_decap_12
XFILLER_26_381 vgnd vpwr scs8hd_decap_12
XFILLER_18_337 vpwr vgnd scs8hd_fill_2
XFILLER_41_384 vgnd vpwr scs8hd_decap_12
XFILLER_14_91 vgnd vpwr scs8hd_fill_1
X_75_ right_width_0_height_0__pin_36_lower right_width_0_height_0__pin_36_upper vgnd
+ vpwr scs8hd_buf_2
XFILLER_36_178 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XFILLER_51_159 vgnd vpwr scs8hd_decap_12
XFILLER_32_384 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_381 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_27_101 vpwr vgnd scs8hd_fill_2
XFILLER_19_47 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_90 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_33_159 vgnd vpwr scs8hd_decap_12
XFILLER_25_90 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XFILLER_44_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _51_/HI vgnd vpwr scs8hd_diode_2
XFILLER_64_273 vgnd vpwr scs8hd_decap_6
XFILLER_49_281 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
X_58_ _58_/HI _58_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_72 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_15 vgnd vpwr scs8hd_decap_12
XFILLER_20_398 vgnd vpwr scs8hd_decap_8
XFILLER_20_321 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_56 vgnd vpwr scs8hd_decap_12
XFILLER_62_44 vgnd vpwr scs8hd_decap_12
XFILLER_30_129 vgnd vpwr scs8hd_decap_12
XFILLER_23_192 vpwr vgnd scs8hd_fill_2
XFILLER_15_137 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_7_314 vpwr vgnd scs8hd_fill_2
XFILLER_7_347 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_11_81 vgnd vpwr scs8hd_decap_12
XFILLER_61_232 vgnd vpwr scs8hd_decap_12
XFILLER_46_273 vpwr vgnd scs8hd_fill_2
XFILLER_46_251 vpwr vgnd scs8hd_fill_2
XFILLER_14_192 vgnd vpwr scs8hd_fill_1
XFILLER_37_240 vpwr vgnd scs8hd_fill_2
XFILLER_52_276 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_16_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_107 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_240 vgnd vpwr scs8hd_decap_4
XPHY_496 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_485 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_474 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_463 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_452 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_441 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_430 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_298 vgnd vpwr scs8hd_fill_1
XFILLER_31_405 vpwr vgnd scs8hd_fill_2
XFILLER_7_111 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_184 vpwr vgnd scs8hd_fill_2
XFILLER_34_210 vpwr vgnd scs8hd_fill_2
XFILLER_19_262 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
+ right_width_0_height_0__pin_1_ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
+ bottom_width_0_height_0__pin_21_ vgnd vpwr scs8hd_diode_2
XFILLER_8_82 vgnd vpwr scs8hd_decap_8
XFILLER_8_93 vgnd vpwr scs8hd_decap_4
XFILLER_57_346 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_213 vgnd vpwr scs8hd_fill_1
XFILLER_40_202 vgnd vpwr scs8hd_decap_8
XFILLER_25_298 vpwr vgnd scs8hd_fill_2
XFILLER_13_405 vpwr vgnd scs8hd_fill_2
XFILLER_4_114 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_48_335 vgnd vpwr scs8hd_fill_1
XFILLER_0_386 vpwr vgnd scs8hd_fill_2
XFILLER_0_342 vpwr vgnd scs8hd_fill_2
XFILLER_16_276 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_31_257 vgnd vpwr scs8hd_decap_12
XPHY_293 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_349 vpwr vgnd scs8hd_fill_2
XFILLER_54_327 vgnd vpwr scs8hd_decap_4
XFILLER_22_235 vgnd vpwr scs8hd_fill_1
XFILLER_22_202 vgnd vpwr scs8hd_decap_12
XFILLER_13_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_110 vgnd vpwr scs8hd_decap_12
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
XFILLER_1_117 vgnd vpwr scs8hd_decap_3
XFILLER_54_56 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_13_202 vpwr vgnd scs8hd_fill_2
XFILLER_13_257 vgnd vpwr scs8hd_decap_4
XFILLER_63_135 vgnd vpwr scs8hd_decap_12
XFILLER_48_154 vgnd vpwr scs8hd_decap_12
XFILLER_29_390 vgnd vpwr scs8hd_decap_12
XFILLER_0_183 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_5_83 vpwr vgnd scs8hd_fill_2
XFILLER_42_308 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_62_190 vgnd vpwr scs8hd_decap_12
XFILLER_50_341 vgnd vpwr scs8hd_decap_8
XFILLER_10_205 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_45_135 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_349 vgnd vpwr scs8hd_decap_12
XFILLER_60_105 vgnd vpwr scs8hd_decap_12
XFILLER_41_330 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_26_393 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_41_396 vgnd vpwr scs8hd_decap_8
XFILLER_14_81 vpwr vgnd scs8hd_fill_2
XFILLER_30_80 vgnd vpwr scs8hd_decap_12
X_74_ right_width_0_height_0__pin_35_lower right_width_0_height_0__pin_35_upper vgnd
+ vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_190 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_1__f_clk/X vgnd vpwr scs8hd_diode_2
XFILLER_32_396 vgnd vpwr scs8hd_fill_1
XFILLER_32_352 vpwr vgnd scs8hd_fill_2
XFILLER_32_341 vgnd vpwr scs8hd_fill_1
XFILLER_17_393 vgnd vpwr scs8hd_decap_12
XFILLER_19_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _53_/HI vgnd vpwr scs8hd_diode_2
XFILLER_42_105 vgnd vpwr scs8hd_decap_12
XFILLER_23_363 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_289 vgnd vpwr scs8hd_fill_1
XFILLER_2_201 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_18_113 vpwr vgnd scs8hd_fill_2
XFILLER_18_102 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_91 vgnd vpwr scs8hd_decap_3
XFILLER_41_171 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_decap_3
XFILLER_26_190 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_84 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_230 vgnd vpwr scs8hd_decap_12
X_57_ _57_/HI _57_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_21_27 vgnd vpwr scs8hd_decap_8
XFILLER_20_366 vpwr vgnd scs8hd_fill_2
XFILLER_20_333 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
+ right_width_0_height_0__pin_15_ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_208 vgnd vpwr scs8hd_decap_12
XFILLER_46_68 vgnd vpwr scs8hd_decap_12
XFILLER_15_116 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ bottom_width_0_height_0__pin_27_ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/A
+ vgnd vpwr scs8hd_or2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_62_56 vgnd vpwr scs8hd_decap_12
XFILLER_23_171 vgnd vpwr scs8hd_decap_12
XFILLER_15_149 vgnd vpwr scs8hd_fill_1
XFILLER_7_304 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_11_322 vpwr vgnd scs8hd_fill_2
XFILLER_11_388 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_14_171 vgnd vpwr scs8hd_decap_8
XFILLER_6_370 vgnd vpwr scs8hd_fill_1
XFILLER_52_288 vgnd vpwr scs8hd_decap_12
XFILLER_40_406 vgnd vpwr scs8hd_fill_1
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
XFILLER_20_141 vgnd vpwr scs8hd_decap_12
XFILLER_16_27 vgnd vpwr scs8hd_decap_4
XFILLER_20_196 vgnd vpwr scs8hd_fill_1
XFILLER_4_329 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_211 vpwr vgnd scs8hd_fill_2
XPHY_497 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_486 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_475 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_464 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_453 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_442 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_431 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_420 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_70 vpwr vgnd scs8hd_fill_2
XFILLER_11_163 vpwr vgnd scs8hd_fill_2
XFILLER_11_174 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_7_167 vgnd vpwr scs8hd_decap_3
XFILLER_19_230 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_22_406 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
+ right_width_0_height_0__pin_0_ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_57_358 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_27_59 vpwr vgnd scs8hd_fill_2
XFILLER_27_15 vgnd vpwr scs8hd_decap_12
XFILLER_25_222 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_25_277 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_137 vpwr vgnd scs8hd_fill_2
XFILLER_63_306 vgnd vpwr scs8hd_decap_12
XFILLER_48_369 vgnd vpwr scs8hd_decap_4
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_81 vpwr vgnd scs8hd_fill_2
XFILLER_16_266 vgnd vpwr scs8hd_fill_1
XFILLER_16_211 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_31_269 vgnd vpwr scs8hd_decap_12
XPHY_294 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_192 vpwr vgnd scs8hd_fill_2
XFILLER_54_306 vgnd vpwr scs8hd_decap_3
XFILLER_39_358 vpwr vgnd scs8hd_fill_2
XFILLER_62_361 vgnd vpwr scs8hd_decap_12
XFILLER_22_247 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_68 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_207 vpwr vgnd scs8hd_fill_2
XFILLER_21_291 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_229 vgnd vpwr scs8hd_fill_1
XFILLER_0_151 vpwr vgnd scs8hd_fill_2
XFILLER_63_147 vgnd vpwr scs8hd_decap_12
XFILLER_48_166 vgnd vpwr scs8hd_decap_12
XFILLER_44_394 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_8_251 vpwr vgnd scs8hd_fill_2
XFILLER_8_284 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
+ prog_clk ccff_head ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_5_95 vpwr vgnd scs8hd_fill_2
XFILLER_24_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_239 vgnd vpwr scs8hd_fill_1
XFILLER_45_147 vgnd vpwr scs8hd_decap_12
XFILLER_60_117 vgnd vpwr scs8hd_decap_12
XFILLER_41_364 vpwr vgnd scs8hd_fill_2
XFILLER_41_320 vpwr vgnd scs8hd_fill_2
XFILLER_26_350 vgnd vpwr scs8hd_decap_4
XFILLER_14_60 vpwr vgnd scs8hd_fill_2
XFILLER_5_221 vpwr vgnd scs8hd_fill_2
XFILLER_5_254 vpwr vgnd scs8hd_fill_2
XFILLER_5_298 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
X_73_ right_width_0_height_0__pin_34_lower right_width_0_height_0__pin_34_upper vgnd
+ vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_361 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_136 vgnd vpwr scs8hd_decap_12
XFILLER_27_114 vpwr vgnd scs8hd_fill_2
XFILLER_19_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_117 vgnd vpwr scs8hd_decap_12
XFILLER_35_59 vpwr vgnd scs8hd_fill_2
XFILLER_2_268 vgnd vpwr scs8hd_decap_4
XFILLER_2_224 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_18_136 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XPHY_92 vgnd vpwr scs8hd_decap_3
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_242 vgnd vpwr scs8hd_decap_6
X_56_ _56_/HI _56_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_96 vpwr vgnd scs8hd_fill_2
XFILLER_2_41 vpwr vgnd scs8hd_fill_2
XFILLER_20_312 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_389 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_55_220 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_11_312 vgnd vpwr scs8hd_fill_1
XFILLER_11_345 vpwr vgnd scs8hd_fill_2
XFILLER_11_356 vgnd vpwr scs8hd_decap_4
XFILLER_11_367 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_61_245 vgnd vpwr scs8hd_decap_12
XFILLER_36_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
+ bottom_width_0_height_0__pin_18_ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xclkbuf_1_0__f_clk clkbuf_0_clk/X clkbuf_1_0__f_clk/X vgnd vpwr scs8hd_clkbuf_16
XFILLER_37_297 vpwr vgnd scs8hd_fill_2
XFILLER_37_231 vpwr vgnd scs8hd_fill_2
X_39_ _39_/HI _39_/LO vgnd vpwr scs8hd_conb_1
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XFILLER_20_164 vpwr vgnd scs8hd_fill_2
XFILLER_20_120 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_ _52_/HI
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ right_width_0_height_0__pin_35_lower vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XPHY_443 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_432 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_421 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_267 vpwr vgnd scs8hd_fill_2
XFILLER_43_245 vgnd vpwr scs8hd_decap_3
XFILLER_43_234 vpwr vgnd scs8hd_fill_2
XPHY_410 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_498 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_487 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_476 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_465 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_454 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_93 vpwr vgnd scs8hd_fill_2
XFILLER_7_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_363 vgnd vpwr scs8hd_decap_3
XFILLER_34_234 vgnd vpwr scs8hd_decap_6
XFILLER_19_253 vgnd vpwr scs8hd_decap_6
XFILLER_19_242 vpwr vgnd scs8hd_fill_2
XFILLER_34_289 vgnd vpwr scs8hd_decap_6
XFILLER_8_51 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_clkbuf_1_0__f_clk_A clkbuf_0_clk/X vgnd vpwr scs8hd_diode_2
XFILLER_6_190 vpwr vgnd scs8hd_fill_2
XFILLER_27_27 vgnd vpwr scs8hd_decap_12
XFILLER_43_15 vgnd vpwr scs8hd_decap_12
XFILLER_40_215 vgnd vpwr scs8hd_decap_3
XFILLER_25_245 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_43_59 vpwr vgnd scs8hd_fill_2
XFILLER_0_333 vpwr vgnd scs8hd_fill_2
XFILLER_0_311 vgnd vpwr scs8hd_decap_3
XFILLER_4_149 vpwr vgnd scs8hd_fill_2
XFILLER_63_318 vgnd vpwr scs8hd_decap_12
XFILLER_48_359 vgnd vpwr scs8hd_fill_1
XFILLER_48_337 vgnd vpwr scs8hd_decap_3
XPHY_295 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_234 vgnd vpwr scs8hd_decap_8
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_ _41_/HI
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ bottom_width_0_height_0__pin_44_lower vgnd vpwr scs8hd_mux2_1
XFILLER_39_326 vgnd vpwr scs8hd_decap_12
XFILLER_39_315 vpwr vgnd scs8hd_fill_2
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XFILLER_62_373 vgnd vpwr scs8hd_decap_12
XFILLER_47_381 vgnd vpwr scs8hd_decap_4
XFILLER_22_215 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_270 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_123 vgnd vpwr scs8hd_decap_12
XFILLER_45_329 vpwr vgnd scs8hd_fill_2
XFILLER_38_15 vgnd vpwr scs8hd_decap_12
XFILLER_53_362 vpwr vgnd scs8hd_fill_2
XFILLER_53_351 vgnd vpwr scs8hd_fill_1
XFILLER_53_340 vgnd vpwr scs8hd_decap_4
XFILLER_9_219 vpwr vgnd scs8hd_fill_2
XFILLER_5_403 vgnd vpwr scs8hd_decap_4
XFILLER_63_159 vgnd vpwr scs8hd_decap_12
XFILLER_48_178 vgnd vpwr scs8hd_decap_12
XFILLER_36_307 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_80 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_5_52 vgnd vpwr scs8hd_decap_3
XFILLER_39_123 vgnd vpwr scs8hd_decap_12
XFILLER_27_329 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _54_/HI vgnd vpwr scs8hd_diode_2
XFILLER_50_398 vgnd vpwr scs8hd_decap_8
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
XFILLER_2_406 vgnd vpwr scs8hd_fill_1
XFILLER_45_159 vgnd vpwr scs8hd_decap_12
XFILLER_26_373 vpwr vgnd scs8hd_fill_2
XFILLER_60_129 vgnd vpwr scs8hd_decap_12
XFILLER_41_376 vpwr vgnd scs8hd_fill_2
XANTENNA__70__A bottom_width_0_height_0__pin_48_lower vgnd vpwr scs8hd_diode_2
XFILLER_30_93 vgnd vpwr scs8hd_decap_12
XFILLER_5_277 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
X_72_ bottom_width_0_height_0__pin_50_ bottom_width_0_height_0__pin_51_ vgnd vpwr
+ scs8hd_buf_2
XFILLER_17_373 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_398 vgnd vpwr scs8hd_decap_8
XFILLER_10_19 vgnd vpwr scs8hd_fill_1
XFILLER_55_402 vgnd vpwr scs8hd_decap_4
XFILLER_35_27 vgnd vpwr scs8hd_decap_12
XFILLER_27_148 vgnd vpwr scs8hd_decap_12
XFILLER_19_39 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XFILLER_51_59 vpwr vgnd scs8hd_fill_2
XFILLER_51_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_129 vgnd vpwr scs8hd_decap_12
XFILLER_23_376 vpwr vgnd scs8hd_fill_2
XFILLER_23_343 vgnd vpwr scs8hd_decap_3
XFILLER_23_310 vgnd vpwr scs8hd_decap_3
XFILLER_2_236 vgnd vpwr scs8hd_decap_3
XFILLER_58_251 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_61_405 vpwr vgnd scs8hd_fill_2
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_60 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA__65__A bottom_width_0_height_0__pin_43_lower vgnd vpwr scs8hd_diode_2
XFILLER_14_310 vpwr vgnd scs8hd_fill_2
XFILLER_14_343 vgnd vpwr scs8hd_fill_1
XPHY_93 vgnd vpwr scs8hd_decap_3
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
XFILLER_14_398 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
X_55_ _55_/HI _55_/LO vgnd vpwr scs8hd_conb_1
XFILLER_20_302 vgnd vpwr scs8hd_decap_4
XFILLER_17_192 vgnd vpwr scs8hd_decap_8
XFILLER_17_170 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_55_232 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_184 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_46_276 vgnd vpwr scs8hd_decap_12
XFILLER_46_243 vgnd vpwr scs8hd_decap_8
XFILLER_61_257 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_14_195 vgnd vpwr scs8hd_fill_1
XFILLER_52_80 vgnd vpwr scs8hd_decap_12
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_52_202 vgnd vpwr scs8hd_decap_12
XFILLER_37_276 vpwr vgnd scs8hd_fill_2
XFILLER_37_254 vpwr vgnd scs8hd_fill_2
XFILLER_25_405 vpwr vgnd scs8hd_fill_2
X_38_ _38_/HI _38_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_20_154 vpwr vgnd scs8hd_fill_2
XFILLER_20_132 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_477 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_466 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_455 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_444 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_433 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_422 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_411 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_400 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_276 vgnd vpwr scs8hd_decap_12
XPHY_499 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_488 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_50 vgnd vpwr scs8hd_fill_1
XFILLER_7_114 vpwr vgnd scs8hd_fill_2
XFILLER_7_136 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
+ right_width_0_height_0__pin_12_ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_353 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_390 vgnd vpwr scs8hd_decap_4
XFILLER_34_202 vgnd vpwr scs8hd_decap_8
XFILLER_19_298 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_27_39 vgnd vpwr scs8hd_decap_12
XFILLER_43_27 vgnd vpwr scs8hd_decap_12
XFILLER_40_227 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_316 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_16_246 vpwr vgnd scs8hd_fill_2
XANTENNA__73__A right_width_0_height_0__pin_34_lower vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_238 vgnd vpwr scs8hd_decap_6
XPHY_296 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_3_161 vgnd vpwr scs8hd_decap_3
XFILLER_39_338 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_62_385 vgnd vpwr scs8hd_decap_12
XFILLER_47_360 vgnd vpwr scs8hd_decap_6
XFILLER_22_238 vgnd vpwr scs8hd_decap_6
XFILLER_22_227 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_109 vpwr vgnd scs8hd_fill_2
XFILLER_57_135 vgnd vpwr scs8hd_decap_12
XFILLER_54_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ right_width_0_height_0__pin_15_ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/A
+ vgnd vpwr scs8hd_or2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA__68__A bottom_width_0_height_0__pin_46_lower vgnd vpwr scs8hd_diode_2
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XFILLER_0_175 vpwr vgnd scs8hd_fill_2
XFILLER_56_190 vgnd vpwr scs8hd_decap_12
XFILLER_44_363 vpwr vgnd scs8hd_fill_2
XFILLER_28_93 vgnd vpwr scs8hd_decap_12
XFILLER_60_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_20 vpwr vgnd scs8hd_fill_2
XFILLER_5_75 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_54_105 vgnd vpwr scs8hd_decap_12
XFILLER_39_135 vgnd vpwr scs8hd_decap_12
XFILLER_35_330 vpwr vgnd scs8hd_fill_2
XFILLER_50_355 vgnd vpwr scs8hd_decap_3
XFILLER_35_363 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_ _34_/HI
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XFILLER_10_219 vgnd vpwr scs8hd_decap_12
XFILLER_49_59 vpwr vgnd scs8hd_fill_2
XFILLER_49_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_53_171 vgnd vpwr scs8hd_decap_12
XFILLER_41_311 vpwr vgnd scs8hd_fill_2
XFILLER_38_190 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_105 vgnd vpwr scs8hd_decap_12
XFILLER_29_190 vgnd vpwr scs8hd_fill_1
X_71_ bottom_width_0_height_0__pin_49_lower bottom_width_0_height_0__pin_49_upper
+ vgnd vpwr scs8hd_buf_2
XFILLER_32_344 vpwr vgnd scs8hd_fill_2
XFILLER_32_333 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_0__f_clk/X vgnd vpwr scs8hd_diode_2
XFILLER_59_208 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_171 vgnd vpwr scs8hd_decap_12
XFILLER_35_39 vgnd vpwr scs8hd_decap_12
XFILLER_51_27 vgnd vpwr scs8hd_decap_12
XFILLER_50_141 vgnd vpwr scs8hd_decap_12
XFILLER_23_388 vpwr vgnd scs8hd_fill_2
XFILLER_23_355 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _39_/HI ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_mux2_1
XFILLER_58_263 vgnd vpwr scs8hd_decap_12
XPHY_94 vgnd vpwr scs8hd_decap_3
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XFILLER_14_366 vgnd vpwr scs8hd_fill_1
XFILLER_14_300 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_196 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_211 vgnd vpwr scs8hd_decap_6
XFILLER_52_406 vgnd vpwr scs8hd_fill_1
XFILLER_49_285 vgnd vpwr scs8hd_fill_1
XFILLER_37_403 vgnd vpwr scs8hd_decap_4
XFILLER_24_108 vgnd vpwr scs8hd_fill_1
XFILLER_2_76 vpwr vgnd scs8hd_fill_2
X_54_ _54_/HI _54_/LO vgnd vpwr scs8hd_conb_1
XFILLER_32_141 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _58_/HI vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_46_27 vgnd vpwr scs8hd_decap_4
XFILLER_62_15 vgnd vpwr scs8hd_decap_12
XFILLER_15_108 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _37_/HI vgnd vpwr scs8hd_diode_2
XFILLER_7_318 vpwr vgnd scs8hd_fill_2
XFILLER_11_41 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_2_3 vgnd vpwr scs8hd_fill_1
XANTENNA__76__A right_width_0_height_0__pin_37_lower vgnd vpwr scs8hd_diode_2
XFILLER_46_288 vgnd vpwr scs8hd_decap_4
XFILLER_34_406 vgnd vpwr scs8hd_fill_1
XFILLER_61_269 vgnd vpwr scs8hd_decap_12
XFILLER_36_93 vgnd vpwr scs8hd_decap_12
XFILLER_6_340 vgnd vpwr scs8hd_decap_12
XFILLER_6_373 vgnd vpwr scs8hd_decap_12
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_37_266 vpwr vgnd scs8hd_fill_2
X_37_ _37_/HI _37_/LO vgnd vpwr scs8hd_conb_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_20_188 vpwr vgnd scs8hd_fill_2
XFILLER_57_15 vgnd vpwr scs8hd_decap_12
XFILLER_57_59 vpwr vgnd scs8hd_fill_2
XFILLER_28_244 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_406 vgnd vpwr scs8hd_fill_1
XPHY_489 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_478 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_467 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_456 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_445 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_434 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_423 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_412 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_401 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_84 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_321 vpwr vgnd scs8hd_fill_2
XFILLER_7_159 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_188 vgnd vpwr scs8hd_decap_4
XFILLER_19_266 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_57_306 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_43_39 vgnd vpwr scs8hd_decap_12
XFILLER_33_291 vgnd vpwr scs8hd_decap_4
XFILLER_25_236 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_368 vpwr vgnd scs8hd_fill_2
XFILLER_0_302 vpwr vgnd scs8hd_fill_2
XFILLER_56_361 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_269 vgnd vpwr scs8hd_decap_6
XFILLER_16_203 vpwr vgnd scs8hd_fill_2
XPHY_297 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_286 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _55_/HI ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_mux2_1
XFILLER_3_184 vpwr vgnd scs8hd_fill_2
XFILLER_58_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_147 vgnd vpwr scs8hd_decap_12
XFILLER_54_27 vgnd vpwr scs8hd_decap_4
XFILLER_53_386 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_187 vgnd vpwr scs8hd_decap_3
XFILLER_44_386 vgnd vpwr scs8hd_decap_8
XFILLER_44_93 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_250 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_5_32 vpwr vgnd scs8hd_fill_2
XFILLER_5_87 vpwr vgnd scs8hd_fill_2
XFILLER_54_117 vgnd vpwr scs8hd_decap_12
XFILLER_39_147 vgnd vpwr scs8hd_decap_12
XFILLER_50_334 vpwr vgnd scs8hd_fill_2
XFILLER_35_397 vgnd vpwr scs8hd_decap_8
XFILLER_35_386 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_27 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_14_85 vgnd vpwr scs8hd_decap_6
XANTENNA__79__A right_width_0_height_0__pin_40_lower vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XFILLER_64_404 vgnd vpwr scs8hd_decap_3
XFILLER_36_117 vgnd vpwr scs8hd_decap_12
X_70_ bottom_width_0_height_0__pin_48_lower bottom_width_0_height_0__pin_48_upper
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_205 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_18_106 vgnd vpwr scs8hd_decap_4
XPHY_95 vgnd vpwr scs8hd_decap_3
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_62 vpwr vgnd scs8hd_fill_2
XFILLER_25_51 vgnd vpwr scs8hd_decap_8
XPHY_40 vgnd vpwr scs8hd_decap_3
XFILLER_14_389 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_323 vpwr vgnd scs8hd_fill_2
XFILLER_49_220 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
X_53_ _53_/HI _53_/LO vgnd vpwr scs8hd_conb_1
XFILLER_49_297 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_2_88 vpwr vgnd scs8hd_fill_2
XFILLER_20_337 vpwr vgnd scs8hd_fill_2
XFILLER_9_360 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_55_245 vgnd vpwr scs8hd_decap_12
XFILLER_62_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_53 vpwr vgnd scs8hd_fill_2
XFILLER_19_404 vgnd vpwr scs8hd_decap_3
XFILLER_46_223 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
+ right_width_0_height_0__pin_9_ vgnd vpwr scs8hd_diode_2
XFILLER_52_93 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_ _32_/HI
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ right_width_0_height_0__pin_41_lower vgnd vpwr scs8hd_mux2_1
XFILLER_6_352 vgnd vpwr scs8hd_decap_12
XFILLER_6_385 vgnd vpwr scs8hd_decap_12
XFILLER_28_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
X_36_ _36_/HI _36_/LO vgnd vpwr scs8hd_conb_1
XFILLER_52_215 vgnd vpwr scs8hd_decap_12
XFILLER_37_289 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_57_27 vgnd vpwr scs8hd_decap_12
XFILLER_28_267 vgnd vpwr scs8hd_decap_8
XPHY_479 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_51_281 vgnd vpwr scs8hd_decap_8
XPHY_468 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_457 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_446 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_435 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_424 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_413 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_402 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_123 vgnd vpwr scs8hd_decap_3
XFILLER_11_156 vgnd vpwr scs8hd_fill_1
XFILLER_11_167 vgnd vpwr scs8hd_decap_3
XFILLER_11_178 vgnd vpwr scs8hd_decap_3
XFILLER_22_74 vgnd vpwr scs8hd_decap_6
XFILLER_19_245 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_8_10 vpwr vgnd scs8hd_fill_2
XFILLER_57_329 vpwr vgnd scs8hd_fill_2
XFILLER_25_226 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _62_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_56_384 vgnd vpwr scs8hd_decap_12
XFILLER_56_351 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _32_/HI vgnd vpwr scs8hd_diode_2
XFILLER_17_85 vpwr vgnd scs8hd_fill_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XFILLER_33_51 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XPHY_298 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_287 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_196 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_62_398 vgnd vpwr scs8hd_decap_8
XFILLER_30_251 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_57_159 vgnd vpwr scs8hd_decap_12
XFILLER_53_354 vpwr vgnd scs8hd_fill_2
XFILLER_53_310 vpwr vgnd scs8hd_fill_2
XFILLER_38_362 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_295 vpwr vgnd scs8hd_fill_2
XFILLER_21_240 vpwr vgnd scs8hd_fill_2
XFILLER_44_332 vpwr vgnd scs8hd_fill_2
XFILLER_29_362 vpwr vgnd scs8hd_fill_2
XFILLER_29_351 vgnd vpwr scs8hd_decap_3
XFILLER_44_398 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_93 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_44 vpwr vgnd scs8hd_fill_2
XFILLER_8_255 vgnd vpwr scs8hd_decap_3
XFILLER_12_295 vgnd vpwr scs8hd_decap_12
XFILLER_39_159 vgnd vpwr scs8hd_decap_12
XFILLER_5_99 vpwr vgnd scs8hd_fill_2
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XFILLER_54_129 vgnd vpwr scs8hd_decap_12
XFILLER_50_313 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_49_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_53_184 vgnd vpwr scs8hd_decap_12
XFILLER_41_324 vgnd vpwr scs8hd_decap_4
XFILLER_41_302 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_26_398 vgnd vpwr scs8hd_decap_8
XFILLER_26_332 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _39_/HI vgnd vpwr scs8hd_diode_2
XFILLER_5_225 vpwr vgnd scs8hd_fill_2
XFILLER_5_236 vpwr vgnd scs8hd_fill_2
XFILLER_5_258 vpwr vgnd scs8hd_fill_2
XFILLER_14_64 vgnd vpwr scs8hd_decap_3
XFILLER_14_97 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_129 vgnd vpwr scs8hd_decap_12
XFILLER_32_313 vgnd vpwr scs8hd_decap_12
XFILLER_17_365 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_32_357 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
+ right_width_0_height_0__pin_3_ vgnd vpwr scs8hd_diode_2
XFILLER_58_3 vgnd vpwr scs8hd_decap_12
XFILLER_4_280 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_154 vgnd vpwr scs8hd_decap_12
XFILLER_35_184 vgnd vpwr scs8hd_decap_12
XFILLER_2_228 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_58_276 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XFILLER_25_85 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_14_335 vgnd vpwr scs8hd_fill_1
XFILLER_14_346 vgnd vpwr scs8hd_decap_3
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
XFILLER_49_232 vgnd vpwr scs8hd_decap_12
XFILLER_2_45 vpwr vgnd scs8hd_fill_2
XFILLER_2_23 vpwr vgnd scs8hd_fill_2
X_52_ _52_/HI _52_/LO vgnd vpwr scs8hd_conb_1
XFILLER_32_154 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_13_390 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_55_257 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ right_width_0_height_0__pin_3_ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ vgnd vpwr scs8hd_or2_1
XFILLER_23_121 vgnd vpwr scs8hd_fill_1
XFILLER_11_349 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_46_202 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_257 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_110 vpwr vgnd scs8hd_fill_2
XFILLER_14_121 vpwr vgnd scs8hd_fill_2
XFILLER_14_154 vpwr vgnd scs8hd_fill_2
XFILLER_10_382 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_6_364 vgnd vpwr scs8hd_decap_6
XFILLER_37_235 vgnd vpwr scs8hd_decap_3
XFILLER_37_213 vpwr vgnd scs8hd_fill_2
X_35_ _35_/HI _35_/LO vgnd vpwr scs8hd_conb_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_227 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_20_168 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XFILLER_57_39 vgnd vpwr scs8hd_decap_12
XFILLER_28_213 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_425 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_238 vgnd vpwr scs8hd_decap_4
XPHY_414 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_403 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_469 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_458 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_447 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_436 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_301 vpwr vgnd scs8hd_fill_2
XFILLER_3_367 vgnd vpwr scs8hd_decap_12
XFILLER_6_150 vgnd vpwr scs8hd_decap_3
XFILLER_6_172 vgnd vpwr scs8hd_decap_3
XFILLER_6_194 vgnd vpwr scs8hd_decap_4
XFILLER_8_55 vpwr vgnd scs8hd_fill_2
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_0_337 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_396 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_31_208 vgnd vpwr scs8hd_decap_12
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_53 vpwr vgnd scs8hd_fill_2
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_33_74 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XPHY_299 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_288 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_120 vpwr vgnd scs8hd_fill_2
XFILLER_39_319 vpwr vgnd scs8hd_fill_2
XFILLER_3_175 vpwr vgnd scs8hd_fill_2
XFILLER_3_131 vgnd vpwr scs8hd_decap_4
XFILLER_62_300 vgnd vpwr scs8hd_decap_12
XFILLER_58_93 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_30_296 vgnd vpwr scs8hd_decap_3
XFILLER_30_274 vgnd vpwr scs8hd_fill_1
XFILLER_30_263 vgnd vpwr scs8hd_decap_4
XFILLER_15_293 vpwr vgnd scs8hd_fill_2
XFILLER_15_271 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_344 vgnd vpwr scs8hd_fill_1
XFILLER_53_300 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_105 vgnd vpwr scs8hd_decap_12
XFILLER_44_322 vgnd vpwr scs8hd_decap_8
XFILLER_44_300 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_8_201 vgnd vpwr scs8hd_decap_12
XFILLER_8_223 vgnd vpwr scs8hd_decap_3
XFILLER_5_78 vgnd vpwr scs8hd_fill_1
XFILLER_8_267 vpwr vgnd scs8hd_fill_2
XFILLER_8_289 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_141 vgnd vpwr scs8hd_decap_12
XFILLER_47_171 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
+ bottom_width_0_height_0__pin_31_ vgnd vpwr scs8hd_diode_2
XFILLER_50_369 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _34_/HI vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_196 vgnd vpwr scs8hd_decap_12
XFILLER_41_358 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_32 vgnd vpwr scs8hd_decap_12
XFILLER_14_76 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_62 vgnd vpwr scs8hd_decap_12
XFILLER_39_51 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_44_141 vgnd vpwr scs8hd_decap_12
XFILLER_32_325 vgnd vpwr scs8hd_decap_8
XFILLER_29_171 vgnd vpwr scs8hd_decap_12
XFILLER_17_377 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_55_406 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_166 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_196 vgnd vpwr scs8hd_decap_8
XFILLER_31_380 vpwr vgnd scs8hd_fill_2
XFILLER_46_406 vgnd vpwr scs8hd_fill_1
XFILLER_58_288 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_152 vgnd vpwr scs8hd_fill_1
XFILLER_26_130 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
+ right_width_0_height_0__pin_6_ vgnd vpwr scs8hd_diode_2
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_97 vgnd vpwr scs8hd_decap_3
XPHY_86 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_369 vgnd vpwr scs8hd_fill_1
XFILLER_14_358 vgnd vpwr scs8hd_decap_8
XFILLER_1_240 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_1_273 vpwr vgnd scs8hd_fill_2
X_51_ _51_/HI _51_/LO vgnd vpwr scs8hd_conb_1
XFILLER_32_166 vgnd vpwr scs8hd_decap_12
XFILLER_20_317 vpwr vgnd scs8hd_fill_2
XFILLER_17_174 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_28_406 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_55_269 vgnd vpwr scs8hd_decap_12
XFILLER_11_306 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_133 vgnd vpwr scs8hd_decap_8
XFILLER_14_188 vgnd vpwr scs8hd_decap_4
XFILLER_10_394 vgnd vpwr scs8hd_decap_3
XFILLER_6_398 vgnd vpwr scs8hd_decap_8
XFILLER_52_239 vgnd vpwr scs8hd_decap_12
XFILLER_37_258 vpwr vgnd scs8hd_fill_2
X_34_ _34_/HI _34_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
+ bottom_width_0_height_0__pin_22_ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_buf_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_20_158 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_247 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_459 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_448 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_437 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_426 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_415 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XPHY_404 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_114 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_32 vgnd vpwr scs8hd_decap_12
XFILLER_7_107 vgnd vpwr scs8hd_decap_4
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_0_3 vgnd vpwr scs8hd_decap_4
XFILLER_3_379 vgnd vpwr scs8hd_decap_12
XFILLER_47_62 vgnd vpwr scs8hd_decap_12
XFILLER_47_51 vgnd vpwr scs8hd_decap_8
XFILLER_19_203 vpwr vgnd scs8hd_fill_2
XFILLER_42_283 vpwr vgnd scs8hd_fill_2
XFILLER_8_23 vpwr vgnd scs8hd_fill_2
XFILLER_8_78 vpwr vgnd scs8hd_fill_2
XFILLER_10_191 vgnd vpwr scs8hd_decap_4
XFILLER_33_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
+ clkbuf_1_1__f_clk/X ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ bottom_width_0_height_0__pin_50_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en vgnd vpwr scs8hd_sdfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_86 vgnd vpwr scs8hd_decap_12
XFILLER_24_272 vgnd vpwr scs8hd_fill_1
XPHY_289 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_47_331 vpwr vgnd scs8hd_fill_2
XFILLER_62_312 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_323 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_117 vgnd vpwr scs8hd_decap_12
XFILLER_0_179 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_29_386 vpwr vgnd scs8hd_fill_2
XFILLER_8_213 vgnd vpwr scs8hd_fill_1
XFILLER_12_253 vgnd vpwr scs8hd_decap_3
XFILLER_5_24 vpwr vgnd scs8hd_fill_2
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XFILLER_35_301 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_326 vgnd vpwr scs8hd_decap_8
XFILLER_35_334 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_315 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_26_356 vpwr vgnd scs8hd_fill_2
XFILLER_26_323 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_14_44 vgnd vpwr scs8hd_decap_12
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_74 vgnd vpwr scs8hd_decap_12
XFILLER_17_301 vpwr vgnd scs8hd_fill_2
XFILLER_55_62 vgnd vpwr scs8hd_decap_12
XFILLER_55_51 vgnd vpwr scs8hd_decap_8
XFILLER_32_348 vpwr vgnd scs8hd_fill_2
XFILLER_32_337 vgnd vpwr scs8hd_decap_4
XFILLER_17_367 vgnd vpwr scs8hd_decap_4
XFILLER_40_381 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_178 vgnd vpwr scs8hd_decap_12
XFILLER_23_359 vgnd vpwr scs8hd_decap_4
XFILLER_23_315 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_98 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_decap_3
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XFILLER_14_337 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_1__f_clk/X vgnd vpwr scs8hd_diode_2
XFILLER_49_245 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_17_153 vpwr vgnd scs8hd_fill_2
XFILLER_17_142 vgnd vpwr scs8hd_decap_6
XFILLER_1_296 vpwr vgnd scs8hd_fill_2
X_50_ _50_/HI _50_/LO vgnd vpwr scs8hd_conb_1
XFILLER_32_178 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XFILLER_63_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_63_281 vgnd vpwr scs8hd_decap_12
XFILLER_23_123 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
+ right_width_0_height_0__pin_0_ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_0__f_clk/X vgnd vpwr scs8hd_diode_2
XFILLER_11_23 vgnd vpwr scs8hd_decap_3
XFILLER_11_318 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _38_/HI vgnd vpwr scs8hd_diode_2
XFILLER_46_215 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_ _44_/HI
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ bottom_width_0_height_0__pin_47_lower vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_145 vgnd vpwr scs8hd_decap_8
XFILLER_37_204 vgnd vpwr scs8hd_decap_3
X_33_ _33_/HI _33_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
+ bottom_width_0_height_0__pin_21_ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_60_251 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_160 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_215 vgnd vpwr scs8hd_decap_6
XPHY_449 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_438 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_427 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_416 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_405 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_159 vpwr vgnd scs8hd_fill_2
XFILLER_59_362 vpwr vgnd scs8hd_fill_2
XFILLER_63_51 vgnd vpwr scs8hd_decap_8
XFILLER_47_74 vgnd vpwr scs8hd_decap_12
XFILLER_19_259 vgnd vpwr scs8hd_fill_1
XFILLER_63_62 vgnd vpwr scs8hd_decap_12
XFILLER_6_163 vgnd vpwr scs8hd_decap_3
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
XFILLER_33_295 vgnd vpwr scs8hd_fill_1
XFILLER_33_240 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_306 vpwr vgnd scs8hd_fill_2
XFILLER_56_398 vgnd vpwr scs8hd_decap_8
XFILLER_16_207 vpwr vgnd scs8hd_fill_2
XFILLER_33_98 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_262 vpwr vgnd scs8hd_fill_2
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_406 vgnd vpwr scs8hd_fill_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_100 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_62_324 vgnd vpwr scs8hd_decap_12
XFILLER_47_387 vgnd vpwr scs8hd_decap_12
XFILLER_30_276 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_398 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_221 vgnd vpwr scs8hd_decap_12
XFILLER_48_129 vgnd vpwr scs8hd_decap_12
XFILLER_29_343 vpwr vgnd scs8hd_fill_2
XFILLER_28_32 vgnd vpwr scs8hd_decap_12
Xclkbuf_1_1__f_clk clkbuf_0_clk/X clkbuf_1_1__f_clk/X vgnd vpwr scs8hd_clkbuf_16
XFILLER_0_125 vgnd vpwr scs8hd_decap_3
XFILLER_0_147 vpwr vgnd scs8hd_fill_2
XFILLER_28_76 vgnd vpwr scs8hd_decap_12
XFILLER_12_210 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _48_/HI vgnd vpwr scs8hd_diode_2
XFILLER_8_247 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_36 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_47_184 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_62_154 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_357 vgnd vpwr scs8hd_decap_4
XFILLER_53_110 vgnd vpwr scs8hd_decap_12
XFILLER_26_346 vpwr vgnd scs8hd_fill_2
XFILLER_26_335 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_5_217 vpwr vgnd scs8hd_fill_2
XFILLER_14_56 vpwr vgnd scs8hd_fill_2
XFILLER_30_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_86 vgnd vpwr scs8hd_decap_12
XFILLER_29_184 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_74 vgnd vpwr scs8hd_decap_12
XFILLER_44_154 vgnd vpwr scs8hd_decap_12
XFILLER_40_360 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_40_393 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_261 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_35_110 vgnd vpwr scs8hd_decap_12
XFILLER_23_338 vgnd vpwr scs8hd_decap_3
XFILLER_31_393 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_209 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_58_202 vgnd vpwr scs8hd_decap_12
XPHY_99 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XPHY_88 vgnd vpwr scs8hd_decap_3
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_154 vgnd vpwr scs8hd_decap_12
XFILLER_22_360 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
+ bottom_width_0_height_0__pin_28_ vgnd vpwr scs8hd_diode_2
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XFILLER_14_327 vgnd vpwr scs8hd_decap_8
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
XFILLER_22_382 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_257 vgnd vpwr scs8hd_decap_12
XFILLER_1_264 vgnd vpwr scs8hd_decap_3
XFILLER_64_249 vgnd vpwr scs8hd_decap_12
XFILLER_57_290 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_40_190 vgnd vpwr scs8hd_decap_12
XFILLER_20_308 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_9_397 vgnd vpwr scs8hd_decap_8
XFILLER_63_293 vgnd vpwr scs8hd_decap_12
XFILLER_48_290 vpwr vgnd scs8hd_fill_2
XFILLER_23_135 vgnd vpwr scs8hd_decap_12
XFILLER_23_113 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_61_208 vgnd vpwr scs8hd_decap_12
XFILLER_46_227 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_10_341 vgnd vpwr scs8hd_fill_1
XFILLER_6_312 vpwr vgnd scs8hd_fill_2
XFILLER_6_334 vpwr vgnd scs8hd_fill_2
X_32_ _32_/HI _32_/LO vgnd vpwr scs8hd_conb_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
+ bottom_width_0_height_0__pin_20_ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_60_263 vgnd vpwr scs8hd_decap_12
XFILLER_33_400 vgnd vpwr scs8hd_decap_6
XFILLER_20_105 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_20_138 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_208 vgnd vpwr scs8hd_fill_1
XPHY_439 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_428 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_417 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_406 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_359 vpwr vgnd scs8hd_fill_2
XFILLER_63_74 vgnd vpwr scs8hd_decap_12
XFILLER_47_86 vgnd vpwr scs8hd_decap_12
XFILLER_42_263 vpwr vgnd scs8hd_fill_2
XFILLER_19_249 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_142 vpwr vgnd scs8hd_fill_2
XFILLER_25_208 vgnd vpwr scs8hd_decap_12
XFILLER_19_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_403 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_24_285 vpwr vgnd scs8hd_fill_2
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _42_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_3_112 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_171 vgnd vpwr scs8hd_decap_12
XFILLER_47_377 vpwr vgnd scs8hd_fill_2
XFILLER_47_399 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _59_/HI vgnd vpwr scs8hd_diode_2
XFILLER_15_285 vpwr vgnd scs8hd_fill_2
XFILLER_15_263 vgnd vpwr scs8hd_decap_4
XFILLER_30_288 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_322 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_ _53_/HI
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ right_width_0_height_0__pin_34_lower vgnd vpwr scs8hd_mux2_1
XFILLER_53_358 vpwr vgnd scs8hd_fill_2
XFILLER_53_347 vgnd vpwr scs8hd_decap_4
XFILLER_38_366 vgnd vpwr scs8hd_fill_1
XFILLER_21_299 vpwr vgnd scs8hd_fill_2
XFILLER_21_233 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_90 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_0_104 vpwr vgnd scs8hd_fill_2
XFILLER_56_141 vgnd vpwr scs8hd_decap_12
XFILLER_28_88 vgnd vpwr scs8hd_decap_4
XFILLER_28_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_32 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_215 vgnd vpwr scs8hd_decap_8
XFILLER_5_48 vpwr vgnd scs8hd_fill_2
XFILLER_62_166 vgnd vpwr scs8hd_decap_12
XFILLER_47_196 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
+ right_width_0_height_0__pin_10_ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_50_317 vgnd vpwr scs8hd_decap_4
XFILLER_43_380 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_406 vgnd vpwr scs8hd_fill_1
XFILLER_38_141 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_41_306 vgnd vpwr scs8hd_decap_3
XFILLER_26_369 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_30_56 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_49_406 vgnd vpwr scs8hd_fill_1
XFILLER_55_86 vgnd vpwr scs8hd_decap_12
XFILLER_39_98 vgnd vpwr scs8hd_decap_12
XFILLER_17_325 vgnd vpwr scs8hd_decap_12
XFILLER_44_166 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_32_306 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_284 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_295 vpwr vgnd scs8hd_fill_2
XFILLER_23_306 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_80 vgnd vpwr scs8hd_decap_12
XPHY_12 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_decap_3
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_26_166 vgnd vpwr scs8hd_decap_12
XFILLER_22_394 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_23 vgnd vpwr scs8hd_decap_3
XFILLER_14_306 vpwr vgnd scs8hd_fill_2
XFILLER_49_269 vgnd vpwr scs8hd_decap_12
XFILLER_2_49 vpwr vgnd scs8hd_fill_2
XFILLER_2_27 vpwr vgnd scs8hd_fill_2
XFILLER_1_221 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_188 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_13_361 vgnd vpwr scs8hd_decap_3
XFILLER_9_321 vgnd vpwr scs8hd_decap_8
XFILLER_49_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_147 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_103 vgnd vpwr scs8hd_fill_1
XFILLER_14_125 vpwr vgnd scs8hd_fill_2
XFILLER_52_32 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
+ clkbuf_1_0__f_clk/X ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en vgnd vpwr scs8hd_sdfxbp_1
XFILLER_6_324 vpwr vgnd scs8hd_fill_2
XFILLER_10_386 vgnd vpwr scs8hd_decap_8
XFILLER_14_158 vpwr vgnd scs8hd_fill_2
XFILLER_37_217 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XFILLER_51_220 vgnd vpwr scs8hd_decap_12
XPHY_407 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_36_261 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_297 vpwr vgnd scs8hd_fill_2
XPHY_429 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_418 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_46 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_349 vpwr vgnd scs8hd_fill_2
XFILLER_59_386 vpwr vgnd scs8hd_fill_2
XFILLER_47_98 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_86 vgnd vpwr scs8hd_decap_12
XFILLER_42_242 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_90 vpwr vgnd scs8hd_fill_2
XFILLER_6_198 vgnd vpwr scs8hd_fill_1
XFILLER_33_264 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_157 vpwr vgnd scs8hd_fill_2
XFILLER_3_135 vgnd vpwr scs8hd_fill_1
XFILLER_62_337 vgnd vpwr scs8hd_decap_12
XFILLER_47_367 vgnd vpwr scs8hd_decap_4
XFILLER_47_323 vgnd vpwr scs8hd_decap_6
XFILLER_47_301 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_267 vgnd vpwr scs8hd_fill_1
XFILLER_15_297 vpwr vgnd scs8hd_fill_2
XFILLER_15_275 vgnd vpwr scs8hd_decap_4
XFILLER_15_242 vpwr vgnd scs8hd_fill_2
XFILLER_38_334 vpwr vgnd scs8hd_fill_2
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
XFILLER_61_381 vgnd vpwr scs8hd_decap_12
XFILLER_53_304 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_389 vgnd vpwr scs8hd_decap_8
XFILLER_0_116 vpwr vgnd scs8hd_fill_2
XFILLER_44_337 vgnd vpwr scs8hd_decap_3
XFILLER_28_56 vgnd vpwr scs8hd_decap_12
XFILLER_52_381 vgnd vpwr scs8hd_decap_12
XFILLER_44_359 vpwr vgnd scs8hd_fill_2
XFILLER_44_44 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_234 vgnd vpwr scs8hd_decap_12
XFILLER_12_267 vgnd vpwr scs8hd_decap_6
XFILLER_60_32 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
+ right_width_0_height_0__pin_9_ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_62_178 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_123 vgnd vpwr scs8hd_decap_12
XFILLER_26_315 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
+ bottom_width_0_height_0__pin_25_ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_30_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_98 vgnd vpwr scs8hd_decap_12
XFILLER_44_178 vgnd vpwr scs8hd_decap_12
XFILLER_17_337 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _46_/HI vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_ _42_/HI
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XFILLER_25_381 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_4_274 vgnd vpwr scs8hd_fill_1
XFILLER_35_123 vgnd vpwr scs8hd_decap_12
XFILLER_31_362 vpwr vgnd scs8hd_fill_2
XFILLER_31_351 vgnd vpwr scs8hd_fill_1
XFILLER_58_215 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_178 vgnd vpwr scs8hd_decap_12
XFILLER_26_134 vgnd vpwr scs8hd_decap_12
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XFILLER_41_159 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_3 vgnd vpwr scs8hd_decap_8
XFILLER_64_218 vgnd vpwr scs8hd_decap_12
XFILLER_57_281 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_1__f_clk/X vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_17_112 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_178 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_340 vpwr vgnd scs8hd_fill_2
XFILLER_9_333 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_ _54_/HI
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XFILLER_23_159 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_0__f_clk/X vgnd vpwr scs8hd_diode_2
XFILLER_11_15 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_54_251 vgnd vpwr scs8hd_decap_12
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_44 vgnd vpwr scs8hd_decap_12
XFILLER_10_321 vgnd vpwr scs8hd_decap_4
XFILLER_10_365 vpwr vgnd scs8hd_fill_2
XFILLER_10_398 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_60_276 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_9_152 vpwr vgnd scs8hd_fill_2
XFILLER_13_181 vpwr vgnd scs8hd_fill_2
XFILLER_61_3 vgnd vpwr scs8hd_decap_12
XFILLER_5_391 vgnd vpwr scs8hd_decap_12
XFILLER_28_207 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_3_71 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_232 vgnd vpwr scs8hd_decap_12
XPHY_419 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_408 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_36_251 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_118 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_310 vpwr vgnd scs8hd_fill_2
XFILLER_3_306 vpwr vgnd scs8hd_fill_2
XFILLER_3_317 vpwr vgnd scs8hd_fill_2
XFILLER_59_398 vpwr vgnd scs8hd_fill_2
XFILLER_27_240 vpwr vgnd scs8hd_fill_2
XFILLER_19_207 vpwr vgnd scs8hd_fill_2
XFILLER_63_98 vgnd vpwr scs8hd_decap_12
XFILLER_42_287 vgnd vpwr scs8hd_decap_4
XFILLER_42_276 vgnd vpwr scs8hd_decap_3
XFILLER_42_210 vgnd vpwr scs8hd_fill_1
XFILLER_27_284 vpwr vgnd scs8hd_fill_2
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
XFILLER_6_177 vpwr vgnd scs8hd_fill_2
XFILLER_10_173 vgnd vpwr scs8hd_decap_3
XFILLER_2_372 vpwr vgnd scs8hd_fill_2
XFILLER_33_221 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_295 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_33_298 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_346 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_210 vgnd vpwr scs8hd_decap_4
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_58_32 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
+ bottom_width_0_height_0__pin_19_ vgnd vpwr scs8hd_diode_2
XFILLER_62_349 vgnd vpwr scs8hd_decap_12
XFILLER_59_184 vgnd vpwr scs8hd_decap_12
XFILLER_47_335 vpwr vgnd scs8hd_fill_2
XFILLER_15_210 vpwr vgnd scs8hd_fill_2
XFILLER_30_202 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_357 vpwr vgnd scs8hd_fill_2
XFILLER_24_3 vgnd vpwr scs8hd_decap_12
XFILLER_61_393 vgnd vpwr scs8hd_decap_12
XFILLER_53_327 vpwr vgnd scs8hd_fill_2
XFILLER_0_72 vpwr vgnd scs8hd_fill_2
XFILLER_0_94 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_81 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_154 vgnd vpwr scs8hd_decap_12
XFILLER_28_68 vgnd vpwr scs8hd_decap_6
XFILLER_60_44 vgnd vpwr scs8hd_decap_12
XFILLER_52_393 vgnd vpwr scs8hd_decap_4
XFILLER_44_56 vgnd vpwr scs8hd_decap_12
XFILLER_12_246 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_110 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
+ right_width_0_height_0__pin_8_ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_283 vpwr vgnd scs8hd_fill_2
XFILLER_53_135 vgnd vpwr scs8hd_decap_12
XFILLER_38_154 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_382 vgnd vpwr scs8hd_decap_12
XFILLER_14_15 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_1_404 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_110 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_25_393 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_17_349 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_52_190 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_135 vgnd vpwr scs8hd_decap_12
XFILLER_50_105 vgnd vpwr scs8hd_decap_12
XFILLER_31_330 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_58_227 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_146 vgnd vpwr scs8hd_decap_6
XFILLER_26_102 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_190 vgnd vpwr scs8hd_decap_12
XFILLER_1_234 vgnd vpwr scs8hd_decap_4
XFILLER_32_105 vgnd vpwr scs8hd_decap_12
XFILLER_17_157 vpwr vgnd scs8hd_fill_2
XFILLER_9_301 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_356 vpwr vgnd scs8hd_fill_2
XFILLER_9_367 vgnd vpwr scs8hd_decap_4
XFILLER_55_208 vgnd vpwr scs8hd_decap_12
XFILLER_31_171 vgnd vpwr scs8hd_decap_12
XFILLER_16_190 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XFILLER_54_263 vgnd vpwr scs8hd_decap_12
XFILLER_52_56 vgnd vpwr scs8hd_decap_12
XFILLER_36_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_10_344 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _50_/HI vgnd vpwr scs8hd_diode_2
XFILLER_45_252 vpwr vgnd scs8hd_fill_2
XFILLER_45_241 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_60_288 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_175 vpwr vgnd scs8hd_fill_2
XFILLER_54_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XPHY_409 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_15 vgnd vpwr scs8hd_decap_12
XFILLER_59_333 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _33_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_406 vgnd vpwr scs8hd_fill_1
XFILLER_6_101 vpwr vgnd scs8hd_fill_2
XFILLER_10_152 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_ top_width_0_height_0__pin_32_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_33_233 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_17_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_24_266 vgnd vpwr scs8hd_decap_6
XFILLER_24_233 vgnd vpwr scs8hd_decap_3
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_406 vgnd vpwr scs8hd_fill_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_3_104 vpwr vgnd scs8hd_fill_2
XFILLER_59_196 vgnd vpwr scs8hd_decap_12
XFILLER_58_44 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
+ clkbuf_1_1__f_clk/X ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 Test_en
+ vgnd vpwr scs8hd_sdfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_ _33_/HI
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ right_width_0_height_0__pin_40_lower vgnd vpwr scs8hd_mux2_1
XFILLER_15_255 vpwr vgnd scs8hd_fill_2
XFILLER_23_91 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_306 vpwr vgnd scs8hd_fill_2
XFILLER_38_369 vgnd vpwr scs8hd_fill_1
XFILLER_17_3 vgnd vpwr scs8hd_decap_12
XFILLER_0_51 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
+ bottom_width_0_height_0__pin_22_ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_303 vpwr vgnd scs8hd_fill_2
XFILLER_56_166 vgnd vpwr scs8hd_decap_12
XFILLER_44_68 vgnd vpwr scs8hd_decap_12
XFILLER_37_391 vgnd vpwr scs8hd_decap_12
XFILLER_29_358 vpwr vgnd scs8hd_fill_2
XFILLER_29_347 vpwr vgnd scs8hd_fill_2
XFILLER_12_203 vgnd vpwr scs8hd_fill_1
XFILLER_60_56 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_91 vgnd vpwr scs8hd_fill_1
XFILLER_7_240 vpwr vgnd scs8hd_fill_2
XFILLER_7_262 vpwr vgnd scs8hd_fill_2
XFILLER_53_147 vgnd vpwr scs8hd_decap_12
XFILLER_38_166 vgnd vpwr scs8hd_decap_12
XFILLER_26_328 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_34_394 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _43_/HI ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_mux2_1
XFILLER_14_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_40_353 vgnd vpwr scs8hd_decap_4
XFILLER_40_320 vgnd vpwr scs8hd_decap_12
XFILLER_32_309 vpwr vgnd scs8hd_fill_2
XFILLER_25_350 vpwr vgnd scs8hd_fill_2
XFILLER_40_364 vgnd vpwr scs8hd_decap_3
XFILLER_4_210 vgnd vpwr scs8hd_decap_4
XFILLER_4_221 vpwr vgnd scs8hd_fill_2
XFILLER_20_81 vgnd vpwr scs8hd_decap_8
XFILLER_4_265 vpwr vgnd scs8hd_fill_2
XFILLER_4_276 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_147 vgnd vpwr scs8hd_decap_12
XFILLER_50_117 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_6_72 vpwr vgnd scs8hd_fill_2
XFILLER_58_239 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
+ clkbuf_1_0__f_clk/X ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en vgnd vpwr scs8hd_sdfxbp_1
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_25_59 vpwr vgnd scs8hd_fill_2
XFILLER_25_15 vgnd vpwr scs8hd_decap_12
XPHY_48 vgnd vpwr scs8hd_decap_3
XFILLER_22_342 vpwr vgnd scs8hd_fill_2
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XFILLER_22_386 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_294 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_117 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_397 vgnd vpwr scs8hd_decap_8
XFILLER_13_386 vpwr vgnd scs8hd_fill_2
XFILLER_13_353 vpwr vgnd scs8hd_fill_2
XFILLER_63_220 vgnd vpwr scs8hd_decap_12
XFILLER_23_117 vgnd vpwr scs8hd_decap_4
XFILLER_11_28 vpwr vgnd scs8hd_fill_2
XFILLER_39_283 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_68 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_14_106 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_316 vpwr vgnd scs8hd_fill_2
XFILLER_37_209 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_45_297 vpwr vgnd scs8hd_fill_2
XFILLER_45_275 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_47_3 vgnd vpwr scs8hd_decap_12
XFILLER_51_289 vpwr vgnd scs8hd_fill_2
XFILLER_51_245 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_345 vpwr vgnd scs8hd_fill_2
XFILLER_59_301 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_9 vpwr vgnd scs8hd_fill_2
XFILLER_42_234 vgnd vpwr scs8hd_decap_8
XFILLER_27_297 vpwr vgnd scs8hd_fill_2
XFILLER_27_264 vgnd vpwr scs8hd_decap_12
XFILLER_15_404 vgnd vpwr scs8hd_decap_3
XFILLER_42_267 vgnd vpwr scs8hd_decap_6
XFILLER_10_142 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _59_/HI ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_2_341 vpwr vgnd scs8hd_fill_2
XFILLER_6_146 vpwr vgnd scs8hd_fill_2
XFILLER_6_168 vpwr vgnd scs8hd_fill_2
XFILLER_10_197 vgnd vpwr scs8hd_decap_3
XFILLER_12_82 vgnd vpwr scs8hd_decap_8
XFILLER_12_93 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_231 vgnd vpwr scs8hd_decap_12
XFILLER_2_396 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_190 vpwr vgnd scs8hd_fill_2
XFILLER_24_245 vpwr vgnd scs8hd_fill_2
XFILLER_17_27 vgnd vpwr scs8hd_decap_12
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_59 vpwr vgnd scs8hd_fill_2
XFILLER_33_15 vgnd vpwr scs8hd_decap_12
XFILLER_24_289 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ top_width_0_height_0__pin_32_ vgnd vpwr scs8hd_diode_2
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_3_127 vpwr vgnd scs8hd_fill_2
XFILLER_3_116 vpwr vgnd scs8hd_fill_2
XFILLER_58_56 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_47_348 vgnd vpwr scs8hd_decap_12
XFILLER_47_315 vpwr vgnd scs8hd_fill_2
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
XFILLER_15_289 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_buf_2
XFILLER_15_245 vgnd vpwr scs8hd_decap_8
XFILLER_15_234 vgnd vpwr scs8hd_decap_8
XFILLER_23_81 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_337 vgnd vpwr scs8hd_decap_12
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
XFILLER_21_237 vgnd vpwr scs8hd_fill_1
XFILLER_0_108 vpwr vgnd scs8hd_fill_2
XFILLER_29_315 vpwr vgnd scs8hd_fill_2
XFILLER_28_15 vgnd vpwr scs8hd_decap_12
XFILLER_56_178 vgnd vpwr scs8hd_decap_12
XFILLER_52_351 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_68 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _60_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_270 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_123 vgnd vpwr scs8hd_decap_12
XFILLER_28_381 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_560 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_362 vpwr vgnd scs8hd_fill_2
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
XFILLER_7_296 vpwr vgnd scs8hd_fill_2
XFILLER_11_270 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
+ bottom_width_0_height_0__pin_16_ vgnd vpwr scs8hd_diode_2
XFILLER_53_159 vgnd vpwr scs8hd_decap_12
XFILLER_38_178 vgnd vpwr scs8hd_decap_12
XFILLER_19_392 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_30_27 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_29_123 vgnd vpwr scs8hd_decap_12
XFILLER_40_332 vpwr vgnd scs8hd_fill_2
XFILLER_25_362 vpwr vgnd scs8hd_fill_2
XFILLER_40_398 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_93 vpwr vgnd scs8hd_fill_2
XFILLER_4_299 vpwr vgnd scs8hd_fill_2
XFILLER_50_129 vgnd vpwr scs8hd_decap_12
XFILLER_35_159 vgnd vpwr scs8hd_decap_12
XPHY_390 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_376 vpwr vgnd scs8hd_fill_2
XFILLER_31_343 vgnd vpwr scs8hd_decap_8
XFILLER_16_395 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ bottom_width_0_height_0__pin_23_ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/A
+ vgnd vpwr scs8hd_or2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_27 vgnd vpwr scs8hd_decap_12
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_22_321 vgnd vpwr scs8hd_decap_12
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XFILLER_22_398 vgnd vpwr scs8hd_decap_8
XFILLER_1_269 vpwr vgnd scs8hd_fill_2
XFILLER_32_129 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_71 vpwr vgnd scs8hd_fill_2
XFILLER_13_310 vgnd vpwr scs8hd_fill_1
XFILLER_48_251 vgnd vpwr scs8hd_decap_12
XFILLER_0_280 vgnd vpwr scs8hd_decap_3
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_63_232 vgnd vpwr scs8hd_decap_12
XFILLER_31_184 vgnd vpwr scs8hd_decap_12
XFILLER_8_380 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_276 vgnd vpwr scs8hd_decap_12
XFILLER_39_262 vpwr vgnd scs8hd_fill_2
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_14_129 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_3 vgnd vpwr scs8hd_decap_4
XFILLER_6_328 vgnd vpwr scs8hd_decap_4
XFILLER_60_202 vgnd vpwr scs8hd_decap_12
XFILLER_45_287 vgnd vpwr scs8hd_decap_3
XFILLER_45_221 vpwr vgnd scs8hd_fill_2
XFILLER_13_140 vpwr vgnd scs8hd_fill_2
XFILLER_42_80 vgnd vpwr scs8hd_decap_12
XFILLER_13_184 vpwr vgnd scs8hd_fill_2
XFILLER_3_52 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_36_276 vgnd vpwr scs8hd_decap_3
XFILLER_51_257 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_246 vpwr vgnd scs8hd_fill_2
XFILLER_42_213 vgnd vpwr scs8hd_fill_1
XFILLER_42_202 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_276 vgnd vpwr scs8hd_decap_6
XFILLER_27_232 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_290 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_6_125 vpwr vgnd scs8hd_fill_2
XFILLER_10_121 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XFILLER_18_265 vpwr vgnd scs8hd_fill_2
XFILLER_18_243 vgnd vpwr scs8hd_decap_3
XFILLER_41_290 vpwr vgnd scs8hd_fill_2
XFILLER_33_268 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_17_39 vgnd vpwr scs8hd_decap_12
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XFILLER_59_110 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_58_68 vgnd vpwr scs8hd_decap_12
XFILLER_30_227 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_38_349 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_28_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_44_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_105 vgnd vpwr scs8hd_decap_12
XFILLER_47_135 vgnd vpwr scs8hd_decap_12
XFILLER_28_393 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_561 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_550 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_50_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_319 vgnd vpwr scs8hd_decap_4
XFILLER_22_3 vgnd vpwr scs8hd_decap_12
XFILLER_61_171 vgnd vpwr scs8hd_decap_12
XFILLER_46_190 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_39_59 vpwr vgnd scs8hd_fill_2
XFILLER_39_15 vgnd vpwr scs8hd_decap_12
XFILLER_44_105 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_135 vgnd vpwr scs8hd_decap_12
XFILLER_4_234 vpwr vgnd scs8hd_fill_2
XFILLER_63_403 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_43_171 vgnd vpwr scs8hd_decap_12
XFILLER_28_190 vgnd vpwr scs8hd_decap_3
XFILLER_16_341 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XPHY_391 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_380 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_6_30 vgnd vpwr scs8hd_fill_1
XFILLER_6_41 vpwr vgnd scs8hd_fill_2
XFILLER_39_400 vgnd vpwr scs8hd_decap_6
XFILLER_19_190 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XFILLER_25_39 vgnd vpwr scs8hd_decap_12
XFILLER_22_355 vgnd vpwr scs8hd_decap_3
XFILLER_22_333 vgnd vpwr scs8hd_fill_1
XFILLER_22_311 vgnd vpwr scs8hd_fill_1
XPHY_39 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_49_208 vgnd vpwr scs8hd_decap_12
XFILLER_60_406 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_182 vgnd vpwr scs8hd_fill_1
XFILLER_40_141 vgnd vpwr scs8hd_decap_12
XANTENNA__71__A bottom_width_0_height_0__pin_49_lower vgnd vpwr scs8hd_diode_2
XFILLER_48_263 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_406 vgnd vpwr scs8hd_fill_1
XFILLER_23_108 vgnd vpwr scs8hd_decap_3
XFILLER_31_196 vgnd vpwr scs8hd_decap_12
XFILLER_39_241 vgnd vpwr scs8hd_decap_3
XFILLER_54_288 vgnd vpwr scs8hd_decap_12
XFILLER_52_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_406 vgnd vpwr scs8hd_fill_1
XFILLER_39_274 vpwr vgnd scs8hd_fill_2
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_10_314 vgnd vpwr scs8hd_decap_4
XFILLER_10_325 vgnd vpwr scs8hd_fill_1
XFILLER_10_369 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA__66__A bottom_width_0_height_0__pin_44_lower vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_406 vgnd vpwr scs8hd_fill_1
XFILLER_26_82 vgnd vpwr scs8hd_decap_8
XFILLER_9_123 vgnd vpwr scs8hd_decap_3
XFILLER_13_152 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_ _56_/HI
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ right_width_0_height_0__pin_37_lower vgnd vpwr scs8hd_mux2_1
XFILLER_9_156 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_1__f_clk/X vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_42 vgnd vpwr scs8hd_fill_1
XFILLER_36_255 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_406 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
+ clkbuf_1_0__f_clk/X ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 Test_en
+ vgnd vpwr scs8hd_sdfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_51_269 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _47_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_59_358 vpwr vgnd scs8hd_fill_2
XFILLER_47_59 vpwr vgnd scs8hd_fill_2
XFILLER_47_15 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
+ clkbuf_1_1__f_clk/X vgnd vpwr scs8hd_diode_2
XFILLER_12_62 vgnd vpwr scs8hd_fill_1
XFILLER_2_398 vgnd vpwr scs8hd_decap_8
XFILLER_2_376 vgnd vpwr scs8hd_decap_12
XFILLER_2_332 vpwr vgnd scs8hd_fill_2
XFILLER_33_236 vpwr vgnd scs8hd_fill_2
XFILLER_33_214 vgnd vpwr scs8hd_fill_1
XFILLER_18_299 vpwr vgnd scs8hd_fill_2
XFILLER_52_3 vgnd vpwr scs8hd_decap_12
XFILLER_56_328 vgnd vpwr scs8hd_decap_6
XFILLER_56_306 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_39 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
X_69_ bottom_width_0_height_0__pin_47_lower bottom_width_0_height_0__pin_47_upper
+ vgnd vpwr scs8hd_buf_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_280 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_ _45_/HI
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ bottom_width_0_height_0__pin_46_lower vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_/QN
+ vgnd vpwr scs8hd_dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_30_239 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _49_/HI vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_140 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_80 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
+ right_width_0_height_0__pin_13_ vgnd vpwr scs8hd_diode_2
XFILLER_2_173 vpwr vgnd scs8hd_fill_2
XFILLER_46_394 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_0_76 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_85 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_180 vgnd vpwr scs8hd_decap_6
XFILLER_60_15 vgnd vpwr scs8hd_decap_12
XFILLER_44_27 vgnd vpwr scs8hd_decap_4
XFILLER_12_206 vpwr vgnd scs8hd_fill_2
XFILLER_62_117 vgnd vpwr scs8hd_decap_12
XANTENNA__74__A right_width_0_height_0__pin_35_lower vgnd vpwr scs8hd_diode_2
XFILLER_47_147 vgnd vpwr scs8hd_decap_12
XFILLER_43_342 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
+ clkbuf_1_0__f_clk/X ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en vgnd vpwr scs8hd_sdfxbp_1
XPHY_562 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_551 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_540 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_254 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_372 vgnd vpwr scs8hd_fill_1
XFILLER_15_3 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_39_27 vgnd vpwr scs8hd_decap_12
XFILLER_55_59 vpwr vgnd scs8hd_fill_2
XFILLER_55_15 vgnd vpwr scs8hd_decap_12
XFILLER_44_117 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_147 vgnd vpwr scs8hd_decap_12
XFILLER_40_345 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_73 vpwr vgnd scs8hd_fill_2
XANTENNA__69__A bottom_width_0_height_0__pin_47_lower vgnd vpwr scs8hd_diode_2
XFILLER_4_202 vgnd vpwr scs8hd_fill_1
XPHY_370 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_375 vgnd vpwr scs8hd_decap_12
XFILLER_16_353 vgnd vpwr scs8hd_decap_12
XFILLER_16_331 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XPHY_392 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_381 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_389 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_97 vpwr vgnd scs8hd_fill_2
XPHY_29 vgnd vpwr scs8hd_decap_3
XPHY_18 vgnd vpwr scs8hd_decap_3
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_57_220 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_51 vgnd vpwr scs8hd_decap_4
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_0_271 vpwr vgnd scs8hd_fill_2
XFILLER_63_245 vgnd vpwr scs8hd_decap_12
XFILLER_56_80 vgnd vpwr scs8hd_decap_12
XFILLER_16_183 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_231 vgnd vpwr scs8hd_decap_4
XFILLER_27_404 vgnd vpwr scs8hd_decap_3
XFILLER_52_27 vgnd vpwr scs8hd_decap_4
XFILLER_39_297 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_22_175 vgnd vpwr scs8hd_decap_6
XFILLER_10_337 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_245 vgnd vpwr scs8hd_decap_4
XFILLER_45_234 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XFILLER_60_215 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_113 vpwr vgnd scs8hd_fill_2
XFILLER_13_175 vgnd vpwr scs8hd_decap_4
XFILLER_42_93 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_341 vpwr vgnd scs8hd_fill_2
XFILLER_5_352 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_168 vgnd vpwr scs8hd_fill_1
XFILLER_9_179 vpwr vgnd scs8hd_fill_2
XFILLER_36_267 vgnd vpwr scs8hd_decap_6
XFILLER_36_234 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
+ right_width_0_height_0__pin_7_ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_337 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_15 vgnd vpwr scs8hd_decap_12
XFILLER_47_27 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_59 vpwr vgnd scs8hd_fill_2
XFILLER_42_259 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_10_178 vpwr vgnd scs8hd_fill_2
XANTENNA__77__A right_width_0_height_0__pin_38_lower vgnd vpwr scs8hd_diode_2
XFILLER_2_388 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ right_width_0_height_0__pin_11_ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_/X
+ vgnd vpwr scs8hd_or2_1
XFILLER_45_3 vgnd vpwr scs8hd_decap_12
X_68_ bottom_width_0_height_0__pin_46_lower bottom_width_0_height_0__pin_46_upper
+ vgnd vpwr scs8hd_buf_2
XFILLER_64_373 vgnd vpwr scs8hd_decap_12
XFILLER_24_215 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_59_123 vgnd vpwr scs8hd_decap_12
XFILLER_58_15 vgnd vpwr scs8hd_decap_12
XFILLER_55_362 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
XFILLER_15_259 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_95 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_152 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_/X
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_365 vgnd vpwr scs8hd_fill_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_0_55 vpwr vgnd scs8hd_fill_2
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_37_362 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_60_27 vgnd vpwr scs8hd_decap_4
XFILLER_52_398 vgnd vpwr scs8hd_decap_8
XFILLER_20_262 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ccff_tail
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_4_406 vgnd vpwr scs8hd_fill_1
XFILLER_47_159 vgnd vpwr scs8hd_decap_12
XPHY_552 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_541 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_62_129 vgnd vpwr scs8hd_decap_12
XPHY_530 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_43_387 vgnd vpwr scs8hd_decap_12
XFILLER_43_376 vpwr vgnd scs8hd_fill_2
XFILLER_43_310 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XPHY_563 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_50_93 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_266 vpwr vgnd scs8hd_fill_2
XFILLER_19_362 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_61_184 vgnd vpwr scs8hd_decap_12
XFILLER_34_398 vgnd vpwr scs8hd_decap_8
XFILLER_34_365 vpwr vgnd scs8hd_fill_2
XFILLER_39_39 vgnd vpwr scs8hd_decap_12
XFILLER_29_159 vgnd vpwr scs8hd_decap_12
XFILLER_55_27 vgnd vpwr scs8hd_decap_12
XFILLER_44_129 vgnd vpwr scs8hd_decap_12
XFILLER_25_332 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_357 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_4_269 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _44_/HI vgnd vpwr scs8hd_diode_2
XFILLER_43_184 vgnd vpwr scs8hd_decap_12
XPHY_393 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_382 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_371 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_360 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_398 vgnd vpwr scs8hd_decap_8
XFILLER_16_387 vgnd vpwr scs8hd_decap_8
XFILLER_16_365 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_107 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_1_217 vpwr vgnd scs8hd_fill_2
XFILLER_57_298 vgnd vpwr scs8hd_fill_1
XFILLER_57_287 vgnd vpwr scs8hd_fill_1
XFILLER_57_232 vgnd vpwr scs8hd_decap_12
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_40_154 vgnd vpwr scs8hd_decap_12
XFILLER_25_184 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_13_313 vpwr vgnd scs8hd_fill_2
XFILLER_13_357 vpwr vgnd scs8hd_fill_2
XFILLER_31_62 vgnd vpwr scs8hd_decap_12
XFILLER_31_51 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_257 vgnd vpwr scs8hd_decap_12
XFILLER_48_276 vgnd vpwr scs8hd_decap_12
XFILLER_31_110 vgnd vpwr scs8hd_decap_12
XFILLER_16_151 vpwr vgnd scs8hd_fill_2
XFILLER_16_195 vpwr vgnd scs8hd_fill_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_54_202 vgnd vpwr scs8hd_decap_12
XFILLER_39_287 vgnd vpwr scs8hd_fill_1
XFILLER_39_210 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ vgnd vpwr scs8hd_mux2_1
XFILLER_22_154 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_227 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_13_132 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_22 vpwr vgnd scs8hd_fill_2
XFILLER_5_364 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_36_202 vgnd vpwr scs8hd_decap_12
XFILLER_3_77 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_27 vgnd vpwr scs8hd_decap_12
XFILLER_47_39 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_10_146 vgnd vpwr scs8hd_decap_6
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_2_345 vpwr vgnd scs8hd_fill_2
XFILLER_2_301 vgnd vpwr scs8hd_decap_4
XFILLER_5_3 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
+ right_width_0_height_0__pin_10_ vgnd vpwr scs8hd_diode_2
XFILLER_18_213 vgnd vpwr scs8hd_fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
+ Test_en vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XFILLER_5_194 vpwr vgnd scs8hd_fill_2
XFILLER_64_385 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
X_67_ bottom_width_0_height_0__pin_45_lower bottom_width_0_height_0__pin_45_upper
+ vgnd vpwr scs8hd_buf_2
XFILLER_32_271 vgnd vpwr scs8hd_fill_1
XFILLER_24_249 vpwr vgnd scs8hd_fill_2
XFILLER_17_290 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XFILLER_59_135 vgnd vpwr scs8hd_decap_12
XFILLER_58_27 vgnd vpwr scs8hd_decap_4
XFILLER_47_319 vpwr vgnd scs8hd_fill_2
XFILLER_55_341 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_buf_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_293 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
+ bottom_width_0_height_0__pin_30_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_/X
+ vgnd vpwr scs8hd_buf_2
XFILLER_7_404 vgnd vpwr scs8hd_decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 vgnd
+ vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_58_190 vgnd vpwr scs8hd_decap_12
XFILLER_48_93 vgnd vpwr scs8hd_decap_12
XFILLER_46_330 vgnd vpwr scs8hd_decap_4
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XFILLER_61_377 vpwr vgnd scs8hd_fill_2
XFILLER_0_89 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ vgnd vpwr scs8hd_diode_2
XFILLER_56_105 vgnd vpwr scs8hd_decap_12
XFILLER_29_319 vgnd vpwr scs8hd_decap_3
XFILLER_52_333 vgnd vpwr scs8hd_decap_3
XFILLER_52_300 vgnd vpwr scs8hd_decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_ prog_clk
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_564 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_553 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_542 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_531 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_520 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_55_171 vgnd vpwr scs8hd_decap_12
XFILLER_43_399 vgnd vpwr scs8hd_decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_223 vpwr vgnd scs8hd_fill_2
XFILLER_11_274 vpwr vgnd scs8hd_fill_2
XFILLER_38_105 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_196 vgnd vpwr scs8hd_decap_12
XFILLER_55_39 vgnd vpwr scs8hd_decap_12
XFILLER_52_141 vgnd vpwr scs8hd_decap_12
XFILLER_40_369 vgnd vpwr scs8hd_decap_3
XFILLER_37_171 vgnd vpwr scs8hd_decap_12
XFILLER_25_377 vpwr vgnd scs8hd_fill_2
XFILLER_25_311 vpwr vgnd scs8hd_fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_/D
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_215 vgnd vpwr scs8hd_decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_29_62 vgnd vpwr scs8hd_decap_12
XFILLER_29_51 vgnd vpwr scs8hd_decap_8
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_196 vgnd vpwr scs8hd_decap_12
XPHY_394 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_383 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_372 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_361 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_350 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_358 vpwr vgnd scs8hd_fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ vgnd vpwr scs8hd_buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_3_281 vgnd vpwr scs8hd_decap_4
XFILLER_6_22 vpwr vgnd scs8hd_fill_2
XFILLER_6_55 vpwr vgnd scs8hd_fill_2
XFILLER_54_406 vgnd vpwr scs8hd_fill_1
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
+ prog_clk vgnd vpwr scs8hd_diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_ _50_/HI
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X ccff_tail
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_mux2_1
XFILLER_34_141 vgnd vpwr scs8hd_decap_12
XFILLER_17_108 vpwr vgnd scs8hd_fill_2
XFILLER_40_166 vgnd vpwr scs8hd_decap_12
XFILLER_25_196 vgnd vpwr scs8hd_decap_12
XFILLER_21_391 vgnd vpwr scs8hd_decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_75 vpwr vgnd scs8hd_fill_2
XFILLER_9_329 vpwr vgnd scs8hd_fill_2
XFILLER_13_336 vpwr vgnd scs8hd_fill_2
XFILLER_31_74 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
+ clkbuf_1_0__f_clk/X ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_/QN
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 Test_en
+ vgnd vpwr scs8hd_sdfxbp_1
XFILLER_36_406 vgnd vpwr scs8hd_fill_1
XFILLER_63_269 vgnd vpwr scs8hd_decap_12
XFILLER_56_93 vgnd vpwr scs8hd_decap_12
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
+ prog_clk ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_/QN
+ vgnd vpwr scs8hd_dfxbp_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_362 vgnd vpwr scs8hd_decap_3
XFILLER_8_384 vpwr vgnd scs8hd_fill_2
.ends

