magic
tech sky130A
magscale 1 2
timestamp 1606931478
<< locali >>
rect 11253 19159 11287 19329
rect 15945 19159 15979 19261
rect 3341 18207 3375 18377
rect 3283 18173 3375 18207
rect 5089 18071 5123 18309
rect 12357 17833 12449 17867
rect 5641 17527 5675 17765
rect 12357 17527 12391 17833
rect 6377 16983 6411 17289
rect 10057 16099 10091 16201
rect 4905 15419 4939 15589
rect 9413 14807 9447 14977
rect 11989 13719 12023 13889
rect 10609 12699 10643 12869
rect 14381 12631 14415 12869
rect 4905 12087 4939 12189
rect 6285 10047 6319 10217
rect 12265 9503 12299 9673
rect 7297 8823 7331 8925
rect 11621 8891 11655 9129
rect 13277 8347 13311 8585
rect 14323 7497 14415 7531
rect 6653 7327 6687 7497
rect 11253 7191 11287 7361
rect 14381 7327 14415 7497
rect 9413 6817 9597 6851
rect 9413 6783 9447 6817
rect 11253 6171 11287 6273
rect 2789 4471 2823 4709
rect 8309 4471 8343 4641
rect 15025 4471 15059 4709
rect 8251 4437 8343 4471
rect 13093 3383 13127 3553
rect 2513 2907 2547 3145
rect 13277 3043 13311 3145
rect 13737 2363 13771 2533
<< viali >>
rect 4537 20009 4571 20043
rect 6561 20009 6595 20043
rect 9229 20009 9263 20043
rect 10701 20009 10735 20043
rect 12817 20009 12851 20043
rect 13369 20009 13403 20043
rect 14381 20009 14415 20043
rect 14933 20009 14967 20043
rect 15669 20009 15703 20043
rect 16221 20009 16255 20043
rect 17233 20009 17267 20043
rect 2513 19941 2547 19975
rect 10793 19941 10827 19975
rect 1685 19873 1719 19907
rect 2237 19873 2271 19907
rect 3065 19873 3099 19907
rect 4445 19873 4479 19907
rect 5448 19873 5482 19907
rect 7656 19873 7690 19907
rect 9045 19873 9079 19907
rect 9781 19873 9815 19907
rect 11345 19873 11379 19907
rect 11621 19873 11655 19907
rect 12633 19873 12667 19907
rect 13185 19873 13219 19907
rect 14197 19873 14231 19907
rect 14749 19873 14783 19907
rect 15485 19873 15519 19907
rect 16037 19873 16071 19907
rect 17049 19873 17083 19907
rect 3249 19805 3283 19839
rect 4721 19805 4755 19839
rect 5181 19805 5215 19839
rect 6929 19805 6963 19839
rect 7389 19805 7423 19839
rect 10977 19805 11011 19839
rect 12081 19805 12115 19839
rect 9965 19737 9999 19771
rect 1869 19669 1903 19703
rect 4077 19669 4111 19703
rect 8769 19669 8803 19703
rect 10333 19669 10367 19703
rect 6469 19465 6503 19499
rect 13829 19465 13863 19499
rect 7389 19329 7423 19363
rect 8033 19329 8067 19363
rect 11253 19329 11287 19363
rect 11897 19329 11931 19363
rect 1593 19261 1627 19295
rect 2145 19261 2179 19295
rect 2973 19261 3007 19295
rect 3240 19261 3274 19295
rect 5089 19261 5123 19295
rect 7297 19261 7331 19295
rect 9689 19261 9723 19295
rect 2421 19193 2455 19227
rect 4629 19193 4663 19227
rect 5356 19193 5390 19227
rect 8300 19193 8334 19227
rect 9956 19193 9990 19227
rect 11713 19261 11747 19295
rect 12449 19261 12483 19295
rect 14105 19261 14139 19295
rect 14933 19261 14967 19295
rect 15945 19261 15979 19295
rect 16037 19261 16071 19295
rect 16589 19261 16623 19295
rect 17141 19261 17175 19295
rect 18061 19261 18095 19295
rect 18613 19261 18647 19295
rect 19441 19261 19475 19295
rect 11805 19193 11839 19227
rect 12716 19193 12750 19227
rect 15577 19193 15611 19227
rect 1777 19125 1811 19159
rect 4353 19125 4387 19159
rect 6837 19125 6871 19159
rect 7205 19125 7239 19159
rect 9413 19125 9447 19159
rect 11069 19125 11103 19159
rect 11253 19125 11287 19159
rect 11345 19125 11379 19159
rect 14289 19125 14323 19159
rect 15945 19125 15979 19159
rect 16221 19125 16255 19159
rect 16773 19125 16807 19159
rect 17325 19125 17359 19159
rect 18245 19125 18279 19159
rect 18797 19125 18831 19159
rect 19625 19125 19659 19159
rect 2973 18921 3007 18955
rect 3341 18921 3375 18955
rect 3433 18921 3467 18955
rect 6561 18921 6595 18955
rect 7021 18921 7055 18955
rect 8861 18921 8895 18955
rect 13369 18921 13403 18955
rect 2421 18853 2455 18887
rect 4537 18853 4571 18887
rect 7748 18853 7782 18887
rect 13921 18853 13955 18887
rect 14657 18853 14691 18887
rect 15577 18853 15611 18887
rect 18797 18853 18831 18887
rect 1409 18785 1443 18819
rect 2329 18785 2363 18819
rect 4445 18785 4479 18819
rect 5448 18785 5482 18819
rect 6837 18785 6871 18819
rect 9137 18785 9171 18819
rect 10057 18785 10091 18819
rect 11345 18785 11379 18819
rect 11437 18785 11471 18819
rect 11989 18785 12023 18819
rect 12256 18785 12290 18819
rect 13645 18785 13679 18819
rect 14381 18785 14415 18819
rect 15301 18785 15335 18819
rect 18521 18785 18555 18819
rect 2605 18717 2639 18751
rect 3617 18717 3651 18751
rect 4721 18717 4755 18751
rect 5181 18717 5215 18751
rect 7481 18717 7515 18751
rect 10149 18717 10183 18751
rect 10241 18717 10275 18751
rect 11621 18717 11655 18751
rect 1593 18649 1627 18683
rect 4077 18649 4111 18683
rect 1961 18581 1995 18615
rect 9689 18581 9723 18615
rect 10977 18581 11011 18615
rect 3341 18377 3375 18411
rect 12449 18377 12483 18411
rect 13461 18377 13495 18411
rect 14657 18377 14691 18411
rect 1685 18309 1719 18343
rect 4905 18309 4939 18343
rect 5089 18309 5123 18343
rect 9045 18309 9079 18343
rect 1501 18173 1535 18207
rect 2053 18173 2087 18207
rect 2789 18173 2823 18207
rect 3249 18173 3283 18207
rect 3525 18173 3559 18207
rect 2329 18105 2363 18139
rect 3065 18105 3099 18139
rect 3792 18105 3826 18139
rect 5733 18241 5767 18275
rect 7481 18241 7515 18275
rect 8401 18241 8435 18275
rect 8585 18241 8619 18275
rect 9597 18241 9631 18275
rect 10241 18241 10275 18275
rect 11529 18241 11563 18275
rect 13001 18241 13035 18275
rect 14013 18241 14047 18275
rect 5641 18173 5675 18207
rect 6193 18173 6227 18207
rect 10057 18173 10091 18207
rect 11897 18173 11931 18207
rect 12817 18173 12851 18207
rect 14473 18173 14507 18207
rect 5549 18105 5583 18139
rect 9413 18105 9447 18139
rect 11345 18105 11379 18139
rect 13829 18105 13863 18139
rect 5089 18037 5123 18071
rect 5181 18037 5215 18071
rect 6377 18037 6411 18071
rect 6837 18037 6871 18071
rect 7205 18037 7239 18071
rect 7297 18037 7331 18071
rect 7941 18037 7975 18071
rect 8309 18037 8343 18071
rect 9505 18037 9539 18071
rect 10885 18037 10919 18071
rect 11253 18037 11287 18071
rect 12909 18037 12943 18071
rect 13921 18037 13955 18071
rect 3341 17833 3375 17867
rect 6469 17833 6503 17867
rect 9137 17833 9171 17867
rect 9689 17833 9723 17867
rect 12449 17833 12483 17867
rect 13921 17833 13955 17867
rect 14473 17833 14507 17867
rect 5641 17765 5675 17799
rect 6009 17765 6043 17799
rect 1501 17697 1535 17731
rect 2237 17697 2271 17731
rect 4077 17697 4111 17731
rect 4344 17697 4378 17731
rect 1685 17629 1719 17663
rect 2421 17629 2455 17663
rect 3433 17629 3467 17663
rect 3617 17629 3651 17663
rect 2973 17561 3007 17595
rect 5457 17561 5491 17595
rect 5733 17697 5767 17731
rect 6837 17697 6871 17731
rect 7748 17697 7782 17731
rect 10057 17697 10091 17731
rect 10149 17697 10183 17731
rect 10885 17697 10919 17731
rect 11152 17697 11186 17731
rect 6929 17629 6963 17663
rect 7021 17629 7055 17663
rect 7481 17629 7515 17663
rect 10333 17629 10367 17663
rect 8861 17561 8895 17595
rect 12808 17765 12842 17799
rect 14289 17697 14323 17731
rect 12541 17629 12575 17663
rect 5641 17493 5675 17527
rect 12265 17493 12299 17527
rect 12357 17493 12391 17527
rect 1777 17289 1811 17323
rect 4905 17289 4939 17323
rect 6377 17289 6411 17323
rect 8217 17289 8251 17323
rect 10057 17289 10091 17323
rect 11713 17289 11747 17323
rect 12449 17289 12483 17323
rect 13645 17289 13679 17323
rect 14197 17289 14231 17323
rect 4629 17221 4663 17255
rect 6101 17221 6135 17255
rect 3249 17153 3283 17187
rect 5365 17153 5399 17187
rect 5457 17153 5491 17187
rect 1593 17085 1627 17119
rect 2155 17085 2189 17119
rect 5917 17085 5951 17119
rect 2421 17017 2455 17051
rect 3516 17017 3550 17051
rect 13001 17153 13035 17187
rect 6653 17085 6687 17119
rect 6837 17085 6871 17119
rect 8677 17085 8711 17119
rect 8944 17085 8978 17119
rect 10333 17085 10367 17119
rect 10589 17085 10623 17119
rect 12173 17085 12207 17119
rect 13461 17085 13495 17119
rect 14013 17085 14047 17119
rect 7093 17017 7127 17051
rect 5273 16949 5307 16983
rect 6377 16949 6411 16983
rect 6469 16949 6503 16983
rect 11989 16949 12023 16983
rect 12817 16949 12851 16983
rect 12909 16949 12943 16983
rect 1869 16745 1903 16779
rect 3433 16745 3467 16779
rect 8125 16745 8159 16779
rect 9137 16745 9171 16779
rect 9965 16745 9999 16779
rect 10333 16745 10367 16779
rect 10977 16745 11011 16779
rect 2513 16677 2547 16711
rect 3341 16677 3375 16711
rect 11345 16677 11379 16711
rect 14565 16677 14599 16711
rect 1685 16609 1719 16643
rect 2237 16609 2271 16643
rect 4077 16609 4111 16643
rect 4629 16609 4663 16643
rect 4896 16609 4930 16643
rect 6285 16609 6319 16643
rect 6552 16609 6586 16643
rect 8493 16609 8527 16643
rect 8585 16609 8619 16643
rect 10425 16609 10459 16643
rect 11989 16609 12023 16643
rect 12633 16609 12667 16643
rect 12900 16609 12934 16643
rect 14289 16609 14323 16643
rect 3617 16541 3651 16575
rect 8677 16541 8711 16575
rect 10517 16541 10551 16575
rect 11437 16541 11471 16575
rect 11621 16541 11655 16575
rect 4261 16473 4295 16507
rect 7665 16473 7699 16507
rect 12173 16473 12207 16507
rect 2973 16405 3007 16439
rect 6009 16405 6043 16439
rect 14013 16405 14047 16439
rect 1961 16201 1995 16235
rect 2513 16201 2547 16235
rect 7941 16201 7975 16235
rect 10057 16201 10091 16235
rect 10149 16201 10183 16235
rect 2973 16133 3007 16167
rect 11161 16133 11195 16167
rect 3617 16065 3651 16099
rect 4629 16065 4663 16099
rect 5825 16065 5859 16099
rect 7481 16065 7515 16099
rect 8401 16065 8435 16099
rect 8585 16065 8619 16099
rect 9689 16065 9723 16099
rect 10057 16065 10091 16099
rect 10609 16065 10643 16099
rect 10793 16065 10827 16099
rect 11713 16065 11747 16099
rect 13277 16065 13311 16099
rect 13829 16065 13863 16099
rect 1777 15997 1811 16031
rect 2329 15997 2363 16031
rect 3433 15997 3467 16031
rect 5641 15997 5675 16031
rect 6218 15997 6252 16031
rect 7205 15997 7239 16031
rect 9505 15997 9539 16031
rect 11529 15997 11563 16031
rect 13645 15997 13679 16031
rect 4353 15929 4387 15963
rect 8309 15929 8343 15963
rect 10517 15929 10551 15963
rect 13093 15929 13127 15963
rect 3341 15861 3375 15895
rect 3985 15861 4019 15895
rect 4445 15861 4479 15895
rect 5181 15861 5215 15895
rect 5549 15861 5583 15895
rect 6377 15861 6411 15895
rect 6837 15861 6871 15895
rect 7297 15861 7331 15895
rect 9137 15861 9171 15895
rect 9597 15861 9631 15895
rect 11621 15861 11655 15895
rect 12633 15861 12667 15895
rect 13001 15861 13035 15895
rect 1593 15657 1627 15691
rect 2329 15657 2363 15691
rect 4077 15657 4111 15691
rect 4537 15657 4571 15691
rect 5457 15657 5491 15691
rect 5549 15657 5583 15691
rect 7113 15657 7147 15691
rect 11621 15657 11655 15691
rect 11989 15657 12023 15691
rect 14289 15657 14323 15691
rect 4905 15589 4939 15623
rect 6469 15589 6503 15623
rect 6561 15589 6595 15623
rect 9934 15589 9968 15623
rect 12081 15589 12115 15623
rect 1409 15521 1443 15555
rect 2421 15521 2455 15555
rect 3341 15521 3375 15555
rect 4445 15521 4479 15555
rect 2605 15453 2639 15487
rect 3433 15453 3467 15487
rect 3617 15453 3651 15487
rect 4721 15453 4755 15487
rect 7757 15521 7791 15555
rect 8197 15521 8231 15555
rect 9689 15521 9723 15555
rect 12633 15521 12667 15555
rect 12900 15521 12934 15555
rect 5733 15453 5767 15487
rect 6745 15453 6779 15487
rect 7941 15453 7975 15487
rect 12265 15453 12299 15487
rect 1961 15385 1995 15419
rect 4905 15385 4939 15419
rect 5089 15385 5123 15419
rect 9321 15385 9355 15419
rect 14013 15385 14047 15419
rect 2973 15317 3007 15351
rect 6101 15317 6135 15351
rect 7573 15317 7607 15351
rect 11069 15317 11103 15351
rect 3433 15113 3467 15147
rect 5733 15113 5767 15147
rect 14013 15113 14047 15147
rect 15025 15113 15059 15147
rect 8217 15045 8251 15079
rect 12817 15045 12851 15079
rect 1685 14977 1719 15011
rect 2881 14977 2915 15011
rect 6193 14977 6227 15011
rect 6377 14977 6411 15011
rect 8953 14977 8987 15011
rect 9045 14977 9079 15011
rect 9413 14977 9447 15011
rect 9505 14977 9539 15011
rect 10333 14977 10367 15011
rect 12449 14977 12483 15011
rect 13461 14977 13495 15011
rect 14473 14977 14507 15011
rect 14565 14977 14599 15011
rect 15669 14977 15703 15011
rect 1511 14909 1545 14943
rect 3249 14909 3283 14943
rect 3985 14909 4019 14943
rect 4252 14909 4286 14943
rect 6837 14909 6871 14943
rect 2605 14841 2639 14875
rect 6101 14841 6135 14875
rect 7104 14841 7138 14875
rect 10241 14909 10275 14943
rect 10600 14909 10634 14943
rect 13921 14909 13955 14943
rect 14381 14909 14415 14943
rect 15485 14909 15519 14943
rect 13277 14841 13311 14875
rect 2237 14773 2271 14807
rect 2697 14773 2731 14807
rect 5365 14773 5399 14807
rect 8493 14773 8527 14807
rect 8861 14773 8895 14807
rect 9413 14773 9447 14807
rect 10057 14773 10091 14807
rect 11713 14773 11747 14807
rect 13185 14773 13219 14807
rect 15393 14773 15427 14807
rect 1685 14569 1719 14603
rect 7481 14569 7515 14603
rect 8677 14569 8711 14603
rect 9321 14569 9355 14603
rect 9689 14569 9723 14603
rect 14197 14569 14231 14603
rect 15301 14569 15335 14603
rect 15669 14569 15703 14603
rect 15761 14569 15795 14603
rect 5549 14501 5583 14535
rect 10057 14501 10091 14535
rect 1501 14433 1535 14467
rect 2053 14433 2087 14467
rect 2309 14433 2343 14467
rect 4997 14433 5031 14467
rect 5457 14433 5491 14467
rect 6101 14433 6135 14467
rect 6745 14433 6779 14467
rect 7849 14433 7883 14467
rect 9505 14433 9539 14467
rect 10149 14433 10183 14467
rect 11161 14433 11195 14467
rect 11428 14433 11462 14467
rect 13084 14433 13118 14467
rect 5641 14365 5675 14399
rect 6837 14365 6871 14399
rect 7021 14365 7055 14399
rect 7941 14365 7975 14399
rect 8125 14365 8159 14399
rect 8769 14365 8803 14399
rect 8861 14365 8895 14399
rect 10333 14365 10367 14399
rect 10701 14365 10735 14399
rect 12817 14365 12851 14399
rect 15853 14365 15887 14399
rect 8309 14297 8343 14331
rect 3433 14229 3467 14263
rect 5089 14229 5123 14263
rect 5917 14229 5951 14263
rect 6377 14229 6411 14263
rect 12541 14229 12575 14263
rect 1501 14025 1535 14059
rect 3893 14025 3927 14059
rect 4905 14025 4939 14059
rect 7573 14025 7607 14059
rect 9413 14025 9447 14059
rect 10241 14025 10275 14059
rect 11069 14025 11103 14059
rect 13829 14025 13863 14059
rect 16129 14025 16163 14059
rect 4077 13957 4111 13991
rect 8585 13957 8619 13991
rect 2145 13889 2179 13923
rect 2513 13889 2547 13923
rect 4629 13889 4663 13923
rect 5365 13889 5399 13923
rect 5457 13889 5491 13923
rect 6285 13889 6319 13923
rect 8125 13889 8159 13923
rect 9229 13889 9263 13923
rect 9965 13889 9999 13923
rect 10701 13889 10735 13923
rect 10885 13889 10919 13923
rect 11529 13889 11563 13923
rect 11713 13889 11747 13923
rect 11989 13889 12023 13923
rect 12449 13889 12483 13923
rect 1961 13821 1995 13855
rect 2780 13821 2814 13855
rect 4445 13821 4479 13855
rect 5273 13821 5307 13855
rect 6193 13821 6227 13855
rect 11437 13821 11471 13855
rect 1869 13753 1903 13787
rect 4537 13753 4571 13787
rect 6837 13753 6871 13787
rect 8033 13753 8067 13787
rect 9045 13753 9079 13787
rect 9781 13753 9815 13787
rect 9873 13753 9907 13787
rect 10609 13753 10643 13787
rect 12265 13821 12299 13855
rect 12705 13821 12739 13855
rect 14749 13821 14783 13855
rect 15016 13821 15050 13855
rect 5733 13685 5767 13719
rect 6101 13685 6135 13719
rect 7941 13685 7975 13719
rect 8953 13685 8987 13719
rect 11989 13685 12023 13719
rect 12081 13685 12115 13719
rect 2145 13481 2179 13515
rect 3341 13481 3375 13515
rect 7113 13481 7147 13515
rect 9689 13481 9723 13515
rect 10057 13481 10091 13515
rect 11069 13481 11103 13515
rect 12081 13481 12115 13515
rect 13369 13481 13403 13515
rect 15301 13481 15335 13515
rect 16313 13481 16347 13515
rect 1685 13413 1719 13447
rect 4344 13413 4378 13447
rect 6000 13413 6034 13447
rect 7634 13413 7668 13447
rect 9321 13413 9355 13447
rect 10149 13413 10183 13447
rect 1409 13345 1443 13379
rect 2513 13345 2547 13379
rect 2605 13345 2639 13379
rect 3157 13345 3191 13379
rect 9045 13345 9079 13379
rect 10977 13345 11011 13379
rect 11989 13345 12023 13379
rect 13277 13345 13311 13379
rect 14289 13345 14323 13379
rect 14381 13345 14415 13379
rect 15669 13345 15703 13379
rect 15761 13345 15795 13379
rect 16681 13345 16715 13379
rect 2697 13277 2731 13311
rect 4077 13277 4111 13311
rect 5733 13277 5767 13311
rect 7389 13277 7423 13311
rect 10333 13277 10367 13311
rect 11161 13277 11195 13311
rect 12265 13277 12299 13311
rect 13461 13277 13495 13311
rect 14473 13277 14507 13311
rect 15853 13277 15887 13311
rect 16773 13277 16807 13311
rect 16865 13277 16899 13311
rect 8769 13209 8803 13243
rect 12909 13209 12943 13243
rect 5457 13141 5491 13175
rect 10609 13141 10643 13175
rect 11621 13141 11655 13175
rect 13921 13141 13955 13175
rect 6837 12937 6871 12971
rect 9689 12937 9723 12971
rect 15577 12937 15611 12971
rect 10609 12869 10643 12903
rect 12081 12869 12115 12903
rect 14381 12869 14415 12903
rect 2237 12801 2271 12835
rect 2421 12801 2455 12835
rect 3433 12801 3467 12835
rect 7389 12801 7423 12835
rect 10333 12801 10367 12835
rect 3249 12733 3283 12767
rect 3801 12733 3835 12767
rect 4721 12733 4755 12767
rect 4988 12733 5022 12767
rect 7297 12733 7331 12767
rect 7941 12733 7975 12767
rect 8208 12733 8242 12767
rect 12449 12801 12483 12835
rect 10701 12733 10735 12767
rect 12909 12733 12943 12767
rect 10057 12665 10091 12699
rect 10609 12665 10643 12699
rect 10968 12665 11002 12699
rect 13176 12665 13210 12699
rect 15117 12801 15151 12835
rect 16129 12801 16163 12835
rect 14933 12733 14967 12767
rect 15025 12733 15059 12767
rect 16037 12665 16071 12699
rect 1777 12597 1811 12631
rect 2145 12597 2179 12631
rect 2789 12597 2823 12631
rect 3157 12597 3191 12631
rect 3985 12597 4019 12631
rect 6101 12597 6135 12631
rect 7205 12597 7239 12631
rect 9321 12597 9355 12631
rect 10149 12597 10183 12631
rect 14289 12597 14323 12631
rect 14381 12597 14415 12631
rect 14565 12597 14599 12631
rect 15945 12597 15979 12631
rect 1777 12393 1811 12427
rect 2237 12393 2271 12427
rect 2789 12393 2823 12427
rect 3157 12393 3191 12427
rect 4537 12393 4571 12427
rect 9689 12393 9723 12427
rect 11621 12393 11655 12427
rect 11897 12393 11931 12427
rect 4445 12325 4479 12359
rect 8493 12325 8527 12359
rect 12265 12325 12299 12359
rect 13728 12325 13762 12359
rect 2145 12257 2179 12291
rect 3249 12257 3283 12291
rect 5089 12257 5123 12291
rect 5917 12257 5951 12291
rect 6184 12257 6218 12291
rect 8401 12257 8435 12291
rect 10508 12257 10542 12291
rect 2421 12189 2455 12223
rect 3433 12189 3467 12223
rect 4721 12189 4755 12223
rect 4905 12189 4939 12223
rect 8585 12189 8619 12223
rect 10241 12189 10275 12223
rect 12357 12189 12391 12223
rect 12449 12189 12483 12223
rect 13461 12189 13495 12223
rect 5273 12121 5307 12155
rect 4077 12053 4111 12087
rect 4905 12053 4939 12087
rect 7297 12053 7331 12087
rect 8033 12053 8067 12087
rect 14841 12053 14875 12087
rect 4997 11849 5031 11883
rect 6837 11849 6871 11883
rect 10885 11849 10919 11883
rect 13829 11849 13863 11883
rect 14105 11849 14139 11883
rect 3709 11781 3743 11815
rect 1869 11713 1903 11747
rect 4537 11713 4571 11747
rect 5457 11713 5491 11747
rect 5549 11713 5583 11747
rect 7389 11713 7423 11747
rect 11437 11713 11471 11747
rect 12449 11713 12483 11747
rect 14657 11713 14691 11747
rect 16957 11713 16991 11747
rect 1593 11645 1627 11679
rect 2329 11645 2363 11679
rect 2596 11645 2630 11679
rect 4353 11645 4387 11679
rect 7205 11645 7239 11679
rect 8401 11645 8435 11679
rect 11253 11645 11287 11679
rect 16681 11645 16715 11679
rect 5365 11577 5399 11611
rect 7297 11577 7331 11611
rect 12694 11577 12728 11611
rect 3985 11509 4019 11543
rect 4445 11509 4479 11543
rect 9689 11509 9723 11543
rect 11345 11509 11379 11543
rect 14473 11509 14507 11543
rect 14565 11509 14599 11543
rect 2789 11305 2823 11339
rect 4077 11305 4111 11339
rect 6929 11305 6963 11339
rect 7297 11305 7331 11339
rect 9321 11305 9355 11339
rect 11069 11305 11103 11339
rect 12817 11305 12851 11339
rect 13093 11305 13127 11339
rect 14105 11305 14139 11339
rect 1676 11237 1710 11271
rect 3341 11237 3375 11271
rect 8208 11237 8242 11271
rect 9934 11237 9968 11271
rect 1409 11169 1443 11203
rect 3065 11169 3099 11203
rect 5080 11169 5114 11203
rect 9689 11169 9723 11203
rect 11704 11169 11738 11203
rect 13461 11169 13495 11203
rect 13553 11169 13587 11203
rect 14473 11169 14507 11203
rect 4813 11101 4847 11135
rect 7389 11101 7423 11135
rect 7573 11101 7607 11135
rect 7941 11101 7975 11135
rect 11437 11101 11471 11135
rect 13645 11101 13679 11135
rect 14565 11101 14599 11135
rect 14657 11101 14691 11135
rect 6193 11033 6227 11067
rect 8953 10761 8987 10795
rect 11069 10761 11103 10795
rect 13277 10761 13311 10795
rect 13461 10761 13495 10795
rect 5825 10693 5859 10727
rect 3709 10625 3743 10659
rect 9229 10625 9263 10659
rect 11805 10625 11839 10659
rect 14013 10625 14047 10659
rect 2053 10557 2087 10591
rect 4445 10557 4479 10591
rect 7573 10557 7607 10591
rect 9689 10557 9723 10591
rect 9956 10557 9990 10591
rect 11621 10557 11655 10591
rect 13921 10557 13955 10591
rect 2320 10489 2354 10523
rect 4712 10489 4746 10523
rect 6101 10489 6135 10523
rect 7840 10489 7874 10523
rect 13829 10489 13863 10523
rect 14473 10489 14507 10523
rect 3433 10421 3467 10455
rect 6837 10421 6871 10455
rect 11161 10421 11195 10455
rect 11529 10421 11563 10455
rect 11989 10421 12023 10455
rect 3709 10217 3743 10251
rect 5549 10217 5583 10251
rect 6285 10217 6319 10251
rect 7757 10217 7791 10251
rect 9873 10217 9907 10251
rect 11989 10217 12023 10251
rect 12449 10217 12483 10251
rect 12909 10217 12943 10251
rect 13277 10217 13311 10251
rect 1869 10149 1903 10183
rect 1593 10081 1627 10115
rect 2596 10081 2630 10115
rect 4445 10081 4479 10115
rect 5457 10081 5491 10115
rect 10876 10149 10910 10183
rect 13645 10149 13679 10183
rect 6377 10081 6411 10115
rect 6633 10081 6667 10115
rect 8585 10081 8619 10115
rect 10057 10081 10091 10115
rect 10609 10081 10643 10115
rect 12817 10081 12851 10115
rect 2329 10013 2363 10047
rect 4537 10013 4571 10047
rect 4721 10013 4755 10047
rect 5733 10013 5767 10047
rect 6285 10013 6319 10047
rect 8677 10013 8711 10047
rect 8769 10013 8803 10047
rect 10149 10013 10183 10047
rect 13093 10013 13127 10047
rect 13737 10013 13771 10047
rect 13921 10013 13955 10047
rect 4077 9877 4111 9911
rect 5089 9877 5123 9911
rect 8217 9877 8251 9911
rect 12265 9673 12299 9707
rect 12449 9673 12483 9707
rect 6469 9605 6503 9639
rect 8125 9605 8159 9639
rect 10609 9605 10643 9639
rect 2605 9537 2639 9571
rect 3525 9537 3559 9571
rect 4537 9537 4571 9571
rect 5089 9537 5123 9571
rect 7297 9537 7331 9571
rect 7389 9537 7423 9571
rect 8677 9537 8711 9571
rect 9137 9537 9171 9571
rect 10149 9537 10183 9571
rect 11161 9537 11195 9571
rect 11989 9537 12023 9571
rect 13001 9537 13035 9571
rect 13737 9537 13771 9571
rect 13829 9537 13863 9571
rect 14657 9537 14691 9571
rect 3433 9469 3467 9503
rect 7205 9469 7239 9503
rect 8033 9469 8067 9503
rect 10057 9469 10091 9503
rect 10977 9469 11011 9503
rect 11805 9469 11839 9503
rect 12265 9469 12299 9503
rect 12817 9469 12851 9503
rect 14473 9469 14507 9503
rect 5356 9401 5390 9435
rect 11897 9401 11931 9435
rect 1961 9333 1995 9367
rect 2329 9333 2363 9367
rect 2421 9333 2455 9367
rect 2973 9333 3007 9367
rect 3341 9333 3375 9367
rect 3985 9333 4019 9367
rect 4353 9333 4387 9367
rect 4445 9333 4479 9367
rect 6837 9333 6871 9367
rect 7849 9333 7883 9367
rect 8493 9333 8527 9367
rect 8585 9333 8619 9367
rect 9597 9333 9631 9367
rect 9965 9333 9999 9367
rect 11069 9333 11103 9367
rect 11437 9333 11471 9367
rect 12909 9333 12943 9367
rect 13277 9333 13311 9367
rect 13645 9333 13679 9367
rect 14105 9333 14139 9367
rect 14565 9333 14599 9367
rect 3709 9129 3743 9163
rect 4445 9129 4479 9163
rect 7481 9129 7515 9163
rect 7849 9129 7883 9163
rect 8861 9129 8895 9163
rect 11621 9129 11655 9163
rect 11713 9129 11747 9163
rect 12725 9129 12759 9163
rect 14105 9129 14139 9163
rect 2320 9061 2354 9095
rect 2053 8993 2087 9027
rect 3893 8993 3927 9027
rect 4813 8993 4847 9027
rect 5825 8993 5859 9027
rect 5917 8993 5951 9027
rect 6837 8993 6871 9027
rect 7941 8993 7975 9027
rect 10057 8993 10091 9027
rect 11069 8993 11103 9027
rect 4905 8925 4939 8959
rect 5089 8925 5123 8959
rect 6009 8925 6043 8959
rect 6929 8925 6963 8959
rect 7113 8925 7147 8959
rect 7297 8925 7331 8959
rect 8033 8925 8067 8959
rect 8953 8925 8987 8959
rect 9045 8925 9079 8959
rect 10149 8925 10183 8959
rect 10241 8925 10275 8959
rect 11161 8925 11195 8959
rect 11253 8925 11287 8959
rect 6469 8857 6503 8891
rect 12173 9061 12207 9095
rect 13185 9061 13219 9095
rect 12081 8993 12115 9027
rect 13093 8993 13127 9027
rect 14197 8993 14231 9027
rect 12265 8925 12299 8959
rect 13369 8925 13403 8959
rect 14289 8925 14323 8959
rect 11621 8857 11655 8891
rect 3433 8789 3467 8823
rect 5457 8789 5491 8823
rect 7297 8789 7331 8823
rect 8493 8789 8527 8823
rect 9689 8789 9723 8823
rect 10701 8789 10735 8823
rect 13737 8789 13771 8823
rect 3065 8585 3099 8619
rect 4077 8585 4111 8619
rect 6469 8585 6503 8619
rect 10057 8585 10091 8619
rect 13277 8585 13311 8619
rect 13461 8585 13495 8619
rect 2789 8517 2823 8551
rect 8401 8517 8435 8551
rect 10333 8517 10367 8551
rect 12081 8517 12115 8551
rect 12449 8517 12483 8551
rect 3525 8449 3559 8483
rect 3617 8449 3651 8483
rect 4537 8449 4571 8483
rect 4721 8449 4755 8483
rect 10701 8449 10735 8483
rect 13001 8449 13035 8483
rect 1409 8381 1443 8415
rect 1676 8381 1710 8415
rect 5089 8381 5123 8415
rect 7021 8381 7055 8415
rect 8677 8381 8711 8415
rect 8944 8381 8978 8415
rect 10517 8381 10551 8415
rect 12909 8381 12943 8415
rect 14473 8517 14507 8551
rect 14013 8449 14047 8483
rect 14933 8449 14967 8483
rect 15025 8449 15059 8483
rect 13829 8381 13863 8415
rect 14841 8381 14875 8415
rect 5356 8313 5390 8347
rect 7288 8313 7322 8347
rect 10968 8313 11002 8347
rect 12817 8313 12851 8347
rect 13277 8313 13311 8347
rect 3433 8245 3467 8279
rect 4445 8245 4479 8279
rect 13921 8245 13955 8279
rect 2145 8041 2179 8075
rect 2513 8041 2547 8075
rect 3157 8041 3191 8075
rect 4261 8041 4295 8075
rect 6377 8041 6411 8075
rect 7389 8041 7423 8075
rect 8585 8041 8619 8075
rect 13093 8041 13127 8075
rect 4629 7973 4663 8007
rect 5825 7973 5859 8007
rect 6745 7973 6779 8007
rect 9956 7973 9990 8007
rect 11980 7973 12014 8007
rect 13614 7973 13648 8007
rect 5733 7905 5767 7939
rect 7757 7905 7791 7939
rect 8953 7905 8987 7939
rect 9689 7905 9723 7939
rect 2605 7837 2639 7871
rect 2697 7837 2731 7871
rect 4721 7837 4755 7871
rect 4905 7837 4939 7871
rect 5917 7837 5951 7871
rect 6837 7837 6871 7871
rect 6929 7837 6963 7871
rect 7849 7837 7883 7871
rect 8033 7837 8067 7871
rect 9045 7837 9079 7871
rect 9229 7837 9263 7871
rect 11713 7837 11747 7871
rect 13369 7837 13403 7871
rect 5365 7701 5399 7735
rect 11069 7701 11103 7735
rect 14749 7701 14783 7735
rect 6285 7497 6319 7531
rect 6653 7497 6687 7531
rect 8585 7497 8619 7531
rect 14289 7497 14323 7531
rect 2513 7361 2547 7395
rect 3525 7361 3559 7395
rect 4169 7361 4203 7395
rect 4629 7361 4663 7395
rect 11345 7429 11379 7463
rect 13461 7429 13495 7463
rect 7389 7361 7423 7395
rect 8125 7361 8159 7395
rect 9045 7361 9079 7395
rect 9229 7361 9263 7395
rect 10057 7361 10091 7395
rect 10241 7361 10275 7395
rect 11253 7361 11287 7395
rect 11989 7361 12023 7395
rect 13001 7361 13035 7395
rect 14013 7361 14047 7395
rect 2329 7293 2363 7327
rect 4896 7293 4930 7327
rect 6469 7293 6503 7327
rect 6653 7293 6687 7327
rect 7205 7293 7239 7327
rect 9965 7293 9999 7327
rect 10793 7293 10827 7327
rect 2421 7225 2455 7259
rect 14933 7361 14967 7395
rect 15025 7361 15059 7395
rect 13921 7293 13955 7327
rect 14381 7293 14415 7327
rect 14841 7293 14875 7327
rect 13829 7225 13863 7259
rect 1961 7157 1995 7191
rect 2973 7157 3007 7191
rect 3341 7157 3375 7191
rect 3433 7157 3467 7191
rect 6009 7157 6043 7191
rect 6837 7157 6871 7191
rect 7297 7157 7331 7191
rect 8953 7157 8987 7191
rect 9597 7157 9631 7191
rect 10609 7157 10643 7191
rect 11253 7157 11287 7191
rect 11713 7157 11747 7191
rect 11805 7157 11839 7191
rect 12449 7157 12483 7191
rect 12817 7157 12851 7191
rect 12909 7157 12943 7191
rect 14473 7157 14507 7191
rect 3065 6953 3099 6987
rect 5457 6953 5491 6987
rect 7941 6953 7975 6987
rect 8585 6953 8619 6987
rect 13001 6953 13035 6987
rect 13645 6953 13679 6987
rect 15669 6953 15703 6987
rect 4344 6885 4378 6919
rect 8953 6885 8987 6919
rect 1685 6817 1719 6851
rect 1952 6817 1986 6851
rect 4077 6817 4111 6851
rect 5917 6817 5951 6851
rect 6184 6817 6218 6851
rect 9597 6817 9631 6851
rect 9945 6817 9979 6851
rect 11888 6817 11922 6851
rect 3341 6749 3375 6783
rect 8033 6749 8067 6783
rect 8125 6749 8159 6783
rect 9045 6749 9079 6783
rect 9229 6749 9263 6783
rect 9413 6749 9447 6783
rect 9689 6749 9723 6783
rect 11621 6749 11655 6783
rect 13737 6749 13771 6783
rect 13921 6749 13955 6783
rect 14749 6749 14783 6783
rect 15761 6749 15795 6783
rect 15853 6749 15887 6783
rect 11069 6681 11103 6715
rect 13277 6681 13311 6715
rect 7297 6613 7331 6647
rect 7573 6613 7607 6647
rect 15301 6613 15335 6647
rect 3249 6409 3283 6443
rect 5733 6409 5767 6443
rect 10057 6409 10091 6443
rect 2973 6341 3007 6375
rect 9229 6341 9263 6375
rect 3801 6273 3835 6307
rect 4905 6273 4939 6307
rect 6285 6273 6319 6307
rect 7389 6273 7423 6307
rect 10701 6273 10735 6307
rect 11253 6273 11287 6307
rect 11989 6273 12023 6307
rect 13093 6273 13127 6307
rect 13553 6273 13587 6307
rect 1593 6205 1627 6239
rect 1860 6205 1894 6239
rect 4721 6205 4755 6239
rect 5457 6205 5491 6239
rect 7205 6205 7239 6239
rect 7849 6205 7883 6239
rect 8116 6205 8150 6239
rect 15209 6205 15243 6239
rect 7297 6137 7331 6171
rect 11253 6137 11287 6171
rect 11713 6137 11747 6171
rect 12817 6137 12851 6171
rect 13820 6137 13854 6171
rect 15454 6137 15488 6171
rect 3617 6069 3651 6103
rect 3709 6069 3743 6103
rect 4261 6069 4295 6103
rect 4629 6069 4663 6103
rect 5273 6069 5307 6103
rect 6101 6069 6135 6103
rect 6193 6069 6227 6103
rect 6837 6069 6871 6103
rect 10425 6069 10459 6103
rect 10517 6069 10551 6103
rect 11345 6069 11379 6103
rect 11805 6069 11839 6103
rect 12449 6069 12483 6103
rect 12909 6069 12943 6103
rect 14933 6069 14967 6103
rect 16589 6069 16623 6103
rect 2053 5865 2087 5899
rect 2605 5865 2639 5899
rect 6101 5865 6135 5899
rect 10609 5865 10643 5899
rect 10977 5865 11011 5899
rect 14565 5865 14599 5899
rect 16681 5865 16715 5899
rect 17417 5865 17451 5899
rect 2973 5797 3007 5831
rect 4988 5797 5022 5831
rect 7564 5797 7598 5831
rect 15568 5797 15602 5831
rect 1961 5729 1995 5763
rect 11888 5729 11922 5763
rect 14657 5729 14691 5763
rect 15301 5729 15335 5763
rect 17325 5729 17359 5763
rect 18889 5729 18923 5763
rect 2237 5661 2271 5695
rect 3065 5661 3099 5695
rect 3249 5661 3283 5695
rect 4721 5661 4755 5695
rect 7297 5661 7331 5695
rect 11069 5661 11103 5695
rect 11253 5661 11287 5695
rect 11621 5661 11655 5695
rect 13277 5661 13311 5695
rect 14841 5661 14875 5695
rect 17509 5661 17543 5695
rect 19165 5661 19199 5695
rect 1593 5593 1627 5627
rect 8677 5525 8711 5559
rect 13001 5525 13035 5559
rect 14197 5525 14231 5559
rect 16957 5525 16991 5559
rect 6009 5321 6043 5355
rect 8493 5321 8527 5355
rect 11345 5321 11379 5355
rect 12541 5321 12575 5355
rect 13461 5321 13495 5355
rect 15209 5253 15243 5287
rect 3893 5185 3927 5219
rect 8953 5185 8987 5219
rect 9137 5185 9171 5219
rect 10517 5185 10551 5219
rect 11989 5185 12023 5219
rect 13001 5185 13035 5219
rect 13185 5185 13219 5219
rect 14749 5185 14783 5219
rect 15761 5185 15795 5219
rect 2053 5117 2087 5151
rect 2320 5117 2354 5151
rect 3709 5117 3743 5151
rect 4629 5117 4663 5151
rect 4896 5117 4930 5151
rect 6837 5117 6871 5151
rect 7104 5117 7138 5151
rect 10333 5117 10367 5151
rect 12909 5117 12943 5151
rect 13553 5117 13587 5151
rect 14565 5117 14599 5151
rect 14657 5117 14691 5151
rect 16957 5117 16991 5151
rect 19809 5117 19843 5151
rect 15577 5049 15611 5083
rect 17233 5049 17267 5083
rect 3433 4981 3467 5015
rect 8217 4981 8251 5015
rect 8861 4981 8895 5015
rect 9873 4981 9907 5015
rect 10241 4981 10275 5015
rect 11713 4981 11747 5015
rect 11805 4981 11839 5015
rect 13737 4981 13771 5015
rect 14197 4981 14231 5015
rect 15669 4981 15703 5015
rect 19993 4981 20027 5015
rect 5549 4777 5583 4811
rect 6193 4777 6227 4811
rect 7389 4777 7423 4811
rect 10149 4777 10183 4811
rect 12909 4777 12943 4811
rect 14657 4777 14691 4811
rect 15669 4777 15703 4811
rect 15761 4777 15795 4811
rect 2789 4709 2823 4743
rect 6561 4709 6595 4743
rect 7757 4709 7791 4743
rect 8769 4709 8803 4743
rect 11520 4709 11554 4743
rect 14565 4709 14599 4743
rect 15025 4709 15059 4743
rect 2237 4641 2271 4675
rect 2329 4641 2363 4675
rect 2421 4573 2455 4607
rect 3249 4641 3283 4675
rect 4169 4641 4203 4675
rect 4436 4641 4470 4675
rect 8309 4641 8343 4675
rect 10057 4641 10091 4675
rect 13277 4641 13311 4675
rect 3341 4573 3375 4607
rect 3433 4573 3467 4607
rect 6653 4573 6687 4607
rect 6837 4573 6871 4607
rect 7849 4573 7883 4607
rect 8033 4573 8067 4607
rect 8861 4573 8895 4607
rect 9045 4573 9079 4607
rect 10241 4573 10275 4607
rect 11253 4573 11287 4607
rect 13369 4573 13403 4607
rect 13553 4573 13587 4607
rect 14841 4573 14875 4607
rect 12633 4505 12667 4539
rect 17877 4641 17911 4675
rect 15853 4573 15887 4607
rect 1869 4437 1903 4471
rect 2789 4437 2823 4471
rect 2881 4437 2915 4471
rect 8217 4437 8251 4471
rect 8401 4437 8435 4471
rect 9689 4437 9723 4471
rect 14197 4437 14231 4471
rect 15025 4437 15059 4471
rect 15301 4437 15335 4471
rect 18061 4437 18095 4471
rect 3157 4233 3191 4267
rect 5641 4233 5675 4267
rect 7113 4233 7147 4267
rect 8125 4233 8159 4267
rect 9321 4233 9355 4267
rect 4813 4165 4847 4199
rect 6285 4097 6319 4131
rect 7665 4097 7699 4131
rect 8677 4097 8711 4131
rect 9781 4097 9815 4131
rect 9965 4097 9999 4131
rect 11529 4097 11563 4131
rect 14657 4097 14691 4131
rect 1777 4029 1811 4063
rect 3433 4029 3467 4063
rect 6101 4029 6135 4063
rect 10333 4029 10367 4063
rect 12449 4029 12483 4063
rect 14473 4029 14507 4063
rect 15117 4029 15151 4063
rect 2044 3961 2078 3995
rect 3678 3961 3712 3995
rect 7573 3961 7607 3995
rect 12716 3961 12750 3995
rect 14565 3961 14599 3995
rect 5181 3893 5215 3927
rect 6009 3893 6043 3927
rect 7481 3893 7515 3927
rect 8493 3893 8527 3927
rect 8585 3893 8619 3927
rect 9689 3893 9723 3927
rect 10517 3893 10551 3927
rect 10885 3893 10919 3927
rect 11253 3893 11287 3927
rect 11345 3893 11379 3927
rect 13829 3893 13863 3927
rect 14105 3893 14139 3927
rect 15301 3893 15335 3927
rect 6193 3689 6227 3723
rect 9137 3689 9171 3723
rect 11253 3689 11287 3723
rect 12909 3689 12943 3723
rect 13185 3689 13219 3723
rect 16221 3689 16255 3723
rect 2044 3621 2078 3655
rect 4436 3621 4470 3655
rect 10140 3621 10174 3655
rect 11774 3621 11808 3655
rect 7380 3553 7414 3587
rect 13093 3553 13127 3587
rect 13553 3553 13587 3587
rect 14197 3553 14231 3587
rect 15301 3553 15335 3587
rect 16037 3553 16071 3587
rect 1777 3485 1811 3519
rect 3433 3485 3467 3519
rect 4169 3485 4203 3519
rect 6285 3485 6319 3519
rect 6377 3485 6411 3519
rect 7113 3485 7147 3519
rect 9873 3485 9907 3519
rect 11529 3485 11563 3519
rect 5549 3417 5583 3451
rect 5825 3417 5859 3451
rect 13645 3485 13679 3519
rect 13737 3485 13771 3519
rect 15577 3485 15611 3519
rect 3157 3349 3191 3383
rect 8493 3349 8527 3383
rect 13093 3349 13127 3383
rect 14381 3349 14415 3383
rect 1685 3145 1719 3179
rect 2513 3145 2547 3179
rect 2697 3145 2731 3179
rect 3709 3145 3743 3179
rect 4721 3145 4755 3179
rect 5733 3145 5767 3179
rect 9597 3145 9631 3179
rect 13277 3145 13311 3179
rect 14381 3145 14415 3179
rect 2329 3009 2363 3043
rect 2053 2941 2087 2975
rect 14933 3077 14967 3111
rect 3341 3009 3375 3043
rect 4169 3009 4203 3043
rect 4353 3009 4387 3043
rect 5273 3009 5307 3043
rect 6377 3009 6411 3043
rect 7757 3009 7791 3043
rect 8217 3009 8251 3043
rect 10425 3009 10459 3043
rect 11437 3009 11471 3043
rect 12909 3009 12943 3043
rect 13093 3009 13127 3043
rect 13277 3009 13311 3043
rect 3157 2941 3191 2975
rect 5181 2941 5215 2975
rect 7481 2941 7515 2975
rect 13461 2941 13495 2975
rect 13737 2941 13771 2975
rect 14197 2941 14231 2975
rect 14749 2941 14783 2975
rect 15301 2941 15335 2975
rect 16129 2941 16163 2975
rect 17049 2941 17083 2975
rect 18337 2941 18371 2975
rect 19165 2941 19199 2975
rect 2145 2873 2179 2907
rect 2513 2873 2547 2907
rect 4077 2873 4111 2907
rect 6101 2873 6135 2907
rect 8462 2873 8496 2907
rect 11345 2873 11379 2907
rect 12817 2873 12851 2907
rect 3065 2805 3099 2839
rect 5089 2805 5123 2839
rect 6193 2805 6227 2839
rect 7113 2805 7147 2839
rect 7573 2805 7607 2839
rect 9873 2805 9907 2839
rect 10241 2805 10275 2839
rect 10333 2805 10367 2839
rect 10885 2805 10919 2839
rect 11253 2805 11287 2839
rect 12449 2805 12483 2839
rect 15485 2805 15519 2839
rect 16313 2805 16347 2839
rect 17233 2805 17267 2839
rect 18521 2805 18555 2839
rect 19349 2805 19383 2839
rect 2329 2601 2363 2635
rect 2697 2601 2731 2635
rect 5365 2601 5399 2635
rect 9045 2601 9079 2635
rect 10149 2601 10183 2635
rect 10241 2601 10275 2635
rect 11161 2601 11195 2635
rect 4721 2533 4755 2567
rect 8125 2533 8159 2567
rect 9137 2533 9171 2567
rect 12081 2533 12115 2567
rect 12909 2533 12943 2567
rect 13737 2533 13771 2567
rect 5733 2465 5767 2499
rect 5825 2465 5859 2499
rect 6929 2465 6963 2499
rect 8033 2465 8067 2499
rect 11805 2465 11839 2499
rect 12643 2465 12677 2499
rect 13369 2465 13403 2499
rect 2789 2397 2823 2431
rect 2973 2397 3007 2431
rect 4813 2397 4847 2431
rect 4997 2397 5031 2431
rect 6009 2397 6043 2431
rect 7205 2397 7239 2431
rect 8217 2397 8251 2431
rect 9321 2397 9355 2431
rect 10333 2397 10367 2431
rect 11253 2397 11287 2431
rect 11437 2397 11471 2431
rect 13921 2465 13955 2499
rect 14749 2465 14783 2499
rect 15669 2465 15703 2499
rect 16589 2465 16623 2499
rect 17509 2465 17543 2499
rect 8677 2329 8711 2363
rect 10793 2329 10827 2363
rect 13553 2329 13587 2363
rect 13737 2329 13771 2363
rect 14105 2329 14139 2363
rect 4353 2261 4387 2295
rect 7665 2261 7699 2295
rect 9781 2261 9815 2295
rect 14933 2261 14967 2295
rect 15853 2261 15887 2295
rect 16773 2261 16807 2295
rect 17693 2261 17727 2295
<< metal1 >>
rect 3694 20816 3700 20868
rect 3752 20856 3758 20868
rect 6914 20856 6920 20868
rect 3752 20828 6920 20856
rect 3752 20816 3758 20828
rect 6914 20816 6920 20828
rect 6972 20816 6978 20868
rect 4062 20272 4068 20324
rect 4120 20312 4126 20324
rect 6362 20312 6368 20324
rect 4120 20284 6368 20312
rect 4120 20272 4126 20284
rect 6362 20272 6368 20284
rect 6420 20272 6426 20324
rect 3694 20204 3700 20256
rect 3752 20244 3758 20256
rect 6730 20244 6736 20256
rect 3752 20216 6736 20244
rect 3752 20204 3758 20216
rect 6730 20204 6736 20216
rect 6788 20204 6794 20256
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 4525 20043 4583 20049
rect 4525 20009 4537 20043
rect 4571 20040 4583 20043
rect 5166 20040 5172 20052
rect 4571 20012 5172 20040
rect 4571 20009 4583 20012
rect 4525 20003 4583 20009
rect 5166 20000 5172 20012
rect 5224 20000 5230 20052
rect 5534 20000 5540 20052
rect 5592 20040 5598 20052
rect 6549 20043 6607 20049
rect 6549 20040 6561 20043
rect 5592 20012 6561 20040
rect 5592 20000 5598 20012
rect 6549 20009 6561 20012
rect 6595 20009 6607 20043
rect 6549 20003 6607 20009
rect 6914 20000 6920 20052
rect 6972 20040 6978 20052
rect 9217 20043 9275 20049
rect 9217 20040 9229 20043
rect 6972 20012 9229 20040
rect 6972 20000 6978 20012
rect 9217 20009 9229 20012
rect 9263 20009 9275 20043
rect 9217 20003 9275 20009
rect 10689 20043 10747 20049
rect 10689 20009 10701 20043
rect 10735 20040 10747 20043
rect 10870 20040 10876 20052
rect 10735 20012 10876 20040
rect 10735 20009 10747 20012
rect 10689 20003 10747 20009
rect 10870 20000 10876 20012
rect 10928 20000 10934 20052
rect 12805 20043 12863 20049
rect 12805 20009 12817 20043
rect 12851 20040 12863 20043
rect 12894 20040 12900 20052
rect 12851 20012 12900 20040
rect 12851 20009 12863 20012
rect 12805 20003 12863 20009
rect 12894 20000 12900 20012
rect 12952 20000 12958 20052
rect 13354 20040 13360 20052
rect 13315 20012 13360 20040
rect 13354 20000 13360 20012
rect 13412 20000 13418 20052
rect 14369 20043 14427 20049
rect 14369 20009 14381 20043
rect 14415 20040 14427 20043
rect 14550 20040 14556 20052
rect 14415 20012 14556 20040
rect 14415 20009 14427 20012
rect 14369 20003 14427 20009
rect 14550 20000 14556 20012
rect 14608 20000 14614 20052
rect 14921 20043 14979 20049
rect 14921 20009 14933 20043
rect 14967 20040 14979 20043
rect 15194 20040 15200 20052
rect 14967 20012 15200 20040
rect 14967 20009 14979 20012
rect 14921 20003 14979 20009
rect 15194 20000 15200 20012
rect 15252 20000 15258 20052
rect 15654 20040 15660 20052
rect 15615 20012 15660 20040
rect 15654 20000 15660 20012
rect 15712 20000 15718 20052
rect 16209 20043 16267 20049
rect 16209 20009 16221 20043
rect 16255 20040 16267 20043
rect 16574 20040 16580 20052
rect 16255 20012 16580 20040
rect 16255 20009 16267 20012
rect 16209 20003 16267 20009
rect 16574 20000 16580 20012
rect 16632 20000 16638 20052
rect 17221 20043 17279 20049
rect 17221 20009 17233 20043
rect 17267 20040 17279 20043
rect 17954 20040 17960 20052
rect 17267 20012 17960 20040
rect 17267 20009 17279 20012
rect 17221 20003 17279 20009
rect 17954 20000 17960 20012
rect 18012 20000 18018 20052
rect 2501 19975 2559 19981
rect 2501 19941 2513 19975
rect 2547 19972 2559 19975
rect 10781 19975 10839 19981
rect 2547 19944 9076 19972
rect 2547 19941 2559 19944
rect 2501 19935 2559 19941
rect 1673 19907 1731 19913
rect 1673 19873 1685 19907
rect 1719 19873 1731 19907
rect 1673 19867 1731 19873
rect 2225 19907 2283 19913
rect 2225 19873 2237 19907
rect 2271 19904 2283 19907
rect 2866 19904 2872 19916
rect 2271 19876 2872 19904
rect 2271 19873 2283 19876
rect 2225 19867 2283 19873
rect 1688 19768 1716 19867
rect 2866 19864 2872 19876
rect 2924 19864 2930 19916
rect 3050 19904 3056 19916
rect 3011 19876 3056 19904
rect 3050 19864 3056 19876
rect 3108 19864 3114 19916
rect 4433 19907 4491 19913
rect 4433 19873 4445 19907
rect 4479 19904 4491 19907
rect 5258 19904 5264 19916
rect 4479 19876 5264 19904
rect 4479 19873 4491 19876
rect 4433 19867 4491 19873
rect 5258 19864 5264 19876
rect 5316 19864 5322 19916
rect 5436 19907 5494 19913
rect 5436 19873 5448 19907
rect 5482 19904 5494 19907
rect 6454 19904 6460 19916
rect 5482 19876 6460 19904
rect 5482 19873 5494 19876
rect 5436 19867 5494 19873
rect 6454 19864 6460 19876
rect 6512 19864 6518 19916
rect 7644 19907 7702 19913
rect 7644 19873 7656 19907
rect 7690 19904 7702 19907
rect 8846 19904 8852 19916
rect 7690 19876 8852 19904
rect 7690 19873 7702 19876
rect 7644 19867 7702 19873
rect 8846 19864 8852 19876
rect 8904 19864 8910 19916
rect 9048 19913 9076 19944
rect 10781 19941 10793 19975
rect 10827 19972 10839 19975
rect 12434 19972 12440 19984
rect 10827 19944 12440 19972
rect 10827 19941 10839 19944
rect 10781 19935 10839 19941
rect 12434 19932 12440 19944
rect 12492 19932 12498 19984
rect 9033 19907 9091 19913
rect 9033 19873 9045 19907
rect 9079 19873 9091 19907
rect 9033 19867 9091 19873
rect 9769 19907 9827 19913
rect 9769 19873 9781 19907
rect 9815 19904 9827 19907
rect 9858 19904 9864 19916
rect 9815 19876 9864 19904
rect 9815 19873 9827 19876
rect 9769 19867 9827 19873
rect 9858 19864 9864 19876
rect 9916 19864 9922 19916
rect 11333 19907 11391 19913
rect 11333 19873 11345 19907
rect 11379 19873 11391 19907
rect 11333 19867 11391 19873
rect 11609 19907 11667 19913
rect 11609 19873 11621 19907
rect 11655 19904 11667 19907
rect 12621 19907 12679 19913
rect 12621 19904 12633 19907
rect 11655 19876 12633 19904
rect 11655 19873 11667 19876
rect 11609 19867 11667 19873
rect 12621 19873 12633 19876
rect 12667 19873 12679 19907
rect 12621 19867 12679 19873
rect 13173 19907 13231 19913
rect 13173 19873 13185 19907
rect 13219 19904 13231 19907
rect 13906 19904 13912 19916
rect 13219 19876 13912 19904
rect 13219 19873 13231 19876
rect 13173 19867 13231 19873
rect 3234 19836 3240 19848
rect 3195 19808 3240 19836
rect 3234 19796 3240 19808
rect 3292 19796 3298 19848
rect 4709 19839 4767 19845
rect 3436 19808 4292 19836
rect 3436 19768 3464 19808
rect 1688 19740 3464 19768
rect 3510 19728 3516 19780
rect 3568 19768 3574 19780
rect 4264 19768 4292 19808
rect 4709 19805 4721 19839
rect 4755 19836 4767 19839
rect 4890 19836 4896 19848
rect 4755 19808 4896 19836
rect 4755 19805 4767 19808
rect 4709 19799 4767 19805
rect 4890 19796 4896 19808
rect 4948 19796 4954 19848
rect 5074 19796 5080 19848
rect 5132 19836 5138 19848
rect 5169 19839 5227 19845
rect 5169 19836 5181 19839
rect 5132 19808 5181 19836
rect 5132 19796 5138 19808
rect 5169 19805 5181 19808
rect 5215 19805 5227 19839
rect 5169 19799 5227 19805
rect 6917 19839 6975 19845
rect 6917 19805 6929 19839
rect 6963 19805 6975 19839
rect 7374 19836 7380 19848
rect 7335 19808 7380 19836
rect 6917 19799 6975 19805
rect 4982 19768 4988 19780
rect 3568 19740 4200 19768
rect 4264 19740 4988 19768
rect 3568 19728 3574 19740
rect 1854 19700 1860 19712
rect 1815 19672 1860 19700
rect 1854 19660 1860 19672
rect 1912 19660 1918 19712
rect 4062 19700 4068 19712
rect 4023 19672 4068 19700
rect 4062 19660 4068 19672
rect 4120 19660 4126 19712
rect 4172 19700 4200 19740
rect 4982 19728 4988 19740
rect 5040 19728 5046 19780
rect 6932 19768 6960 19799
rect 7374 19796 7380 19808
rect 7432 19796 7438 19848
rect 10962 19836 10968 19848
rect 10923 19808 10968 19836
rect 10962 19796 10968 19808
rect 11020 19796 11026 19848
rect 11348 19836 11376 19867
rect 13906 19864 13912 19876
rect 13964 19864 13970 19916
rect 14182 19904 14188 19916
rect 14143 19876 14188 19904
rect 14182 19864 14188 19876
rect 14240 19864 14246 19916
rect 14458 19864 14464 19916
rect 14516 19904 14522 19916
rect 14737 19907 14795 19913
rect 14737 19904 14749 19907
rect 14516 19876 14749 19904
rect 14516 19864 14522 19876
rect 14737 19873 14749 19876
rect 14783 19873 14795 19907
rect 15470 19904 15476 19916
rect 15431 19876 15476 19904
rect 14737 19867 14795 19873
rect 15470 19864 15476 19876
rect 15528 19864 15534 19916
rect 15562 19864 15568 19916
rect 15620 19904 15626 19916
rect 16025 19907 16083 19913
rect 16025 19904 16037 19907
rect 15620 19876 16037 19904
rect 15620 19864 15626 19876
rect 16025 19873 16037 19876
rect 16071 19873 16083 19907
rect 17034 19904 17040 19916
rect 16995 19876 17040 19904
rect 16025 19867 16083 19873
rect 17034 19864 17040 19876
rect 17092 19864 17098 19916
rect 11698 19836 11704 19848
rect 11348 19808 11704 19836
rect 11698 19796 11704 19808
rect 11756 19796 11762 19848
rect 12066 19836 12072 19848
rect 12027 19808 12072 19836
rect 12066 19796 12072 19808
rect 12124 19796 12130 19848
rect 6104 19740 6960 19768
rect 9953 19771 10011 19777
rect 6104 19700 6132 19740
rect 9953 19737 9965 19771
rect 9999 19768 10011 19771
rect 19794 19768 19800 19780
rect 9999 19740 19800 19768
rect 9999 19737 10011 19740
rect 9953 19731 10011 19737
rect 19794 19728 19800 19740
rect 19852 19728 19858 19780
rect 4172 19672 6132 19700
rect 6914 19660 6920 19712
rect 6972 19700 6978 19712
rect 8757 19703 8815 19709
rect 8757 19700 8769 19703
rect 6972 19672 8769 19700
rect 6972 19660 6978 19672
rect 8757 19669 8769 19672
rect 8803 19669 8815 19703
rect 8757 19663 8815 19669
rect 10321 19703 10379 19709
rect 10321 19669 10333 19703
rect 10367 19700 10379 19703
rect 11790 19700 11796 19712
rect 10367 19672 11796 19700
rect 10367 19669 10379 19672
rect 10321 19663 10379 19669
rect 11790 19660 11796 19672
rect 11848 19660 11854 19712
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 3234 19456 3240 19508
rect 3292 19496 3298 19508
rect 5810 19496 5816 19508
rect 3292 19468 5816 19496
rect 3292 19456 3298 19468
rect 5810 19456 5816 19468
rect 5868 19456 5874 19508
rect 6454 19496 6460 19508
rect 6415 19468 6460 19496
rect 6454 19456 6460 19468
rect 6512 19456 6518 19508
rect 7374 19456 7380 19508
rect 7432 19456 7438 19508
rect 10962 19456 10968 19508
rect 11020 19496 11026 19508
rect 13817 19499 13875 19505
rect 13817 19496 13829 19499
rect 11020 19468 13829 19496
rect 11020 19456 11026 19468
rect 13817 19465 13829 19468
rect 13863 19465 13875 19499
rect 13817 19459 13875 19465
rect 3970 19320 3976 19372
rect 4028 19360 4034 19372
rect 6472 19360 6500 19456
rect 7392 19428 7420 19456
rect 7392 19400 8064 19428
rect 8036 19369 8064 19400
rect 7377 19363 7435 19369
rect 7377 19360 7389 19363
rect 4028 19332 5212 19360
rect 6472 19332 7389 19360
rect 4028 19320 4034 19332
rect 1581 19295 1639 19301
rect 1581 19261 1593 19295
rect 1627 19261 1639 19295
rect 2130 19292 2136 19304
rect 2091 19264 2136 19292
rect 1581 19255 1639 19261
rect 1596 19224 1624 19255
rect 2130 19252 2136 19264
rect 2188 19252 2194 19304
rect 2961 19295 3019 19301
rect 2961 19261 2973 19295
rect 3007 19261 3019 19295
rect 2961 19255 3019 19261
rect 3228 19295 3286 19301
rect 3228 19261 3240 19295
rect 3274 19292 3286 19295
rect 4890 19292 4896 19304
rect 3274 19264 4896 19292
rect 3274 19261 3286 19264
rect 3228 19255 3286 19261
rect 2222 19224 2228 19236
rect 1596 19196 2228 19224
rect 2222 19184 2228 19196
rect 2280 19184 2286 19236
rect 2409 19227 2467 19233
rect 2409 19193 2421 19227
rect 2455 19224 2467 19227
rect 2590 19224 2596 19236
rect 2455 19196 2596 19224
rect 2455 19193 2467 19196
rect 2409 19187 2467 19193
rect 2590 19184 2596 19196
rect 2648 19184 2654 19236
rect 1762 19156 1768 19168
rect 1723 19128 1768 19156
rect 1762 19116 1768 19128
rect 1820 19116 1826 19168
rect 2976 19156 3004 19255
rect 4890 19252 4896 19264
rect 4948 19252 4954 19304
rect 5074 19292 5080 19304
rect 5035 19264 5080 19292
rect 5074 19252 5080 19264
rect 5132 19252 5138 19304
rect 5184 19292 5212 19332
rect 7377 19329 7389 19332
rect 7423 19329 7435 19363
rect 7377 19323 7435 19329
rect 8021 19363 8079 19369
rect 8021 19329 8033 19363
rect 8067 19329 8079 19363
rect 8021 19323 8079 19329
rect 11241 19363 11299 19369
rect 11241 19329 11253 19363
rect 11287 19360 11299 19363
rect 11885 19363 11943 19369
rect 11885 19360 11897 19363
rect 11287 19332 11897 19360
rect 11287 19329 11299 19332
rect 11241 19323 11299 19329
rect 11885 19329 11897 19332
rect 11931 19329 11943 19363
rect 11885 19323 11943 19329
rect 5184 19264 7052 19292
rect 4246 19184 4252 19236
rect 4304 19224 4310 19236
rect 4617 19227 4675 19233
rect 4617 19224 4629 19227
rect 4304 19196 4629 19224
rect 4304 19184 4310 19196
rect 4617 19193 4629 19196
rect 4663 19193 4675 19227
rect 4617 19187 4675 19193
rect 5344 19227 5402 19233
rect 5344 19193 5356 19227
rect 5390 19224 5402 19227
rect 5718 19224 5724 19236
rect 5390 19196 5724 19224
rect 5390 19193 5402 19196
rect 5344 19187 5402 19193
rect 5718 19184 5724 19196
rect 5776 19184 5782 19236
rect 5810 19184 5816 19236
rect 5868 19224 5874 19236
rect 6914 19224 6920 19236
rect 5868 19196 6920 19224
rect 5868 19184 5874 19196
rect 6914 19184 6920 19196
rect 6972 19184 6978 19236
rect 7024 19224 7052 19264
rect 7098 19252 7104 19304
rect 7156 19292 7162 19304
rect 7285 19295 7343 19301
rect 7285 19292 7297 19295
rect 7156 19264 7297 19292
rect 7156 19252 7162 19264
rect 7285 19261 7297 19264
rect 7331 19261 7343 19295
rect 8754 19292 8760 19304
rect 7285 19255 7343 19261
rect 8128 19264 8760 19292
rect 8128 19224 8156 19264
rect 8754 19252 8760 19264
rect 8812 19252 8818 19304
rect 9677 19295 9735 19301
rect 9677 19261 9689 19295
rect 9723 19292 9735 19295
rect 10318 19292 10324 19304
rect 9723 19264 10324 19292
rect 9723 19261 9735 19264
rect 9677 19255 9735 19261
rect 10318 19252 10324 19264
rect 10376 19252 10382 19304
rect 11701 19295 11759 19301
rect 11701 19261 11713 19295
rect 11747 19292 11759 19295
rect 12066 19292 12072 19304
rect 11747 19264 12072 19292
rect 11747 19261 11759 19264
rect 11701 19255 11759 19261
rect 12066 19252 12072 19264
rect 12124 19252 12130 19304
rect 12158 19252 12164 19304
rect 12216 19292 12222 19304
rect 12437 19295 12495 19301
rect 12437 19292 12449 19295
rect 12216 19264 12449 19292
rect 12216 19252 12222 19264
rect 12437 19261 12449 19264
rect 12483 19261 12495 19295
rect 14090 19292 14096 19304
rect 14051 19264 14096 19292
rect 12437 19255 12495 19261
rect 14090 19252 14096 19264
rect 14148 19252 14154 19304
rect 14921 19295 14979 19301
rect 14921 19261 14933 19295
rect 14967 19292 14979 19295
rect 15933 19295 15991 19301
rect 14967 19264 15884 19292
rect 14967 19261 14979 19264
rect 14921 19255 14979 19261
rect 7024 19196 8156 19224
rect 8288 19227 8346 19233
rect 8288 19193 8300 19227
rect 8334 19224 8346 19227
rect 9944 19227 10002 19233
rect 8334 19196 9904 19224
rect 8334 19193 8346 19196
rect 8288 19187 8346 19193
rect 3234 19156 3240 19168
rect 2976 19128 3240 19156
rect 3234 19116 3240 19128
rect 3292 19116 3298 19168
rect 3326 19116 3332 19168
rect 3384 19156 3390 19168
rect 3510 19156 3516 19168
rect 3384 19128 3516 19156
rect 3384 19116 3390 19128
rect 3510 19116 3516 19128
rect 3568 19116 3574 19168
rect 3602 19116 3608 19168
rect 3660 19156 3666 19168
rect 4341 19159 4399 19165
rect 4341 19156 4353 19159
rect 3660 19128 4353 19156
rect 3660 19116 3666 19128
rect 4341 19125 4353 19128
rect 4387 19125 4399 19159
rect 4341 19119 4399 19125
rect 4430 19116 4436 19168
rect 4488 19156 4494 19168
rect 5828 19156 5856 19184
rect 4488 19128 5856 19156
rect 4488 19116 4494 19128
rect 6638 19116 6644 19168
rect 6696 19156 6702 19168
rect 6825 19159 6883 19165
rect 6825 19156 6837 19159
rect 6696 19128 6837 19156
rect 6696 19116 6702 19128
rect 6825 19125 6837 19128
rect 6871 19125 6883 19159
rect 6825 19119 6883 19125
rect 7006 19116 7012 19168
rect 7064 19156 7070 19168
rect 7193 19159 7251 19165
rect 7193 19156 7205 19159
rect 7064 19128 7205 19156
rect 7064 19116 7070 19128
rect 7193 19125 7205 19128
rect 7239 19125 7251 19159
rect 7193 19119 7251 19125
rect 8386 19116 8392 19168
rect 8444 19156 8450 19168
rect 9030 19156 9036 19168
rect 8444 19128 9036 19156
rect 8444 19116 8450 19128
rect 9030 19116 9036 19128
rect 9088 19116 9094 19168
rect 9398 19156 9404 19168
rect 9359 19128 9404 19156
rect 9398 19116 9404 19128
rect 9456 19116 9462 19168
rect 9876 19156 9904 19196
rect 9944 19193 9956 19227
rect 9990 19224 10002 19227
rect 10962 19224 10968 19236
rect 9990 19196 10968 19224
rect 9990 19193 10002 19196
rect 9944 19187 10002 19193
rect 10962 19184 10968 19196
rect 11020 19184 11026 19236
rect 11790 19224 11796 19236
rect 11751 19196 11796 19224
rect 11790 19184 11796 19196
rect 11848 19184 11854 19236
rect 12710 19233 12716 19236
rect 12704 19224 12716 19233
rect 12671 19196 12716 19224
rect 12704 19187 12716 19196
rect 12710 19184 12716 19187
rect 12768 19184 12774 19236
rect 13722 19184 13728 19236
rect 13780 19224 13786 19236
rect 15565 19227 15623 19233
rect 15565 19224 15577 19227
rect 13780 19196 15577 19224
rect 13780 19184 13786 19196
rect 15565 19193 15577 19196
rect 15611 19193 15623 19227
rect 15856 19224 15884 19264
rect 15933 19261 15945 19295
rect 15979 19292 15991 19295
rect 16025 19295 16083 19301
rect 16025 19292 16037 19295
rect 15979 19264 16037 19292
rect 15979 19261 15991 19264
rect 15933 19255 15991 19261
rect 16025 19261 16037 19264
rect 16071 19261 16083 19295
rect 16574 19292 16580 19304
rect 16535 19264 16580 19292
rect 16025 19255 16083 19261
rect 16574 19252 16580 19264
rect 16632 19252 16638 19304
rect 17126 19292 17132 19304
rect 17087 19264 17132 19292
rect 17126 19252 17132 19264
rect 17184 19252 17190 19304
rect 17218 19252 17224 19304
rect 17276 19292 17282 19304
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 17276 19264 18061 19292
rect 17276 19252 17282 19264
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18598 19292 18604 19304
rect 18559 19264 18604 19292
rect 18049 19255 18107 19261
rect 18598 19252 18604 19264
rect 18656 19252 18662 19304
rect 18782 19252 18788 19304
rect 18840 19292 18846 19304
rect 19429 19295 19487 19301
rect 19429 19292 19441 19295
rect 18840 19264 19441 19292
rect 18840 19252 18846 19264
rect 19429 19261 19441 19264
rect 19475 19261 19487 19295
rect 19429 19255 19487 19261
rect 22094 19224 22100 19236
rect 15856 19196 22100 19224
rect 15565 19187 15623 19193
rect 22094 19184 22100 19196
rect 22152 19184 22158 19236
rect 11057 19159 11115 19165
rect 11057 19156 11069 19159
rect 9876 19128 11069 19156
rect 11057 19125 11069 19128
rect 11103 19156 11115 19159
rect 11241 19159 11299 19165
rect 11241 19156 11253 19159
rect 11103 19128 11253 19156
rect 11103 19125 11115 19128
rect 11057 19119 11115 19125
rect 11241 19125 11253 19128
rect 11287 19125 11299 19159
rect 11241 19119 11299 19125
rect 11333 19159 11391 19165
rect 11333 19125 11345 19159
rect 11379 19156 11391 19159
rect 11422 19156 11428 19168
rect 11379 19128 11428 19156
rect 11379 19125 11391 19128
rect 11333 19119 11391 19125
rect 11422 19116 11428 19128
rect 11480 19116 11486 19168
rect 14274 19156 14280 19168
rect 14235 19128 14280 19156
rect 14274 19116 14280 19128
rect 14332 19116 14338 19168
rect 15102 19116 15108 19168
rect 15160 19156 15166 19168
rect 15933 19159 15991 19165
rect 15933 19156 15945 19159
rect 15160 19128 15945 19156
rect 15160 19116 15166 19128
rect 15933 19125 15945 19128
rect 15979 19125 15991 19159
rect 15933 19119 15991 19125
rect 16114 19116 16120 19168
rect 16172 19156 16178 19168
rect 16209 19159 16267 19165
rect 16209 19156 16221 19159
rect 16172 19128 16221 19156
rect 16172 19116 16178 19128
rect 16209 19125 16221 19128
rect 16255 19125 16267 19159
rect 16209 19119 16267 19125
rect 16761 19159 16819 19165
rect 16761 19125 16773 19159
rect 16807 19156 16819 19159
rect 16942 19156 16948 19168
rect 16807 19128 16948 19156
rect 16807 19125 16819 19128
rect 16761 19119 16819 19125
rect 16942 19116 16948 19128
rect 17000 19116 17006 19168
rect 17313 19159 17371 19165
rect 17313 19125 17325 19159
rect 17359 19156 17371 19159
rect 17494 19156 17500 19168
rect 17359 19128 17500 19156
rect 17359 19125 17371 19128
rect 17313 19119 17371 19125
rect 17494 19116 17500 19128
rect 17552 19116 17558 19168
rect 18233 19159 18291 19165
rect 18233 19125 18245 19159
rect 18279 19156 18291 19159
rect 18506 19156 18512 19168
rect 18279 19128 18512 19156
rect 18279 19125 18291 19128
rect 18233 19119 18291 19125
rect 18506 19116 18512 19128
rect 18564 19116 18570 19168
rect 18785 19159 18843 19165
rect 18785 19125 18797 19159
rect 18831 19156 18843 19159
rect 18874 19156 18880 19168
rect 18831 19128 18880 19156
rect 18831 19125 18843 19128
rect 18785 19119 18843 19125
rect 18874 19116 18880 19128
rect 18932 19116 18938 19168
rect 19613 19159 19671 19165
rect 19613 19125 19625 19159
rect 19659 19156 19671 19159
rect 20254 19156 20260 19168
rect 19659 19128 20260 19156
rect 19659 19125 19671 19128
rect 19613 19119 19671 19125
rect 20254 19116 20260 19128
rect 20312 19116 20318 19168
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 1486 18912 1492 18964
rect 1544 18952 1550 18964
rect 2498 18952 2504 18964
rect 1544 18924 2504 18952
rect 1544 18912 1550 18924
rect 2498 18912 2504 18924
rect 2556 18912 2562 18964
rect 2866 18912 2872 18964
rect 2924 18952 2930 18964
rect 2961 18955 3019 18961
rect 2961 18952 2973 18955
rect 2924 18924 2973 18952
rect 2924 18912 2930 18924
rect 2961 18921 2973 18924
rect 3007 18921 3019 18955
rect 3326 18952 3332 18964
rect 3287 18924 3332 18952
rect 2961 18915 3019 18921
rect 3326 18912 3332 18924
rect 3384 18912 3390 18964
rect 3421 18955 3479 18961
rect 3421 18921 3433 18955
rect 3467 18952 3479 18955
rect 4062 18952 4068 18964
rect 3467 18924 4068 18952
rect 3467 18921 3479 18924
rect 3421 18915 3479 18921
rect 4062 18912 4068 18924
rect 4120 18912 4126 18964
rect 4338 18912 4344 18964
rect 4396 18952 4402 18964
rect 5166 18952 5172 18964
rect 4396 18924 5172 18952
rect 4396 18912 4402 18924
rect 5166 18912 5172 18924
rect 5224 18912 5230 18964
rect 5534 18952 5540 18964
rect 5276 18924 5540 18952
rect 2409 18887 2467 18893
rect 2409 18853 2421 18887
rect 2455 18884 2467 18887
rect 3970 18884 3976 18896
rect 2455 18856 3976 18884
rect 2455 18853 2467 18856
rect 2409 18847 2467 18853
rect 3970 18844 3976 18856
rect 4028 18844 4034 18896
rect 4522 18884 4528 18896
rect 4483 18856 4528 18884
rect 4522 18844 4528 18856
rect 4580 18844 4586 18896
rect 5276 18884 5304 18924
rect 5534 18912 5540 18924
rect 5592 18912 5598 18964
rect 5718 18912 5724 18964
rect 5776 18952 5782 18964
rect 6549 18955 6607 18961
rect 6549 18952 6561 18955
rect 5776 18924 6561 18952
rect 5776 18912 5782 18924
rect 6549 18921 6561 18924
rect 6595 18921 6607 18955
rect 6549 18915 6607 18921
rect 6730 18912 6736 18964
rect 6788 18952 6794 18964
rect 7009 18955 7067 18961
rect 7009 18952 7021 18955
rect 6788 18924 7021 18952
rect 6788 18912 6794 18924
rect 7009 18921 7021 18924
rect 7055 18921 7067 18955
rect 8846 18952 8852 18964
rect 8807 18924 8852 18952
rect 7009 18915 7067 18921
rect 8846 18912 8852 18924
rect 8904 18912 8910 18964
rect 9306 18912 9312 18964
rect 9364 18952 9370 18964
rect 11882 18952 11888 18964
rect 9364 18924 10272 18952
rect 9364 18912 9370 18924
rect 7374 18884 7380 18896
rect 4724 18856 5304 18884
rect 5368 18856 7380 18884
rect 1394 18816 1400 18828
rect 1355 18788 1400 18816
rect 1394 18776 1400 18788
rect 1452 18776 1458 18828
rect 2317 18819 2375 18825
rect 2317 18785 2329 18819
rect 2363 18816 2375 18819
rect 3326 18816 3332 18828
rect 2363 18788 3332 18816
rect 2363 18785 2375 18788
rect 2317 18779 2375 18785
rect 3326 18776 3332 18788
rect 3384 18776 3390 18828
rect 4338 18816 4344 18828
rect 3436 18788 4344 18816
rect 198 18708 204 18760
rect 256 18748 262 18760
rect 2593 18751 2651 18757
rect 256 18720 1716 18748
rect 256 18708 262 18720
rect 1578 18680 1584 18692
rect 1539 18652 1584 18680
rect 1578 18640 1584 18652
rect 1636 18640 1642 18692
rect 1688 18680 1716 18720
rect 2593 18717 2605 18751
rect 2639 18748 2651 18751
rect 3436 18748 3464 18788
rect 4338 18776 4344 18788
rect 4396 18776 4402 18828
rect 4433 18819 4491 18825
rect 4433 18785 4445 18819
rect 4479 18785 4491 18819
rect 4433 18779 4491 18785
rect 3602 18748 3608 18760
rect 2639 18720 3464 18748
rect 3563 18720 3608 18748
rect 2639 18717 2651 18720
rect 2593 18711 2651 18717
rect 3602 18708 3608 18720
rect 3660 18708 3666 18760
rect 4448 18748 4476 18779
rect 4724 18757 4752 18856
rect 5368 18816 5396 18856
rect 7374 18844 7380 18856
rect 7432 18844 7438 18896
rect 7736 18887 7794 18893
rect 7736 18853 7748 18887
rect 7782 18884 7794 18887
rect 9398 18884 9404 18896
rect 7782 18856 9404 18884
rect 7782 18853 7794 18856
rect 7736 18847 7794 18853
rect 9398 18844 9404 18856
rect 9456 18884 9462 18896
rect 10244 18884 10272 18924
rect 11808 18924 11888 18952
rect 11808 18884 11836 18924
rect 11882 18912 11888 18924
rect 11940 18912 11946 18964
rect 12710 18952 12716 18964
rect 11992 18924 12716 18952
rect 11992 18884 12020 18924
rect 12710 18912 12716 18924
rect 12768 18952 12774 18964
rect 13357 18955 13415 18961
rect 13357 18952 13369 18955
rect 12768 18924 13369 18952
rect 12768 18912 12774 18924
rect 13357 18921 13369 18924
rect 13403 18921 13415 18955
rect 13357 18915 13415 18921
rect 19334 18912 19340 18964
rect 19392 18952 19398 18964
rect 21174 18952 21180 18964
rect 19392 18924 21180 18952
rect 19392 18912 19398 18924
rect 21174 18912 21180 18924
rect 21232 18912 21238 18964
rect 9456 18856 10180 18884
rect 10244 18856 11836 18884
rect 11900 18856 12020 18884
rect 9456 18844 9462 18856
rect 5276 18788 5396 18816
rect 5436 18819 5494 18825
rect 4709 18751 4767 18757
rect 4448 18720 4660 18748
rect 2774 18680 2780 18692
rect 1688 18652 2780 18680
rect 2774 18640 2780 18652
rect 2832 18640 2838 18692
rect 3050 18640 3056 18692
rect 3108 18680 3114 18692
rect 4065 18683 4123 18689
rect 4065 18680 4077 18683
rect 3108 18652 4077 18680
rect 3108 18640 3114 18652
rect 4065 18649 4077 18652
rect 4111 18649 4123 18683
rect 4065 18643 4123 18649
rect 1949 18615 2007 18621
rect 1949 18581 1961 18615
rect 1995 18612 2007 18615
rect 4154 18612 4160 18624
rect 1995 18584 4160 18612
rect 1995 18581 2007 18584
rect 1949 18575 2007 18581
rect 4154 18572 4160 18584
rect 4212 18572 4218 18624
rect 4632 18612 4660 18720
rect 4709 18717 4721 18751
rect 4755 18748 4767 18751
rect 4798 18748 4804 18760
rect 4755 18720 4804 18748
rect 4755 18717 4767 18720
rect 4709 18711 4767 18717
rect 4798 18708 4804 18720
rect 4856 18708 4862 18760
rect 5074 18708 5080 18760
rect 5132 18748 5138 18760
rect 5169 18751 5227 18757
rect 5169 18748 5181 18751
rect 5132 18720 5181 18748
rect 5132 18708 5138 18720
rect 5169 18717 5181 18720
rect 5215 18748 5227 18751
rect 5276 18748 5304 18788
rect 5436 18785 5448 18819
rect 5482 18816 5494 18819
rect 5810 18816 5816 18828
rect 5482 18788 5816 18816
rect 5482 18785 5494 18788
rect 5436 18779 5494 18785
rect 5810 18776 5816 18788
rect 5868 18776 5874 18828
rect 5994 18776 6000 18828
rect 6052 18816 6058 18828
rect 6825 18819 6883 18825
rect 6825 18816 6837 18819
rect 6052 18788 6837 18816
rect 6052 18776 6058 18788
rect 6825 18785 6837 18788
rect 6871 18785 6883 18819
rect 9125 18819 9183 18825
rect 9125 18816 9137 18819
rect 6825 18779 6883 18785
rect 7300 18788 9137 18816
rect 5215 18720 5304 18748
rect 5215 18717 5227 18720
rect 5169 18711 5227 18717
rect 7300 18612 7328 18788
rect 9125 18785 9137 18788
rect 9171 18785 9183 18819
rect 10045 18819 10103 18825
rect 10045 18816 10057 18819
rect 9125 18779 9183 18785
rect 9968 18788 10057 18816
rect 7374 18708 7380 18760
rect 7432 18748 7438 18760
rect 7469 18751 7527 18757
rect 7469 18748 7481 18751
rect 7432 18720 7481 18748
rect 7432 18708 7438 18720
rect 7469 18717 7481 18720
rect 7515 18717 7527 18751
rect 7469 18711 7527 18717
rect 4632 18584 7328 18612
rect 8386 18572 8392 18624
rect 8444 18612 8450 18624
rect 9677 18615 9735 18621
rect 9677 18612 9689 18615
rect 8444 18584 9689 18612
rect 8444 18572 8450 18584
rect 9677 18581 9689 18584
rect 9723 18581 9735 18615
rect 9968 18612 9996 18788
rect 10045 18785 10057 18788
rect 10091 18785 10103 18819
rect 10152 18816 10180 18856
rect 11330 18816 11336 18828
rect 10152 18788 10272 18816
rect 11291 18788 11336 18816
rect 10045 18779 10103 18785
rect 10134 18748 10140 18760
rect 10095 18720 10140 18748
rect 10134 18708 10140 18720
rect 10192 18708 10198 18760
rect 10244 18757 10272 18788
rect 11330 18776 11336 18788
rect 11388 18776 11394 18828
rect 11425 18819 11483 18825
rect 11425 18785 11437 18819
rect 11471 18816 11483 18819
rect 11790 18816 11796 18828
rect 11471 18788 11796 18816
rect 11471 18785 11483 18788
rect 11425 18779 11483 18785
rect 11790 18776 11796 18788
rect 11848 18776 11854 18828
rect 10229 18751 10287 18757
rect 10229 18717 10241 18751
rect 10275 18717 10287 18751
rect 10229 18711 10287 18717
rect 11609 18751 11667 18757
rect 11609 18717 11621 18751
rect 11655 18748 11667 18751
rect 11900 18748 11928 18856
rect 12342 18844 12348 18896
rect 12400 18884 12406 18896
rect 13906 18884 13912 18896
rect 12400 18856 13676 18884
rect 13867 18856 13912 18884
rect 12400 18844 12406 18856
rect 11977 18819 12035 18825
rect 11977 18785 11989 18819
rect 12023 18816 12035 18819
rect 12066 18816 12072 18828
rect 12023 18788 12072 18816
rect 12023 18785 12035 18788
rect 11977 18779 12035 18785
rect 12066 18776 12072 18788
rect 12124 18776 12130 18828
rect 12244 18819 12302 18825
rect 12244 18785 12256 18819
rect 12290 18816 12302 18819
rect 12986 18816 12992 18828
rect 12290 18788 12992 18816
rect 12290 18785 12302 18788
rect 12244 18779 12302 18785
rect 12986 18776 12992 18788
rect 13044 18776 13050 18828
rect 13648 18825 13676 18856
rect 13906 18844 13912 18856
rect 13964 18844 13970 18896
rect 14182 18844 14188 18896
rect 14240 18884 14246 18896
rect 14645 18887 14703 18893
rect 14645 18884 14657 18887
rect 14240 18856 14657 18884
rect 14240 18844 14246 18856
rect 14645 18853 14657 18856
rect 14691 18853 14703 18887
rect 15562 18884 15568 18896
rect 15523 18856 15568 18884
rect 14645 18847 14703 18853
rect 15562 18844 15568 18856
rect 15620 18844 15626 18896
rect 18782 18884 18788 18896
rect 18743 18856 18788 18884
rect 18782 18844 18788 18856
rect 18840 18844 18846 18896
rect 13633 18819 13691 18825
rect 13633 18785 13645 18819
rect 13679 18785 13691 18819
rect 13633 18779 13691 18785
rect 14369 18819 14427 18825
rect 14369 18785 14381 18819
rect 14415 18785 14427 18819
rect 14369 18779 14427 18785
rect 11655 18720 11928 18748
rect 14384 18748 14412 18779
rect 15194 18776 15200 18828
rect 15252 18816 15258 18828
rect 15289 18819 15347 18825
rect 15289 18816 15301 18819
rect 15252 18788 15301 18816
rect 15252 18776 15258 18788
rect 15289 18785 15301 18788
rect 15335 18785 15347 18819
rect 18506 18816 18512 18828
rect 18467 18788 18512 18816
rect 15289 18779 15347 18785
rect 18506 18776 18512 18788
rect 18564 18776 18570 18828
rect 15562 18748 15568 18760
rect 14384 18720 15568 18748
rect 11655 18717 11667 18720
rect 11609 18711 11667 18717
rect 15562 18708 15568 18720
rect 15620 18708 15626 18760
rect 10686 18612 10692 18624
rect 9968 18584 10692 18612
rect 9677 18575 9735 18581
rect 10686 18572 10692 18584
rect 10744 18572 10750 18624
rect 10962 18612 10968 18624
rect 10923 18584 10968 18612
rect 10962 18572 10968 18584
rect 11020 18572 11026 18624
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 1026 18368 1032 18420
rect 1084 18408 1090 18420
rect 2590 18408 2596 18420
rect 1084 18380 2596 18408
rect 1084 18368 1090 18380
rect 2590 18368 2596 18380
rect 2648 18368 2654 18420
rect 2774 18368 2780 18420
rect 2832 18408 2838 18420
rect 3050 18408 3056 18420
rect 2832 18380 3056 18408
rect 2832 18368 2838 18380
rect 3050 18368 3056 18380
rect 3108 18368 3114 18420
rect 3329 18411 3387 18417
rect 3329 18377 3341 18411
rect 3375 18408 3387 18411
rect 10962 18408 10968 18420
rect 3375 18380 10968 18408
rect 3375 18377 3387 18380
rect 3329 18371 3387 18377
rect 10962 18368 10968 18380
rect 11020 18368 11026 18420
rect 11790 18368 11796 18420
rect 11848 18408 11854 18420
rect 12437 18411 12495 18417
rect 12437 18408 12449 18411
rect 11848 18380 12449 18408
rect 11848 18368 11854 18380
rect 12437 18377 12449 18380
rect 12483 18377 12495 18411
rect 13446 18408 13452 18420
rect 13407 18380 13452 18408
rect 12437 18371 12495 18377
rect 13446 18368 13452 18380
rect 13504 18368 13510 18420
rect 14645 18411 14703 18417
rect 14645 18377 14657 18411
rect 14691 18408 14703 18411
rect 21634 18408 21640 18420
rect 14691 18380 21640 18408
rect 14691 18377 14703 18380
rect 14645 18371 14703 18377
rect 21634 18368 21640 18380
rect 21692 18368 21698 18420
rect 1670 18340 1676 18352
rect 1631 18312 1676 18340
rect 1670 18300 1676 18312
rect 1728 18300 1734 18352
rect 4890 18340 4896 18352
rect 4851 18312 4896 18340
rect 4890 18300 4896 18312
rect 4948 18300 4954 18352
rect 5077 18343 5135 18349
rect 5077 18309 5089 18343
rect 5123 18340 5135 18343
rect 9033 18343 9091 18349
rect 9033 18340 9045 18343
rect 5123 18312 9045 18340
rect 5123 18309 5135 18312
rect 5077 18303 5135 18309
rect 9033 18309 9045 18312
rect 9079 18309 9091 18343
rect 10042 18340 10048 18352
rect 9033 18303 9091 18309
rect 9600 18312 10048 18340
rect 5718 18272 5724 18284
rect 2056 18244 3372 18272
rect 5679 18244 5724 18272
rect 2056 18213 2084 18244
rect 1489 18207 1547 18213
rect 1489 18173 1501 18207
rect 1535 18173 1547 18207
rect 1489 18167 1547 18173
rect 2041 18207 2099 18213
rect 2041 18173 2053 18207
rect 2087 18173 2099 18207
rect 2041 18167 2099 18173
rect 1504 18136 1532 18167
rect 2222 18164 2228 18216
rect 2280 18204 2286 18216
rect 2777 18207 2835 18213
rect 2280 18176 2452 18204
rect 2280 18164 2286 18176
rect 2317 18139 2375 18145
rect 2317 18136 2329 18139
rect 1504 18108 2329 18136
rect 2317 18105 2329 18108
rect 2363 18105 2375 18139
rect 2424 18136 2452 18176
rect 2777 18173 2789 18207
rect 2823 18204 2835 18207
rect 3237 18207 3295 18213
rect 3237 18204 3249 18207
rect 2823 18176 3249 18204
rect 2823 18173 2835 18176
rect 2777 18167 2835 18173
rect 3237 18173 3249 18176
rect 3283 18173 3295 18207
rect 3237 18167 3295 18173
rect 3053 18139 3111 18145
rect 3053 18136 3065 18139
rect 2424 18108 3065 18136
rect 2317 18099 2375 18105
rect 3053 18105 3065 18108
rect 3099 18105 3111 18139
rect 3053 18099 3111 18105
rect 566 18028 572 18080
rect 624 18068 630 18080
rect 2682 18068 2688 18080
rect 624 18040 2688 18068
rect 624 18028 630 18040
rect 2682 18028 2688 18040
rect 2740 18028 2746 18080
rect 3344 18068 3372 18244
rect 5718 18232 5724 18244
rect 5776 18232 5782 18284
rect 7469 18275 7527 18281
rect 7469 18241 7481 18275
rect 7515 18272 7527 18275
rect 8110 18272 8116 18284
rect 7515 18244 8116 18272
rect 7515 18241 7527 18244
rect 7469 18235 7527 18241
rect 8110 18232 8116 18244
rect 8168 18232 8174 18284
rect 8386 18272 8392 18284
rect 8347 18244 8392 18272
rect 8386 18232 8392 18244
rect 8444 18232 8450 18284
rect 8573 18275 8631 18281
rect 8573 18241 8585 18275
rect 8619 18272 8631 18275
rect 8846 18272 8852 18284
rect 8619 18244 8852 18272
rect 8619 18241 8631 18244
rect 8573 18235 8631 18241
rect 8846 18232 8852 18244
rect 8904 18232 8910 18284
rect 9600 18281 9628 18312
rect 10042 18300 10048 18312
rect 10100 18300 10106 18352
rect 11606 18300 11612 18352
rect 11664 18340 11670 18352
rect 13078 18340 13084 18352
rect 11664 18312 13084 18340
rect 11664 18300 11670 18312
rect 13078 18300 13084 18312
rect 13136 18300 13142 18352
rect 9585 18275 9643 18281
rect 9585 18241 9597 18275
rect 9631 18241 9643 18275
rect 10229 18275 10287 18281
rect 10229 18272 10241 18275
rect 9585 18235 9643 18241
rect 9692 18244 10241 18272
rect 3513 18207 3571 18213
rect 3513 18173 3525 18207
rect 3559 18204 3571 18207
rect 4062 18204 4068 18216
rect 3559 18176 4068 18204
rect 3559 18173 3571 18176
rect 3513 18167 3571 18173
rect 4062 18164 4068 18176
rect 4120 18164 4126 18216
rect 4154 18164 4160 18216
rect 4212 18204 4218 18216
rect 5629 18207 5687 18213
rect 5629 18204 5641 18207
rect 4212 18176 5641 18204
rect 4212 18164 4218 18176
rect 5629 18173 5641 18176
rect 5675 18173 5687 18207
rect 5629 18167 5687 18173
rect 6181 18207 6239 18213
rect 6181 18173 6193 18207
rect 6227 18204 6239 18207
rect 9692 18204 9720 18244
rect 10229 18241 10241 18244
rect 10275 18241 10287 18275
rect 10229 18235 10287 18241
rect 11146 18232 11152 18284
rect 11204 18232 11210 18284
rect 11517 18275 11575 18281
rect 11517 18241 11529 18275
rect 11563 18272 11575 18275
rect 11790 18272 11796 18284
rect 11563 18244 11796 18272
rect 11563 18241 11575 18244
rect 11517 18235 11575 18241
rect 11790 18232 11796 18244
rect 11848 18232 11854 18284
rect 12986 18272 12992 18284
rect 12947 18244 12992 18272
rect 12986 18232 12992 18244
rect 13044 18272 13050 18284
rect 13906 18272 13912 18284
rect 13044 18244 13912 18272
rect 13044 18232 13050 18244
rect 13906 18232 13912 18244
rect 13964 18272 13970 18284
rect 14001 18275 14059 18281
rect 14001 18272 14013 18275
rect 13964 18244 14013 18272
rect 13964 18232 13970 18244
rect 14001 18241 14013 18244
rect 14047 18241 14059 18275
rect 14001 18235 14059 18241
rect 6227 18176 9720 18204
rect 10045 18207 10103 18213
rect 6227 18173 6239 18176
rect 6181 18167 6239 18173
rect 10045 18173 10057 18207
rect 10091 18204 10103 18207
rect 11164 18204 11192 18232
rect 10091 18176 11192 18204
rect 11885 18207 11943 18213
rect 10091 18173 10103 18176
rect 10045 18167 10103 18173
rect 11885 18173 11897 18207
rect 11931 18204 11943 18207
rect 12805 18207 12863 18213
rect 11931 18176 12296 18204
rect 11931 18173 11943 18176
rect 11885 18167 11943 18173
rect 3780 18139 3838 18145
rect 3780 18105 3792 18139
rect 3826 18136 3838 18139
rect 4798 18136 4804 18148
rect 3826 18108 4804 18136
rect 3826 18105 3838 18108
rect 3780 18099 3838 18105
rect 4798 18096 4804 18108
rect 4856 18096 4862 18148
rect 4890 18096 4896 18148
rect 4948 18136 4954 18148
rect 5537 18139 5595 18145
rect 4948 18108 5212 18136
rect 4948 18096 4954 18108
rect 5184 18077 5212 18108
rect 5537 18105 5549 18139
rect 5583 18136 5595 18139
rect 9122 18136 9128 18148
rect 5583 18108 9128 18136
rect 5583 18105 5595 18108
rect 5537 18099 5595 18105
rect 9122 18096 9128 18108
rect 9180 18096 9186 18148
rect 9401 18139 9459 18145
rect 9401 18105 9413 18139
rect 9447 18136 9459 18139
rect 9674 18136 9680 18148
rect 9447 18108 9680 18136
rect 9447 18105 9459 18108
rect 9401 18099 9459 18105
rect 9674 18096 9680 18108
rect 9732 18096 9738 18148
rect 11333 18139 11391 18145
rect 11333 18105 11345 18139
rect 11379 18136 11391 18139
rect 12268 18136 12296 18176
rect 12805 18173 12817 18207
rect 12851 18204 12863 18207
rect 13170 18204 13176 18216
rect 12851 18176 13176 18204
rect 12851 18173 12863 18176
rect 12805 18167 12863 18173
rect 13170 18164 13176 18176
rect 13228 18204 13234 18216
rect 14461 18207 14519 18213
rect 14461 18204 14473 18207
rect 13228 18176 14473 18204
rect 13228 18164 13234 18176
rect 14461 18173 14473 18176
rect 14507 18173 14519 18207
rect 14461 18167 14519 18173
rect 13817 18139 13875 18145
rect 13817 18136 13829 18139
rect 11379 18108 12112 18136
rect 12268 18108 12664 18136
rect 11379 18105 11391 18108
rect 11333 18099 11391 18105
rect 5077 18071 5135 18077
rect 5077 18068 5089 18071
rect 3344 18040 5089 18068
rect 5077 18037 5089 18040
rect 5123 18037 5135 18071
rect 5077 18031 5135 18037
rect 5169 18071 5227 18077
rect 5169 18037 5181 18071
rect 5215 18037 5227 18071
rect 6362 18068 6368 18080
rect 6323 18040 6368 18068
rect 5169 18031 5227 18037
rect 6362 18028 6368 18040
rect 6420 18028 6426 18080
rect 6454 18028 6460 18080
rect 6512 18068 6518 18080
rect 6825 18071 6883 18077
rect 6825 18068 6837 18071
rect 6512 18040 6837 18068
rect 6512 18028 6518 18040
rect 6825 18037 6837 18040
rect 6871 18037 6883 18071
rect 7190 18068 7196 18080
rect 7151 18040 7196 18068
rect 6825 18031 6883 18037
rect 7190 18028 7196 18040
rect 7248 18028 7254 18080
rect 7282 18028 7288 18080
rect 7340 18068 7346 18080
rect 7340 18040 7385 18068
rect 7340 18028 7346 18040
rect 7466 18028 7472 18080
rect 7524 18068 7530 18080
rect 7929 18071 7987 18077
rect 7929 18068 7941 18071
rect 7524 18040 7941 18068
rect 7524 18028 7530 18040
rect 7929 18037 7941 18040
rect 7975 18037 7987 18071
rect 8294 18068 8300 18080
rect 8255 18040 8300 18068
rect 7929 18031 7987 18037
rect 8294 18028 8300 18040
rect 8352 18028 8358 18080
rect 9493 18071 9551 18077
rect 9493 18037 9505 18071
rect 9539 18068 9551 18071
rect 9950 18068 9956 18080
rect 9539 18040 9956 18068
rect 9539 18037 9551 18040
rect 9493 18031 9551 18037
rect 9950 18028 9956 18040
rect 10008 18028 10014 18080
rect 10870 18068 10876 18080
rect 10831 18040 10876 18068
rect 10870 18028 10876 18040
rect 10928 18028 10934 18080
rect 11054 18028 11060 18080
rect 11112 18068 11118 18080
rect 11241 18071 11299 18077
rect 11241 18068 11253 18071
rect 11112 18040 11253 18068
rect 11112 18028 11118 18040
rect 11241 18037 11253 18040
rect 11287 18037 11299 18071
rect 12084 18068 12112 18108
rect 12434 18068 12440 18080
rect 12084 18040 12440 18068
rect 11241 18031 11299 18037
rect 12434 18028 12440 18040
rect 12492 18028 12498 18080
rect 12636 18068 12664 18108
rect 12789 18108 13829 18136
rect 12789 18068 12817 18108
rect 13817 18105 13829 18108
rect 13863 18105 13875 18139
rect 13817 18099 13875 18105
rect 12636 18040 12817 18068
rect 12894 18028 12900 18080
rect 12952 18068 12958 18080
rect 13538 18068 13544 18080
rect 12952 18040 13544 18068
rect 12952 18028 12958 18040
rect 13538 18028 13544 18040
rect 13596 18028 13602 18080
rect 13909 18071 13967 18077
rect 13909 18037 13921 18071
rect 13955 18068 13967 18071
rect 13998 18068 14004 18080
rect 13955 18040 14004 18068
rect 13955 18037 13967 18040
rect 13909 18031 13967 18037
rect 13998 18028 14004 18040
rect 14056 18028 14062 18080
rect 19518 18028 19524 18080
rect 19576 18068 19582 18080
rect 22554 18068 22560 18080
rect 19576 18040 22560 18068
rect 19576 18028 19582 18040
rect 22554 18028 22560 18040
rect 22612 18028 22618 18080
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 3329 17867 3387 17873
rect 3329 17833 3341 17867
rect 3375 17864 3387 17867
rect 4246 17864 4252 17876
rect 3375 17836 4252 17864
rect 3375 17833 3387 17836
rect 3329 17827 3387 17833
rect 4246 17824 4252 17836
rect 4304 17824 4310 17876
rect 6457 17867 6515 17873
rect 6457 17833 6469 17867
rect 6503 17864 6515 17867
rect 7190 17864 7196 17876
rect 6503 17836 7196 17864
rect 6503 17833 6515 17836
rect 6457 17827 6515 17833
rect 7190 17824 7196 17836
rect 7248 17824 7254 17876
rect 9122 17864 9128 17876
rect 9083 17836 9128 17864
rect 9122 17824 9128 17836
rect 9180 17824 9186 17876
rect 9674 17864 9680 17876
rect 9635 17836 9680 17864
rect 9674 17824 9680 17836
rect 9732 17824 9738 17876
rect 12437 17867 12495 17873
rect 12437 17833 12449 17867
rect 12483 17864 12495 17867
rect 13906 17864 13912 17876
rect 12483 17836 12848 17864
rect 13867 17836 13912 17864
rect 12483 17833 12495 17836
rect 12437 17827 12495 17833
rect 5629 17799 5687 17805
rect 5629 17796 5641 17799
rect 1504 17768 5641 17796
rect 1504 17737 1532 17768
rect 5629 17765 5641 17768
rect 5675 17765 5687 17799
rect 5994 17796 6000 17808
rect 5955 17768 6000 17796
rect 5629 17759 5687 17765
rect 5994 17756 6000 17768
rect 6052 17756 6058 17808
rect 7466 17796 7472 17808
rect 6196 17768 7472 17796
rect 1489 17731 1547 17737
rect 1489 17697 1501 17731
rect 1535 17697 1547 17731
rect 1489 17691 1547 17697
rect 2225 17731 2283 17737
rect 2225 17697 2237 17731
rect 2271 17728 2283 17731
rect 2271 17700 2636 17728
rect 2271 17697 2283 17700
rect 2225 17691 2283 17697
rect 1394 17620 1400 17672
rect 1452 17660 1458 17672
rect 1673 17663 1731 17669
rect 1673 17660 1685 17663
rect 1452 17632 1685 17660
rect 1452 17620 1458 17632
rect 1673 17629 1685 17632
rect 1719 17629 1731 17663
rect 1673 17623 1731 17629
rect 2409 17663 2467 17669
rect 2409 17629 2421 17663
rect 2455 17629 2467 17663
rect 2608 17660 2636 17700
rect 3234 17688 3240 17740
rect 3292 17728 3298 17740
rect 4062 17728 4068 17740
rect 3292 17700 4068 17728
rect 3292 17688 3298 17700
rect 4062 17688 4068 17700
rect 4120 17688 4126 17740
rect 4332 17731 4390 17737
rect 4332 17697 4344 17731
rect 4378 17728 4390 17731
rect 4706 17728 4712 17740
rect 4378 17700 4712 17728
rect 4378 17697 4390 17700
rect 4332 17691 4390 17697
rect 4706 17688 4712 17700
rect 4764 17688 4770 17740
rect 5721 17731 5779 17737
rect 5721 17697 5733 17731
rect 5767 17728 5779 17731
rect 6196 17728 6224 17768
rect 7466 17756 7472 17768
rect 7524 17756 7530 17808
rect 12158 17796 12164 17808
rect 7576 17768 12164 17796
rect 5767 17700 6224 17728
rect 6825 17731 6883 17737
rect 5767 17697 5779 17700
rect 5721 17691 5779 17697
rect 6825 17697 6837 17731
rect 6871 17728 6883 17731
rect 7098 17728 7104 17740
rect 6871 17700 7104 17728
rect 6871 17697 6883 17700
rect 6825 17691 6883 17697
rect 7098 17688 7104 17700
rect 7156 17688 7162 17740
rect 7576 17728 7604 17768
rect 12158 17756 12164 17768
rect 12216 17756 12222 17808
rect 12820 17805 12848 17836
rect 13906 17824 13912 17836
rect 13964 17824 13970 17876
rect 14461 17867 14519 17873
rect 14461 17833 14473 17867
rect 14507 17864 14519 17867
rect 20622 17864 20628 17876
rect 14507 17836 20628 17864
rect 14507 17833 14519 17836
rect 14461 17827 14519 17833
rect 20622 17824 20628 17836
rect 20680 17824 20686 17876
rect 12796 17799 12854 17805
rect 12796 17765 12808 17799
rect 12842 17765 12854 17799
rect 12796 17759 12854 17765
rect 7208 17700 7604 17728
rect 7736 17731 7794 17737
rect 3418 17660 3424 17672
rect 2608 17632 3004 17660
rect 3379 17632 3424 17660
rect 2409 17623 2467 17629
rect 2424 17524 2452 17623
rect 2976 17601 3004 17632
rect 3418 17620 3424 17632
rect 3476 17620 3482 17672
rect 3605 17663 3663 17669
rect 3605 17629 3617 17663
rect 3651 17660 3663 17663
rect 3651 17632 4108 17660
rect 3651 17629 3663 17632
rect 3605 17623 3663 17629
rect 2961 17595 3019 17601
rect 2961 17561 2973 17595
rect 3007 17561 3019 17595
rect 2961 17555 3019 17561
rect 3970 17524 3976 17536
rect 2424 17496 3976 17524
rect 3970 17484 3976 17496
rect 4028 17484 4034 17536
rect 4080 17524 4108 17632
rect 5810 17620 5816 17672
rect 5868 17660 5874 17672
rect 6730 17660 6736 17672
rect 5868 17632 6736 17660
rect 5868 17620 5874 17632
rect 6730 17620 6736 17632
rect 6788 17660 6794 17672
rect 6917 17663 6975 17669
rect 6917 17660 6929 17663
rect 6788 17632 6929 17660
rect 6788 17620 6794 17632
rect 6917 17629 6929 17632
rect 6963 17629 6975 17663
rect 6917 17623 6975 17629
rect 7006 17620 7012 17672
rect 7064 17660 7070 17672
rect 7064 17632 7109 17660
rect 7064 17620 7070 17632
rect 5445 17595 5503 17601
rect 5445 17561 5457 17595
rect 5491 17592 5503 17595
rect 7208 17592 7236 17700
rect 7736 17697 7748 17731
rect 7782 17728 7794 17731
rect 8202 17728 8208 17740
rect 7782 17700 8208 17728
rect 7782 17697 7794 17700
rect 7736 17691 7794 17697
rect 8202 17688 8208 17700
rect 8260 17688 8266 17740
rect 9490 17688 9496 17740
rect 9548 17728 9554 17740
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 9548 17700 10057 17728
rect 9548 17688 9554 17700
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 10045 17691 10103 17697
rect 10134 17688 10140 17740
rect 10192 17728 10198 17740
rect 10192 17700 10237 17728
rect 10192 17688 10198 17700
rect 10410 17688 10416 17740
rect 10468 17728 10474 17740
rect 10873 17731 10931 17737
rect 10873 17728 10885 17731
rect 10468 17700 10885 17728
rect 10468 17688 10474 17700
rect 10873 17697 10885 17700
rect 10919 17697 10931 17731
rect 10873 17691 10931 17697
rect 11140 17731 11198 17737
rect 11140 17697 11152 17731
rect 11186 17728 11198 17731
rect 11698 17728 11704 17740
rect 11186 17700 11704 17728
rect 11186 17697 11198 17700
rect 11140 17691 11198 17697
rect 11698 17688 11704 17700
rect 11756 17688 11762 17740
rect 11974 17688 11980 17740
rect 12032 17728 12038 17740
rect 14277 17731 14335 17737
rect 14277 17728 14289 17731
rect 12032 17700 14289 17728
rect 12032 17688 12038 17700
rect 14277 17697 14289 17700
rect 14323 17697 14335 17731
rect 14277 17691 14335 17697
rect 7466 17660 7472 17672
rect 7427 17632 7472 17660
rect 7466 17620 7472 17632
rect 7524 17620 7530 17672
rect 8478 17620 8484 17672
rect 8536 17660 8542 17672
rect 9858 17660 9864 17672
rect 8536 17632 9864 17660
rect 8536 17620 8542 17632
rect 9858 17620 9864 17632
rect 9916 17620 9922 17672
rect 10321 17663 10379 17669
rect 10321 17629 10333 17663
rect 10367 17660 10379 17663
rect 10502 17660 10508 17672
rect 10367 17632 10508 17660
rect 10367 17629 10379 17632
rect 10321 17623 10379 17629
rect 5491 17564 7236 17592
rect 8849 17595 8907 17601
rect 5491 17561 5503 17564
rect 5445 17555 5503 17561
rect 8849 17561 8861 17595
rect 8895 17592 8907 17595
rect 9674 17592 9680 17604
rect 8895 17564 9680 17592
rect 8895 17561 8907 17564
rect 8849 17555 8907 17561
rect 5460 17524 5488 17555
rect 9674 17552 9680 17564
rect 9732 17592 9738 17604
rect 10336 17592 10364 17623
rect 10502 17620 10508 17632
rect 10560 17620 10566 17672
rect 12066 17620 12072 17672
rect 12124 17660 12130 17672
rect 12526 17660 12532 17672
rect 12124 17632 12532 17660
rect 12124 17620 12130 17632
rect 12526 17620 12532 17632
rect 12584 17620 12590 17672
rect 9732 17564 10364 17592
rect 9732 17552 9738 17564
rect 4080 17496 5488 17524
rect 5629 17527 5687 17533
rect 5629 17493 5641 17527
rect 5675 17524 5687 17527
rect 10870 17524 10876 17536
rect 5675 17496 10876 17524
rect 5675 17493 5687 17496
rect 5629 17487 5687 17493
rect 10870 17484 10876 17496
rect 10928 17484 10934 17536
rect 11790 17484 11796 17536
rect 11848 17524 11854 17536
rect 12253 17527 12311 17533
rect 12253 17524 12265 17527
rect 11848 17496 12265 17524
rect 11848 17484 11854 17496
rect 12253 17493 12265 17496
rect 12299 17524 12311 17527
rect 12345 17527 12403 17533
rect 12345 17524 12357 17527
rect 12299 17496 12357 17524
rect 12299 17493 12311 17496
rect 12253 17487 12311 17493
rect 12345 17493 12357 17496
rect 12391 17493 12403 17527
rect 12345 17487 12403 17493
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 1762 17320 1768 17332
rect 1723 17292 1768 17320
rect 1762 17280 1768 17292
rect 1820 17280 1826 17332
rect 3418 17280 3424 17332
rect 3476 17320 3482 17332
rect 4893 17323 4951 17329
rect 4893 17320 4905 17323
rect 3476 17292 4905 17320
rect 3476 17280 3482 17292
rect 4893 17289 4905 17292
rect 4939 17289 4951 17323
rect 4893 17283 4951 17289
rect 5626 17280 5632 17332
rect 5684 17320 5690 17332
rect 6270 17320 6276 17332
rect 5684 17292 6276 17320
rect 5684 17280 5690 17292
rect 6270 17280 6276 17292
rect 6328 17280 6334 17332
rect 6365 17323 6423 17329
rect 6365 17289 6377 17323
rect 6411 17320 6423 17323
rect 8202 17320 8208 17332
rect 6411 17292 7779 17320
rect 8163 17292 8208 17320
rect 6411 17289 6423 17292
rect 6365 17283 6423 17289
rect 4617 17255 4675 17261
rect 4617 17221 4629 17255
rect 4663 17252 4675 17255
rect 4706 17252 4712 17264
rect 4663 17224 4712 17252
rect 4663 17221 4675 17224
rect 4617 17215 4675 17221
rect 4706 17212 4712 17224
rect 4764 17252 4770 17264
rect 4764 17224 5488 17252
rect 4764 17212 4770 17224
rect 3234 17184 3240 17196
rect 2148 17156 2728 17184
rect 3195 17156 3240 17184
rect 1578 17116 1584 17128
rect 1539 17088 1584 17116
rect 1578 17076 1584 17088
rect 1636 17076 1642 17128
rect 2148 17125 2176 17156
rect 2143 17119 2201 17125
rect 2143 17085 2155 17119
rect 2189 17085 2201 17119
rect 2143 17079 2201 17085
rect 2314 17008 2320 17060
rect 2372 17048 2378 17060
rect 2409 17051 2467 17057
rect 2409 17048 2421 17051
rect 2372 17020 2421 17048
rect 2372 17008 2378 17020
rect 2409 17017 2421 17020
rect 2455 17017 2467 17051
rect 2700 17048 2728 17156
rect 3234 17144 3240 17156
rect 3292 17144 3298 17196
rect 5166 17144 5172 17196
rect 5224 17184 5230 17196
rect 5460 17193 5488 17224
rect 5534 17212 5540 17264
rect 5592 17252 5598 17264
rect 6089 17255 6147 17261
rect 6089 17252 6101 17255
rect 5592 17224 6101 17252
rect 5592 17212 5598 17224
rect 6089 17221 6101 17224
rect 6135 17221 6147 17255
rect 7751 17252 7779 17292
rect 8202 17280 8208 17292
rect 8260 17280 8266 17332
rect 10042 17320 10048 17332
rect 8680 17292 9628 17320
rect 10003 17292 10048 17320
rect 8680 17252 8708 17292
rect 7751 17224 8708 17252
rect 9600 17252 9628 17292
rect 10042 17280 10048 17292
rect 10100 17280 10106 17332
rect 11698 17320 11704 17332
rect 10152 17292 11468 17320
rect 11659 17292 11704 17320
rect 10152 17252 10180 17292
rect 11440 17264 11468 17292
rect 11698 17280 11704 17292
rect 11756 17280 11762 17332
rect 12434 17280 12440 17332
rect 12492 17320 12498 17332
rect 13633 17323 13691 17329
rect 12492 17292 12537 17320
rect 12492 17280 12498 17292
rect 13633 17289 13645 17323
rect 13679 17320 13691 17323
rect 13814 17320 13820 17332
rect 13679 17292 13820 17320
rect 13679 17289 13691 17292
rect 13633 17283 13691 17289
rect 13814 17280 13820 17292
rect 13872 17280 13878 17332
rect 14185 17323 14243 17329
rect 14185 17289 14197 17323
rect 14231 17320 14243 17323
rect 19334 17320 19340 17332
rect 14231 17292 19340 17320
rect 14231 17289 14243 17292
rect 14185 17283 14243 17289
rect 19334 17280 19340 17292
rect 19392 17280 19398 17332
rect 9600 17224 10180 17252
rect 6089 17215 6147 17221
rect 11422 17212 11428 17264
rect 11480 17212 11486 17264
rect 5353 17187 5411 17193
rect 5353 17184 5365 17187
rect 5224 17156 5365 17184
rect 5224 17144 5230 17156
rect 5353 17153 5365 17156
rect 5399 17153 5411 17187
rect 5353 17147 5411 17153
rect 5445 17187 5503 17193
rect 5445 17153 5457 17187
rect 5491 17153 5503 17187
rect 6454 17184 6460 17196
rect 5445 17147 5503 17153
rect 5552 17156 6460 17184
rect 5552 17116 5580 17156
rect 6454 17144 6460 17156
rect 6512 17144 6518 17196
rect 10042 17144 10048 17196
rect 10100 17184 10106 17196
rect 10100 17156 10456 17184
rect 10100 17144 10106 17156
rect 5902 17116 5908 17128
rect 3436 17088 5580 17116
rect 5863 17088 5908 17116
rect 3436 17048 3464 17088
rect 5902 17076 5908 17088
rect 5960 17076 5966 17128
rect 6641 17119 6699 17125
rect 6641 17085 6653 17119
rect 6687 17116 6699 17119
rect 6730 17116 6736 17128
rect 6687 17088 6736 17116
rect 6687 17085 6699 17088
rect 6641 17079 6699 17085
rect 6730 17076 6736 17088
rect 6788 17076 6794 17128
rect 6822 17076 6828 17128
rect 6880 17116 6886 17128
rect 7466 17116 7472 17128
rect 6880 17088 7472 17116
rect 6880 17076 6886 17088
rect 7466 17076 7472 17088
rect 7524 17116 7530 17128
rect 8662 17116 8668 17128
rect 7524 17088 8668 17116
rect 7524 17076 7530 17088
rect 8662 17076 8668 17088
rect 8720 17076 8726 17128
rect 8932 17119 8990 17125
rect 8932 17085 8944 17119
rect 8978 17116 8990 17119
rect 9674 17116 9680 17128
rect 8978 17088 9680 17116
rect 8978 17085 8990 17088
rect 8932 17079 8990 17085
rect 9674 17076 9680 17088
rect 9732 17076 9738 17128
rect 10318 17116 10324 17128
rect 10279 17088 10324 17116
rect 10318 17076 10324 17088
rect 10376 17076 10382 17128
rect 10428 17116 10456 17156
rect 11698 17144 11704 17196
rect 11756 17184 11762 17196
rect 12989 17187 13047 17193
rect 12989 17184 13001 17187
rect 11756 17156 13001 17184
rect 11756 17144 11762 17156
rect 12989 17153 13001 17156
rect 13035 17153 13047 17187
rect 12989 17147 13047 17153
rect 13372 17156 14044 17184
rect 10577 17119 10635 17125
rect 10577 17116 10589 17119
rect 10428 17088 10589 17116
rect 10577 17085 10589 17088
rect 10623 17085 10635 17119
rect 10577 17079 10635 17085
rect 10870 17076 10876 17128
rect 10928 17116 10934 17128
rect 11974 17116 11980 17128
rect 10928 17088 11980 17116
rect 10928 17076 10934 17088
rect 11974 17076 11980 17088
rect 12032 17076 12038 17128
rect 12158 17116 12164 17128
rect 12119 17088 12164 17116
rect 12158 17076 12164 17088
rect 12216 17076 12222 17128
rect 12802 17076 12808 17128
rect 12860 17116 12866 17128
rect 13372 17116 13400 17156
rect 14016 17125 14044 17156
rect 12860 17088 13400 17116
rect 13449 17119 13507 17125
rect 12860 17076 12866 17088
rect 13449 17085 13461 17119
rect 13495 17085 13507 17119
rect 13449 17079 13507 17085
rect 14001 17119 14059 17125
rect 14001 17085 14013 17119
rect 14047 17085 14059 17119
rect 14001 17079 14059 17085
rect 2700 17020 3464 17048
rect 3504 17051 3562 17057
rect 2409 17011 2467 17017
rect 3504 17017 3516 17051
rect 3550 17048 3562 17051
rect 3602 17048 3608 17060
rect 3550 17020 3608 17048
rect 3550 17017 3562 17020
rect 3504 17011 3562 17017
rect 3602 17008 3608 17020
rect 3660 17008 3666 17060
rect 3786 17008 3792 17060
rect 3844 17048 3850 17060
rect 4798 17048 4804 17060
rect 3844 17020 4804 17048
rect 3844 17008 3850 17020
rect 4798 17008 4804 17020
rect 4856 17008 4862 17060
rect 7081 17051 7139 17057
rect 5184 17020 6960 17048
rect 1670 16940 1676 16992
rect 1728 16980 1734 16992
rect 5184 16980 5212 17020
rect 1728 16952 5212 16980
rect 1728 16940 1734 16952
rect 5258 16940 5264 16992
rect 5316 16980 5322 16992
rect 6365 16983 6423 16989
rect 6365 16980 6377 16983
rect 5316 16952 6377 16980
rect 5316 16940 5322 16952
rect 6365 16949 6377 16952
rect 6411 16949 6423 16983
rect 6365 16943 6423 16949
rect 6457 16983 6515 16989
rect 6457 16949 6469 16983
rect 6503 16980 6515 16983
rect 6822 16980 6828 16992
rect 6503 16952 6828 16980
rect 6503 16949 6515 16952
rect 6457 16943 6515 16949
rect 6822 16940 6828 16952
rect 6880 16940 6886 16992
rect 6932 16980 6960 17020
rect 7081 17017 7093 17051
rect 7127 17048 7139 17051
rect 7374 17048 7380 17060
rect 7127 17020 7380 17048
rect 7127 17017 7139 17020
rect 7081 17011 7139 17017
rect 7374 17008 7380 17020
rect 7432 17008 7438 17060
rect 12250 17048 12256 17060
rect 7751 17020 12256 17048
rect 7751 16980 7779 17020
rect 12250 17008 12256 17020
rect 12308 17008 12314 17060
rect 13464 17048 13492 17079
rect 14550 17048 14556 17060
rect 13464 17020 14556 17048
rect 14550 17008 14556 17020
rect 14608 17008 14614 17060
rect 6932 16952 7779 16980
rect 8202 16940 8208 16992
rect 8260 16980 8266 16992
rect 9674 16980 9680 16992
rect 8260 16952 9680 16980
rect 8260 16940 8266 16952
rect 9674 16940 9680 16952
rect 9732 16940 9738 16992
rect 10318 16940 10324 16992
rect 10376 16980 10382 16992
rect 11977 16983 12035 16989
rect 11977 16980 11989 16983
rect 10376 16952 11989 16980
rect 10376 16940 10382 16952
rect 11977 16949 11989 16952
rect 12023 16980 12035 16983
rect 12066 16980 12072 16992
rect 12023 16952 12072 16980
rect 12023 16949 12035 16952
rect 11977 16943 12035 16949
rect 12066 16940 12072 16952
rect 12124 16940 12130 16992
rect 12802 16980 12808 16992
rect 12763 16952 12808 16980
rect 12802 16940 12808 16952
rect 12860 16940 12866 16992
rect 12897 16983 12955 16989
rect 12897 16949 12909 16983
rect 12943 16980 12955 16983
rect 13078 16980 13084 16992
rect 12943 16952 13084 16980
rect 12943 16949 12955 16952
rect 12897 16943 12955 16949
rect 13078 16940 13084 16952
rect 13136 16940 13142 16992
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 1854 16776 1860 16788
rect 1815 16748 1860 16776
rect 1854 16736 1860 16748
rect 1912 16736 1918 16788
rect 2958 16736 2964 16788
rect 3016 16776 3022 16788
rect 3418 16776 3424 16788
rect 3016 16748 3424 16776
rect 3016 16736 3022 16748
rect 3418 16736 3424 16748
rect 3476 16736 3482 16788
rect 3970 16736 3976 16788
rect 4028 16776 4034 16788
rect 6178 16776 6184 16788
rect 4028 16748 6184 16776
rect 4028 16736 4034 16748
rect 6178 16736 6184 16748
rect 6236 16736 6242 16788
rect 7282 16736 7288 16788
rect 7340 16776 7346 16788
rect 8113 16779 8171 16785
rect 8113 16776 8125 16779
rect 7340 16748 8125 16776
rect 7340 16736 7346 16748
rect 8113 16745 8125 16748
rect 8159 16745 8171 16779
rect 8113 16739 8171 16745
rect 8294 16736 8300 16788
rect 8352 16776 8358 16788
rect 9125 16779 9183 16785
rect 9125 16776 9137 16779
rect 8352 16748 9137 16776
rect 8352 16736 8358 16748
rect 9125 16745 9137 16748
rect 9171 16745 9183 16779
rect 9950 16776 9956 16788
rect 9911 16748 9956 16776
rect 9125 16739 9183 16745
rect 9950 16736 9956 16748
rect 10008 16736 10014 16788
rect 10321 16779 10379 16785
rect 10321 16745 10333 16779
rect 10367 16776 10379 16779
rect 10870 16776 10876 16788
rect 10367 16748 10876 16776
rect 10367 16745 10379 16748
rect 10321 16739 10379 16745
rect 10870 16736 10876 16748
rect 10928 16736 10934 16788
rect 10965 16779 11023 16785
rect 10965 16745 10977 16779
rect 11011 16776 11023 16779
rect 11054 16776 11060 16788
rect 11011 16748 11060 16776
rect 11011 16745 11023 16748
rect 10965 16739 11023 16745
rect 11054 16736 11060 16748
rect 11112 16736 11118 16788
rect 11164 16748 14320 16776
rect 1578 16668 1584 16720
rect 1636 16708 1642 16720
rect 2501 16711 2559 16717
rect 2501 16708 2513 16711
rect 1636 16680 2513 16708
rect 1636 16668 1642 16680
rect 2501 16677 2513 16680
rect 2547 16677 2559 16711
rect 2501 16671 2559 16677
rect 3142 16668 3148 16720
rect 3200 16708 3206 16720
rect 3329 16711 3387 16717
rect 3329 16708 3341 16711
rect 3200 16680 3341 16708
rect 3200 16668 3206 16680
rect 3329 16677 3341 16680
rect 3375 16677 3387 16711
rect 3329 16671 3387 16677
rect 3510 16668 3516 16720
rect 3568 16708 3574 16720
rect 6822 16708 6828 16720
rect 3568 16680 4108 16708
rect 3568 16668 3574 16680
rect 1670 16640 1676 16652
rect 1631 16612 1676 16640
rect 1670 16600 1676 16612
rect 1728 16600 1734 16652
rect 4080 16649 4108 16680
rect 6288 16680 6828 16708
rect 2225 16643 2283 16649
rect 2225 16609 2237 16643
rect 2271 16609 2283 16643
rect 2225 16603 2283 16609
rect 4065 16643 4123 16649
rect 4065 16609 4077 16643
rect 4111 16609 4123 16643
rect 4065 16603 4123 16609
rect 2240 16504 2268 16603
rect 4246 16600 4252 16652
rect 4304 16640 4310 16652
rect 4617 16643 4675 16649
rect 4617 16640 4629 16643
rect 4304 16612 4629 16640
rect 4304 16600 4310 16612
rect 4617 16609 4629 16612
rect 4663 16609 4675 16643
rect 4617 16603 4675 16609
rect 4884 16643 4942 16649
rect 4884 16609 4896 16643
rect 4930 16640 4942 16643
rect 5810 16640 5816 16652
rect 4930 16612 5816 16640
rect 4930 16609 4942 16612
rect 4884 16603 4942 16609
rect 5810 16600 5816 16612
rect 5868 16600 5874 16652
rect 6288 16649 6316 16680
rect 6822 16668 6828 16680
rect 6880 16668 6886 16720
rect 7190 16668 7196 16720
rect 7248 16708 7254 16720
rect 7248 16680 10088 16708
rect 7248 16668 7254 16680
rect 6546 16649 6552 16652
rect 6273 16643 6331 16649
rect 6273 16609 6285 16643
rect 6319 16609 6331 16643
rect 6540 16640 6552 16649
rect 6507 16612 6552 16640
rect 6273 16603 6331 16609
rect 6540 16603 6552 16612
rect 6546 16600 6552 16603
rect 6604 16600 6610 16652
rect 7006 16600 7012 16652
rect 7064 16640 7070 16652
rect 7374 16640 7380 16652
rect 7064 16612 7380 16640
rect 7064 16600 7070 16612
rect 7374 16600 7380 16612
rect 7432 16640 7438 16652
rect 8478 16640 8484 16652
rect 7432 16612 7779 16640
rect 8439 16612 8484 16640
rect 7432 16600 7438 16612
rect 2682 16532 2688 16584
rect 2740 16572 2746 16584
rect 3234 16572 3240 16584
rect 2740 16544 3240 16572
rect 2740 16532 2746 16544
rect 3234 16532 3240 16544
rect 3292 16532 3298 16584
rect 3605 16575 3663 16581
rect 3605 16541 3617 16575
rect 3651 16572 3663 16575
rect 3786 16572 3792 16584
rect 3651 16544 3792 16572
rect 3651 16541 3663 16544
rect 3605 16535 3663 16541
rect 3786 16532 3792 16544
rect 3844 16532 3850 16584
rect 3418 16504 3424 16516
rect 2240 16476 3424 16504
rect 3418 16464 3424 16476
rect 3476 16464 3482 16516
rect 3694 16464 3700 16516
rect 3752 16504 3758 16516
rect 7637 16513 7665 16612
rect 7751 16572 7779 16612
rect 8478 16600 8484 16612
rect 8536 16600 8542 16652
rect 8573 16643 8631 16649
rect 8573 16609 8585 16643
rect 8619 16640 8631 16643
rect 9950 16640 9956 16652
rect 8619 16612 9956 16640
rect 8619 16609 8631 16612
rect 8573 16603 8631 16609
rect 9950 16600 9956 16612
rect 10008 16600 10014 16652
rect 10060 16640 10088 16680
rect 10134 16668 10140 16720
rect 10192 16708 10198 16720
rect 11164 16708 11192 16748
rect 10192 16680 11192 16708
rect 11333 16711 11391 16717
rect 10192 16668 10198 16680
rect 11333 16677 11345 16711
rect 11379 16708 11391 16711
rect 12066 16708 12072 16720
rect 11379 16680 12072 16708
rect 11379 16677 11391 16680
rect 11333 16671 11391 16677
rect 12066 16668 12072 16680
rect 12124 16668 12130 16720
rect 12176 16680 14228 16708
rect 10413 16643 10471 16649
rect 10060 16612 10364 16640
rect 8665 16575 8723 16581
rect 8665 16572 8677 16575
rect 7751 16544 8677 16572
rect 8665 16541 8677 16544
rect 8711 16541 8723 16575
rect 8665 16535 8723 16541
rect 9674 16532 9680 16584
rect 9732 16572 9738 16584
rect 9732 16544 9904 16572
rect 9732 16532 9738 16544
rect 4249 16507 4307 16513
rect 4249 16504 4261 16507
rect 3752 16476 4261 16504
rect 3752 16464 3758 16476
rect 4249 16473 4261 16476
rect 4295 16473 4307 16507
rect 7637 16507 7711 16513
rect 7637 16476 7665 16507
rect 4249 16467 4307 16473
rect 7653 16473 7665 16476
rect 7699 16473 7711 16507
rect 7653 16467 7711 16473
rect 8846 16464 8852 16516
rect 8904 16504 8910 16516
rect 9766 16504 9772 16516
rect 8904 16476 9772 16504
rect 8904 16464 8910 16476
rect 9766 16464 9772 16476
rect 9824 16464 9830 16516
rect 9876 16504 9904 16544
rect 10336 16504 10364 16612
rect 10413 16609 10425 16643
rect 10459 16640 10471 16643
rect 11146 16640 11152 16652
rect 10459 16612 11152 16640
rect 10459 16609 10471 16612
rect 10413 16603 10471 16609
rect 11146 16600 11152 16612
rect 11204 16640 11210 16652
rect 11790 16640 11796 16652
rect 11204 16612 11796 16640
rect 11204 16600 11210 16612
rect 11790 16600 11796 16612
rect 11848 16600 11854 16652
rect 11977 16643 12035 16649
rect 11977 16640 11989 16643
rect 11900 16612 11989 16640
rect 10502 16572 10508 16584
rect 10463 16544 10508 16572
rect 10502 16532 10508 16544
rect 10560 16532 10566 16584
rect 11422 16572 11428 16584
rect 11383 16544 11428 16572
rect 11422 16532 11428 16544
rect 11480 16532 11486 16584
rect 11609 16575 11667 16581
rect 11609 16541 11621 16575
rect 11655 16572 11667 16575
rect 11698 16572 11704 16584
rect 11655 16544 11704 16572
rect 11655 16541 11667 16544
rect 11609 16535 11667 16541
rect 11698 16532 11704 16544
rect 11756 16532 11762 16584
rect 11900 16504 11928 16612
rect 11977 16609 11989 16612
rect 12023 16609 12035 16643
rect 11977 16603 12035 16609
rect 12176 16513 12204 16680
rect 12526 16600 12532 16652
rect 12584 16640 12590 16652
rect 12894 16649 12900 16652
rect 12621 16643 12679 16649
rect 12621 16640 12633 16643
rect 12584 16612 12633 16640
rect 12584 16600 12590 16612
rect 12621 16609 12633 16612
rect 12667 16609 12679 16643
rect 12888 16640 12900 16649
rect 12855 16612 12900 16640
rect 12621 16603 12679 16609
rect 12888 16603 12900 16612
rect 12894 16600 12900 16603
rect 12952 16600 12958 16652
rect 14200 16572 14228 16680
rect 14292 16649 14320 16748
rect 14550 16708 14556 16720
rect 14511 16680 14556 16708
rect 14550 16668 14556 16680
rect 14608 16668 14614 16720
rect 14277 16643 14335 16649
rect 14277 16609 14289 16643
rect 14323 16609 14335 16643
rect 19426 16640 19432 16652
rect 14277 16603 14335 16609
rect 19260 16612 19432 16640
rect 19260 16572 19288 16612
rect 19426 16600 19432 16612
rect 19484 16600 19490 16652
rect 14200 16544 19288 16572
rect 9876 16476 10088 16504
rect 10336 16476 11928 16504
rect 12161 16507 12219 16513
rect 2958 16436 2964 16448
rect 2919 16408 2964 16436
rect 2958 16396 2964 16408
rect 3016 16396 3022 16448
rect 3326 16396 3332 16448
rect 3384 16436 3390 16448
rect 5258 16436 5264 16448
rect 3384 16408 5264 16436
rect 3384 16396 3390 16408
rect 5258 16396 5264 16408
rect 5316 16396 5322 16448
rect 5994 16436 6000 16448
rect 5955 16408 6000 16436
rect 5994 16396 6000 16408
rect 6052 16396 6058 16448
rect 6454 16396 6460 16448
rect 6512 16436 6518 16448
rect 9950 16436 9956 16448
rect 6512 16408 9956 16436
rect 6512 16396 6518 16408
rect 9950 16396 9956 16408
rect 10008 16396 10014 16448
rect 10060 16436 10088 16476
rect 12161 16473 12173 16507
rect 12207 16473 12219 16507
rect 12161 16467 12219 16473
rect 14001 16439 14059 16445
rect 14001 16436 14013 16439
rect 10060 16408 14013 16436
rect 14001 16405 14013 16408
rect 14047 16405 14059 16439
rect 14001 16399 14059 16405
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 1946 16232 1952 16244
rect 1907 16204 1952 16232
rect 1946 16192 1952 16204
rect 2004 16192 2010 16244
rect 2501 16235 2559 16241
rect 2501 16201 2513 16235
rect 2547 16232 2559 16235
rect 2774 16232 2780 16244
rect 2547 16204 2780 16232
rect 2547 16201 2559 16204
rect 2501 16195 2559 16201
rect 2774 16192 2780 16204
rect 2832 16192 2838 16244
rect 3050 16192 3056 16244
rect 3108 16232 3114 16244
rect 3510 16232 3516 16244
rect 3108 16204 3516 16232
rect 3108 16192 3114 16204
rect 3510 16192 3516 16204
rect 3568 16192 3574 16244
rect 3694 16192 3700 16244
rect 3752 16232 3758 16244
rect 6454 16232 6460 16244
rect 3752 16204 6460 16232
rect 3752 16192 3758 16204
rect 6454 16192 6460 16204
rect 6512 16192 6518 16244
rect 7929 16235 7987 16241
rect 7929 16201 7941 16235
rect 7975 16232 7987 16235
rect 10045 16235 10103 16241
rect 10045 16232 10057 16235
rect 7975 16204 10057 16232
rect 7975 16201 7987 16204
rect 7929 16195 7987 16201
rect 10045 16201 10057 16204
rect 10091 16201 10103 16235
rect 10045 16195 10103 16201
rect 10134 16192 10140 16244
rect 10192 16232 10198 16244
rect 10192 16204 10237 16232
rect 10192 16192 10198 16204
rect 2961 16167 3019 16173
rect 2961 16133 2973 16167
rect 3007 16164 3019 16167
rect 6822 16164 6828 16176
rect 3007 16136 6828 16164
rect 3007 16133 3019 16136
rect 2961 16127 3019 16133
rect 6822 16124 6828 16136
rect 6880 16124 6886 16176
rect 11149 16167 11207 16173
rect 11149 16164 11161 16167
rect 8404 16136 11161 16164
rect 3605 16099 3663 16105
rect 3605 16065 3617 16099
rect 3651 16096 3663 16099
rect 3786 16096 3792 16108
rect 3651 16068 3792 16096
rect 3651 16065 3663 16068
rect 3605 16059 3663 16065
rect 3786 16056 3792 16068
rect 3844 16056 3850 16108
rect 4062 16056 4068 16108
rect 4120 16096 4126 16108
rect 4522 16096 4528 16108
rect 4120 16068 4528 16096
rect 4120 16056 4126 16068
rect 4522 16056 4528 16068
rect 4580 16056 4586 16108
rect 4617 16099 4675 16105
rect 4617 16065 4629 16099
rect 4663 16096 4675 16099
rect 5350 16096 5356 16108
rect 4663 16068 5356 16096
rect 4663 16065 4675 16068
rect 4617 16059 4675 16065
rect 5350 16056 5356 16068
rect 5408 16056 5414 16108
rect 5810 16096 5816 16108
rect 5723 16068 5816 16096
rect 5810 16056 5816 16068
rect 5868 16096 5874 16108
rect 7469 16099 7527 16105
rect 7469 16096 7481 16099
rect 5868 16068 7481 16096
rect 5868 16056 5874 16068
rect 7469 16065 7481 16068
rect 7515 16096 7527 16099
rect 8202 16096 8208 16108
rect 7515 16068 8208 16096
rect 7515 16065 7527 16068
rect 7469 16059 7527 16065
rect 8202 16056 8208 16068
rect 8260 16056 8266 16108
rect 8404 16105 8432 16136
rect 11149 16133 11161 16136
rect 11195 16133 11207 16167
rect 14182 16164 14188 16176
rect 11149 16127 11207 16133
rect 13280 16136 14188 16164
rect 8389 16099 8447 16105
rect 8389 16065 8401 16099
rect 8435 16065 8447 16099
rect 8389 16059 8447 16065
rect 8573 16099 8631 16105
rect 8573 16065 8585 16099
rect 8619 16096 8631 16099
rect 9306 16096 9312 16108
rect 8619 16068 9312 16096
rect 8619 16065 8631 16068
rect 8573 16059 8631 16065
rect 9306 16056 9312 16068
rect 9364 16096 9370 16108
rect 9677 16099 9735 16105
rect 9677 16096 9689 16099
rect 9364 16068 9689 16096
rect 9364 16056 9370 16068
rect 9677 16065 9689 16068
rect 9723 16065 9735 16099
rect 9677 16059 9735 16065
rect 10045 16099 10103 16105
rect 10045 16065 10057 16099
rect 10091 16096 10103 16099
rect 10597 16099 10655 16105
rect 10597 16096 10609 16099
rect 10091 16068 10609 16096
rect 10091 16065 10103 16068
rect 10045 16059 10103 16065
rect 10597 16065 10609 16068
rect 10643 16065 10655 16099
rect 10597 16059 10655 16065
rect 10781 16099 10839 16105
rect 10781 16065 10793 16099
rect 10827 16096 10839 16099
rect 10962 16096 10968 16108
rect 10827 16068 10968 16096
rect 10827 16065 10839 16068
rect 10781 16059 10839 16065
rect 10962 16056 10968 16068
rect 11020 16056 11026 16108
rect 11701 16099 11759 16105
rect 11701 16096 11713 16099
rect 11072 16068 11713 16096
rect 1762 16028 1768 16040
rect 1723 16000 1768 16028
rect 1762 15988 1768 16000
rect 1820 15988 1826 16040
rect 2314 16028 2320 16040
rect 2275 16000 2320 16028
rect 2314 15988 2320 16000
rect 2372 15988 2378 16040
rect 3421 16031 3479 16037
rect 3421 15997 3433 16031
rect 3467 16028 3479 16031
rect 4982 16028 4988 16040
rect 3467 16000 4988 16028
rect 3467 15997 3479 16000
rect 3421 15991 3479 15997
rect 2590 15920 2596 15972
rect 2648 15960 2654 15972
rect 3436 15960 3464 15991
rect 4982 15988 4988 16000
rect 5040 15988 5046 16040
rect 5258 15988 5264 16040
rect 5316 16028 5322 16040
rect 5629 16031 5687 16037
rect 5629 16028 5641 16031
rect 5316 16000 5641 16028
rect 5316 15988 5322 16000
rect 5629 15997 5641 16000
rect 5675 15997 5687 16031
rect 5629 15991 5687 15997
rect 6206 16031 6264 16037
rect 6206 15997 6218 16031
rect 6252 16028 6264 16031
rect 6454 16028 6460 16040
rect 6252 16000 6460 16028
rect 6252 15997 6264 16000
rect 6206 15991 6264 15997
rect 6454 15988 6460 16000
rect 6512 15988 6518 16040
rect 7190 16028 7196 16040
rect 7151 16000 7196 16028
rect 7190 15988 7196 16000
rect 7248 15988 7254 16040
rect 9493 16031 9551 16037
rect 9493 15997 9505 16031
rect 9539 16028 9551 16031
rect 9766 16028 9772 16040
rect 9539 16000 9772 16028
rect 9539 15997 9551 16000
rect 9493 15991 9551 15997
rect 9766 15988 9772 16000
rect 9824 15988 9830 16040
rect 9950 15988 9956 16040
rect 10008 16028 10014 16040
rect 10008 16000 10620 16028
rect 10008 15988 10014 16000
rect 2648 15932 3464 15960
rect 2648 15920 2654 15932
rect 3510 15920 3516 15972
rect 3568 15960 3574 15972
rect 4062 15960 4068 15972
rect 3568 15932 4068 15960
rect 3568 15920 3574 15932
rect 4062 15920 4068 15932
rect 4120 15920 4126 15972
rect 4341 15963 4399 15969
rect 4341 15929 4353 15963
rect 4387 15960 4399 15963
rect 5810 15960 5816 15972
rect 4387 15932 5816 15960
rect 4387 15929 4399 15932
rect 4341 15923 4399 15929
rect 5810 15920 5816 15932
rect 5868 15920 5874 15972
rect 8297 15963 8355 15969
rect 8297 15960 8309 15963
rect 5920 15932 8309 15960
rect 2498 15852 2504 15904
rect 2556 15892 2562 15904
rect 3329 15895 3387 15901
rect 3329 15892 3341 15895
rect 2556 15864 3341 15892
rect 2556 15852 2562 15864
rect 3329 15861 3341 15864
rect 3375 15892 3387 15895
rect 3602 15892 3608 15904
rect 3375 15864 3608 15892
rect 3375 15861 3387 15864
rect 3329 15855 3387 15861
rect 3602 15852 3608 15864
rect 3660 15852 3666 15904
rect 3973 15895 4031 15901
rect 3973 15861 3985 15895
rect 4019 15892 4031 15895
rect 4246 15892 4252 15904
rect 4019 15864 4252 15892
rect 4019 15861 4031 15864
rect 3973 15855 4031 15861
rect 4246 15852 4252 15864
rect 4304 15852 4310 15904
rect 4430 15892 4436 15904
rect 4391 15864 4436 15892
rect 4430 15852 4436 15864
rect 4488 15852 4494 15904
rect 5169 15895 5227 15901
rect 5169 15861 5181 15895
rect 5215 15892 5227 15895
rect 5258 15892 5264 15904
rect 5215 15864 5264 15892
rect 5215 15861 5227 15864
rect 5169 15855 5227 15861
rect 5258 15852 5264 15864
rect 5316 15852 5322 15904
rect 5534 15892 5540 15904
rect 5495 15864 5540 15892
rect 5534 15852 5540 15864
rect 5592 15852 5598 15904
rect 5718 15852 5724 15904
rect 5776 15892 5782 15904
rect 5920 15892 5948 15932
rect 8297 15929 8309 15932
rect 8343 15929 8355 15963
rect 10505 15963 10563 15969
rect 10505 15960 10517 15963
rect 8297 15923 8355 15929
rect 9140 15932 10517 15960
rect 5776 15864 5948 15892
rect 5776 15852 5782 15864
rect 6178 15852 6184 15904
rect 6236 15892 6242 15904
rect 6365 15895 6423 15901
rect 6365 15892 6377 15895
rect 6236 15864 6377 15892
rect 6236 15852 6242 15864
rect 6365 15861 6377 15864
rect 6411 15861 6423 15895
rect 6822 15892 6828 15904
rect 6783 15864 6828 15892
rect 6365 15855 6423 15861
rect 6822 15852 6828 15864
rect 6880 15852 6886 15904
rect 7285 15895 7343 15901
rect 7285 15861 7297 15895
rect 7331 15892 7343 15895
rect 8846 15892 8852 15904
rect 7331 15864 8852 15892
rect 7331 15861 7343 15864
rect 7285 15855 7343 15861
rect 8846 15852 8852 15864
rect 8904 15852 8910 15904
rect 9140 15901 9168 15932
rect 10505 15929 10517 15932
rect 10551 15929 10563 15963
rect 10505 15923 10563 15929
rect 9125 15895 9183 15901
rect 9125 15861 9137 15895
rect 9171 15861 9183 15895
rect 9125 15855 9183 15861
rect 9585 15895 9643 15901
rect 9585 15861 9597 15895
rect 9631 15892 9643 15895
rect 10042 15892 10048 15904
rect 9631 15864 10048 15892
rect 9631 15861 9643 15864
rect 9585 15855 9643 15861
rect 10042 15852 10048 15864
rect 10100 15852 10106 15904
rect 10592 15892 10620 16000
rect 10870 15988 10876 16040
rect 10928 16028 10934 16040
rect 11072 16028 11100 16068
rect 11701 16065 11713 16068
rect 11747 16065 11759 16099
rect 11701 16059 11759 16065
rect 12066 16056 12072 16108
rect 12124 16096 12130 16108
rect 12434 16096 12440 16108
rect 12124 16068 12440 16096
rect 12124 16056 12130 16068
rect 12434 16056 12440 16068
rect 12492 16056 12498 16108
rect 13280 16105 13308 16136
rect 14182 16124 14188 16136
rect 14240 16124 14246 16176
rect 13265 16099 13323 16105
rect 13265 16065 13277 16099
rect 13311 16065 13323 16099
rect 13814 16096 13820 16108
rect 13775 16068 13820 16096
rect 13265 16059 13323 16065
rect 13814 16056 13820 16068
rect 13872 16056 13878 16108
rect 11514 16028 11520 16040
rect 10928 16000 11100 16028
rect 11475 16000 11520 16028
rect 10928 15988 10934 16000
rect 11514 15988 11520 16000
rect 11572 15988 11578 16040
rect 11606 15988 11612 16040
rect 11664 16028 11670 16040
rect 13633 16031 13691 16037
rect 13633 16028 13645 16031
rect 11664 16000 13645 16028
rect 11664 15988 11670 16000
rect 13633 15997 13645 16000
rect 13679 15997 13691 16031
rect 13633 15991 13691 15997
rect 10686 15920 10692 15972
rect 10744 15960 10750 15972
rect 13081 15963 13139 15969
rect 13081 15960 13093 15963
rect 10744 15932 13093 15960
rect 10744 15920 10750 15932
rect 13081 15929 13093 15932
rect 13127 15929 13139 15963
rect 13081 15923 13139 15929
rect 11609 15895 11667 15901
rect 11609 15892 11621 15895
rect 10592 15864 11621 15892
rect 11609 15861 11621 15864
rect 11655 15861 11667 15895
rect 11609 15855 11667 15861
rect 11974 15852 11980 15904
rect 12032 15892 12038 15904
rect 12621 15895 12679 15901
rect 12621 15892 12633 15895
rect 12032 15864 12633 15892
rect 12032 15852 12038 15864
rect 12621 15861 12633 15864
rect 12667 15861 12679 15895
rect 12986 15892 12992 15904
rect 12947 15864 12992 15892
rect 12621 15855 12679 15861
rect 12986 15852 12992 15864
rect 13044 15852 13050 15904
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 1578 15688 1584 15700
rect 1539 15660 1584 15688
rect 1578 15648 1584 15660
rect 1636 15648 1642 15700
rect 2317 15691 2375 15697
rect 2317 15657 2329 15691
rect 2363 15688 2375 15691
rect 2958 15688 2964 15700
rect 2363 15660 2964 15688
rect 2363 15657 2375 15660
rect 2317 15651 2375 15657
rect 2958 15648 2964 15660
rect 3016 15648 3022 15700
rect 4065 15691 4123 15697
rect 4065 15657 4077 15691
rect 4111 15688 4123 15691
rect 4430 15688 4436 15700
rect 4111 15660 4436 15688
rect 4111 15657 4123 15660
rect 4065 15651 4123 15657
rect 4430 15648 4436 15660
rect 4488 15648 4494 15700
rect 4522 15648 4528 15700
rect 4580 15688 4586 15700
rect 4580 15660 5212 15688
rect 4580 15648 4586 15660
rect 3418 15580 3424 15632
rect 3476 15620 3482 15632
rect 4893 15623 4951 15629
rect 4893 15620 4905 15623
rect 3476 15592 4905 15620
rect 3476 15580 3482 15592
rect 4893 15589 4905 15592
rect 4939 15589 4951 15623
rect 5184 15620 5212 15660
rect 5258 15648 5264 15700
rect 5316 15688 5322 15700
rect 5445 15691 5503 15697
rect 5445 15688 5457 15691
rect 5316 15660 5457 15688
rect 5316 15648 5322 15660
rect 5445 15657 5457 15660
rect 5491 15657 5503 15691
rect 5445 15651 5503 15657
rect 5537 15691 5595 15697
rect 5537 15657 5549 15691
rect 5583 15688 5595 15691
rect 6822 15688 6828 15700
rect 5583 15660 6828 15688
rect 5583 15657 5595 15660
rect 5537 15651 5595 15657
rect 6822 15648 6828 15660
rect 6880 15648 6886 15700
rect 7098 15688 7104 15700
rect 7059 15660 7104 15688
rect 7098 15648 7104 15660
rect 7156 15648 7162 15700
rect 11146 15688 11152 15700
rect 7668 15660 11152 15688
rect 6178 15620 6184 15632
rect 5184 15592 6184 15620
rect 4893 15583 4951 15589
rect 6178 15580 6184 15592
rect 6236 15580 6242 15632
rect 6362 15580 6368 15632
rect 6420 15620 6426 15632
rect 6457 15623 6515 15629
rect 6457 15620 6469 15623
rect 6420 15592 6469 15620
rect 6420 15580 6426 15592
rect 6457 15589 6469 15592
rect 6503 15589 6515 15623
rect 6457 15583 6515 15589
rect 6546 15580 6552 15632
rect 6604 15620 6610 15632
rect 7668 15620 7696 15660
rect 11146 15648 11152 15660
rect 11204 15688 11210 15700
rect 11422 15688 11428 15700
rect 11204 15660 11428 15688
rect 11204 15648 11210 15660
rect 11422 15648 11428 15660
rect 11480 15648 11486 15700
rect 11606 15688 11612 15700
rect 11567 15660 11612 15688
rect 11606 15648 11612 15660
rect 11664 15648 11670 15700
rect 11974 15688 11980 15700
rect 11935 15660 11980 15688
rect 11974 15648 11980 15660
rect 12032 15648 12038 15700
rect 12986 15648 12992 15700
rect 13044 15688 13050 15700
rect 14277 15691 14335 15697
rect 14277 15688 14289 15691
rect 13044 15660 14289 15688
rect 13044 15648 13050 15660
rect 14277 15657 14289 15660
rect 14323 15657 14335 15691
rect 14277 15651 14335 15657
rect 9214 15620 9220 15632
rect 6604 15592 7696 15620
rect 7760 15592 9220 15620
rect 6604 15580 6610 15592
rect 1397 15555 1455 15561
rect 1397 15521 1409 15555
rect 1443 15552 1455 15555
rect 1670 15552 1676 15564
rect 1443 15524 1676 15552
rect 1443 15521 1455 15524
rect 1397 15515 1455 15521
rect 1670 15512 1676 15524
rect 1728 15512 1734 15564
rect 2406 15552 2412 15564
rect 2367 15524 2412 15552
rect 2406 15512 2412 15524
rect 2464 15512 2470 15564
rect 3234 15512 3240 15564
rect 3292 15552 3298 15564
rect 3329 15555 3387 15561
rect 3329 15552 3341 15555
rect 3292 15524 3341 15552
rect 3292 15512 3298 15524
rect 3329 15521 3341 15524
rect 3375 15552 3387 15555
rect 3786 15552 3792 15564
rect 3375 15524 3792 15552
rect 3375 15521 3387 15524
rect 3329 15515 3387 15521
rect 3786 15512 3792 15524
rect 3844 15512 3850 15564
rect 4433 15555 4491 15561
rect 4433 15521 4445 15555
rect 4479 15552 4491 15555
rect 4982 15552 4988 15564
rect 4479 15524 4988 15552
rect 4479 15521 4491 15524
rect 4433 15515 4491 15521
rect 4982 15512 4988 15524
rect 5040 15512 5046 15564
rect 7760 15561 7788 15592
rect 9214 15580 9220 15592
rect 9272 15580 9278 15632
rect 9306 15580 9312 15632
rect 9364 15620 9370 15632
rect 9922 15623 9980 15629
rect 9922 15620 9934 15623
rect 9364 15592 9934 15620
rect 9364 15580 9370 15592
rect 9922 15589 9934 15592
rect 9968 15589 9980 15623
rect 9922 15583 9980 15589
rect 10226 15580 10232 15632
rect 10284 15620 10290 15632
rect 11698 15620 11704 15632
rect 10284 15592 11704 15620
rect 10284 15580 10290 15592
rect 11698 15580 11704 15592
rect 11756 15580 11762 15632
rect 12069 15623 12127 15629
rect 12069 15589 12081 15623
rect 12115 15620 12127 15623
rect 13998 15620 14004 15632
rect 12115 15592 14004 15620
rect 12115 15589 12127 15592
rect 12069 15583 12127 15589
rect 13998 15580 14004 15592
rect 14056 15580 14062 15632
rect 7745 15555 7803 15561
rect 7745 15521 7757 15555
rect 7791 15521 7803 15555
rect 7745 15515 7803 15521
rect 8018 15512 8024 15564
rect 8076 15552 8082 15564
rect 8185 15555 8243 15561
rect 8185 15552 8197 15555
rect 8076 15524 8197 15552
rect 8076 15512 8082 15524
rect 8185 15521 8197 15524
rect 8231 15552 8243 15555
rect 9677 15555 9735 15561
rect 8231 15524 8975 15552
rect 8231 15521 8243 15524
rect 8185 15515 8243 15521
rect 2590 15484 2596 15496
rect 2551 15456 2596 15484
rect 2590 15444 2596 15456
rect 2648 15444 2654 15496
rect 3421 15487 3479 15493
rect 3421 15453 3433 15487
rect 3467 15484 3479 15487
rect 3510 15484 3516 15496
rect 3467 15456 3516 15484
rect 3467 15453 3479 15456
rect 3421 15447 3479 15453
rect 3510 15444 3516 15456
rect 3568 15444 3574 15496
rect 3605 15487 3663 15493
rect 3605 15453 3617 15487
rect 3651 15484 3663 15487
rect 3970 15484 3976 15496
rect 3651 15456 3976 15484
rect 3651 15453 3663 15456
rect 3605 15447 3663 15453
rect 3970 15444 3976 15456
rect 4028 15444 4034 15496
rect 4706 15484 4712 15496
rect 4619 15456 4712 15484
rect 4706 15444 4712 15456
rect 4764 15484 4770 15496
rect 5721 15487 5779 15493
rect 4764 15456 5672 15484
rect 4764 15444 4770 15456
rect 1949 15419 2007 15425
rect 1949 15385 1961 15419
rect 1995 15416 2007 15419
rect 4893 15419 4951 15425
rect 1995 15388 4568 15416
rect 1995 15385 2007 15388
rect 1949 15379 2007 15385
rect 2961 15351 3019 15357
rect 2961 15317 2973 15351
rect 3007 15348 3019 15351
rect 3694 15348 3700 15360
rect 3007 15320 3700 15348
rect 3007 15317 3019 15320
rect 2961 15311 3019 15317
rect 3694 15308 3700 15320
rect 3752 15308 3758 15360
rect 4540 15348 4568 15388
rect 4893 15385 4905 15419
rect 4939 15416 4951 15419
rect 5077 15419 5135 15425
rect 5077 15416 5089 15419
rect 4939 15388 5089 15416
rect 4939 15385 4951 15388
rect 4893 15379 4951 15385
rect 5077 15385 5089 15388
rect 5123 15385 5135 15419
rect 5644 15416 5672 15456
rect 5721 15453 5733 15487
rect 5767 15484 5779 15487
rect 5994 15484 6000 15496
rect 5767 15456 6000 15484
rect 5767 15453 5779 15456
rect 5721 15447 5779 15453
rect 5994 15444 6000 15456
rect 6052 15444 6058 15496
rect 6733 15487 6791 15493
rect 6733 15453 6745 15487
rect 6779 15484 6791 15487
rect 7374 15484 7380 15496
rect 6779 15456 7380 15484
rect 6779 15453 6791 15456
rect 6733 15447 6791 15453
rect 6748 15416 6776 15447
rect 7374 15444 7380 15456
rect 7432 15444 7438 15496
rect 7929 15487 7987 15493
rect 7929 15453 7941 15487
rect 7975 15453 7987 15487
rect 7929 15447 7987 15453
rect 5644 15388 6776 15416
rect 5077 15379 5135 15385
rect 5718 15348 5724 15360
rect 4540 15320 5724 15348
rect 5718 15308 5724 15320
rect 5776 15308 5782 15360
rect 5810 15308 5816 15360
rect 5868 15348 5874 15360
rect 6089 15351 6147 15357
rect 6089 15348 6101 15351
rect 5868 15320 6101 15348
rect 5868 15308 5874 15320
rect 6089 15317 6101 15320
rect 6135 15317 6147 15351
rect 6089 15311 6147 15317
rect 6546 15308 6552 15360
rect 6604 15348 6610 15360
rect 6730 15348 6736 15360
rect 6604 15320 6736 15348
rect 6604 15308 6610 15320
rect 6730 15308 6736 15320
rect 6788 15348 6794 15360
rect 7561 15351 7619 15357
rect 7561 15348 7573 15351
rect 6788 15320 7573 15348
rect 6788 15308 6794 15320
rect 7561 15317 7573 15320
rect 7607 15317 7619 15351
rect 7944 15348 7972 15447
rect 8662 15348 8668 15360
rect 7944 15320 8668 15348
rect 7561 15311 7619 15317
rect 8662 15308 8668 15320
rect 8720 15308 8726 15360
rect 8947 15348 8975 15524
rect 9677 15521 9689 15555
rect 9723 15552 9735 15555
rect 10318 15552 10324 15564
rect 9723 15524 10324 15552
rect 9723 15521 9735 15524
rect 9677 15515 9735 15521
rect 10318 15512 10324 15524
rect 10376 15512 10382 15564
rect 12526 15512 12532 15564
rect 12584 15552 12590 15564
rect 12621 15555 12679 15561
rect 12621 15552 12633 15555
rect 12584 15524 12633 15552
rect 12584 15512 12590 15524
rect 12621 15521 12633 15524
rect 12667 15521 12679 15555
rect 12621 15515 12679 15521
rect 12888 15555 12946 15561
rect 12888 15521 12900 15555
rect 12934 15552 12946 15555
rect 14182 15552 14188 15564
rect 12934 15524 14188 15552
rect 12934 15521 12946 15524
rect 12888 15515 12946 15521
rect 14182 15512 14188 15524
rect 14240 15512 14246 15564
rect 12250 15484 12256 15496
rect 12211 15456 12256 15484
rect 12250 15444 12256 15456
rect 12308 15444 12314 15496
rect 9306 15416 9312 15428
rect 9267 15388 9312 15416
rect 9306 15376 9312 15388
rect 9364 15376 9370 15428
rect 13630 15376 13636 15428
rect 13688 15416 13694 15428
rect 14001 15419 14059 15425
rect 14001 15416 14013 15419
rect 13688 15388 14013 15416
rect 13688 15376 13694 15388
rect 14001 15385 14013 15388
rect 14047 15385 14059 15419
rect 14001 15379 14059 15385
rect 10870 15348 10876 15360
rect 8947 15320 10876 15348
rect 10870 15308 10876 15320
rect 10928 15308 10934 15360
rect 10962 15308 10968 15360
rect 11020 15348 11026 15360
rect 11057 15351 11115 15357
rect 11057 15348 11069 15351
rect 11020 15320 11069 15348
rect 11020 15308 11026 15320
rect 11057 15317 11069 15320
rect 11103 15317 11115 15351
rect 11057 15311 11115 15317
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 3418 15144 3424 15156
rect 3379 15116 3424 15144
rect 3418 15104 3424 15116
rect 3476 15104 3482 15156
rect 5721 15147 5779 15153
rect 5721 15113 5733 15147
rect 5767 15144 5779 15147
rect 8754 15144 8760 15156
rect 5767 15116 8760 15144
rect 5767 15113 5779 15116
rect 5721 15107 5779 15113
rect 8754 15104 8760 15116
rect 8812 15104 8818 15156
rect 13722 15144 13728 15156
rect 8956 15116 13728 15144
rect 1504 15048 2728 15076
rect 1504 14949 1532 15048
rect 1670 15008 1676 15020
rect 1631 14980 1676 15008
rect 1670 14968 1676 14980
rect 1728 14968 1734 15020
rect 1499 14943 1557 14949
rect 1499 14909 1511 14943
rect 1545 14909 1557 14943
rect 1499 14903 1557 14909
rect 1762 14832 1768 14884
rect 1820 14872 1826 14884
rect 2593 14875 2651 14881
rect 2593 14872 2605 14875
rect 1820 14844 2605 14872
rect 1820 14832 1826 14844
rect 2593 14841 2605 14844
rect 2639 14841 2651 14875
rect 2700 14872 2728 15048
rect 8018 15036 8024 15088
rect 8076 15076 8082 15088
rect 8205 15079 8263 15085
rect 8205 15076 8217 15079
rect 8076 15048 8217 15076
rect 8076 15036 8082 15048
rect 8205 15045 8217 15048
rect 8251 15045 8263 15079
rect 8205 15039 8263 15045
rect 2869 15011 2927 15017
rect 2869 14977 2881 15011
rect 2915 15008 2927 15011
rect 3510 15008 3516 15020
rect 2915 14980 3516 15008
rect 2915 14977 2927 14980
rect 2869 14971 2927 14977
rect 3510 14968 3516 14980
rect 3568 14968 3574 15020
rect 4982 14968 4988 15020
rect 5040 15008 5046 15020
rect 8956 15017 8984 15116
rect 13722 15104 13728 15116
rect 13780 15104 13786 15156
rect 13998 15144 14004 15156
rect 13959 15116 14004 15144
rect 13998 15104 14004 15116
rect 14056 15104 14062 15156
rect 14182 15104 14188 15156
rect 14240 15144 14246 15156
rect 15010 15144 15016 15156
rect 14240 15116 14596 15144
rect 14971 15116 15016 15144
rect 14240 15104 14246 15116
rect 9048 15048 9260 15076
rect 9048 15017 9076 15048
rect 6181 15011 6239 15017
rect 6181 15008 6193 15011
rect 5040 14980 6193 15008
rect 5040 14968 5046 14980
rect 6181 14977 6193 14980
rect 6227 14977 6239 15011
rect 6181 14971 6239 14977
rect 6365 15011 6423 15017
rect 6365 14977 6377 15011
rect 6411 15008 6423 15011
rect 8941 15011 8999 15017
rect 6411 14980 6960 15008
rect 6411 14977 6423 14980
rect 6365 14971 6423 14977
rect 3234 14940 3240 14952
rect 3195 14912 3240 14940
rect 3234 14900 3240 14912
rect 3292 14900 3298 14952
rect 3694 14900 3700 14952
rect 3752 14940 3758 14952
rect 3878 14940 3884 14952
rect 3752 14912 3884 14940
rect 3752 14900 3758 14912
rect 3878 14900 3884 14912
rect 3936 14940 3942 14952
rect 3973 14943 4031 14949
rect 3973 14940 3985 14943
rect 3936 14912 3985 14940
rect 3936 14900 3942 14912
rect 3973 14909 3985 14912
rect 4019 14909 4031 14943
rect 3973 14903 4031 14909
rect 4240 14943 4298 14949
rect 4240 14909 4252 14943
rect 4286 14940 4298 14943
rect 4706 14940 4712 14952
rect 4286 14912 4712 14940
rect 4286 14909 4298 14912
rect 4240 14903 4298 14909
rect 4706 14900 4712 14912
rect 4764 14900 4770 14952
rect 5902 14900 5908 14952
rect 5960 14940 5966 14952
rect 6825 14943 6883 14949
rect 6825 14940 6837 14943
rect 5960 14912 6837 14940
rect 5960 14900 5966 14912
rect 6825 14909 6837 14912
rect 6871 14909 6883 14943
rect 6932 14940 6960 14980
rect 8941 14977 8953 15011
rect 8987 14977 8999 15011
rect 8941 14971 8999 14977
rect 9033 15011 9091 15017
rect 9033 14977 9045 15011
rect 9079 14977 9091 15011
rect 9232 15008 9260 15048
rect 9306 15036 9312 15088
rect 9364 15076 9370 15088
rect 10226 15076 10232 15088
rect 9364 15048 10232 15076
rect 9364 15036 9370 15048
rect 10226 15036 10232 15048
rect 10284 15036 10290 15088
rect 11606 15036 11612 15088
rect 11664 15076 11670 15088
rect 12805 15079 12863 15085
rect 11664 15048 12756 15076
rect 11664 15036 11670 15048
rect 9401 15011 9459 15017
rect 9401 15008 9413 15011
rect 9232 14980 9413 15008
rect 9033 14971 9091 14977
rect 9401 14977 9413 14980
rect 9447 14977 9459 15011
rect 9401 14971 9459 14977
rect 9490 14968 9496 15020
rect 9548 15008 9554 15020
rect 10318 15008 10324 15020
rect 9548 14980 9593 15008
rect 10279 14980 10324 15008
rect 9548 14968 9554 14980
rect 10318 14968 10324 14980
rect 10376 14968 10382 15020
rect 12434 15008 12440 15020
rect 12395 14980 12440 15008
rect 12434 14968 12440 14980
rect 12492 14968 12498 15020
rect 12728 15008 12756 15048
rect 12805 15045 12817 15079
rect 12851 15076 12863 15079
rect 12851 15048 14504 15076
rect 12851 15045 12863 15048
rect 12805 15039 12863 15045
rect 13449 15011 13507 15017
rect 12728 14980 13400 15008
rect 6932 14912 7236 14940
rect 6825 14903 6883 14909
rect 7208 14884 7236 14912
rect 9582 14900 9588 14952
rect 9640 14940 9646 14952
rect 10229 14943 10287 14949
rect 10229 14940 10241 14943
rect 9640 14912 10241 14940
rect 9640 14900 9646 14912
rect 10229 14909 10241 14912
rect 10275 14909 10287 14943
rect 10229 14903 10287 14909
rect 10588 14943 10646 14949
rect 10588 14909 10600 14943
rect 10634 14940 10646 14943
rect 10962 14940 10968 14952
rect 10634 14912 10968 14940
rect 10634 14909 10646 14912
rect 10588 14903 10646 14909
rect 10962 14900 10968 14912
rect 11020 14900 11026 14952
rect 11054 14900 11060 14952
rect 11112 14940 11118 14952
rect 12158 14940 12164 14952
rect 11112 14912 12164 14940
rect 11112 14900 11118 14912
rect 12158 14900 12164 14912
rect 12216 14900 12222 14952
rect 5442 14872 5448 14884
rect 2700 14844 5448 14872
rect 2593 14835 2651 14841
rect 5442 14832 5448 14844
rect 5500 14832 5506 14884
rect 6089 14875 6147 14881
rect 6089 14841 6101 14875
rect 6135 14872 6147 14875
rect 6362 14872 6368 14884
rect 6135 14844 6368 14872
rect 6135 14841 6147 14844
rect 6089 14835 6147 14841
rect 6362 14832 6368 14844
rect 6420 14832 6426 14884
rect 7098 14881 7104 14884
rect 7092 14872 7104 14881
rect 7059 14844 7104 14872
rect 7092 14835 7104 14844
rect 7098 14832 7104 14835
rect 7156 14832 7162 14884
rect 7190 14832 7196 14884
rect 7248 14832 7254 14884
rect 7374 14832 7380 14884
rect 7432 14872 7438 14884
rect 12710 14872 12716 14884
rect 7432 14844 9076 14872
rect 7432 14832 7438 14844
rect 2222 14804 2228 14816
rect 2183 14776 2228 14804
rect 2222 14764 2228 14776
rect 2280 14764 2286 14816
rect 2682 14804 2688 14816
rect 2643 14776 2688 14804
rect 2682 14764 2688 14776
rect 2740 14764 2746 14816
rect 3050 14764 3056 14816
rect 3108 14804 3114 14816
rect 3326 14804 3332 14816
rect 3108 14776 3332 14804
rect 3108 14764 3114 14776
rect 3326 14764 3332 14776
rect 3384 14764 3390 14816
rect 5350 14804 5356 14816
rect 5311 14776 5356 14804
rect 5350 14764 5356 14776
rect 5408 14764 5414 14816
rect 8478 14804 8484 14816
rect 8439 14776 8484 14804
rect 8478 14764 8484 14776
rect 8536 14764 8542 14816
rect 8849 14807 8907 14813
rect 8849 14773 8861 14807
rect 8895 14804 8907 14807
rect 8938 14804 8944 14816
rect 8895 14776 8944 14804
rect 8895 14773 8907 14776
rect 8849 14767 8907 14773
rect 8938 14764 8944 14776
rect 8996 14764 9002 14816
rect 9048 14804 9076 14844
rect 9968 14844 12716 14872
rect 9401 14807 9459 14813
rect 9401 14804 9413 14807
rect 9048 14776 9413 14804
rect 9401 14773 9413 14776
rect 9447 14804 9459 14807
rect 9968 14804 9996 14844
rect 12710 14832 12716 14844
rect 12768 14832 12774 14884
rect 13265 14875 13323 14881
rect 13265 14872 13277 14875
rect 12820 14844 13277 14872
rect 9447 14776 9996 14804
rect 10045 14807 10103 14813
rect 9447 14773 9459 14776
rect 9401 14767 9459 14773
rect 10045 14773 10057 14807
rect 10091 14804 10103 14807
rect 11054 14804 11060 14816
rect 10091 14776 11060 14804
rect 10091 14773 10103 14776
rect 10045 14767 10103 14773
rect 11054 14764 11060 14776
rect 11112 14764 11118 14816
rect 11422 14764 11428 14816
rect 11480 14804 11486 14816
rect 11701 14807 11759 14813
rect 11701 14804 11713 14807
rect 11480 14776 11713 14804
rect 11480 14764 11486 14776
rect 11701 14773 11713 14776
rect 11747 14773 11759 14807
rect 11701 14767 11759 14773
rect 11882 14764 11888 14816
rect 11940 14804 11946 14816
rect 12820 14804 12848 14844
rect 13265 14841 13277 14844
rect 13311 14841 13323 14875
rect 13372 14872 13400 14980
rect 13449 14977 13461 15011
rect 13495 15008 13507 15011
rect 13814 15008 13820 15020
rect 13495 14980 13820 15008
rect 13495 14977 13507 14980
rect 13449 14971 13507 14977
rect 13814 14968 13820 14980
rect 13872 14968 13878 15020
rect 14476 15017 14504 15048
rect 14568 15017 14596 15116
rect 15010 15104 15016 15116
rect 15068 15104 15074 15156
rect 14461 15011 14519 15017
rect 14461 14977 14473 15011
rect 14507 14977 14519 15011
rect 14461 14971 14519 14977
rect 14553 15011 14611 15017
rect 14553 14977 14565 15011
rect 14599 14977 14611 15011
rect 14553 14971 14611 14977
rect 15657 15011 15715 15017
rect 15657 14977 15669 15011
rect 15703 15008 15715 15011
rect 15838 15008 15844 15020
rect 15703 14980 15844 15008
rect 15703 14977 15715 14980
rect 15657 14971 15715 14977
rect 15838 14968 15844 14980
rect 15896 14968 15902 15020
rect 13909 14943 13967 14949
rect 13909 14909 13921 14943
rect 13955 14940 13967 14943
rect 14366 14940 14372 14952
rect 13955 14912 14372 14940
rect 13955 14909 13967 14912
rect 13909 14903 13967 14909
rect 14366 14900 14372 14912
rect 14424 14900 14430 14952
rect 15473 14943 15531 14949
rect 15473 14940 15485 14943
rect 14476 14912 15485 14940
rect 14476 14872 14504 14912
rect 15473 14909 15485 14912
rect 15519 14909 15531 14943
rect 15473 14903 15531 14909
rect 18598 14872 18604 14884
rect 13372 14844 14504 14872
rect 14752 14844 18604 14872
rect 13265 14835 13323 14841
rect 11940 14776 12848 14804
rect 11940 14764 11946 14776
rect 12986 14764 12992 14816
rect 13044 14804 13050 14816
rect 13173 14807 13231 14813
rect 13173 14804 13185 14807
rect 13044 14776 13185 14804
rect 13044 14764 13050 14776
rect 13173 14773 13185 14776
rect 13219 14804 13231 14807
rect 14752 14804 14780 14844
rect 18598 14832 18604 14844
rect 18656 14832 18662 14884
rect 15378 14804 15384 14816
rect 13219 14776 14780 14804
rect 15339 14776 15384 14804
rect 13219 14773 13231 14776
rect 13173 14767 13231 14773
rect 15378 14764 15384 14776
rect 15436 14764 15442 14816
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 1670 14600 1676 14612
rect 1631 14572 1676 14600
rect 1670 14560 1676 14572
rect 1728 14560 1734 14612
rect 2222 14560 2228 14612
rect 2280 14600 2286 14612
rect 5258 14600 5264 14612
rect 2280 14572 5264 14600
rect 2280 14560 2286 14572
rect 5258 14560 5264 14572
rect 5316 14560 5322 14612
rect 7469 14603 7527 14609
rect 7469 14569 7481 14603
rect 7515 14600 7527 14603
rect 8665 14603 8723 14609
rect 8665 14600 8677 14603
rect 7515 14572 8677 14600
rect 7515 14569 7527 14572
rect 7469 14563 7527 14569
rect 8665 14569 8677 14572
rect 8711 14569 8723 14603
rect 8665 14563 8723 14569
rect 9214 14560 9220 14612
rect 9272 14600 9278 14612
rect 9309 14603 9367 14609
rect 9309 14600 9321 14603
rect 9272 14572 9321 14600
rect 9272 14560 9278 14572
rect 9309 14569 9321 14572
rect 9355 14600 9367 14603
rect 9490 14600 9496 14612
rect 9355 14572 9496 14600
rect 9355 14569 9367 14572
rect 9309 14563 9367 14569
rect 9490 14560 9496 14572
rect 9548 14560 9554 14612
rect 9677 14603 9735 14609
rect 9677 14569 9689 14603
rect 9723 14600 9735 14603
rect 13998 14600 14004 14612
rect 9723 14572 14004 14600
rect 9723 14569 9735 14572
rect 9677 14563 9735 14569
rect 13998 14560 14004 14572
rect 14056 14560 14062 14612
rect 14182 14600 14188 14612
rect 14143 14572 14188 14600
rect 14182 14560 14188 14572
rect 14240 14560 14246 14612
rect 15289 14603 15347 14609
rect 15289 14569 15301 14603
rect 15335 14569 15347 14603
rect 15289 14563 15347 14569
rect 2056 14504 2452 14532
rect 1486 14464 1492 14476
rect 1447 14436 1492 14464
rect 1486 14424 1492 14436
rect 1544 14424 1550 14476
rect 2056 14473 2084 14504
rect 2041 14467 2099 14473
rect 2041 14433 2053 14467
rect 2087 14433 2099 14467
rect 2041 14427 2099 14433
rect 2130 14424 2136 14476
rect 2188 14464 2194 14476
rect 2314 14473 2320 14476
rect 2297 14467 2320 14473
rect 2297 14464 2309 14467
rect 2188 14436 2309 14464
rect 2188 14424 2194 14436
rect 2297 14433 2309 14436
rect 2297 14427 2320 14433
rect 2314 14424 2320 14427
rect 2372 14424 2378 14476
rect 2424 14464 2452 14504
rect 2590 14492 2596 14544
rect 2648 14532 2654 14544
rect 5350 14532 5356 14544
rect 2648 14504 5356 14532
rect 2648 14492 2654 14504
rect 2774 14464 2780 14476
rect 2424 14436 2780 14464
rect 2774 14424 2780 14436
rect 2832 14424 2838 14476
rect 4908 14396 4936 14504
rect 5350 14492 5356 14504
rect 5408 14492 5414 14544
rect 5537 14535 5595 14541
rect 5537 14501 5549 14535
rect 5583 14532 5595 14535
rect 8478 14532 8484 14544
rect 5583 14504 8484 14532
rect 5583 14501 5595 14504
rect 5537 14495 5595 14501
rect 8478 14492 8484 14504
rect 8536 14492 8542 14544
rect 8754 14492 8760 14544
rect 8812 14532 8818 14544
rect 10045 14535 10103 14541
rect 8812 14504 9628 14532
rect 8812 14492 8818 14504
rect 4985 14467 5043 14473
rect 4985 14433 4997 14467
rect 5031 14464 5043 14467
rect 5445 14467 5503 14473
rect 5445 14464 5457 14467
rect 5031 14436 5457 14464
rect 5031 14433 5043 14436
rect 4985 14427 5043 14433
rect 5445 14433 5457 14436
rect 5491 14464 5503 14467
rect 5810 14464 5816 14476
rect 5491 14436 5816 14464
rect 5491 14433 5503 14436
rect 5445 14427 5503 14433
rect 5810 14424 5816 14436
rect 5868 14424 5874 14476
rect 6089 14467 6147 14473
rect 6089 14433 6101 14467
rect 6135 14464 6147 14467
rect 6546 14464 6552 14476
rect 6135 14436 6552 14464
rect 6135 14433 6147 14436
rect 6089 14427 6147 14433
rect 6546 14424 6552 14436
rect 6604 14424 6610 14476
rect 6730 14464 6736 14476
rect 6691 14436 6736 14464
rect 6730 14424 6736 14436
rect 6788 14424 6794 14476
rect 7834 14464 7840 14476
rect 7795 14436 7840 14464
rect 7834 14424 7840 14436
rect 7892 14424 7898 14476
rect 8036 14436 8892 14464
rect 5629 14399 5687 14405
rect 5629 14396 5641 14399
rect 4908 14368 5641 14396
rect 5629 14365 5641 14368
rect 5675 14365 5687 14399
rect 5629 14359 5687 14365
rect 5718 14356 5724 14408
rect 5776 14396 5782 14408
rect 6825 14399 6883 14405
rect 6825 14396 6837 14399
rect 5776 14368 6837 14396
rect 5776 14356 5782 14368
rect 6825 14365 6837 14368
rect 6871 14365 6883 14399
rect 6825 14359 6883 14365
rect 7009 14399 7067 14405
rect 7009 14365 7021 14399
rect 7055 14365 7067 14399
rect 7009 14359 7067 14365
rect 3786 14288 3792 14340
rect 3844 14328 3850 14340
rect 7024 14328 7052 14359
rect 7466 14356 7472 14408
rect 7524 14396 7530 14408
rect 7929 14399 7987 14405
rect 7929 14396 7941 14399
rect 7524 14368 7941 14396
rect 7524 14356 7530 14368
rect 7929 14365 7941 14368
rect 7975 14365 7987 14399
rect 7929 14359 7987 14365
rect 7098 14328 7104 14340
rect 3844 14300 6960 14328
rect 7011 14300 7104 14328
rect 3844 14288 3850 14300
rect 3421 14263 3479 14269
rect 3421 14229 3433 14263
rect 3467 14260 3479 14263
rect 3510 14260 3516 14272
rect 3467 14232 3516 14260
rect 3467 14229 3479 14232
rect 3421 14223 3479 14229
rect 3510 14220 3516 14232
rect 3568 14220 3574 14272
rect 5074 14260 5080 14272
rect 5035 14232 5080 14260
rect 5074 14220 5080 14232
rect 5132 14220 5138 14272
rect 5902 14260 5908 14272
rect 5863 14232 5908 14260
rect 5902 14220 5908 14232
rect 5960 14220 5966 14272
rect 6362 14260 6368 14272
rect 6323 14232 6368 14260
rect 6362 14220 6368 14232
rect 6420 14220 6426 14272
rect 6932 14260 6960 14300
rect 7098 14288 7104 14300
rect 7156 14328 7162 14340
rect 8036 14328 8064 14436
rect 8113 14399 8171 14405
rect 8113 14365 8125 14399
rect 8159 14396 8171 14399
rect 8202 14396 8208 14408
rect 8159 14368 8208 14396
rect 8159 14365 8171 14368
rect 8113 14359 8171 14365
rect 8202 14356 8208 14368
rect 8260 14356 8266 14408
rect 8754 14396 8760 14408
rect 8715 14368 8760 14396
rect 8754 14356 8760 14368
rect 8812 14356 8818 14408
rect 8864 14405 8892 14436
rect 9398 14424 9404 14476
rect 9456 14464 9462 14476
rect 9493 14467 9551 14473
rect 9493 14464 9505 14467
rect 9456 14436 9505 14464
rect 9456 14424 9462 14436
rect 9493 14433 9505 14436
rect 9539 14433 9551 14467
rect 9600 14464 9628 14504
rect 10045 14501 10057 14535
rect 10091 14532 10103 14535
rect 10091 14504 11560 14532
rect 10091 14501 10103 14504
rect 10045 14495 10103 14501
rect 10137 14467 10195 14473
rect 10137 14464 10149 14467
rect 9600 14436 10149 14464
rect 9493 14427 9551 14433
rect 10137 14433 10149 14436
rect 10183 14433 10195 14467
rect 10137 14427 10195 14433
rect 10410 14424 10416 14476
rect 10468 14464 10474 14476
rect 11422 14473 11428 14476
rect 11149 14467 11207 14473
rect 11149 14464 11161 14467
rect 10468 14436 11161 14464
rect 10468 14424 10474 14436
rect 11149 14433 11161 14436
rect 11195 14433 11207 14467
rect 11416 14464 11428 14473
rect 11383 14436 11428 14464
rect 11149 14427 11207 14433
rect 11416 14427 11428 14436
rect 11422 14424 11428 14427
rect 11480 14424 11486 14476
rect 11532 14464 11560 14504
rect 11882 14492 11888 14544
rect 11940 14532 11946 14544
rect 15304 14532 15332 14563
rect 15470 14560 15476 14612
rect 15528 14600 15534 14612
rect 15654 14600 15660 14612
rect 15528 14572 15660 14600
rect 15528 14560 15534 14572
rect 15654 14560 15660 14572
rect 15712 14560 15718 14612
rect 15749 14603 15807 14609
rect 15749 14569 15761 14603
rect 15795 14600 15807 14603
rect 19518 14600 19524 14612
rect 15795 14572 19524 14600
rect 15795 14569 15807 14572
rect 15749 14563 15807 14569
rect 11940 14504 15332 14532
rect 11940 14492 11946 14504
rect 12894 14464 12900 14476
rect 11532 14436 12900 14464
rect 12894 14424 12900 14436
rect 12952 14424 12958 14476
rect 13072 14467 13130 14473
rect 13072 14433 13084 14467
rect 13118 14464 13130 14467
rect 13814 14464 13820 14476
rect 13118 14436 13820 14464
rect 13118 14433 13130 14436
rect 13072 14427 13130 14433
rect 13814 14424 13820 14436
rect 13872 14424 13878 14476
rect 15764 14464 15792 14563
rect 19518 14560 19524 14572
rect 19576 14560 19582 14612
rect 13924 14436 15792 14464
rect 8849 14399 8907 14405
rect 8849 14365 8861 14399
rect 8895 14365 8907 14399
rect 8849 14359 8907 14365
rect 9674 14356 9680 14408
rect 9732 14356 9738 14408
rect 10321 14399 10379 14405
rect 10321 14365 10333 14399
rect 10367 14396 10379 14399
rect 10502 14396 10508 14408
rect 10367 14368 10508 14396
rect 10367 14365 10379 14368
rect 10321 14359 10379 14365
rect 10502 14356 10508 14368
rect 10560 14356 10566 14408
rect 10686 14396 10692 14408
rect 10647 14368 10692 14396
rect 10686 14356 10692 14368
rect 10744 14356 10750 14408
rect 12250 14356 12256 14408
rect 12308 14396 12314 14408
rect 12805 14399 12863 14405
rect 12805 14396 12817 14399
rect 12308 14368 12817 14396
rect 12308 14356 12314 14368
rect 12805 14365 12817 14368
rect 12851 14365 12863 14399
rect 12805 14359 12863 14365
rect 7156 14300 8064 14328
rect 8297 14331 8355 14337
rect 7156 14288 7162 14300
rect 8297 14297 8309 14331
rect 8343 14328 8355 14331
rect 9692 14328 9720 14356
rect 8343 14300 9720 14328
rect 8343 14297 8355 14300
rect 8297 14291 8355 14297
rect 7006 14260 7012 14272
rect 6932 14232 7012 14260
rect 7006 14220 7012 14232
rect 7064 14220 7070 14272
rect 7834 14220 7840 14272
rect 7892 14260 7898 14272
rect 9306 14260 9312 14272
rect 7892 14232 9312 14260
rect 7892 14220 7898 14232
rect 9306 14220 9312 14232
rect 9364 14220 9370 14272
rect 9490 14220 9496 14272
rect 9548 14260 9554 14272
rect 12342 14260 12348 14272
rect 9548 14232 12348 14260
rect 9548 14220 9554 14232
rect 12342 14220 12348 14232
rect 12400 14220 12406 14272
rect 12526 14260 12532 14272
rect 12487 14232 12532 14260
rect 12526 14220 12532 14232
rect 12584 14220 12590 14272
rect 13722 14220 13728 14272
rect 13780 14260 13786 14272
rect 13924 14260 13952 14436
rect 15838 14396 15844 14408
rect 15799 14368 15844 14396
rect 15838 14356 15844 14368
rect 15896 14356 15902 14408
rect 13780 14232 13952 14260
rect 13780 14220 13786 14232
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 1489 14059 1547 14065
rect 1489 14025 1501 14059
rect 1535 14056 1547 14059
rect 1762 14056 1768 14068
rect 1535 14028 1768 14056
rect 1535 14025 1547 14028
rect 1489 14019 1547 14025
rect 1762 14016 1768 14028
rect 1820 14016 1826 14068
rect 2774 14056 2780 14068
rect 2516 14028 2780 14056
rect 2130 13920 2136 13932
rect 2091 13892 2136 13920
rect 2130 13880 2136 13892
rect 2188 13880 2194 13932
rect 2516 13929 2544 14028
rect 2774 14016 2780 14028
rect 2832 14056 2838 14068
rect 3694 14056 3700 14068
rect 2832 14028 3700 14056
rect 2832 14016 2838 14028
rect 3694 14016 3700 14028
rect 3752 14016 3758 14068
rect 3881 14059 3939 14065
rect 3881 14025 3893 14059
rect 3927 14056 3939 14059
rect 4154 14056 4160 14068
rect 3927 14028 4160 14056
rect 3927 14025 3939 14028
rect 3881 14019 3939 14025
rect 4154 14016 4160 14028
rect 4212 14016 4218 14068
rect 4893 14059 4951 14065
rect 4893 14025 4905 14059
rect 4939 14056 4951 14059
rect 5442 14056 5448 14068
rect 4939 14028 5448 14056
rect 4939 14025 4951 14028
rect 4893 14019 4951 14025
rect 5442 14016 5448 14028
rect 5500 14016 5506 14068
rect 7561 14059 7619 14065
rect 7561 14025 7573 14059
rect 7607 14056 7619 14059
rect 8754 14056 8760 14068
rect 7607 14028 8760 14056
rect 7607 14025 7619 14028
rect 7561 14019 7619 14025
rect 8754 14016 8760 14028
rect 8812 14016 8818 14068
rect 9401 14059 9459 14065
rect 9401 14025 9413 14059
rect 9447 14056 9459 14059
rect 9490 14056 9496 14068
rect 9447 14028 9496 14056
rect 9447 14025 9459 14028
rect 9401 14019 9459 14025
rect 9490 14016 9496 14028
rect 9548 14016 9554 14068
rect 10042 14016 10048 14068
rect 10100 14056 10106 14068
rect 10229 14059 10287 14065
rect 10229 14056 10241 14059
rect 10100 14028 10241 14056
rect 10100 14016 10106 14028
rect 10229 14025 10241 14028
rect 10275 14025 10287 14059
rect 10229 14019 10287 14025
rect 11057 14059 11115 14065
rect 11057 14025 11069 14059
rect 11103 14056 11115 14059
rect 12434 14056 12440 14068
rect 11103 14028 12440 14056
rect 11103 14025 11115 14028
rect 11057 14019 11115 14025
rect 12434 14016 12440 14028
rect 12492 14016 12498 14068
rect 12710 14016 12716 14068
rect 12768 14056 12774 14068
rect 13814 14056 13820 14068
rect 12768 14028 13400 14056
rect 13775 14028 13820 14056
rect 12768 14016 12774 14028
rect 4065 13991 4123 13997
rect 4065 13957 4077 13991
rect 4111 13988 4123 13991
rect 4111 13960 5396 13988
rect 4111 13957 4123 13960
rect 4065 13951 4123 13957
rect 2501 13923 2559 13929
rect 2501 13889 2513 13923
rect 2547 13889 2559 13923
rect 2501 13883 2559 13889
rect 3510 13880 3516 13932
rect 3568 13920 3574 13932
rect 5368 13929 5396 13960
rect 5810 13948 5816 14000
rect 5868 13988 5874 14000
rect 8573 13991 8631 13997
rect 5868 13960 8248 13988
rect 5868 13948 5874 13960
rect 4617 13923 4675 13929
rect 4617 13920 4629 13923
rect 3568 13892 4629 13920
rect 3568 13880 3574 13892
rect 4617 13889 4629 13892
rect 4663 13889 4675 13923
rect 4617 13883 4675 13889
rect 5353 13923 5411 13929
rect 5353 13889 5365 13923
rect 5399 13889 5411 13923
rect 5353 13883 5411 13889
rect 5442 13880 5448 13932
rect 5500 13920 5506 13932
rect 6273 13923 6331 13929
rect 5500 13892 5545 13920
rect 5500 13880 5506 13892
rect 6273 13889 6285 13923
rect 6319 13920 6331 13923
rect 6914 13920 6920 13932
rect 6319 13892 6920 13920
rect 6319 13889 6331 13892
rect 6273 13883 6331 13889
rect 6914 13880 6920 13892
rect 6972 13920 6978 13932
rect 8110 13920 8116 13932
rect 6972 13892 8116 13920
rect 6972 13880 6978 13892
rect 8110 13880 8116 13892
rect 8168 13880 8174 13932
rect 8220 13920 8248 13960
rect 8573 13957 8585 13991
rect 8619 13988 8631 13991
rect 11882 13988 11888 14000
rect 8619 13960 10272 13988
rect 8619 13957 8631 13960
rect 8573 13951 8631 13957
rect 10244 13932 10272 13960
rect 10704 13960 11888 13988
rect 8938 13920 8944 13932
rect 8220 13892 8944 13920
rect 8938 13880 8944 13892
rect 8996 13880 9002 13932
rect 9217 13923 9275 13929
rect 9217 13889 9229 13923
rect 9263 13920 9275 13923
rect 9858 13920 9864 13932
rect 9263 13892 9864 13920
rect 9263 13889 9275 13892
rect 9217 13883 9275 13889
rect 9858 13880 9864 13892
rect 9916 13880 9922 13932
rect 9950 13880 9956 13932
rect 10008 13920 10014 13932
rect 10008 13892 10053 13920
rect 10008 13880 10014 13892
rect 10226 13880 10232 13932
rect 10284 13880 10290 13932
rect 10704 13929 10732 13960
rect 11882 13948 11888 13960
rect 11940 13948 11946 14000
rect 12250 13948 12256 14000
rect 12308 13948 12314 14000
rect 13372 13988 13400 14028
rect 13814 14016 13820 14028
rect 13872 14016 13878 14068
rect 16117 14059 16175 14065
rect 16117 14056 16129 14059
rect 13924 14028 16129 14056
rect 13924 13988 13952 14028
rect 16117 14025 16129 14028
rect 16163 14025 16175 14059
rect 16117 14019 16175 14025
rect 13372 13960 13952 13988
rect 10689 13923 10747 13929
rect 10689 13889 10701 13923
rect 10735 13889 10747 13923
rect 10870 13920 10876 13932
rect 10831 13892 10876 13920
rect 10689 13883 10747 13889
rect 10870 13880 10876 13892
rect 10928 13880 10934 13932
rect 11054 13880 11060 13932
rect 11112 13920 11118 13932
rect 11517 13923 11575 13929
rect 11517 13920 11529 13923
rect 11112 13892 11529 13920
rect 11112 13880 11118 13892
rect 11517 13889 11529 13892
rect 11563 13889 11575 13923
rect 11701 13923 11759 13929
rect 11701 13920 11713 13923
rect 11517 13883 11575 13889
rect 11624 13892 11713 13920
rect 1394 13812 1400 13864
rect 1452 13852 1458 13864
rect 1949 13855 2007 13861
rect 1949 13852 1961 13855
rect 1452 13824 1961 13852
rect 1452 13812 1458 13824
rect 1949 13821 1961 13824
rect 1995 13821 2007 13855
rect 1949 13815 2007 13821
rect 2768 13855 2826 13861
rect 2768 13821 2780 13855
rect 2814 13852 2826 13855
rect 3528 13852 3556 13880
rect 11624 13864 11652 13892
rect 11701 13889 11713 13892
rect 11747 13889 11759 13923
rect 11701 13883 11759 13889
rect 11977 13923 12035 13929
rect 11977 13889 11989 13923
rect 12023 13920 12035 13923
rect 12268 13920 12296 13948
rect 12437 13923 12495 13929
rect 12437 13920 12449 13923
rect 12023 13892 12449 13920
rect 12023 13889 12035 13892
rect 11977 13883 12035 13889
rect 12437 13889 12449 13892
rect 12483 13889 12495 13923
rect 12437 13883 12495 13889
rect 2814 13824 3556 13852
rect 2814 13821 2826 13824
rect 2768 13815 2826 13821
rect 4246 13812 4252 13864
rect 4304 13852 4310 13864
rect 4433 13855 4491 13861
rect 4304 13824 4384 13852
rect 4304 13812 4310 13824
rect 1857 13787 1915 13793
rect 1857 13753 1869 13787
rect 1903 13784 1915 13787
rect 3418 13784 3424 13796
rect 1903 13756 3424 13784
rect 1903 13753 1915 13756
rect 1857 13747 1915 13753
rect 3418 13744 3424 13756
rect 3476 13744 3482 13796
rect 4356 13784 4384 13824
rect 4433 13821 4445 13855
rect 4479 13852 4491 13855
rect 5074 13852 5080 13864
rect 4479 13824 5080 13852
rect 4479 13821 4491 13824
rect 4433 13815 4491 13821
rect 5074 13812 5080 13824
rect 5132 13812 5138 13864
rect 5258 13852 5264 13864
rect 5219 13824 5264 13852
rect 5258 13812 5264 13824
rect 5316 13812 5322 13864
rect 6178 13852 6184 13864
rect 6139 13824 6184 13852
rect 6178 13812 6184 13824
rect 6236 13812 6242 13864
rect 6362 13812 6368 13864
rect 6420 13852 6426 13864
rect 6420 13824 9904 13852
rect 6420 13812 6426 13824
rect 4525 13787 4583 13793
rect 4525 13784 4537 13787
rect 4356 13756 4537 13784
rect 4525 13753 4537 13756
rect 4571 13753 4583 13787
rect 4525 13747 4583 13753
rect 5534 13744 5540 13796
rect 5592 13784 5598 13796
rect 6825 13787 6883 13793
rect 6825 13784 6837 13787
rect 5592 13756 6837 13784
rect 5592 13744 5598 13756
rect 6825 13753 6837 13756
rect 6871 13753 6883 13787
rect 6825 13747 6883 13753
rect 7282 13744 7288 13796
rect 7340 13784 7346 13796
rect 8021 13787 8079 13793
rect 8021 13784 8033 13787
rect 7340 13756 8033 13784
rect 7340 13744 7346 13756
rect 8021 13753 8033 13756
rect 8067 13753 8079 13787
rect 8021 13747 8079 13753
rect 8202 13744 8208 13796
rect 8260 13784 8266 13796
rect 9033 13787 9091 13793
rect 9033 13784 9045 13787
rect 8260 13756 9045 13784
rect 8260 13744 8266 13756
rect 9033 13753 9045 13756
rect 9079 13753 9091 13787
rect 9033 13747 9091 13753
rect 9674 13744 9680 13796
rect 9732 13784 9738 13796
rect 9876 13793 9904 13824
rect 11146 13812 11152 13864
rect 11204 13852 11210 13864
rect 11425 13855 11483 13861
rect 11425 13852 11437 13855
rect 11204 13824 11437 13852
rect 11204 13812 11210 13824
rect 11425 13821 11437 13824
rect 11471 13821 11483 13855
rect 11425 13815 11483 13821
rect 11606 13812 11612 13864
rect 11664 13812 11670 13864
rect 12158 13812 12164 13864
rect 12216 13852 12222 13864
rect 12253 13855 12311 13861
rect 12253 13852 12265 13855
rect 12216 13824 12265 13852
rect 12216 13812 12222 13824
rect 12253 13821 12265 13824
rect 12299 13821 12311 13855
rect 12253 13815 12311 13821
rect 12342 13812 12348 13864
rect 12400 13852 12406 13864
rect 12693 13855 12751 13861
rect 12693 13852 12705 13855
rect 12400 13824 12705 13852
rect 12400 13812 12406 13824
rect 12693 13821 12705 13824
rect 12739 13821 12751 13855
rect 12693 13815 12751 13821
rect 13538 13812 13544 13864
rect 13596 13852 13602 13864
rect 14182 13852 14188 13864
rect 13596 13824 14188 13852
rect 13596 13812 13602 13824
rect 14182 13812 14188 13824
rect 14240 13812 14246 13864
rect 14737 13855 14795 13861
rect 14737 13852 14749 13855
rect 14292 13824 14749 13852
rect 9769 13787 9827 13793
rect 9769 13784 9781 13787
rect 9732 13756 9781 13784
rect 9732 13744 9738 13756
rect 9769 13753 9781 13756
rect 9815 13753 9827 13787
rect 9769 13747 9827 13753
rect 9861 13787 9919 13793
rect 9861 13753 9873 13787
rect 9907 13753 9919 13787
rect 9861 13747 9919 13753
rect 10597 13787 10655 13793
rect 10597 13753 10609 13787
rect 10643 13784 10655 13787
rect 13814 13784 13820 13796
rect 10643 13756 13820 13784
rect 10643 13753 10655 13756
rect 10597 13747 10655 13753
rect 13814 13744 13820 13756
rect 13872 13744 13878 13796
rect 3510 13676 3516 13728
rect 3568 13716 3574 13728
rect 4706 13716 4712 13728
rect 3568 13688 4712 13716
rect 3568 13676 3574 13688
rect 4706 13676 4712 13688
rect 4764 13676 4770 13728
rect 5718 13716 5724 13728
rect 5679 13688 5724 13716
rect 5718 13676 5724 13688
rect 5776 13676 5782 13728
rect 5994 13676 6000 13728
rect 6052 13716 6058 13728
rect 6089 13719 6147 13725
rect 6089 13716 6101 13719
rect 6052 13688 6101 13716
rect 6052 13676 6058 13688
rect 6089 13685 6101 13688
rect 6135 13685 6147 13719
rect 6089 13679 6147 13685
rect 7650 13676 7656 13728
rect 7708 13716 7714 13728
rect 7929 13719 7987 13725
rect 7929 13716 7941 13719
rect 7708 13688 7941 13716
rect 7708 13676 7714 13688
rect 7929 13685 7941 13688
rect 7975 13685 7987 13719
rect 7929 13679 7987 13685
rect 8754 13676 8760 13728
rect 8812 13716 8818 13728
rect 8941 13719 8999 13725
rect 8941 13716 8953 13719
rect 8812 13688 8953 13716
rect 8812 13676 8818 13688
rect 8941 13685 8953 13688
rect 8987 13685 8999 13719
rect 8941 13679 8999 13685
rect 9122 13676 9128 13728
rect 9180 13716 9186 13728
rect 11146 13716 11152 13728
rect 9180 13688 11152 13716
rect 9180 13676 9186 13688
rect 11146 13676 11152 13688
rect 11204 13676 11210 13728
rect 11698 13676 11704 13728
rect 11756 13716 11762 13728
rect 11977 13719 12035 13725
rect 11977 13716 11989 13719
rect 11756 13688 11989 13716
rect 11756 13676 11762 13688
rect 11977 13685 11989 13688
rect 12023 13716 12035 13719
rect 12069 13719 12127 13725
rect 12069 13716 12081 13719
rect 12023 13688 12081 13716
rect 12023 13685 12035 13688
rect 11977 13679 12035 13685
rect 12069 13685 12081 13688
rect 12115 13716 12127 13719
rect 14292 13716 14320 13824
rect 14737 13821 14749 13824
rect 14783 13821 14795 13855
rect 14737 13815 14795 13821
rect 15004 13855 15062 13861
rect 15004 13821 15016 13855
rect 15050 13852 15062 13855
rect 18690 13852 18696 13864
rect 15050 13824 18696 13852
rect 15050 13821 15062 13824
rect 15004 13815 15062 13821
rect 18690 13812 18696 13824
rect 18748 13812 18754 13864
rect 12115 13688 14320 13716
rect 12115 13685 12127 13688
rect 12069 13679 12127 13685
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 2133 13515 2191 13521
rect 2133 13481 2145 13515
rect 2179 13512 2191 13515
rect 2682 13512 2688 13524
rect 2179 13484 2688 13512
rect 2179 13481 2191 13484
rect 2133 13475 2191 13481
rect 2682 13472 2688 13484
rect 2740 13472 2746 13524
rect 3326 13512 3332 13524
rect 3287 13484 3332 13512
rect 3326 13472 3332 13484
rect 3384 13472 3390 13524
rect 3602 13472 3608 13524
rect 3660 13512 3666 13524
rect 6362 13512 6368 13524
rect 3660 13484 6368 13512
rect 3660 13472 3666 13484
rect 6362 13472 6368 13484
rect 6420 13472 6426 13524
rect 7098 13512 7104 13524
rect 7059 13484 7104 13512
rect 7098 13472 7104 13484
rect 7156 13472 7162 13524
rect 8754 13472 8760 13524
rect 8812 13512 8818 13524
rect 9677 13515 9735 13521
rect 8812 13484 9444 13512
rect 8812 13472 8818 13484
rect 1486 13404 1492 13456
rect 1544 13444 1550 13456
rect 1673 13447 1731 13453
rect 1673 13444 1685 13447
rect 1544 13416 1685 13444
rect 1544 13404 1550 13416
rect 1673 13413 1685 13416
rect 1719 13413 1731 13447
rect 1673 13407 1731 13413
rect 2056 13416 4108 13444
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 2056 13376 2084 13416
rect 2498 13376 2504 13388
rect 1443 13348 2084 13376
rect 2459 13348 2504 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 2498 13336 2504 13348
rect 2556 13336 2562 13388
rect 2593 13379 2651 13385
rect 2593 13345 2605 13379
rect 2639 13376 2651 13379
rect 2866 13376 2872 13388
rect 2639 13348 2872 13376
rect 2639 13345 2651 13348
rect 2593 13339 2651 13345
rect 2866 13336 2872 13348
rect 2924 13336 2930 13388
rect 3145 13379 3203 13385
rect 3145 13345 3157 13379
rect 3191 13376 3203 13379
rect 3878 13376 3884 13388
rect 3191 13348 3884 13376
rect 3191 13345 3203 13348
rect 3145 13339 3203 13345
rect 3878 13336 3884 13348
rect 3936 13336 3942 13388
rect 4080 13376 4108 13416
rect 4154 13404 4160 13456
rect 4212 13444 4218 13456
rect 4332 13447 4390 13453
rect 4332 13444 4344 13447
rect 4212 13416 4344 13444
rect 4212 13404 4218 13416
rect 4332 13413 4344 13416
rect 4378 13444 4390 13447
rect 5442 13444 5448 13456
rect 4378 13416 5448 13444
rect 4378 13413 4390 13416
rect 4332 13407 4390 13413
rect 5442 13404 5448 13416
rect 5500 13404 5506 13456
rect 5988 13447 6046 13453
rect 5988 13413 6000 13447
rect 6034 13444 6046 13447
rect 6914 13444 6920 13456
rect 6034 13416 6920 13444
rect 6034 13413 6046 13416
rect 5988 13407 6046 13413
rect 6914 13404 6920 13416
rect 6972 13404 6978 13456
rect 7116 13444 7144 13472
rect 7622 13447 7680 13453
rect 7622 13444 7634 13447
rect 7116 13416 7634 13444
rect 7622 13413 7634 13416
rect 7668 13413 7680 13447
rect 7622 13407 7680 13413
rect 8294 13404 8300 13456
rect 8352 13444 8358 13456
rect 9309 13447 9367 13453
rect 9309 13444 9321 13447
rect 8352 13416 9321 13444
rect 8352 13404 8358 13416
rect 9309 13413 9321 13416
rect 9355 13413 9367 13447
rect 9416 13444 9444 13484
rect 9677 13481 9689 13515
rect 9723 13512 9735 13515
rect 9766 13512 9772 13524
rect 9723 13484 9772 13512
rect 9723 13481 9735 13484
rect 9677 13475 9735 13481
rect 9766 13472 9772 13484
rect 9824 13472 9830 13524
rect 10045 13515 10103 13521
rect 10045 13481 10057 13515
rect 10091 13512 10103 13515
rect 10686 13512 10692 13524
rect 10091 13484 10692 13512
rect 10091 13481 10103 13484
rect 10045 13475 10103 13481
rect 10686 13472 10692 13484
rect 10744 13472 10750 13524
rect 10778 13472 10784 13524
rect 10836 13512 10842 13524
rect 11057 13515 11115 13521
rect 11057 13512 11069 13515
rect 10836 13484 11069 13512
rect 10836 13472 10842 13484
rect 11057 13481 11069 13484
rect 11103 13481 11115 13515
rect 11057 13475 11115 13481
rect 11146 13472 11152 13524
rect 11204 13512 11210 13524
rect 12069 13515 12127 13521
rect 12069 13512 12081 13515
rect 11204 13484 12081 13512
rect 11204 13472 11210 13484
rect 12069 13481 12081 13484
rect 12115 13481 12127 13515
rect 12069 13475 12127 13481
rect 12434 13472 12440 13524
rect 12492 13512 12498 13524
rect 13357 13515 13415 13521
rect 13357 13512 13369 13515
rect 12492 13484 13369 13512
rect 12492 13472 12498 13484
rect 13357 13481 13369 13484
rect 13403 13481 13415 13515
rect 13357 13475 13415 13481
rect 13814 13472 13820 13524
rect 13872 13512 13878 13524
rect 15289 13515 15347 13521
rect 15289 13512 15301 13515
rect 13872 13484 15301 13512
rect 13872 13472 13878 13484
rect 15289 13481 15301 13484
rect 15335 13481 15347 13515
rect 15289 13475 15347 13481
rect 16301 13515 16359 13521
rect 16301 13481 16313 13515
rect 16347 13481 16359 13515
rect 16301 13475 16359 13481
rect 10137 13447 10195 13453
rect 9416 13416 10088 13444
rect 9309 13407 9367 13413
rect 6546 13376 6552 13388
rect 4080 13348 6552 13376
rect 6546 13336 6552 13348
rect 6604 13336 6610 13388
rect 7006 13336 7012 13388
rect 7064 13376 7070 13388
rect 8202 13376 8208 13388
rect 7064 13348 8208 13376
rect 7064 13336 7070 13348
rect 8202 13336 8208 13348
rect 8260 13336 8266 13388
rect 9033 13379 9091 13385
rect 9033 13345 9045 13379
rect 9079 13376 9091 13379
rect 9674 13376 9680 13388
rect 9079 13348 9680 13376
rect 9079 13345 9091 13348
rect 9033 13339 9091 13345
rect 9674 13336 9680 13348
rect 9732 13336 9738 13388
rect 10060 13376 10088 13416
rect 10137 13413 10149 13447
rect 10183 13444 10195 13447
rect 16316 13444 16344 13475
rect 10183 13416 16344 13444
rect 10183 13413 10195 13416
rect 10137 13407 10195 13413
rect 10410 13376 10416 13388
rect 10060 13348 10416 13376
rect 10410 13336 10416 13348
rect 10468 13336 10474 13388
rect 10965 13379 11023 13385
rect 10965 13345 10977 13379
rect 11011 13345 11023 13379
rect 10965 13339 11023 13345
rect 2130 13268 2136 13320
rect 2188 13308 2194 13320
rect 2685 13311 2743 13317
rect 2685 13308 2697 13311
rect 2188 13280 2697 13308
rect 2188 13268 2194 13280
rect 2685 13277 2697 13280
rect 2731 13277 2743 13311
rect 2685 13271 2743 13277
rect 3694 13268 3700 13320
rect 3752 13308 3758 13320
rect 4065 13311 4123 13317
rect 4065 13308 4077 13311
rect 3752 13280 4077 13308
rect 3752 13268 3758 13280
rect 4065 13277 4077 13280
rect 4111 13277 4123 13311
rect 5718 13308 5724 13320
rect 5679 13280 5724 13308
rect 4065 13271 4123 13277
rect 5718 13268 5724 13280
rect 5776 13268 5782 13320
rect 7374 13308 7380 13320
rect 7335 13280 7380 13308
rect 7374 13268 7380 13280
rect 7432 13268 7438 13320
rect 8478 13268 8484 13320
rect 8536 13308 8542 13320
rect 9766 13308 9772 13320
rect 8536 13280 9772 13308
rect 8536 13268 8542 13280
rect 9766 13268 9772 13280
rect 9824 13268 9830 13320
rect 10321 13311 10379 13317
rect 10321 13277 10333 13311
rect 10367 13308 10379 13311
rect 10870 13308 10876 13320
rect 10367 13280 10876 13308
rect 10367 13277 10379 13280
rect 10321 13271 10379 13277
rect 10870 13268 10876 13280
rect 10928 13268 10934 13320
rect 10980 13308 11008 13339
rect 11330 13336 11336 13388
rect 11388 13376 11394 13388
rect 11977 13379 12035 13385
rect 11977 13376 11989 13379
rect 11388 13348 11989 13376
rect 11388 13336 11394 13348
rect 11977 13345 11989 13348
rect 12023 13345 12035 13379
rect 12986 13376 12992 13388
rect 11977 13339 12035 13345
rect 12452 13348 12992 13376
rect 11054 13308 11060 13320
rect 10980 13280 11060 13308
rect 11054 13268 11060 13280
rect 11112 13268 11118 13320
rect 11146 13268 11152 13320
rect 11204 13308 11210 13320
rect 12250 13308 12256 13320
rect 11204 13280 11249 13308
rect 12211 13280 12256 13308
rect 11204 13268 11210 13280
rect 12250 13268 12256 13280
rect 12308 13268 12314 13320
rect 8757 13243 8815 13249
rect 8757 13209 8769 13243
rect 8803 13240 8815 13243
rect 9950 13240 9956 13252
rect 8803 13212 9956 13240
rect 8803 13209 8815 13212
rect 8757 13203 8815 13209
rect 9950 13200 9956 13212
rect 10008 13200 10014 13252
rect 12452 13240 12480 13348
rect 12986 13336 12992 13348
rect 13044 13336 13050 13388
rect 13265 13379 13323 13385
rect 13265 13345 13277 13379
rect 13311 13376 13323 13379
rect 13722 13376 13728 13388
rect 13311 13348 13728 13376
rect 13311 13345 13323 13348
rect 13265 13339 13323 13345
rect 13722 13336 13728 13348
rect 13780 13336 13786 13388
rect 14274 13376 14280 13388
rect 14235 13348 14280 13376
rect 14274 13336 14280 13348
rect 14332 13336 14338 13388
rect 14369 13379 14427 13385
rect 14369 13345 14381 13379
rect 14415 13376 14427 13379
rect 14826 13376 14832 13388
rect 14415 13348 14832 13376
rect 14415 13345 14427 13348
rect 14369 13339 14427 13345
rect 14826 13336 14832 13348
rect 14884 13376 14890 13388
rect 15102 13376 15108 13388
rect 14884 13348 15108 13376
rect 14884 13336 14890 13348
rect 15102 13336 15108 13348
rect 15160 13336 15166 13388
rect 15286 13336 15292 13388
rect 15344 13376 15350 13388
rect 15657 13379 15715 13385
rect 15657 13376 15669 13379
rect 15344 13348 15669 13376
rect 15344 13336 15350 13348
rect 15657 13345 15669 13348
rect 15703 13345 15715 13379
rect 15657 13339 15715 13345
rect 15746 13336 15752 13388
rect 15804 13376 15810 13388
rect 16669 13379 16727 13385
rect 16669 13376 16681 13379
rect 15804 13348 15849 13376
rect 15948 13348 16681 13376
rect 15804 13336 15810 13348
rect 12526 13268 12532 13320
rect 12584 13308 12590 13320
rect 13449 13311 13507 13317
rect 13449 13308 13461 13311
rect 12584 13280 13461 13308
rect 12584 13268 12590 13280
rect 13449 13277 13461 13280
rect 13495 13308 13507 13311
rect 14461 13311 14519 13317
rect 14461 13308 14473 13311
rect 13495 13280 14473 13308
rect 13495 13277 13507 13280
rect 13449 13271 13507 13277
rect 14461 13277 14473 13280
rect 14507 13277 14519 13311
rect 14461 13271 14519 13277
rect 14642 13268 14648 13320
rect 14700 13308 14706 13320
rect 15838 13308 15844 13320
rect 14700 13280 15148 13308
rect 15799 13280 15844 13308
rect 14700 13268 14706 13280
rect 10060 13212 12480 13240
rect 12897 13243 12955 13249
rect 3418 13132 3424 13184
rect 3476 13172 3482 13184
rect 4062 13172 4068 13184
rect 3476 13144 4068 13172
rect 3476 13132 3482 13144
rect 4062 13132 4068 13144
rect 4120 13132 4126 13184
rect 5445 13175 5503 13181
rect 5445 13141 5457 13175
rect 5491 13172 5503 13175
rect 5718 13172 5724 13184
rect 5491 13144 5724 13172
rect 5491 13141 5503 13144
rect 5445 13135 5503 13141
rect 5718 13132 5724 13144
rect 5776 13132 5782 13184
rect 5902 13132 5908 13184
rect 5960 13172 5966 13184
rect 10060 13172 10088 13212
rect 12897 13209 12909 13243
rect 12943 13240 12955 13243
rect 15010 13240 15016 13252
rect 12943 13212 15016 13240
rect 12943 13209 12955 13212
rect 12897 13203 12955 13209
rect 15010 13200 15016 13212
rect 15068 13200 15074 13252
rect 15120 13240 15148 13280
rect 15838 13268 15844 13280
rect 15896 13268 15902 13320
rect 15948 13240 15976 13348
rect 16669 13345 16681 13348
rect 16715 13345 16727 13379
rect 16669 13339 16727 13345
rect 16758 13308 16764 13320
rect 16719 13280 16764 13308
rect 16758 13268 16764 13280
rect 16816 13268 16822 13320
rect 16853 13311 16911 13317
rect 16853 13277 16865 13311
rect 16899 13277 16911 13311
rect 16853 13271 16911 13277
rect 16868 13240 16896 13271
rect 15120 13212 15976 13240
rect 16776 13212 16896 13240
rect 5960 13144 10088 13172
rect 5960 13132 5966 13144
rect 10318 13132 10324 13184
rect 10376 13172 10382 13184
rect 10597 13175 10655 13181
rect 10597 13172 10609 13175
rect 10376 13144 10609 13172
rect 10376 13132 10382 13144
rect 10597 13141 10609 13144
rect 10643 13141 10655 13175
rect 10597 13135 10655 13141
rect 11609 13175 11667 13181
rect 11609 13141 11621 13175
rect 11655 13172 11667 13175
rect 13538 13172 13544 13184
rect 11655 13144 13544 13172
rect 11655 13141 11667 13144
rect 11609 13135 11667 13141
rect 13538 13132 13544 13144
rect 13596 13132 13602 13184
rect 13909 13175 13967 13181
rect 13909 13141 13921 13175
rect 13955 13172 13967 13175
rect 14918 13172 14924 13184
rect 13955 13144 14924 13172
rect 13955 13141 13967 13144
rect 13909 13135 13967 13141
rect 14918 13132 14924 13144
rect 14976 13132 14982 13184
rect 15838 13132 15844 13184
rect 15896 13172 15902 13184
rect 16776 13172 16804 13212
rect 15896 13144 16804 13172
rect 15896 13132 15902 13144
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 3142 12928 3148 12980
rect 3200 12968 3206 12980
rect 5994 12968 6000 12980
rect 3200 12940 6000 12968
rect 3200 12928 3206 12940
rect 5994 12928 6000 12940
rect 6052 12928 6058 12980
rect 6178 12928 6184 12980
rect 6236 12968 6242 12980
rect 6825 12971 6883 12977
rect 6825 12968 6837 12971
rect 6236 12940 6837 12968
rect 6236 12928 6242 12940
rect 6825 12937 6837 12940
rect 6871 12937 6883 12971
rect 6825 12931 6883 12937
rect 7282 12928 7288 12980
rect 7340 12968 7346 12980
rect 7650 12968 7656 12980
rect 7340 12940 7656 12968
rect 7340 12928 7346 12940
rect 7650 12928 7656 12940
rect 7708 12928 7714 12980
rect 9674 12968 9680 12980
rect 9635 12940 9680 12968
rect 9674 12928 9680 12940
rect 9732 12928 9738 12980
rect 10704 12940 12112 12968
rect 4154 12900 4160 12912
rect 2240 12872 4160 12900
rect 2240 12841 2268 12872
rect 4154 12860 4160 12872
rect 4212 12860 4218 12912
rect 9306 12860 9312 12912
rect 9364 12900 9370 12912
rect 9858 12900 9864 12912
rect 9364 12872 9864 12900
rect 9364 12860 9370 12872
rect 9858 12860 9864 12872
rect 9916 12860 9922 12912
rect 10597 12903 10655 12909
rect 10597 12900 10609 12903
rect 9968 12872 10609 12900
rect 2225 12835 2283 12841
rect 2225 12801 2237 12835
rect 2271 12801 2283 12835
rect 2406 12832 2412 12844
rect 2367 12804 2412 12832
rect 2225 12795 2283 12801
rect 2406 12792 2412 12804
rect 2464 12792 2470 12844
rect 3418 12832 3424 12844
rect 3379 12804 3424 12832
rect 3418 12792 3424 12804
rect 3476 12792 3482 12844
rect 3694 12792 3700 12844
rect 3752 12832 3758 12844
rect 3752 12804 3924 12832
rect 3752 12792 3758 12804
rect 3237 12767 3295 12773
rect 3237 12733 3249 12767
rect 3283 12764 3295 12767
rect 3326 12764 3332 12776
rect 3283 12736 3332 12764
rect 3283 12733 3295 12736
rect 3237 12727 3295 12733
rect 3326 12724 3332 12736
rect 3384 12764 3390 12776
rect 3510 12764 3516 12776
rect 3384 12736 3516 12764
rect 3384 12724 3390 12736
rect 3510 12724 3516 12736
rect 3568 12724 3574 12776
rect 3786 12764 3792 12776
rect 3747 12736 3792 12764
rect 3786 12724 3792 12736
rect 3844 12724 3850 12776
rect 3896 12764 3924 12804
rect 3970 12792 3976 12844
rect 4028 12832 4034 12844
rect 4028 12804 4844 12832
rect 4028 12792 4034 12804
rect 4709 12767 4767 12773
rect 4709 12764 4721 12767
rect 3896 12736 4721 12764
rect 4709 12733 4721 12736
rect 4755 12733 4767 12767
rect 4709 12727 4767 12733
rect 2958 12656 2964 12708
rect 3016 12696 3022 12708
rect 3016 12668 4016 12696
rect 3016 12656 3022 12668
rect 1578 12588 1584 12640
rect 1636 12628 1642 12640
rect 1765 12631 1823 12637
rect 1765 12628 1777 12631
rect 1636 12600 1777 12628
rect 1636 12588 1642 12600
rect 1765 12597 1777 12600
rect 1811 12597 1823 12631
rect 2130 12628 2136 12640
rect 2091 12600 2136 12628
rect 1765 12591 1823 12597
rect 2130 12588 2136 12600
rect 2188 12588 2194 12640
rect 2774 12588 2780 12640
rect 2832 12628 2838 12640
rect 3142 12628 3148 12640
rect 2832 12600 2877 12628
rect 3103 12600 3148 12628
rect 2832 12588 2838 12600
rect 3142 12588 3148 12600
rect 3200 12588 3206 12640
rect 3988 12637 4016 12668
rect 3973 12631 4031 12637
rect 3973 12597 3985 12631
rect 4019 12597 4031 12631
rect 4724 12628 4752 12727
rect 4816 12696 4844 12804
rect 5718 12792 5724 12844
rect 5776 12832 5782 12844
rect 7377 12835 7435 12841
rect 7377 12832 7389 12835
rect 5776 12804 6132 12832
rect 5776 12792 5782 12804
rect 4976 12767 5034 12773
rect 4976 12733 4988 12767
rect 5022 12764 5034 12767
rect 5736 12764 5764 12792
rect 5022 12736 5764 12764
rect 5022 12733 5034 12736
rect 4976 12727 5034 12733
rect 5810 12724 5816 12776
rect 5868 12764 5874 12776
rect 6104 12764 6132 12804
rect 6932 12804 7389 12832
rect 6932 12764 6960 12804
rect 7377 12801 7389 12804
rect 7423 12801 7435 12835
rect 7377 12795 7435 12801
rect 9030 12792 9036 12844
rect 9088 12832 9094 12844
rect 9490 12832 9496 12844
rect 9088 12804 9496 12832
rect 9088 12792 9094 12804
rect 9490 12792 9496 12804
rect 9548 12832 9554 12844
rect 9968 12832 9996 12872
rect 10597 12869 10609 12872
rect 10643 12869 10655 12903
rect 10597 12863 10655 12869
rect 9548 12804 9996 12832
rect 10321 12835 10379 12841
rect 9548 12792 9554 12804
rect 10321 12801 10333 12835
rect 10367 12832 10379 12835
rect 10704 12832 10732 12940
rect 12084 12909 12112 12940
rect 12158 12928 12164 12980
rect 12216 12968 12222 12980
rect 14274 12968 14280 12980
rect 12216 12940 14280 12968
rect 12216 12928 12222 12940
rect 14274 12928 14280 12940
rect 14332 12928 14338 12980
rect 15562 12968 15568 12980
rect 15523 12940 15568 12968
rect 15562 12928 15568 12940
rect 15620 12928 15626 12980
rect 12069 12903 12127 12909
rect 12069 12869 12081 12903
rect 12115 12900 12127 12903
rect 12342 12900 12348 12912
rect 12115 12872 12348 12900
rect 12115 12869 12127 12872
rect 12069 12863 12127 12869
rect 12342 12860 12348 12872
rect 12400 12860 12406 12912
rect 14369 12903 14427 12909
rect 14369 12869 14381 12903
rect 14415 12900 14427 12903
rect 14415 12872 16160 12900
rect 14415 12869 14427 12872
rect 14369 12863 14427 12869
rect 12434 12832 12440 12844
rect 10367 12804 10732 12832
rect 12395 12804 12440 12832
rect 10367 12801 10379 12804
rect 10321 12795 10379 12801
rect 12434 12792 12440 12804
rect 12492 12792 12498 12844
rect 15102 12832 15108 12844
rect 15063 12804 15108 12832
rect 15102 12792 15108 12804
rect 15160 12792 15166 12844
rect 16132 12841 16160 12872
rect 16117 12835 16175 12841
rect 16117 12801 16129 12835
rect 16163 12801 16175 12835
rect 16117 12795 16175 12801
rect 5868 12736 6040 12764
rect 6104 12736 6960 12764
rect 5868 12724 5874 12736
rect 5902 12696 5908 12708
rect 4816 12668 5908 12696
rect 5902 12656 5908 12668
rect 5960 12656 5966 12708
rect 6012 12696 6040 12736
rect 7006 12724 7012 12776
rect 7064 12764 7070 12776
rect 7285 12767 7343 12773
rect 7285 12764 7297 12767
rect 7064 12736 7297 12764
rect 7064 12724 7070 12736
rect 7285 12733 7297 12736
rect 7331 12733 7343 12767
rect 7285 12727 7343 12733
rect 7929 12767 7987 12773
rect 7929 12733 7941 12767
rect 7975 12733 7987 12767
rect 7929 12727 7987 12733
rect 8196 12767 8254 12773
rect 8196 12733 8208 12767
rect 8242 12764 8254 12767
rect 9950 12764 9956 12776
rect 8242 12736 9956 12764
rect 8242 12733 8254 12736
rect 8196 12727 8254 12733
rect 7374 12696 7380 12708
rect 6012 12668 7380 12696
rect 5534 12628 5540 12640
rect 4724 12600 5540 12628
rect 3973 12591 4031 12597
rect 5534 12588 5540 12600
rect 5592 12628 5598 12640
rect 6012 12628 6040 12668
rect 7374 12656 7380 12668
rect 7432 12696 7438 12708
rect 7944 12696 7972 12727
rect 9950 12724 9956 12736
rect 10008 12724 10014 12776
rect 10410 12724 10416 12776
rect 10468 12764 10474 12776
rect 10689 12767 10747 12773
rect 10689 12764 10701 12767
rect 10468 12736 10701 12764
rect 10468 12724 10474 12736
rect 10689 12733 10701 12736
rect 10735 12733 10747 12767
rect 12710 12764 12716 12776
rect 10689 12727 10747 12733
rect 10796 12736 12716 12764
rect 7432 12668 7972 12696
rect 10045 12699 10103 12705
rect 7432 12656 7438 12668
rect 10045 12665 10057 12699
rect 10091 12696 10103 12699
rect 10318 12696 10324 12708
rect 10091 12668 10324 12696
rect 10091 12665 10103 12668
rect 10045 12659 10103 12665
rect 10318 12656 10324 12668
rect 10376 12656 10382 12708
rect 10597 12699 10655 12705
rect 10597 12665 10609 12699
rect 10643 12696 10655 12699
rect 10796 12696 10824 12736
rect 12710 12724 12716 12736
rect 12768 12724 12774 12776
rect 12897 12767 12955 12773
rect 12897 12733 12909 12767
rect 12943 12733 12955 12767
rect 14642 12764 14648 12776
rect 12897 12727 12955 12733
rect 14108 12736 14648 12764
rect 10643 12668 10824 12696
rect 10956 12699 11014 12705
rect 10643 12665 10655 12668
rect 10597 12659 10655 12665
rect 10956 12665 10968 12699
rect 11002 12696 11014 12699
rect 11146 12696 11152 12708
rect 11002 12668 11152 12696
rect 11002 12665 11014 12668
rect 10956 12659 11014 12665
rect 11146 12656 11152 12668
rect 11204 12696 11210 12708
rect 11606 12696 11612 12708
rect 11204 12668 11612 12696
rect 11204 12656 11210 12668
rect 11606 12656 11612 12668
rect 11664 12656 11670 12708
rect 11698 12656 11704 12708
rect 11756 12696 11762 12708
rect 12434 12696 12440 12708
rect 11756 12668 12440 12696
rect 11756 12656 11762 12668
rect 12434 12656 12440 12668
rect 12492 12696 12498 12708
rect 12912 12696 12940 12727
rect 12492 12668 12940 12696
rect 13164 12699 13222 12705
rect 12492 12656 12498 12668
rect 13164 12665 13176 12699
rect 13210 12696 13222 12699
rect 13814 12696 13820 12708
rect 13210 12668 13820 12696
rect 13210 12665 13222 12668
rect 13164 12659 13222 12665
rect 13814 12656 13820 12668
rect 13872 12656 13878 12708
rect 5592 12600 6040 12628
rect 6089 12631 6147 12637
rect 5592 12588 5598 12600
rect 6089 12597 6101 12631
rect 6135 12628 6147 12631
rect 6178 12628 6184 12640
rect 6135 12600 6184 12628
rect 6135 12597 6147 12600
rect 6089 12591 6147 12597
rect 6178 12588 6184 12600
rect 6236 12588 6242 12640
rect 6362 12588 6368 12640
rect 6420 12628 6426 12640
rect 7193 12631 7251 12637
rect 7193 12628 7205 12631
rect 6420 12600 7205 12628
rect 6420 12588 6426 12600
rect 7193 12597 7205 12600
rect 7239 12628 7251 12631
rect 9122 12628 9128 12640
rect 7239 12600 9128 12628
rect 7239 12597 7251 12600
rect 7193 12591 7251 12597
rect 9122 12588 9128 12600
rect 9180 12588 9186 12640
rect 9309 12631 9367 12637
rect 9309 12597 9321 12631
rect 9355 12628 9367 12631
rect 9490 12628 9496 12640
rect 9355 12600 9496 12628
rect 9355 12597 9367 12600
rect 9309 12591 9367 12597
rect 9490 12588 9496 12600
rect 9548 12588 9554 12640
rect 10137 12631 10195 12637
rect 10137 12597 10149 12631
rect 10183 12628 10195 12631
rect 11882 12628 11888 12640
rect 10183 12600 11888 12628
rect 10183 12597 10195 12600
rect 10137 12591 10195 12597
rect 11882 12588 11888 12600
rect 11940 12588 11946 12640
rect 12066 12588 12072 12640
rect 12124 12628 12130 12640
rect 14108 12628 14136 12736
rect 14642 12724 14648 12736
rect 14700 12724 14706 12776
rect 14918 12764 14924 12776
rect 14879 12736 14924 12764
rect 14918 12724 14924 12736
rect 14976 12724 14982 12776
rect 15010 12724 15016 12776
rect 15068 12764 15074 12776
rect 15068 12736 15113 12764
rect 15068 12724 15074 12736
rect 16025 12699 16083 12705
rect 16025 12696 16037 12699
rect 14568 12668 16037 12696
rect 14274 12628 14280 12640
rect 12124 12600 14136 12628
rect 14187 12600 14280 12628
rect 12124 12588 12130 12600
rect 14274 12588 14280 12600
rect 14332 12628 14338 12640
rect 14568 12637 14596 12668
rect 16025 12665 16037 12668
rect 16071 12665 16083 12699
rect 16025 12659 16083 12665
rect 14369 12631 14427 12637
rect 14369 12628 14381 12631
rect 14332 12600 14381 12628
rect 14332 12588 14338 12600
rect 14369 12597 14381 12600
rect 14415 12597 14427 12631
rect 14369 12591 14427 12597
rect 14553 12631 14611 12637
rect 14553 12597 14565 12631
rect 14599 12597 14611 12631
rect 15930 12628 15936 12640
rect 15891 12600 15936 12628
rect 14553 12591 14611 12597
rect 15930 12588 15936 12600
rect 15988 12588 15994 12640
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 1765 12427 1823 12433
rect 1765 12393 1777 12427
rect 1811 12424 1823 12427
rect 2130 12424 2136 12436
rect 1811 12396 2136 12424
rect 1811 12393 1823 12396
rect 1765 12387 1823 12393
rect 2130 12384 2136 12396
rect 2188 12384 2194 12436
rect 2225 12427 2283 12433
rect 2225 12393 2237 12427
rect 2271 12424 2283 12427
rect 2777 12427 2835 12433
rect 2777 12424 2789 12427
rect 2271 12396 2789 12424
rect 2271 12393 2283 12396
rect 2225 12387 2283 12393
rect 2777 12393 2789 12396
rect 2823 12393 2835 12427
rect 2777 12387 2835 12393
rect 3050 12384 3056 12436
rect 3108 12424 3114 12436
rect 3145 12427 3203 12433
rect 3145 12424 3157 12427
rect 3108 12396 3157 12424
rect 3108 12384 3114 12396
rect 3145 12393 3157 12396
rect 3191 12393 3203 12427
rect 3145 12387 3203 12393
rect 4525 12427 4583 12433
rect 4525 12393 4537 12427
rect 4571 12424 4583 12427
rect 4798 12424 4804 12436
rect 4571 12396 4804 12424
rect 4571 12393 4583 12396
rect 4525 12387 4583 12393
rect 4798 12384 4804 12396
rect 4856 12384 4862 12436
rect 9677 12427 9735 12433
rect 9677 12393 9689 12427
rect 9723 12424 9735 12427
rect 9858 12424 9864 12436
rect 9723 12396 9864 12424
rect 9723 12393 9735 12396
rect 9677 12387 9735 12393
rect 9858 12384 9864 12396
rect 9916 12384 9922 12436
rect 10778 12424 10784 12436
rect 10152 12396 10784 12424
rect 4430 12356 4436 12368
rect 4391 12328 4436 12356
rect 4430 12316 4436 12328
rect 4488 12316 4494 12368
rect 4982 12316 4988 12368
rect 5040 12356 5046 12368
rect 8481 12359 8539 12365
rect 8481 12356 8493 12359
rect 5040 12328 8493 12356
rect 5040 12316 5046 12328
rect 8481 12325 8493 12328
rect 8527 12325 8539 12359
rect 8481 12319 8539 12325
rect 8754 12316 8760 12368
rect 8812 12356 8818 12368
rect 10152 12356 10180 12396
rect 10778 12384 10784 12396
rect 10836 12384 10842 12436
rect 10962 12384 10968 12436
rect 11020 12424 11026 12436
rect 11606 12424 11612 12436
rect 11020 12396 11284 12424
rect 11567 12396 11612 12424
rect 11020 12384 11026 12396
rect 10410 12356 10416 12368
rect 8812 12328 10180 12356
rect 10244 12328 10416 12356
rect 8812 12316 8818 12328
rect 2133 12291 2191 12297
rect 2133 12257 2145 12291
rect 2179 12288 2191 12291
rect 2774 12288 2780 12300
rect 2179 12260 2780 12288
rect 2179 12257 2191 12260
rect 2133 12251 2191 12257
rect 2774 12248 2780 12260
rect 2832 12248 2838 12300
rect 3237 12291 3295 12297
rect 3237 12257 3249 12291
rect 3283 12288 3295 12291
rect 3510 12288 3516 12300
rect 3283 12260 3516 12288
rect 3283 12257 3295 12260
rect 3237 12251 3295 12257
rect 3510 12248 3516 12260
rect 3568 12248 3574 12300
rect 5077 12291 5135 12297
rect 5077 12288 5089 12291
rect 4540 12260 5089 12288
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12189 2467 12223
rect 3418 12220 3424 12232
rect 3379 12192 3424 12220
rect 2409 12183 2467 12189
rect 1670 12112 1676 12164
rect 1728 12152 1734 12164
rect 2424 12152 2452 12183
rect 3418 12180 3424 12192
rect 3476 12180 3482 12232
rect 3970 12180 3976 12232
rect 4028 12220 4034 12232
rect 4540 12220 4568 12260
rect 5077 12257 5089 12260
rect 5123 12257 5135 12291
rect 5077 12251 5135 12257
rect 5534 12248 5540 12300
rect 5592 12288 5598 12300
rect 6178 12297 6184 12300
rect 5905 12291 5963 12297
rect 5905 12288 5917 12291
rect 5592 12260 5917 12288
rect 5592 12248 5598 12260
rect 5905 12257 5917 12260
rect 5951 12257 5963 12291
rect 6172 12288 6184 12297
rect 6139 12260 6184 12288
rect 5905 12251 5963 12257
rect 6172 12251 6184 12260
rect 6178 12248 6184 12251
rect 6236 12248 6242 12300
rect 7098 12248 7104 12300
rect 7156 12288 7162 12300
rect 7558 12288 7564 12300
rect 7156 12260 7564 12288
rect 7156 12248 7162 12260
rect 7558 12248 7564 12260
rect 7616 12248 7622 12300
rect 8389 12291 8447 12297
rect 8389 12257 8401 12291
rect 8435 12288 8447 12291
rect 9214 12288 9220 12300
rect 8435 12260 9220 12288
rect 8435 12257 8447 12260
rect 8389 12251 8447 12257
rect 9214 12248 9220 12260
rect 9272 12248 9278 12300
rect 4028 12192 4568 12220
rect 4709 12223 4767 12229
rect 4028 12180 4034 12192
rect 4709 12189 4721 12223
rect 4755 12220 4767 12223
rect 4798 12220 4804 12232
rect 4755 12192 4804 12220
rect 4755 12189 4767 12192
rect 4709 12183 4767 12189
rect 4798 12180 4804 12192
rect 4856 12180 4862 12232
rect 4893 12223 4951 12229
rect 4893 12189 4905 12223
rect 4939 12220 4951 12223
rect 5166 12220 5172 12232
rect 4939 12192 5172 12220
rect 4939 12189 4951 12192
rect 4893 12183 4951 12189
rect 5166 12180 5172 12192
rect 5224 12180 5230 12232
rect 8570 12180 8576 12232
rect 8628 12220 8634 12232
rect 8628 12192 8673 12220
rect 8628 12180 8634 12192
rect 9858 12180 9864 12232
rect 9916 12220 9922 12232
rect 10244 12229 10272 12328
rect 10410 12316 10416 12328
rect 10468 12316 10474 12368
rect 10686 12316 10692 12368
rect 10744 12356 10750 12368
rect 11256 12356 11284 12396
rect 11606 12384 11612 12396
rect 11664 12384 11670 12436
rect 11882 12424 11888 12436
rect 11843 12396 11888 12424
rect 11882 12384 11888 12396
rect 11940 12384 11946 12436
rect 13814 12384 13820 12436
rect 13872 12424 13878 12436
rect 15102 12424 15108 12436
rect 13872 12396 15108 12424
rect 13872 12384 13878 12396
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 12253 12359 12311 12365
rect 12253 12356 12265 12359
rect 10744 12328 11183 12356
rect 11256 12328 12265 12356
rect 10744 12316 10750 12328
rect 10496 12291 10554 12297
rect 10496 12257 10508 12291
rect 10542 12288 10554 12291
rect 11054 12288 11060 12300
rect 10542 12260 11060 12288
rect 10542 12257 10554 12260
rect 10496 12251 10554 12257
rect 11054 12248 11060 12260
rect 11112 12248 11118 12300
rect 11155 12288 11183 12328
rect 12253 12325 12265 12328
rect 12299 12325 12311 12359
rect 12253 12319 12311 12325
rect 13716 12359 13774 12365
rect 13716 12325 13728 12359
rect 13762 12356 13774 12359
rect 14274 12356 14280 12368
rect 13762 12328 14280 12356
rect 13762 12325 13774 12328
rect 13716 12319 13774 12325
rect 14274 12316 14280 12328
rect 14332 12316 14338 12368
rect 14550 12288 14556 12300
rect 11155 12260 14556 12288
rect 14550 12248 14556 12260
rect 14608 12248 14614 12300
rect 10229 12223 10287 12229
rect 10229 12220 10241 12223
rect 9916 12192 10241 12220
rect 9916 12180 9922 12192
rect 10229 12189 10241 12192
rect 10275 12189 10287 12223
rect 12342 12220 12348 12232
rect 12303 12192 12348 12220
rect 10229 12183 10287 12189
rect 12342 12180 12348 12192
rect 12400 12180 12406 12232
rect 12437 12223 12495 12229
rect 12437 12189 12449 12223
rect 12483 12189 12495 12223
rect 12437 12183 12495 12189
rect 3694 12152 3700 12164
rect 1728 12124 3700 12152
rect 1728 12112 1734 12124
rect 3694 12112 3700 12124
rect 3752 12112 3758 12164
rect 4246 12112 4252 12164
rect 4304 12152 4310 12164
rect 5261 12155 5319 12161
rect 5261 12152 5273 12155
rect 4304 12124 5273 12152
rect 4304 12112 4310 12124
rect 5261 12121 5273 12124
rect 5307 12121 5319 12155
rect 5261 12115 5319 12121
rect 7190 12112 7196 12164
rect 7248 12152 7254 12164
rect 7558 12152 7564 12164
rect 7248 12124 7564 12152
rect 7248 12112 7254 12124
rect 7558 12112 7564 12124
rect 7616 12152 7622 12164
rect 7616 12124 8156 12152
rect 7616 12112 7622 12124
rect 4065 12087 4123 12093
rect 4065 12053 4077 12087
rect 4111 12084 4123 12087
rect 4893 12087 4951 12093
rect 4893 12084 4905 12087
rect 4111 12056 4905 12084
rect 4111 12053 4123 12056
rect 4065 12047 4123 12053
rect 4893 12053 4905 12056
rect 4939 12053 4951 12087
rect 7282 12084 7288 12096
rect 7243 12056 7288 12084
rect 4893 12047 4951 12053
rect 7282 12044 7288 12056
rect 7340 12044 7346 12096
rect 7374 12044 7380 12096
rect 7432 12084 7438 12096
rect 8021 12087 8079 12093
rect 8021 12084 8033 12087
rect 7432 12056 8033 12084
rect 7432 12044 7438 12056
rect 8021 12053 8033 12056
rect 8067 12053 8079 12087
rect 8128 12084 8156 12124
rect 11606 12112 11612 12164
rect 11664 12152 11670 12164
rect 12452 12152 12480 12183
rect 12526 12180 12532 12232
rect 12584 12220 12590 12232
rect 13449 12223 13507 12229
rect 13449 12220 13461 12223
rect 12584 12192 13461 12220
rect 12584 12180 12590 12192
rect 13449 12189 13461 12192
rect 13495 12189 13507 12223
rect 13449 12183 13507 12189
rect 11664 12124 12480 12152
rect 11664 12112 11670 12124
rect 11698 12084 11704 12096
rect 8128 12056 11704 12084
rect 8021 12047 8079 12053
rect 11698 12044 11704 12056
rect 11756 12044 11762 12096
rect 14458 12044 14464 12096
rect 14516 12084 14522 12096
rect 14829 12087 14887 12093
rect 14829 12084 14841 12087
rect 14516 12056 14841 12084
rect 14516 12044 14522 12056
rect 14829 12053 14841 12056
rect 14875 12053 14887 12087
rect 14829 12047 14887 12053
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 3970 11880 3976 11892
rect 1872 11852 3976 11880
rect 1872 11753 1900 11852
rect 3970 11840 3976 11852
rect 4028 11840 4034 11892
rect 4154 11840 4160 11892
rect 4212 11880 4218 11892
rect 4985 11883 5043 11889
rect 4985 11880 4997 11883
rect 4212 11852 4997 11880
rect 4212 11840 4218 11852
rect 4985 11849 4997 11852
rect 5031 11849 5043 11883
rect 4985 11843 5043 11849
rect 6730 11840 6736 11892
rect 6788 11880 6794 11892
rect 6825 11883 6883 11889
rect 6825 11880 6837 11883
rect 6788 11852 6837 11880
rect 6788 11840 6794 11852
rect 6825 11849 6837 11852
rect 6871 11849 6883 11883
rect 6825 11843 6883 11849
rect 7006 11840 7012 11892
rect 7064 11880 7070 11892
rect 7466 11880 7472 11892
rect 7064 11852 7472 11880
rect 7064 11840 7070 11852
rect 7466 11840 7472 11852
rect 7524 11840 7530 11892
rect 10042 11840 10048 11892
rect 10100 11880 10106 11892
rect 10594 11880 10600 11892
rect 10100 11852 10600 11880
rect 10100 11840 10106 11852
rect 10594 11840 10600 11852
rect 10652 11840 10658 11892
rect 10686 11840 10692 11892
rect 10744 11840 10750 11892
rect 10873 11883 10931 11889
rect 10873 11849 10885 11883
rect 10919 11880 10931 11883
rect 12342 11880 12348 11892
rect 10919 11852 12348 11880
rect 10919 11849 10931 11852
rect 10873 11843 10931 11849
rect 12342 11840 12348 11852
rect 12400 11840 12406 11892
rect 13630 11880 13636 11892
rect 12452 11852 13636 11880
rect 3418 11772 3424 11824
rect 3476 11772 3482 11824
rect 3694 11812 3700 11824
rect 3607 11784 3700 11812
rect 3694 11772 3700 11784
rect 3752 11812 3758 11824
rect 3752 11784 5580 11812
rect 3752 11772 3758 11784
rect 1857 11747 1915 11753
rect 1857 11713 1869 11747
rect 1903 11713 1915 11747
rect 1857 11707 1915 11713
rect 3436 11744 3464 11772
rect 4525 11747 4583 11753
rect 4525 11744 4537 11747
rect 3436 11716 4537 11744
rect 1578 11676 1584 11688
rect 1539 11648 1584 11676
rect 1578 11636 1584 11648
rect 1636 11636 1642 11688
rect 2222 11636 2228 11688
rect 2280 11676 2286 11688
rect 2317 11679 2375 11685
rect 2317 11676 2329 11679
rect 2280 11648 2329 11676
rect 2280 11636 2286 11648
rect 2317 11645 2329 11648
rect 2363 11645 2375 11679
rect 2317 11639 2375 11645
rect 2584 11679 2642 11685
rect 2584 11645 2596 11679
rect 2630 11676 2642 11679
rect 3436 11676 3464 11716
rect 4525 11713 4537 11716
rect 4571 11744 4583 11747
rect 4798 11744 4804 11756
rect 4571 11716 4804 11744
rect 4571 11713 4583 11716
rect 4525 11707 4583 11713
rect 4798 11704 4804 11716
rect 4856 11704 4862 11756
rect 5166 11704 5172 11756
rect 5224 11744 5230 11756
rect 5552 11753 5580 11784
rect 7098 11772 7104 11824
rect 7156 11812 7162 11824
rect 7742 11812 7748 11824
rect 7156 11784 7748 11812
rect 7156 11772 7162 11784
rect 7742 11772 7748 11784
rect 7800 11772 7806 11824
rect 10704 11812 10732 11840
rect 12452 11812 12480 11852
rect 13630 11840 13636 11852
rect 13688 11840 13694 11892
rect 13814 11880 13820 11892
rect 13775 11852 13820 11880
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 14093 11883 14151 11889
rect 14093 11849 14105 11883
rect 14139 11880 14151 11883
rect 15930 11880 15936 11892
rect 14139 11852 15936 11880
rect 14139 11849 14151 11852
rect 14093 11843 14151 11849
rect 15930 11840 15936 11852
rect 15988 11840 15994 11892
rect 7843 11784 10732 11812
rect 10980 11784 12480 11812
rect 5445 11747 5503 11753
rect 5445 11744 5457 11747
rect 5224 11716 5457 11744
rect 5224 11704 5230 11716
rect 5445 11713 5457 11716
rect 5491 11713 5503 11747
rect 5445 11707 5503 11713
rect 5537 11747 5595 11753
rect 5537 11713 5549 11747
rect 5583 11713 5595 11747
rect 5537 11707 5595 11713
rect 6914 11704 6920 11756
rect 6972 11744 6978 11756
rect 7377 11747 7435 11753
rect 7377 11744 7389 11747
rect 6972 11716 7389 11744
rect 6972 11704 6978 11716
rect 7377 11713 7389 11716
rect 7423 11713 7435 11747
rect 7377 11707 7435 11713
rect 2630 11648 3464 11676
rect 2630 11645 2642 11648
rect 2584 11639 2642 11645
rect 3694 11636 3700 11688
rect 3752 11676 3758 11688
rect 4341 11679 4399 11685
rect 4341 11676 4353 11679
rect 3752 11648 4353 11676
rect 3752 11636 3758 11648
rect 4341 11645 4353 11648
rect 4387 11645 4399 11679
rect 4341 11639 4399 11645
rect 5902 11636 5908 11688
rect 5960 11676 5966 11688
rect 7193 11679 7251 11685
rect 7193 11676 7205 11679
rect 5960 11648 7205 11676
rect 5960 11636 5966 11648
rect 7193 11645 7205 11648
rect 7239 11676 7251 11679
rect 7843 11676 7871 11784
rect 8478 11744 8484 11756
rect 7239 11648 7871 11676
rect 8220 11716 8484 11744
rect 7239 11645 7251 11648
rect 7193 11639 7251 11645
rect 5353 11611 5411 11617
rect 5353 11608 5365 11611
rect 3988 11580 5365 11608
rect 3988 11549 4016 11580
rect 5353 11577 5365 11580
rect 5399 11577 5411 11611
rect 5353 11571 5411 11577
rect 5994 11568 6000 11620
rect 6052 11608 6058 11620
rect 7285 11611 7343 11617
rect 7285 11608 7297 11611
rect 6052 11580 7297 11608
rect 6052 11568 6058 11580
rect 7285 11577 7297 11580
rect 7331 11608 7343 11611
rect 8220 11608 8248 11716
rect 8478 11704 8484 11716
rect 8536 11704 8542 11756
rect 9582 11704 9588 11756
rect 9640 11744 9646 11756
rect 10318 11744 10324 11756
rect 9640 11716 10324 11744
rect 9640 11704 9646 11716
rect 10318 11704 10324 11716
rect 10376 11704 10382 11756
rect 8389 11679 8447 11685
rect 8389 11645 8401 11679
rect 8435 11676 8447 11679
rect 10980 11676 11008 11784
rect 11054 11704 11060 11756
rect 11112 11744 11118 11756
rect 11425 11747 11483 11753
rect 11425 11744 11437 11747
rect 11112 11716 11437 11744
rect 11112 11704 11118 11716
rect 11425 11713 11437 11716
rect 11471 11713 11483 11747
rect 12434 11744 12440 11756
rect 12395 11716 12440 11744
rect 11425 11707 11483 11713
rect 12434 11704 12440 11716
rect 12492 11704 12498 11756
rect 13814 11704 13820 11756
rect 13872 11744 13878 11756
rect 14645 11747 14703 11753
rect 14645 11744 14657 11747
rect 13872 11716 14657 11744
rect 13872 11704 13878 11716
rect 14645 11713 14657 11716
rect 14691 11713 14703 11747
rect 14645 11707 14703 11713
rect 16945 11747 17003 11753
rect 16945 11713 16957 11747
rect 16991 11744 17003 11747
rect 17218 11744 17224 11756
rect 16991 11716 17224 11744
rect 16991 11713 17003 11716
rect 16945 11707 17003 11713
rect 17218 11704 17224 11716
rect 17276 11704 17282 11756
rect 8435 11648 11008 11676
rect 11241 11679 11299 11685
rect 8435 11645 8447 11648
rect 8389 11639 8447 11645
rect 11241 11645 11253 11679
rect 11287 11676 11299 11679
rect 12342 11676 12348 11688
rect 11287 11648 12348 11676
rect 11287 11645 11299 11648
rect 11241 11639 11299 11645
rect 12342 11636 12348 11648
rect 12400 11676 12406 11688
rect 12400 11648 13584 11676
rect 12400 11636 12406 11648
rect 7331 11580 8248 11608
rect 7331 11577 7343 11580
rect 7285 11571 7343 11577
rect 8478 11568 8484 11620
rect 8536 11608 8542 11620
rect 8536 11580 11836 11608
rect 8536 11568 8542 11580
rect 3973 11543 4031 11549
rect 3973 11509 3985 11543
rect 4019 11509 4031 11543
rect 3973 11503 4031 11509
rect 4433 11543 4491 11549
rect 4433 11509 4445 11543
rect 4479 11540 4491 11543
rect 5442 11540 5448 11552
rect 4479 11512 5448 11540
rect 4479 11509 4491 11512
rect 4433 11503 4491 11509
rect 5442 11500 5448 11512
rect 5500 11540 5506 11552
rect 6454 11540 6460 11552
rect 5500 11512 6460 11540
rect 5500 11500 5506 11512
rect 6454 11500 6460 11512
rect 6512 11500 6518 11552
rect 7466 11500 7472 11552
rect 7524 11540 7530 11552
rect 9306 11540 9312 11552
rect 7524 11512 9312 11540
rect 7524 11500 7530 11512
rect 9306 11500 9312 11512
rect 9364 11500 9370 11552
rect 9398 11500 9404 11552
rect 9456 11540 9462 11552
rect 9677 11543 9735 11549
rect 9677 11540 9689 11543
rect 9456 11512 9689 11540
rect 9456 11500 9462 11512
rect 9677 11509 9689 11512
rect 9723 11509 9735 11543
rect 9677 11503 9735 11509
rect 10318 11500 10324 11552
rect 10376 11540 10382 11552
rect 11333 11543 11391 11549
rect 11333 11540 11345 11543
rect 10376 11512 11345 11540
rect 10376 11500 10382 11512
rect 11333 11509 11345 11512
rect 11379 11509 11391 11543
rect 11808 11540 11836 11580
rect 12618 11568 12624 11620
rect 12676 11617 12682 11620
rect 12676 11611 12740 11617
rect 12676 11577 12694 11611
rect 12728 11608 12740 11611
rect 13354 11608 13360 11620
rect 12728 11580 13360 11608
rect 12728 11577 12740 11580
rect 12676 11571 12740 11577
rect 12676 11568 12682 11571
rect 13354 11568 13360 11580
rect 13412 11568 13418 11620
rect 13556 11608 13584 11648
rect 14090 11636 14096 11688
rect 14148 11676 14154 11688
rect 16669 11679 16727 11685
rect 16669 11676 16681 11679
rect 14148 11648 16681 11676
rect 14148 11636 14154 11648
rect 16669 11645 16681 11648
rect 16715 11645 16727 11679
rect 16669 11639 16727 11645
rect 17034 11608 17040 11620
rect 13556 11580 17040 11608
rect 17034 11568 17040 11580
rect 17092 11568 17098 11620
rect 13906 11540 13912 11552
rect 11808 11512 13912 11540
rect 11333 11503 11391 11509
rect 13906 11500 13912 11512
rect 13964 11500 13970 11552
rect 14274 11500 14280 11552
rect 14332 11540 14338 11552
rect 14461 11543 14519 11549
rect 14461 11540 14473 11543
rect 14332 11512 14473 11540
rect 14332 11500 14338 11512
rect 14461 11509 14473 11512
rect 14507 11509 14519 11543
rect 14461 11503 14519 11509
rect 14553 11543 14611 11549
rect 14553 11509 14565 11543
rect 14599 11540 14611 11543
rect 15102 11540 15108 11552
rect 14599 11512 15108 11540
rect 14599 11509 14611 11512
rect 14553 11503 14611 11509
rect 15102 11500 15108 11512
rect 15160 11500 15166 11552
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 2406 11296 2412 11348
rect 2464 11336 2470 11348
rect 2777 11339 2835 11345
rect 2777 11336 2789 11339
rect 2464 11308 2789 11336
rect 2464 11296 2470 11308
rect 2777 11305 2789 11308
rect 2823 11305 2835 11339
rect 4062 11336 4068 11348
rect 4023 11308 4068 11336
rect 2777 11299 2835 11305
rect 4062 11296 4068 11308
rect 4120 11296 4126 11348
rect 5350 11296 5356 11348
rect 5408 11336 5414 11348
rect 6917 11339 6975 11345
rect 6917 11336 6929 11339
rect 5408 11308 6929 11336
rect 5408 11296 5414 11308
rect 6917 11305 6929 11308
rect 6963 11305 6975 11339
rect 6917 11299 6975 11305
rect 7285 11339 7343 11345
rect 7285 11305 7297 11339
rect 7331 11336 7343 11339
rect 7374 11336 7380 11348
rect 7331 11308 7380 11336
rect 7331 11305 7343 11308
rect 7285 11299 7343 11305
rect 7374 11296 7380 11308
rect 7432 11296 7438 11348
rect 9309 11339 9367 11345
rect 9309 11336 9321 11339
rect 7576 11308 9321 11336
rect 1670 11277 1676 11280
rect 1664 11268 1676 11277
rect 1631 11240 1676 11268
rect 1664 11231 1676 11240
rect 1670 11228 1676 11231
rect 1728 11228 1734 11280
rect 3329 11271 3387 11277
rect 3329 11237 3341 11271
rect 3375 11268 3387 11271
rect 3786 11268 3792 11280
rect 3375 11240 3792 11268
rect 3375 11237 3387 11240
rect 3329 11231 3387 11237
rect 3786 11228 3792 11240
rect 3844 11228 3850 11280
rect 7466 11268 7472 11280
rect 5000 11240 7472 11268
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11200 1455 11203
rect 2222 11200 2228 11212
rect 1443 11172 2228 11200
rect 1443 11169 1455 11172
rect 1397 11163 1455 11169
rect 2222 11160 2228 11172
rect 2280 11160 2286 11212
rect 3050 11200 3056 11212
rect 3011 11172 3056 11200
rect 3050 11160 3056 11172
rect 3108 11160 3114 11212
rect 3602 11160 3608 11212
rect 3660 11200 3666 11212
rect 5000 11200 5028 11240
rect 7466 11228 7472 11240
rect 7524 11228 7530 11280
rect 3660 11172 5028 11200
rect 5068 11203 5126 11209
rect 3660 11160 3666 11172
rect 5068 11169 5080 11203
rect 5114 11200 5126 11203
rect 5810 11200 5816 11212
rect 5114 11172 5816 11200
rect 5114 11169 5126 11172
rect 5068 11163 5126 11169
rect 5810 11160 5816 11172
rect 5868 11160 5874 11212
rect 4246 11092 4252 11144
rect 4304 11132 4310 11144
rect 7576 11141 7604 11308
rect 9309 11305 9321 11308
rect 9355 11336 9367 11339
rect 9582 11336 9588 11348
rect 9355 11308 9588 11336
rect 9355 11305 9367 11308
rect 9309 11299 9367 11305
rect 9582 11296 9588 11308
rect 9640 11296 9646 11348
rect 9674 11296 9680 11348
rect 9732 11296 9738 11348
rect 11054 11336 11060 11348
rect 11015 11308 11060 11336
rect 11054 11296 11060 11308
rect 11112 11296 11118 11348
rect 11698 11296 11704 11348
rect 11756 11336 11762 11348
rect 12710 11336 12716 11348
rect 11756 11308 12716 11336
rect 11756 11296 11762 11308
rect 12710 11296 12716 11308
rect 12768 11336 12774 11348
rect 12805 11339 12863 11345
rect 12805 11336 12817 11339
rect 12768 11308 12817 11336
rect 12768 11296 12774 11308
rect 12805 11305 12817 11308
rect 12851 11305 12863 11339
rect 12805 11299 12863 11305
rect 12894 11296 12900 11348
rect 12952 11336 12958 11348
rect 13081 11339 13139 11345
rect 13081 11336 13093 11339
rect 12952 11308 13093 11336
rect 12952 11296 12958 11308
rect 13081 11305 13093 11308
rect 13127 11305 13139 11339
rect 14090 11336 14096 11348
rect 14051 11308 14096 11336
rect 13081 11299 13139 11305
rect 14090 11296 14096 11308
rect 14148 11296 14154 11348
rect 8196 11271 8254 11277
rect 8196 11237 8208 11271
rect 8242 11268 8254 11271
rect 8570 11268 8576 11280
rect 8242 11240 8576 11268
rect 8242 11237 8254 11240
rect 8196 11231 8254 11237
rect 8570 11228 8576 11240
rect 8628 11228 8634 11280
rect 9692 11268 9720 11296
rect 9922 11271 9980 11277
rect 9922 11268 9934 11271
rect 9692 11240 9934 11268
rect 9922 11237 9934 11240
rect 9968 11237 9980 11271
rect 9922 11231 9980 11237
rect 8754 11200 8760 11212
rect 7852 11172 8760 11200
rect 4801 11135 4859 11141
rect 4801 11132 4813 11135
rect 4304 11104 4813 11132
rect 4304 11092 4310 11104
rect 4801 11101 4813 11104
rect 4847 11101 4859 11135
rect 4801 11095 4859 11101
rect 7377 11135 7435 11141
rect 7377 11101 7389 11135
rect 7423 11101 7435 11135
rect 7377 11095 7435 11101
rect 7561 11135 7619 11141
rect 7561 11101 7573 11135
rect 7607 11101 7619 11135
rect 7561 11095 7619 11101
rect 6178 11064 6184 11076
rect 6091 11036 6184 11064
rect 6178 11024 6184 11036
rect 6236 11064 6242 11076
rect 7392 11064 7420 11095
rect 7742 11064 7748 11076
rect 6236 11036 7328 11064
rect 7392 11036 7748 11064
rect 6236 11024 6242 11036
rect 3970 10956 3976 11008
rect 4028 10996 4034 11008
rect 7006 10996 7012 11008
rect 4028 10968 7012 10996
rect 4028 10956 4034 10968
rect 7006 10956 7012 10968
rect 7064 10956 7070 11008
rect 7300 10996 7328 11036
rect 7742 11024 7748 11036
rect 7800 11024 7806 11076
rect 7852 10996 7880 11172
rect 8754 11160 8760 11172
rect 8812 11160 8818 11212
rect 9582 11160 9588 11212
rect 9640 11200 9646 11212
rect 11698 11209 11704 11212
rect 9677 11203 9735 11209
rect 9677 11200 9689 11203
rect 9640 11172 9689 11200
rect 9640 11160 9646 11172
rect 9677 11169 9689 11172
rect 9723 11169 9735 11203
rect 9677 11163 9735 11169
rect 11692 11163 11704 11209
rect 11756 11200 11762 11212
rect 11756 11172 11792 11200
rect 11698 11160 11704 11163
rect 11756 11160 11762 11172
rect 12434 11160 12440 11212
rect 12492 11200 12498 11212
rect 13170 11200 13176 11212
rect 12492 11172 13176 11200
rect 12492 11160 12498 11172
rect 13170 11160 13176 11172
rect 13228 11200 13234 11212
rect 13449 11203 13507 11209
rect 13449 11200 13461 11203
rect 13228 11172 13461 11200
rect 13228 11160 13234 11172
rect 13449 11169 13461 11172
rect 13495 11169 13507 11203
rect 13449 11163 13507 11169
rect 13541 11203 13599 11209
rect 13541 11169 13553 11203
rect 13587 11200 13599 11203
rect 13587 11172 13768 11200
rect 13587 11169 13599 11172
rect 13541 11163 13599 11169
rect 7929 11135 7987 11141
rect 7929 11101 7941 11135
rect 7975 11101 7987 11135
rect 7929 11095 7987 11101
rect 7300 10968 7880 10996
rect 7944 10996 7972 11095
rect 11054 11092 11060 11144
rect 11112 11132 11118 11144
rect 11425 11135 11483 11141
rect 11425 11132 11437 11135
rect 11112 11104 11437 11132
rect 11112 11092 11118 11104
rect 11425 11101 11437 11104
rect 11471 11101 11483 11135
rect 13630 11132 13636 11144
rect 13591 11104 13636 11132
rect 11425 11095 11483 11101
rect 13630 11092 13636 11104
rect 13688 11092 13694 11144
rect 13740 11132 13768 11172
rect 13814 11160 13820 11212
rect 13872 11200 13878 11212
rect 14461 11203 14519 11209
rect 14461 11200 14473 11203
rect 13872 11172 14473 11200
rect 13872 11160 13878 11172
rect 14461 11169 14473 11172
rect 14507 11169 14519 11203
rect 14461 11163 14519 11169
rect 13740 11104 13952 11132
rect 12710 11024 12716 11076
rect 12768 11064 12774 11076
rect 13924 11064 13952 11104
rect 13998 11092 14004 11144
rect 14056 11132 14062 11144
rect 14553 11135 14611 11141
rect 14553 11132 14565 11135
rect 14056 11104 14565 11132
rect 14056 11092 14062 11104
rect 14553 11101 14565 11104
rect 14599 11101 14611 11135
rect 14553 11095 14611 11101
rect 14642 11092 14648 11144
rect 14700 11132 14706 11144
rect 14700 11104 14745 11132
rect 14700 11092 14706 11104
rect 17126 11064 17132 11076
rect 12768 11036 17132 11064
rect 12768 11024 12774 11036
rect 17126 11024 17132 11036
rect 17184 11024 17190 11076
rect 8662 10996 8668 11008
rect 7944 10968 8668 10996
rect 8662 10956 8668 10968
rect 8720 10956 8726 11008
rect 10870 10956 10876 11008
rect 10928 10996 10934 11008
rect 11606 10996 11612 11008
rect 10928 10968 11612 10996
rect 10928 10956 10934 10968
rect 11606 10956 11612 10968
rect 11664 10996 11670 11008
rect 16758 10996 16764 11008
rect 11664 10968 16764 10996
rect 11664 10956 11670 10968
rect 16758 10956 16764 10968
rect 16816 10956 16822 11008
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 4062 10752 4068 10804
rect 4120 10792 4126 10804
rect 4120 10764 8524 10792
rect 4120 10752 4126 10764
rect 5810 10724 5816 10736
rect 5723 10696 5816 10724
rect 5810 10684 5816 10696
rect 5868 10684 5874 10736
rect 6914 10684 6920 10736
rect 6972 10724 6978 10736
rect 7190 10724 7196 10736
rect 6972 10696 7196 10724
rect 6972 10684 6978 10696
rect 7190 10684 7196 10696
rect 7248 10684 7254 10736
rect 8496 10724 8524 10764
rect 8570 10752 8576 10804
rect 8628 10792 8634 10804
rect 8754 10792 8760 10804
rect 8628 10764 8760 10792
rect 8628 10752 8634 10764
rect 8754 10752 8760 10764
rect 8812 10792 8818 10804
rect 8941 10795 8999 10801
rect 8941 10792 8953 10795
rect 8812 10764 8953 10792
rect 8812 10752 8818 10764
rect 8941 10761 8953 10764
rect 8987 10761 8999 10795
rect 10870 10792 10876 10804
rect 8941 10755 8999 10761
rect 9692 10764 10876 10792
rect 9692 10724 9720 10764
rect 10870 10752 10876 10764
rect 10928 10752 10934 10804
rect 11057 10795 11115 10801
rect 11057 10761 11069 10795
rect 11103 10792 11115 10795
rect 11103 10764 11183 10792
rect 11103 10761 11115 10764
rect 11057 10755 11115 10761
rect 8496 10696 9720 10724
rect 11155 10724 11183 10764
rect 12986 10752 12992 10804
rect 13044 10792 13050 10804
rect 13265 10795 13323 10801
rect 13265 10792 13277 10795
rect 13044 10764 13277 10792
rect 13044 10752 13050 10764
rect 13265 10761 13277 10764
rect 13311 10761 13323 10795
rect 13265 10755 13323 10761
rect 13449 10795 13507 10801
rect 13449 10761 13461 10795
rect 13495 10792 13507 10795
rect 14274 10792 14280 10804
rect 13495 10764 14280 10792
rect 13495 10761 13507 10764
rect 13449 10755 13507 10761
rect 11155 10696 11284 10724
rect 3142 10616 3148 10668
rect 3200 10656 3206 10668
rect 3697 10659 3755 10665
rect 3697 10656 3709 10659
rect 3200 10628 3709 10656
rect 3200 10616 3206 10628
rect 3697 10625 3709 10628
rect 3743 10625 3755 10659
rect 5828 10656 5856 10684
rect 11256 10668 11284 10696
rect 12802 10684 12808 10736
rect 12860 10724 12866 10736
rect 13078 10724 13084 10736
rect 12860 10696 13084 10724
rect 12860 10684 12866 10696
rect 13078 10684 13084 10696
rect 13136 10684 13142 10736
rect 5828 10628 7696 10656
rect 3697 10619 3755 10625
rect 2041 10591 2099 10597
rect 2041 10557 2053 10591
rect 2087 10588 2099 10591
rect 2130 10588 2136 10600
rect 2087 10560 2136 10588
rect 2087 10557 2099 10560
rect 2041 10551 2099 10557
rect 2130 10548 2136 10560
rect 2188 10548 2194 10600
rect 4246 10548 4252 10600
rect 4304 10588 4310 10600
rect 4433 10591 4491 10597
rect 4433 10588 4445 10591
rect 4304 10560 4445 10588
rect 4304 10548 4310 10560
rect 4433 10557 4445 10560
rect 4479 10588 4491 10591
rect 6362 10588 6368 10600
rect 4479 10560 6368 10588
rect 4479 10557 4491 10560
rect 4433 10551 4491 10557
rect 6362 10548 6368 10560
rect 6420 10588 6426 10600
rect 7561 10591 7619 10597
rect 7561 10588 7573 10591
rect 6420 10560 7573 10588
rect 6420 10548 6426 10560
rect 7561 10557 7573 10560
rect 7607 10557 7619 10591
rect 7668 10588 7696 10628
rect 8662 10616 8668 10668
rect 8720 10656 8726 10668
rect 9214 10656 9220 10668
rect 8720 10628 9076 10656
rect 9175 10628 9220 10656
rect 8720 10616 8726 10628
rect 8570 10588 8576 10600
rect 7668 10560 8576 10588
rect 7561 10551 7619 10557
rect 8570 10548 8576 10560
rect 8628 10548 8634 10600
rect 9048 10588 9076 10628
rect 9214 10616 9220 10628
rect 9272 10616 9278 10668
rect 11238 10616 11244 10668
rect 11296 10656 11302 10668
rect 11793 10659 11851 10665
rect 11793 10656 11805 10659
rect 11296 10628 11805 10656
rect 11296 10616 11302 10628
rect 11793 10625 11805 10628
rect 11839 10656 11851 10659
rect 12986 10656 12992 10668
rect 11839 10628 12992 10656
rect 11839 10625 11851 10628
rect 11793 10619 11851 10625
rect 12986 10616 12992 10628
rect 13044 10616 13050 10668
rect 9674 10588 9680 10600
rect 9048 10560 9680 10588
rect 9674 10548 9680 10560
rect 9732 10548 9738 10600
rect 9950 10597 9956 10600
rect 9944 10588 9956 10597
rect 9911 10560 9956 10588
rect 9944 10551 9956 10560
rect 9950 10548 9956 10551
rect 10008 10548 10014 10600
rect 10226 10548 10232 10600
rect 10284 10588 10290 10600
rect 11609 10591 11667 10597
rect 11609 10588 11621 10591
rect 10284 10560 11621 10588
rect 10284 10548 10290 10560
rect 11609 10557 11621 10560
rect 11655 10557 11667 10591
rect 13280 10588 13308 10755
rect 14274 10752 14280 10764
rect 14332 10752 14338 10804
rect 13354 10616 13360 10668
rect 13412 10656 13418 10668
rect 13998 10656 14004 10668
rect 13412 10628 14004 10656
rect 13412 10616 13418 10628
rect 13998 10616 14004 10628
rect 14056 10616 14062 10668
rect 13446 10588 13452 10600
rect 13280 10560 13452 10588
rect 11609 10551 11667 10557
rect 13446 10548 13452 10560
rect 13504 10588 13510 10600
rect 13909 10591 13967 10597
rect 13909 10588 13921 10591
rect 13504 10560 13921 10588
rect 13504 10548 13510 10560
rect 13909 10557 13921 10560
rect 13955 10557 13967 10591
rect 13909 10551 13967 10557
rect 2308 10523 2366 10529
rect 2308 10489 2320 10523
rect 2354 10520 2366 10523
rect 2406 10520 2412 10532
rect 2354 10492 2412 10520
rect 2354 10489 2366 10492
rect 2308 10483 2366 10489
rect 2406 10480 2412 10492
rect 2464 10480 2470 10532
rect 4700 10523 4758 10529
rect 4700 10489 4712 10523
rect 4746 10520 4758 10523
rect 5718 10520 5724 10532
rect 4746 10492 5724 10520
rect 4746 10489 4758 10492
rect 4700 10483 4758 10489
rect 5718 10480 5724 10492
rect 5776 10480 5782 10532
rect 6089 10523 6147 10529
rect 6089 10489 6101 10523
rect 6135 10520 6147 10523
rect 7650 10520 7656 10532
rect 6135 10492 7656 10520
rect 6135 10489 6147 10492
rect 6089 10483 6147 10489
rect 7650 10480 7656 10492
rect 7708 10480 7714 10532
rect 7828 10523 7886 10529
rect 7828 10489 7840 10523
rect 7874 10520 7886 10523
rect 8662 10520 8668 10532
rect 7874 10492 8668 10520
rect 7874 10489 7886 10492
rect 7828 10483 7886 10489
rect 8662 10480 8668 10492
rect 8720 10480 8726 10532
rect 13817 10523 13875 10529
rect 13817 10489 13829 10523
rect 13863 10520 13875 10523
rect 14461 10523 14519 10529
rect 14461 10520 14473 10523
rect 13863 10492 14473 10520
rect 13863 10489 13875 10492
rect 13817 10483 13875 10489
rect 14461 10489 14473 10492
rect 14507 10489 14519 10523
rect 14461 10483 14519 10489
rect 3421 10455 3479 10461
rect 3421 10421 3433 10455
rect 3467 10452 3479 10455
rect 4982 10452 4988 10464
rect 3467 10424 4988 10452
rect 3467 10421 3479 10424
rect 3421 10415 3479 10421
rect 4982 10412 4988 10424
rect 5040 10412 5046 10464
rect 6825 10455 6883 10461
rect 6825 10421 6837 10455
rect 6871 10452 6883 10455
rect 7190 10452 7196 10464
rect 6871 10424 7196 10452
rect 6871 10421 6883 10424
rect 6825 10415 6883 10421
rect 7190 10412 7196 10424
rect 7248 10412 7254 10464
rect 7282 10412 7288 10464
rect 7340 10452 7346 10464
rect 8202 10452 8208 10464
rect 7340 10424 8208 10452
rect 7340 10412 7346 10424
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 8846 10412 8852 10464
rect 8904 10452 8910 10464
rect 9214 10452 9220 10464
rect 8904 10424 9220 10452
rect 8904 10412 8910 10424
rect 9214 10412 9220 10424
rect 9272 10412 9278 10464
rect 9766 10412 9772 10464
rect 9824 10452 9830 10464
rect 9950 10452 9956 10464
rect 9824 10424 9956 10452
rect 9824 10412 9830 10424
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 11146 10452 11152 10464
rect 11107 10424 11152 10452
rect 11146 10412 11152 10424
rect 11204 10412 11210 10464
rect 11514 10452 11520 10464
rect 11475 10424 11520 10452
rect 11514 10412 11520 10424
rect 11572 10412 11578 10464
rect 11974 10452 11980 10464
rect 11935 10424 11980 10452
rect 11974 10412 11980 10424
rect 12032 10412 12038 10464
rect 12894 10412 12900 10464
rect 12952 10452 12958 10464
rect 16574 10452 16580 10464
rect 12952 10424 16580 10452
rect 12952 10412 12958 10424
rect 16574 10412 16580 10424
rect 16632 10412 16638 10464
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 1596 10220 3372 10248
rect 1596 10121 1624 10220
rect 1857 10183 1915 10189
rect 1857 10149 1869 10183
rect 1903 10180 1915 10183
rect 3234 10180 3240 10192
rect 1903 10152 3240 10180
rect 1903 10149 1915 10152
rect 1857 10143 1915 10149
rect 3234 10140 3240 10152
rect 3292 10140 3298 10192
rect 3344 10180 3372 10220
rect 3418 10208 3424 10260
rect 3476 10248 3482 10260
rect 3697 10251 3755 10257
rect 3697 10248 3709 10251
rect 3476 10220 3709 10248
rect 3476 10208 3482 10220
rect 3697 10217 3709 10220
rect 3743 10217 3755 10251
rect 3697 10211 3755 10217
rect 4706 10208 4712 10260
rect 4764 10248 4770 10260
rect 5537 10251 5595 10257
rect 5537 10248 5549 10251
rect 4764 10220 5549 10248
rect 4764 10208 4770 10220
rect 5537 10217 5549 10220
rect 5583 10217 5595 10251
rect 5537 10211 5595 10217
rect 6273 10251 6331 10257
rect 6273 10217 6285 10251
rect 6319 10248 6331 10251
rect 7466 10248 7472 10260
rect 6319 10220 7472 10248
rect 6319 10217 6331 10220
rect 6273 10211 6331 10217
rect 7466 10208 7472 10220
rect 7524 10208 7530 10260
rect 7745 10251 7803 10257
rect 7745 10217 7757 10251
rect 7791 10248 7803 10251
rect 8662 10248 8668 10260
rect 7791 10220 8668 10248
rect 7791 10217 7803 10220
rect 7745 10211 7803 10217
rect 8662 10208 8668 10220
rect 8720 10208 8726 10260
rect 9674 10208 9680 10260
rect 9732 10248 9738 10260
rect 9861 10251 9919 10257
rect 9861 10248 9873 10251
rect 9732 10220 9873 10248
rect 9732 10208 9738 10220
rect 9861 10217 9873 10220
rect 9907 10248 9919 10251
rect 11054 10248 11060 10260
rect 9907 10220 11060 10248
rect 9907 10217 9919 10220
rect 9861 10211 9919 10217
rect 7374 10180 7380 10192
rect 3344 10152 7380 10180
rect 7374 10140 7380 10152
rect 7432 10140 7438 10192
rect 8202 10140 8208 10192
rect 8260 10180 8266 10192
rect 10502 10180 10508 10192
rect 8260 10152 10508 10180
rect 8260 10140 8266 10152
rect 10502 10140 10508 10152
rect 10560 10140 10566 10192
rect 10612 10124 10640 10220
rect 11054 10208 11060 10220
rect 11112 10208 11118 10260
rect 11698 10208 11704 10260
rect 11756 10248 11762 10260
rect 11977 10251 12035 10257
rect 11977 10248 11989 10251
rect 11756 10220 11989 10248
rect 11756 10208 11762 10220
rect 11977 10217 11989 10220
rect 12023 10217 12035 10251
rect 11977 10211 12035 10217
rect 12437 10251 12495 10257
rect 12437 10217 12449 10251
rect 12483 10217 12495 10251
rect 12894 10248 12900 10260
rect 12855 10220 12900 10248
rect 12437 10211 12495 10217
rect 10864 10183 10922 10189
rect 10864 10149 10876 10183
rect 10910 10180 10922 10183
rect 11238 10180 11244 10192
rect 10910 10152 11244 10180
rect 10910 10149 10922 10152
rect 10864 10143 10922 10149
rect 11238 10140 11244 10152
rect 11296 10140 11302 10192
rect 11514 10140 11520 10192
rect 11572 10180 11578 10192
rect 12452 10180 12480 10211
rect 12894 10208 12900 10220
rect 12952 10208 12958 10260
rect 13265 10251 13323 10257
rect 13265 10217 13277 10251
rect 13311 10248 13323 10251
rect 15102 10248 15108 10260
rect 13311 10220 15108 10248
rect 13311 10217 13323 10220
rect 13265 10211 13323 10217
rect 15102 10208 15108 10220
rect 15160 10208 15166 10260
rect 11572 10152 12480 10180
rect 11572 10140 11578 10152
rect 12526 10140 12532 10192
rect 12584 10180 12590 10192
rect 13633 10183 13691 10189
rect 13633 10180 13645 10183
rect 12584 10152 13645 10180
rect 12584 10140 12590 10152
rect 13633 10149 13645 10152
rect 13679 10149 13691 10183
rect 13633 10143 13691 10149
rect 1581 10115 1639 10121
rect 1581 10081 1593 10115
rect 1627 10081 1639 10115
rect 1581 10075 1639 10081
rect 2584 10115 2642 10121
rect 2584 10081 2596 10115
rect 2630 10112 2642 10115
rect 2866 10112 2872 10124
rect 2630 10084 2872 10112
rect 2630 10081 2642 10084
rect 2584 10075 2642 10081
rect 2866 10072 2872 10084
rect 2924 10072 2930 10124
rect 3418 10072 3424 10124
rect 3476 10112 3482 10124
rect 3694 10112 3700 10124
rect 3476 10084 3700 10112
rect 3476 10072 3482 10084
rect 3694 10072 3700 10084
rect 3752 10072 3758 10124
rect 4433 10115 4491 10121
rect 4433 10081 4445 10115
rect 4479 10112 4491 10115
rect 4798 10112 4804 10124
rect 4479 10084 4804 10112
rect 4479 10081 4491 10084
rect 4433 10075 4491 10081
rect 4798 10072 4804 10084
rect 4856 10072 4862 10124
rect 5074 10072 5080 10124
rect 5132 10112 5138 10124
rect 5445 10115 5503 10121
rect 5445 10112 5457 10115
rect 5132 10084 5457 10112
rect 5132 10072 5138 10084
rect 5445 10081 5457 10084
rect 5491 10081 5503 10115
rect 6362 10112 6368 10124
rect 6323 10084 6368 10112
rect 5445 10075 5503 10081
rect 6362 10072 6368 10084
rect 6420 10072 6426 10124
rect 6454 10072 6460 10124
rect 6512 10112 6518 10124
rect 6621 10115 6679 10121
rect 6621 10112 6633 10115
rect 6512 10084 6633 10112
rect 6512 10072 6518 10084
rect 6621 10081 6633 10084
rect 6667 10081 6679 10115
rect 6621 10075 6679 10081
rect 8573 10115 8631 10121
rect 8573 10081 8585 10115
rect 8619 10112 8631 10115
rect 8846 10112 8852 10124
rect 8619 10084 8852 10112
rect 8619 10081 8631 10084
rect 8573 10075 8631 10081
rect 8846 10072 8852 10084
rect 8904 10072 8910 10124
rect 10045 10115 10103 10121
rect 10045 10081 10057 10115
rect 10091 10112 10103 10115
rect 10318 10112 10324 10124
rect 10091 10084 10324 10112
rect 10091 10081 10103 10084
rect 10045 10075 10103 10081
rect 10318 10072 10324 10084
rect 10376 10072 10382 10124
rect 10594 10112 10600 10124
rect 10507 10084 10600 10112
rect 10594 10072 10600 10084
rect 10652 10072 10658 10124
rect 10686 10072 10692 10124
rect 10744 10112 10750 10124
rect 10744 10084 11652 10112
rect 10744 10072 10750 10084
rect 2222 10004 2228 10056
rect 2280 10044 2286 10056
rect 2317 10047 2375 10053
rect 2317 10044 2329 10047
rect 2280 10016 2329 10044
rect 2280 10004 2286 10016
rect 2317 10013 2329 10016
rect 2363 10013 2375 10047
rect 2317 10007 2375 10013
rect 4525 10047 4583 10053
rect 4525 10013 4537 10047
rect 4571 10013 4583 10047
rect 4525 10007 4583 10013
rect 4709 10047 4767 10053
rect 4709 10013 4721 10047
rect 4755 10044 4767 10047
rect 4982 10044 4988 10056
rect 4755 10016 4988 10044
rect 4755 10013 4767 10016
rect 4709 10007 4767 10013
rect 4540 9976 4568 10007
rect 4982 10004 4988 10016
rect 5040 10004 5046 10056
rect 5718 10044 5724 10056
rect 5631 10016 5724 10044
rect 5718 10004 5724 10016
rect 5776 10044 5782 10056
rect 6273 10047 6331 10053
rect 6273 10044 6285 10047
rect 5776 10016 6285 10044
rect 5776 10004 5782 10016
rect 6273 10013 6285 10016
rect 6319 10013 6331 10047
rect 6273 10007 6331 10013
rect 8294 10004 8300 10056
rect 8352 10044 8358 10056
rect 8665 10047 8723 10053
rect 8665 10044 8677 10047
rect 8352 10016 8677 10044
rect 8352 10004 8358 10016
rect 8665 10013 8677 10016
rect 8711 10013 8723 10047
rect 8665 10007 8723 10013
rect 8754 10004 8760 10056
rect 8812 10044 8818 10056
rect 10137 10047 10195 10053
rect 8812 10016 8857 10044
rect 8812 10004 8818 10016
rect 10137 10013 10149 10047
rect 10183 10044 10195 10047
rect 10502 10044 10508 10056
rect 10183 10016 10508 10044
rect 10183 10013 10195 10016
rect 10137 10007 10195 10013
rect 10502 10004 10508 10016
rect 10560 10004 10566 10056
rect 11624 10044 11652 10084
rect 12618 10072 12624 10124
rect 12676 10112 12682 10124
rect 12805 10115 12863 10121
rect 12805 10112 12817 10115
rect 12676 10084 12817 10112
rect 12676 10072 12682 10084
rect 12805 10081 12817 10084
rect 12851 10081 12863 10115
rect 14458 10112 14464 10124
rect 12805 10075 12863 10081
rect 13096 10084 14464 10112
rect 13096 10053 13124 10084
rect 14458 10072 14464 10084
rect 14516 10072 14522 10124
rect 13081 10047 13139 10053
rect 13081 10044 13093 10047
rect 11624 10016 13093 10044
rect 13081 10013 13093 10016
rect 13127 10013 13139 10047
rect 13722 10044 13728 10056
rect 13683 10016 13728 10044
rect 13081 10007 13139 10013
rect 13722 10004 13728 10016
rect 13780 10004 13786 10056
rect 13909 10047 13967 10053
rect 13909 10013 13921 10047
rect 13955 10044 13967 10047
rect 13998 10044 14004 10056
rect 13955 10016 14004 10044
rect 13955 10013 13967 10016
rect 13909 10007 13967 10013
rect 13998 10004 14004 10016
rect 14056 10004 14062 10056
rect 5810 9976 5816 9988
rect 4540 9948 5816 9976
rect 5810 9936 5816 9948
rect 5868 9936 5874 9988
rect 7668 9948 9996 9976
rect 3786 9868 3792 9920
rect 3844 9908 3850 9920
rect 4065 9911 4123 9917
rect 4065 9908 4077 9911
rect 3844 9880 4077 9908
rect 3844 9868 3850 9880
rect 4065 9877 4077 9880
rect 4111 9877 4123 9911
rect 4065 9871 4123 9877
rect 5077 9911 5135 9917
rect 5077 9877 5089 9911
rect 5123 9908 5135 9911
rect 7668 9908 7696 9948
rect 5123 9880 7696 9908
rect 5123 9877 5135 9880
rect 5077 9871 5135 9877
rect 7742 9868 7748 9920
rect 7800 9908 7806 9920
rect 8205 9911 8263 9917
rect 8205 9908 8217 9911
rect 7800 9880 8217 9908
rect 7800 9868 7806 9880
rect 8205 9877 8217 9880
rect 8251 9877 8263 9911
rect 9968 9908 9996 9948
rect 12066 9936 12072 9988
rect 12124 9976 12130 9988
rect 12250 9976 12256 9988
rect 12124 9948 12256 9976
rect 12124 9936 12130 9948
rect 12250 9936 12256 9948
rect 12308 9936 12314 9988
rect 13078 9908 13084 9920
rect 9968 9880 13084 9908
rect 8205 9871 8263 9877
rect 13078 9868 13084 9880
rect 13136 9868 13142 9920
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 5258 9704 5264 9716
rect 5092 9676 5264 9704
rect 4338 9596 4344 9648
rect 4396 9636 4402 9648
rect 5092 9636 5120 9676
rect 5258 9664 5264 9676
rect 5316 9704 5322 9716
rect 6362 9704 6368 9716
rect 5316 9676 6368 9704
rect 5316 9664 5322 9676
rect 6362 9664 6368 9676
rect 6420 9664 6426 9716
rect 12253 9707 12311 9713
rect 10520 9676 12204 9704
rect 6454 9636 6460 9648
rect 4396 9608 5120 9636
rect 6367 9608 6460 9636
rect 4396 9596 4402 9608
rect 2590 9568 2596 9580
rect 2551 9540 2596 9568
rect 2590 9528 2596 9540
rect 2648 9528 2654 9580
rect 2682 9528 2688 9580
rect 2740 9568 2746 9580
rect 3513 9571 3571 9577
rect 3513 9568 3525 9571
rect 2740 9540 3525 9568
rect 2740 9528 2746 9540
rect 3513 9537 3525 9540
rect 3559 9568 3571 9571
rect 4525 9571 4583 9577
rect 4525 9568 4537 9571
rect 3559 9540 4537 9568
rect 3559 9537 3571 9540
rect 3513 9531 3571 9537
rect 4525 9537 4537 9540
rect 4571 9568 4583 9571
rect 4982 9568 4988 9580
rect 4571 9540 4988 9568
rect 4571 9537 4583 9540
rect 4525 9531 4583 9537
rect 4982 9528 4988 9540
rect 5040 9528 5046 9580
rect 5092 9577 5120 9608
rect 6454 9596 6460 9608
rect 6512 9636 6518 9648
rect 8113 9639 8171 9645
rect 6512 9608 7512 9636
rect 6512 9596 6518 9608
rect 5077 9571 5135 9577
rect 5077 9537 5089 9571
rect 5123 9537 5135 9571
rect 7285 9571 7343 9577
rect 7285 9568 7297 9571
rect 5077 9531 5135 9537
rect 6104 9540 7297 9568
rect 3421 9503 3479 9509
rect 3421 9469 3433 9503
rect 3467 9500 3479 9503
rect 3694 9500 3700 9512
rect 3467 9472 3700 9500
rect 3467 9469 3479 9472
rect 3421 9463 3479 9469
rect 3694 9460 3700 9472
rect 3752 9500 3758 9512
rect 4890 9500 4896 9512
rect 3752 9472 4896 9500
rect 3752 9460 3758 9472
rect 4890 9460 4896 9472
rect 4948 9460 4954 9512
rect 6104 9500 6132 9540
rect 7285 9537 7297 9540
rect 7331 9537 7343 9571
rect 7285 9531 7343 9537
rect 7377 9571 7435 9577
rect 7377 9537 7389 9571
rect 7423 9537 7435 9571
rect 7484 9568 7512 9608
rect 8113 9605 8125 9639
rect 8159 9636 8171 9639
rect 8294 9636 8300 9648
rect 8159 9608 8300 9636
rect 8159 9605 8171 9608
rect 8113 9599 8171 9605
rect 8294 9596 8300 9608
rect 8352 9596 8358 9648
rect 10520 9636 10548 9676
rect 9140 9608 10548 9636
rect 10597 9639 10655 9645
rect 8202 9568 8208 9580
rect 7484 9540 8208 9568
rect 7377 9531 7435 9537
rect 7190 9500 7196 9512
rect 5184 9472 6132 9500
rect 7151 9472 7196 9500
rect 3050 9432 3056 9444
rect 1964 9404 3056 9432
rect 1964 9373 1992 9404
rect 3050 9392 3056 9404
rect 3108 9392 3114 9444
rect 4154 9392 4160 9444
rect 4212 9432 4218 9444
rect 5184 9432 5212 9472
rect 7190 9460 7196 9472
rect 7248 9460 7254 9512
rect 7392 9500 7420 9531
rect 8202 9528 8208 9540
rect 8260 9528 8266 9580
rect 8662 9568 8668 9580
rect 8623 9540 8668 9568
rect 8662 9528 8668 9540
rect 8720 9528 8726 9580
rect 9140 9577 9168 9608
rect 10597 9605 10609 9639
rect 10643 9636 10655 9639
rect 12176 9636 12204 9676
rect 12253 9673 12265 9707
rect 12299 9704 12311 9707
rect 12437 9707 12495 9713
rect 12437 9704 12449 9707
rect 12299 9676 12449 9704
rect 12299 9673 12311 9676
rect 12253 9667 12311 9673
rect 12437 9673 12449 9676
rect 12483 9673 12495 9707
rect 12437 9667 12495 9673
rect 10643 9608 12112 9636
rect 12176 9608 14504 9636
rect 10643 9605 10655 9608
rect 10597 9599 10655 9605
rect 9125 9571 9183 9577
rect 9125 9537 9137 9571
rect 9171 9537 9183 9571
rect 9125 9531 9183 9537
rect 9766 9528 9772 9580
rect 9824 9568 9830 9580
rect 10137 9571 10195 9577
rect 10137 9568 10149 9571
rect 9824 9540 10149 9568
rect 9824 9528 9830 9540
rect 10137 9537 10149 9540
rect 10183 9568 10195 9571
rect 10686 9568 10692 9580
rect 10183 9540 10692 9568
rect 10183 9537 10195 9540
rect 10137 9531 10195 9537
rect 10686 9528 10692 9540
rect 10744 9568 10750 9580
rect 11149 9571 11207 9577
rect 11149 9568 11161 9571
rect 10744 9540 11161 9568
rect 10744 9528 10750 9540
rect 11149 9537 11161 9540
rect 11195 9537 11207 9571
rect 11149 9531 11207 9537
rect 11238 9528 11244 9580
rect 11296 9568 11302 9580
rect 11296 9540 11652 9568
rect 11296 9528 11302 9540
rect 7466 9500 7472 9512
rect 7392 9472 7472 9500
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 8021 9503 8079 9509
rect 8021 9469 8033 9503
rect 8067 9500 8079 9503
rect 9398 9500 9404 9512
rect 8067 9472 9404 9500
rect 8067 9469 8079 9472
rect 8021 9463 8079 9469
rect 9398 9460 9404 9472
rect 9456 9460 9462 9512
rect 9582 9460 9588 9512
rect 9640 9500 9646 9512
rect 10045 9503 10103 9509
rect 10045 9500 10057 9503
rect 9640 9472 10057 9500
rect 9640 9460 9646 9472
rect 10045 9469 10057 9472
rect 10091 9469 10103 9503
rect 10045 9463 10103 9469
rect 10502 9460 10508 9512
rect 10560 9500 10566 9512
rect 10965 9503 11023 9509
rect 10965 9500 10977 9503
rect 10560 9472 10977 9500
rect 10560 9460 10566 9472
rect 10965 9469 10977 9472
rect 11011 9469 11023 9503
rect 10965 9463 11023 9469
rect 11072 9472 11560 9500
rect 4212 9404 5212 9432
rect 5344 9435 5402 9441
rect 4212 9392 4218 9404
rect 5344 9401 5356 9435
rect 5390 9432 5402 9435
rect 6454 9432 6460 9444
rect 5390 9404 6460 9432
rect 5390 9401 5402 9404
rect 5344 9395 5402 9401
rect 6454 9392 6460 9404
rect 6512 9392 6518 9444
rect 9490 9432 9496 9444
rect 6840 9404 9496 9432
rect 1949 9367 2007 9373
rect 1949 9333 1961 9367
rect 1995 9333 2007 9367
rect 2314 9364 2320 9376
rect 2275 9336 2320 9364
rect 1949 9327 2007 9333
rect 2314 9324 2320 9336
rect 2372 9324 2378 9376
rect 2406 9324 2412 9376
rect 2464 9364 2470 9376
rect 2958 9364 2964 9376
rect 2464 9336 2509 9364
rect 2919 9336 2964 9364
rect 2464 9324 2470 9336
rect 2958 9324 2964 9336
rect 3016 9324 3022 9376
rect 3326 9364 3332 9376
rect 3287 9336 3332 9364
rect 3326 9324 3332 9336
rect 3384 9324 3390 9376
rect 3510 9324 3516 9376
rect 3568 9364 3574 9376
rect 3973 9367 4031 9373
rect 3973 9364 3985 9367
rect 3568 9336 3985 9364
rect 3568 9324 3574 9336
rect 3973 9333 3985 9336
rect 4019 9333 4031 9367
rect 3973 9327 4031 9333
rect 4246 9324 4252 9376
rect 4304 9364 4310 9376
rect 4341 9367 4399 9373
rect 4341 9364 4353 9367
rect 4304 9336 4353 9364
rect 4304 9324 4310 9336
rect 4341 9333 4353 9336
rect 4387 9333 4399 9367
rect 4341 9327 4399 9333
rect 4433 9367 4491 9373
rect 4433 9333 4445 9367
rect 4479 9364 4491 9367
rect 6270 9364 6276 9376
rect 4479 9336 6276 9364
rect 4479 9333 4491 9336
rect 4433 9327 4491 9333
rect 6270 9324 6276 9336
rect 6328 9324 6334 9376
rect 6840 9373 6868 9404
rect 9490 9392 9496 9404
rect 9548 9392 9554 9444
rect 11072 9432 11100 9472
rect 9600 9404 11100 9432
rect 6825 9367 6883 9373
rect 6825 9333 6837 9367
rect 6871 9333 6883 9367
rect 6825 9327 6883 9333
rect 7006 9324 7012 9376
rect 7064 9364 7070 9376
rect 7190 9364 7196 9376
rect 7064 9336 7196 9364
rect 7064 9324 7070 9336
rect 7190 9324 7196 9336
rect 7248 9324 7254 9376
rect 7742 9324 7748 9376
rect 7800 9364 7806 9376
rect 7837 9367 7895 9373
rect 7837 9364 7849 9367
rect 7800 9336 7849 9364
rect 7800 9324 7806 9336
rect 7837 9333 7849 9336
rect 7883 9333 7895 9367
rect 7837 9327 7895 9333
rect 8294 9324 8300 9376
rect 8352 9364 8358 9376
rect 8481 9367 8539 9373
rect 8481 9364 8493 9367
rect 8352 9336 8493 9364
rect 8352 9324 8358 9336
rect 8481 9333 8493 9336
rect 8527 9333 8539 9367
rect 8481 9327 8539 9333
rect 8570 9324 8576 9376
rect 8628 9364 8634 9376
rect 9398 9364 9404 9376
rect 8628 9336 9404 9364
rect 8628 9324 8634 9336
rect 9398 9324 9404 9336
rect 9456 9324 9462 9376
rect 9600 9373 9628 9404
rect 9585 9367 9643 9373
rect 9585 9333 9597 9367
rect 9631 9333 9643 9367
rect 9585 9327 9643 9333
rect 9674 9324 9680 9376
rect 9732 9364 9738 9376
rect 9953 9367 10011 9373
rect 9953 9364 9965 9367
rect 9732 9336 9965 9364
rect 9732 9324 9738 9336
rect 9953 9333 9965 9336
rect 9999 9333 10011 9367
rect 9953 9327 10011 9333
rect 10042 9324 10048 9376
rect 10100 9364 10106 9376
rect 11057 9367 11115 9373
rect 11057 9364 11069 9367
rect 10100 9336 11069 9364
rect 10100 9324 10106 9336
rect 11057 9333 11069 9336
rect 11103 9333 11115 9367
rect 11422 9364 11428 9376
rect 11383 9336 11428 9364
rect 11057 9327 11115 9333
rect 11422 9324 11428 9336
rect 11480 9324 11486 9376
rect 11532 9364 11560 9472
rect 11624 9432 11652 9540
rect 11698 9528 11704 9580
rect 11756 9568 11762 9580
rect 11977 9571 12035 9577
rect 11977 9568 11989 9571
rect 11756 9540 11989 9568
rect 11756 9528 11762 9540
rect 11977 9537 11989 9540
rect 12023 9537 12035 9571
rect 12084 9568 12112 9608
rect 12986 9568 12992 9580
rect 12084 9540 12848 9568
rect 12947 9540 12992 9568
rect 11977 9531 12035 9537
rect 12820 9509 12848 9540
rect 12986 9528 12992 9540
rect 13044 9528 13050 9580
rect 13078 9528 13084 9580
rect 13136 9568 13142 9580
rect 13725 9571 13783 9577
rect 13725 9568 13737 9571
rect 13136 9540 13737 9568
rect 13136 9528 13142 9540
rect 13725 9537 13737 9540
rect 13771 9537 13783 9571
rect 13725 9531 13783 9537
rect 13817 9571 13875 9577
rect 13817 9537 13829 9571
rect 13863 9537 13875 9571
rect 13817 9531 13875 9537
rect 11793 9503 11851 9509
rect 11793 9469 11805 9503
rect 11839 9500 11851 9503
rect 12253 9503 12311 9509
rect 12253 9500 12265 9503
rect 11839 9472 12265 9500
rect 11839 9469 11851 9472
rect 11793 9463 11851 9469
rect 12253 9469 12265 9472
rect 12299 9469 12311 9503
rect 12253 9463 12311 9469
rect 12805 9503 12863 9509
rect 12805 9469 12817 9503
rect 12851 9469 12863 9503
rect 12805 9463 12863 9469
rect 13170 9460 13176 9512
rect 13228 9500 13234 9512
rect 13832 9500 13860 9531
rect 14476 9509 14504 9608
rect 14645 9571 14703 9577
rect 14645 9568 14657 9571
rect 14568 9540 14657 9568
rect 13228 9472 13860 9500
rect 14461 9503 14519 9509
rect 13228 9460 13234 9472
rect 14461 9469 14473 9503
rect 14507 9469 14519 9503
rect 14461 9463 14519 9469
rect 11885 9435 11943 9441
rect 11885 9432 11897 9435
rect 11624 9404 11897 9432
rect 11885 9401 11897 9404
rect 11931 9401 11943 9435
rect 13814 9432 13820 9444
rect 11885 9395 11943 9401
rect 13464 9404 13820 9432
rect 12897 9367 12955 9373
rect 12897 9364 12909 9367
rect 11532 9336 12909 9364
rect 12897 9333 12909 9336
rect 12943 9333 12955 9367
rect 12897 9327 12955 9333
rect 13265 9367 13323 9373
rect 13265 9333 13277 9367
rect 13311 9364 13323 9367
rect 13464 9364 13492 9404
rect 13814 9392 13820 9404
rect 13872 9392 13878 9444
rect 14274 9392 14280 9444
rect 14332 9432 14338 9444
rect 14568 9432 14596 9540
rect 14645 9537 14657 9540
rect 14691 9537 14703 9571
rect 14645 9531 14703 9537
rect 14332 9404 14596 9432
rect 14332 9392 14338 9404
rect 13630 9364 13636 9376
rect 13311 9336 13492 9364
rect 13591 9336 13636 9364
rect 13311 9333 13323 9336
rect 13265 9327 13323 9333
rect 13630 9324 13636 9336
rect 13688 9324 13694 9376
rect 14090 9364 14096 9376
rect 14051 9336 14096 9364
rect 14090 9324 14096 9336
rect 14148 9324 14154 9376
rect 14550 9364 14556 9376
rect 14511 9336 14556 9364
rect 14550 9324 14556 9336
rect 14608 9324 14614 9376
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 2222 9120 2228 9172
rect 2280 9160 2286 9172
rect 3697 9163 3755 9169
rect 3697 9160 3709 9163
rect 2280 9132 3709 9160
rect 2280 9120 2286 9132
rect 3697 9129 3709 9132
rect 3743 9160 3755 9163
rect 4338 9160 4344 9172
rect 3743 9132 4344 9160
rect 3743 9129 3755 9132
rect 3697 9123 3755 9129
rect 4338 9120 4344 9132
rect 4396 9120 4402 9172
rect 4433 9163 4491 9169
rect 4433 9129 4445 9163
rect 4479 9160 4491 9163
rect 6822 9160 6828 9172
rect 4479 9132 6828 9160
rect 4479 9129 4491 9132
rect 4433 9123 4491 9129
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 7466 9160 7472 9172
rect 7427 9132 7472 9160
rect 7466 9120 7472 9132
rect 7524 9120 7530 9172
rect 7837 9163 7895 9169
rect 7837 9160 7849 9163
rect 7576 9132 7849 9160
rect 1486 8984 1492 9036
rect 1544 9024 1550 9036
rect 2041 9027 2099 9033
rect 2041 9024 2053 9027
rect 1544 8996 2053 9024
rect 1544 8984 1550 8996
rect 2041 8993 2053 8996
rect 2087 9024 2099 9027
rect 2240 9024 2268 9120
rect 2308 9095 2366 9101
rect 2308 9061 2320 9095
rect 2354 9092 2366 9095
rect 2682 9092 2688 9104
rect 2354 9064 2688 9092
rect 2354 9061 2366 9064
rect 2308 9055 2366 9061
rect 2682 9052 2688 9064
rect 2740 9052 2746 9104
rect 3050 9052 3056 9104
rect 3108 9092 3114 9104
rect 3418 9092 3424 9104
rect 3108 9064 3424 9092
rect 3108 9052 3114 9064
rect 3418 9052 3424 9064
rect 3476 9052 3482 9104
rect 2087 8996 2268 9024
rect 3881 9027 3939 9033
rect 2087 8993 2099 8996
rect 2041 8987 2099 8993
rect 3881 8993 3893 9027
rect 3927 8993 3939 9027
rect 3881 8987 3939 8993
rect 3896 8888 3924 8987
rect 4062 8984 4068 9036
rect 4120 9024 4126 9036
rect 4801 9027 4859 9033
rect 4801 9024 4813 9027
rect 4120 8996 4813 9024
rect 4120 8984 4126 8996
rect 4801 8993 4813 8996
rect 4847 8993 4859 9027
rect 4801 8987 4859 8993
rect 5626 8984 5632 9036
rect 5684 9024 5690 9036
rect 5813 9027 5871 9033
rect 5813 9024 5825 9027
rect 5684 8996 5825 9024
rect 5684 8984 5690 8996
rect 5813 8993 5825 8996
rect 5859 8993 5871 9027
rect 5813 8987 5871 8993
rect 5905 9027 5963 9033
rect 5905 8993 5917 9027
rect 5951 9024 5963 9027
rect 6730 9024 6736 9036
rect 5951 8996 6736 9024
rect 5951 8993 5963 8996
rect 5905 8987 5963 8993
rect 6730 8984 6736 8996
rect 6788 8984 6794 9036
rect 6825 9027 6883 9033
rect 6825 8993 6837 9027
rect 6871 9024 6883 9027
rect 7466 9024 7472 9036
rect 6871 8996 7472 9024
rect 6871 8993 6883 8996
rect 6825 8987 6883 8993
rect 7466 8984 7472 8996
rect 7524 8984 7530 9036
rect 7576 9024 7604 9132
rect 7837 9129 7849 9132
rect 7883 9129 7895 9163
rect 8849 9163 8907 9169
rect 8849 9160 8861 9163
rect 7837 9123 7895 9129
rect 8036 9132 8861 9160
rect 7650 9024 7656 9036
rect 7576 8996 7656 9024
rect 7650 8984 7656 8996
rect 7708 8984 7714 9036
rect 7926 9024 7932 9036
rect 7887 8996 7932 9024
rect 7926 8984 7932 8996
rect 7984 8984 7990 9036
rect 8036 9024 8064 9132
rect 8849 9129 8861 9132
rect 8895 9129 8907 9163
rect 8849 9123 8907 9129
rect 9490 9120 9496 9172
rect 9548 9160 9554 9172
rect 11609 9163 11667 9169
rect 11609 9160 11621 9163
rect 9548 9132 11621 9160
rect 9548 9120 9554 9132
rect 11609 9129 11621 9132
rect 11655 9129 11667 9163
rect 11609 9123 11667 9129
rect 11698 9120 11704 9172
rect 11756 9160 11762 9172
rect 12713 9163 12771 9169
rect 11756 9132 11801 9160
rect 11756 9120 11762 9132
rect 12713 9129 12725 9163
rect 12759 9160 12771 9163
rect 14093 9163 14151 9169
rect 14093 9160 14105 9163
rect 12759 9132 14105 9160
rect 12759 9129 12771 9132
rect 12713 9123 12771 9129
rect 14093 9129 14105 9132
rect 14139 9129 14151 9163
rect 14093 9123 14151 9129
rect 8386 9052 8392 9104
rect 8444 9092 8450 9104
rect 11514 9092 11520 9104
rect 8444 9064 11520 9092
rect 8444 9052 8450 9064
rect 11514 9052 11520 9064
rect 11572 9052 11578 9104
rect 12161 9095 12219 9101
rect 12161 9061 12173 9095
rect 12207 9092 12219 9095
rect 12250 9092 12256 9104
rect 12207 9064 12256 9092
rect 12207 9061 12219 9064
rect 12161 9055 12219 9061
rect 12250 9052 12256 9064
rect 12308 9052 12314 9104
rect 13173 9095 13231 9101
rect 13173 9092 13185 9095
rect 12452 9064 13185 9092
rect 8110 9024 8116 9036
rect 8036 8996 8116 9024
rect 8110 8984 8116 8996
rect 8168 8984 8174 9036
rect 8202 8984 8208 9036
rect 8260 9024 8266 9036
rect 8260 8996 9076 9024
rect 8260 8984 8266 8996
rect 4890 8916 4896 8968
rect 4948 8956 4954 8968
rect 5077 8959 5135 8965
rect 4948 8928 4993 8956
rect 4948 8916 4954 8928
rect 5077 8925 5089 8959
rect 5123 8956 5135 8959
rect 5166 8956 5172 8968
rect 5123 8928 5172 8956
rect 5123 8925 5135 8928
rect 5077 8919 5135 8925
rect 5166 8916 5172 8928
rect 5224 8916 5230 8968
rect 5994 8956 6000 8968
rect 5955 8928 6000 8956
rect 5994 8916 6000 8928
rect 6052 8916 6058 8968
rect 6914 8956 6920 8968
rect 6875 8928 6920 8956
rect 6914 8916 6920 8928
rect 6972 8916 6978 8968
rect 9048 8965 9076 8996
rect 9306 8984 9312 9036
rect 9364 9024 9370 9036
rect 10042 9024 10048 9036
rect 9364 8996 10048 9024
rect 9364 8984 9370 8996
rect 10042 8984 10048 8996
rect 10100 8984 10106 9036
rect 11057 9027 11115 9033
rect 11057 8993 11069 9027
rect 11103 9024 11115 9027
rect 11606 9024 11612 9036
rect 11103 8996 11612 9024
rect 11103 8993 11115 8996
rect 11057 8987 11115 8993
rect 11606 8984 11612 8996
rect 11664 8984 11670 9036
rect 11974 8984 11980 9036
rect 12032 9024 12038 9036
rect 12069 9027 12127 9033
rect 12069 9024 12081 9027
rect 12032 8996 12081 9024
rect 12032 8984 12038 8996
rect 12069 8993 12081 8996
rect 12115 8993 12127 9027
rect 12069 8987 12127 8993
rect 12342 8984 12348 9036
rect 12400 9024 12406 9036
rect 12452 9024 12480 9064
rect 13173 9061 13185 9064
rect 13219 9061 13231 9095
rect 13630 9092 13636 9104
rect 13173 9055 13231 9061
rect 13280 9064 13636 9092
rect 13078 9024 13084 9036
rect 12400 8996 12480 9024
rect 13039 8996 13084 9024
rect 12400 8984 12406 8996
rect 13078 8984 13084 8996
rect 13136 8984 13142 9036
rect 7101 8959 7159 8965
rect 7101 8925 7113 8959
rect 7147 8956 7159 8959
rect 7285 8959 7343 8965
rect 7285 8956 7297 8959
rect 7147 8928 7297 8956
rect 7147 8925 7159 8928
rect 7101 8919 7159 8925
rect 7285 8925 7297 8928
rect 7331 8956 7343 8959
rect 8021 8959 8079 8965
rect 8021 8956 8033 8959
rect 7331 8928 8033 8956
rect 7331 8925 7343 8928
rect 7285 8919 7343 8925
rect 8021 8925 8033 8928
rect 8067 8925 8079 8959
rect 8021 8919 8079 8925
rect 8941 8959 8999 8965
rect 8941 8925 8953 8959
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 9033 8959 9091 8965
rect 9033 8925 9045 8959
rect 9079 8925 9091 8959
rect 9033 8919 9091 8925
rect 5350 8888 5356 8900
rect 3896 8860 5356 8888
rect 5350 8848 5356 8860
rect 5408 8848 5414 8900
rect 6457 8891 6515 8897
rect 6457 8857 6469 8891
rect 6503 8888 6515 8891
rect 8956 8888 8984 8919
rect 9674 8916 9680 8968
rect 9732 8956 9738 8968
rect 10137 8959 10195 8965
rect 10137 8956 10149 8959
rect 9732 8928 10149 8956
rect 9732 8916 9738 8928
rect 10137 8925 10149 8928
rect 10183 8925 10195 8959
rect 10137 8919 10195 8925
rect 10226 8916 10232 8968
rect 10284 8956 10290 8968
rect 11149 8959 11207 8965
rect 10284 8928 10329 8956
rect 10284 8916 10290 8928
rect 11149 8925 11161 8959
rect 11195 8925 11207 8959
rect 11149 8919 11207 8925
rect 6503 8860 8984 8888
rect 6503 8857 6515 8860
rect 6457 8851 6515 8857
rect 10778 8848 10784 8900
rect 10836 8888 10842 8900
rect 11164 8888 11192 8919
rect 11238 8916 11244 8968
rect 11296 8956 11302 8968
rect 12253 8959 12311 8965
rect 12253 8956 12265 8959
rect 11296 8928 12265 8956
rect 11296 8916 11302 8928
rect 12253 8925 12265 8928
rect 12299 8925 12311 8959
rect 13280 8956 13308 9064
rect 13630 9052 13636 9064
rect 13688 9052 13694 9104
rect 13814 9052 13820 9104
rect 13872 9092 13878 9104
rect 15102 9092 15108 9104
rect 13872 9064 15108 9092
rect 13872 9052 13878 9064
rect 15102 9052 15108 9064
rect 15160 9052 15166 9104
rect 13538 8984 13544 9036
rect 13596 9024 13602 9036
rect 14185 9027 14243 9033
rect 14185 9024 14197 9027
rect 13596 8996 14197 9024
rect 13596 8984 13602 8996
rect 14185 8993 14197 8996
rect 14231 8993 14243 9027
rect 14185 8987 14243 8993
rect 12253 8919 12311 8925
rect 12360 8928 13308 8956
rect 13357 8959 13415 8965
rect 10836 8860 11192 8888
rect 10836 8848 10842 8860
rect 3418 8820 3424 8832
rect 3379 8792 3424 8820
rect 3418 8780 3424 8792
rect 3476 8780 3482 8832
rect 5442 8820 5448 8832
rect 5403 8792 5448 8820
rect 5442 8780 5448 8792
rect 5500 8780 5506 8832
rect 6362 8780 6368 8832
rect 6420 8820 6426 8832
rect 7285 8823 7343 8829
rect 7285 8820 7297 8823
rect 6420 8792 7297 8820
rect 6420 8780 6426 8792
rect 7285 8789 7297 8792
rect 7331 8789 7343 8823
rect 7285 8783 7343 8789
rect 7374 8780 7380 8832
rect 7432 8820 7438 8832
rect 8481 8823 8539 8829
rect 8481 8820 8493 8823
rect 7432 8792 8493 8820
rect 7432 8780 7438 8792
rect 8481 8789 8493 8792
rect 8527 8789 8539 8823
rect 8481 8783 8539 8789
rect 8754 8780 8760 8832
rect 8812 8820 8818 8832
rect 9582 8820 9588 8832
rect 8812 8792 9588 8820
rect 8812 8780 8818 8792
rect 9582 8780 9588 8792
rect 9640 8780 9646 8832
rect 9677 8823 9735 8829
rect 9677 8789 9689 8823
rect 9723 8820 9735 8823
rect 10042 8820 10048 8832
rect 9723 8792 10048 8820
rect 9723 8789 9735 8792
rect 9677 8783 9735 8789
rect 10042 8780 10048 8792
rect 10100 8780 10106 8832
rect 10686 8820 10692 8832
rect 10647 8792 10692 8820
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 11164 8820 11192 8860
rect 11609 8891 11667 8897
rect 11609 8857 11621 8891
rect 11655 8888 11667 8891
rect 12360 8888 12388 8928
rect 13357 8925 13369 8959
rect 13403 8925 13415 8959
rect 14274 8956 14280 8968
rect 14235 8928 14280 8956
rect 13357 8919 13415 8925
rect 11655 8860 12388 8888
rect 11655 8857 11667 8860
rect 11609 8851 11667 8857
rect 13262 8848 13268 8900
rect 13320 8888 13326 8900
rect 13372 8888 13400 8919
rect 14274 8916 14280 8928
rect 14332 8916 14338 8968
rect 15286 8888 15292 8900
rect 13320 8860 13400 8888
rect 13464 8860 15292 8888
rect 13320 8848 13326 8860
rect 13464 8820 13492 8860
rect 15286 8848 15292 8860
rect 15344 8848 15350 8900
rect 11164 8792 13492 8820
rect 13725 8823 13783 8829
rect 13725 8789 13737 8823
rect 13771 8820 13783 8823
rect 14918 8820 14924 8832
rect 13771 8792 14924 8820
rect 13771 8789 13783 8792
rect 13725 8783 13783 8789
rect 14918 8780 14924 8792
rect 14976 8780 14982 8832
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 2406 8576 2412 8628
rect 2464 8616 2470 8628
rect 3053 8619 3111 8625
rect 3053 8616 3065 8619
rect 2464 8588 3065 8616
rect 2464 8576 2470 8588
rect 3053 8585 3065 8588
rect 3099 8585 3111 8619
rect 4062 8616 4068 8628
rect 4023 8588 4068 8616
rect 3053 8579 3111 8585
rect 4062 8576 4068 8588
rect 4120 8576 4126 8628
rect 6454 8616 6460 8628
rect 5092 8588 6316 8616
rect 6415 8588 6460 8616
rect 2590 8508 2596 8560
rect 2648 8548 2654 8560
rect 2777 8551 2835 8557
rect 2777 8548 2789 8551
rect 2648 8520 2789 8548
rect 2648 8508 2654 8520
rect 2777 8517 2789 8520
rect 2823 8517 2835 8551
rect 2777 8511 2835 8517
rect 3970 8508 3976 8560
rect 4028 8548 4034 8560
rect 5092 8548 5120 8588
rect 4028 8520 5120 8548
rect 6288 8548 6316 8588
rect 6454 8576 6460 8588
rect 6512 8576 6518 8628
rect 9674 8616 9680 8628
rect 7024 8588 9680 8616
rect 7024 8548 7052 8588
rect 9674 8576 9680 8588
rect 9732 8576 9738 8628
rect 9950 8576 9956 8628
rect 10008 8616 10014 8628
rect 10045 8619 10103 8625
rect 10045 8616 10057 8619
rect 10008 8588 10057 8616
rect 10008 8576 10014 8588
rect 10045 8585 10057 8588
rect 10091 8616 10103 8619
rect 13265 8619 13323 8625
rect 13265 8616 13277 8619
rect 10091 8588 13277 8616
rect 10091 8585 10103 8588
rect 10045 8579 10103 8585
rect 13265 8585 13277 8588
rect 13311 8585 13323 8619
rect 13265 8579 13323 8585
rect 13449 8619 13507 8625
rect 13449 8585 13461 8619
rect 13495 8616 13507 8619
rect 14550 8616 14556 8628
rect 13495 8588 14556 8616
rect 13495 8585 13507 8588
rect 13449 8579 13507 8585
rect 14550 8576 14556 8588
rect 14608 8576 14614 8628
rect 6288 8520 7052 8548
rect 8389 8551 8447 8557
rect 4028 8508 4034 8520
rect 8389 8517 8401 8551
rect 8435 8517 8447 8551
rect 10318 8548 10324 8560
rect 10279 8520 10324 8548
rect 8389 8511 8447 8517
rect 3510 8480 3516 8492
rect 3471 8452 3516 8480
rect 3510 8440 3516 8452
rect 3568 8440 3574 8492
rect 3605 8483 3663 8489
rect 3605 8449 3617 8483
rect 3651 8449 3663 8483
rect 3605 8443 3663 8449
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 1486 8412 1492 8424
rect 1443 8384 1492 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 1486 8372 1492 8384
rect 1544 8372 1550 8424
rect 1664 8415 1722 8421
rect 1664 8381 1676 8415
rect 1710 8412 1722 8415
rect 2682 8412 2688 8424
rect 1710 8384 2688 8412
rect 1710 8381 1722 8384
rect 1664 8375 1722 8381
rect 2682 8372 2688 8384
rect 2740 8412 2746 8424
rect 3418 8412 3424 8424
rect 2740 8384 3424 8412
rect 2740 8372 2746 8384
rect 3418 8372 3424 8384
rect 3476 8412 3482 8424
rect 3620 8412 3648 8443
rect 4154 8440 4160 8492
rect 4212 8480 4218 8492
rect 4525 8483 4583 8489
rect 4525 8480 4537 8483
rect 4212 8452 4537 8480
rect 4212 8440 4218 8452
rect 4525 8449 4537 8452
rect 4571 8449 4583 8483
rect 4525 8443 4583 8449
rect 4709 8483 4767 8489
rect 4709 8449 4721 8483
rect 4755 8480 4767 8483
rect 4798 8480 4804 8492
rect 4755 8452 4804 8480
rect 4755 8449 4767 8452
rect 4709 8443 4767 8449
rect 4798 8440 4804 8452
rect 4856 8440 4862 8492
rect 8404 8480 8432 8511
rect 10318 8508 10324 8520
rect 10376 8508 10382 8560
rect 12069 8551 12127 8557
rect 12069 8517 12081 8551
rect 12115 8517 12127 8551
rect 12069 8511 12127 8517
rect 12437 8551 12495 8557
rect 12437 8517 12449 8551
rect 12483 8548 12495 8551
rect 13814 8548 13820 8560
rect 12483 8520 13820 8548
rect 12483 8517 12495 8520
rect 12437 8511 12495 8517
rect 8404 8452 8800 8480
rect 3476 8384 3648 8412
rect 5077 8415 5135 8421
rect 3476 8372 3482 8384
rect 5077 8381 5089 8415
rect 5123 8412 5135 8415
rect 7009 8415 7067 8421
rect 5123 8384 5304 8412
rect 5123 8381 5135 8384
rect 5077 8375 5135 8381
rect 3786 8344 3792 8356
rect 3436 8316 3792 8344
rect 3436 8285 3464 8316
rect 3786 8304 3792 8316
rect 3844 8304 3850 8356
rect 5276 8288 5304 8384
rect 7009 8381 7021 8415
rect 7055 8412 7067 8415
rect 8662 8412 8668 8424
rect 7055 8384 8668 8412
rect 7055 8381 7067 8384
rect 7009 8375 7067 8381
rect 8662 8372 8668 8384
rect 8720 8372 8726 8424
rect 8772 8412 8800 8452
rect 9766 8440 9772 8492
rect 9824 8480 9830 8492
rect 10594 8480 10600 8492
rect 9824 8452 10600 8480
rect 9824 8440 9830 8452
rect 10594 8440 10600 8452
rect 10652 8480 10658 8492
rect 10689 8483 10747 8489
rect 10689 8480 10701 8483
rect 10652 8452 10701 8480
rect 10652 8440 10658 8452
rect 10689 8449 10701 8452
rect 10735 8449 10747 8483
rect 10689 8443 10747 8449
rect 11974 8440 11980 8492
rect 12032 8480 12038 8492
rect 12084 8480 12112 8511
rect 13814 8508 13820 8520
rect 13872 8508 13878 8560
rect 14461 8551 14519 8557
rect 14461 8517 14473 8551
rect 14507 8548 14519 8551
rect 18506 8548 18512 8560
rect 14507 8520 18512 8548
rect 14507 8517 14519 8520
rect 14461 8511 14519 8517
rect 18506 8508 18512 8520
rect 18564 8508 18570 8560
rect 12989 8483 13047 8489
rect 12989 8480 13001 8483
rect 12032 8452 13001 8480
rect 12032 8440 12038 8452
rect 12989 8449 13001 8452
rect 13035 8449 13047 8483
rect 12989 8443 13047 8449
rect 13262 8440 13268 8492
rect 13320 8480 13326 8492
rect 14001 8483 14059 8489
rect 14001 8480 14013 8483
rect 13320 8452 14013 8480
rect 13320 8440 13326 8452
rect 14001 8449 14013 8452
rect 14047 8449 14059 8483
rect 14918 8480 14924 8492
rect 14879 8452 14924 8480
rect 14001 8443 14059 8449
rect 14918 8440 14924 8452
rect 14976 8440 14982 8492
rect 15013 8483 15071 8489
rect 15013 8449 15025 8483
rect 15059 8449 15071 8483
rect 15013 8443 15071 8449
rect 8932 8415 8990 8421
rect 8932 8412 8944 8415
rect 8772 8384 8944 8412
rect 8932 8381 8944 8384
rect 8978 8412 8990 8415
rect 9674 8412 9680 8424
rect 8978 8384 9680 8412
rect 8978 8381 8990 8384
rect 8932 8375 8990 8381
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 10505 8415 10563 8421
rect 10505 8412 10517 8415
rect 9968 8384 10517 8412
rect 5344 8347 5402 8353
rect 5344 8313 5356 8347
rect 5390 8344 5402 8347
rect 5718 8344 5724 8356
rect 5390 8316 5724 8344
rect 5390 8313 5402 8316
rect 5344 8307 5402 8313
rect 5718 8304 5724 8316
rect 5776 8304 5782 8356
rect 7282 8353 7288 8356
rect 7276 8307 7288 8353
rect 7340 8344 7346 8356
rect 7340 8316 7376 8344
rect 7282 8304 7288 8307
rect 7340 8304 7346 8316
rect 7742 8304 7748 8356
rect 7800 8344 7806 8356
rect 9968 8344 9996 8384
rect 10505 8381 10517 8384
rect 10551 8381 10563 8415
rect 12897 8415 12955 8421
rect 12897 8412 12909 8415
rect 10505 8375 10563 8381
rect 10704 8384 12909 8412
rect 10704 8356 10732 8384
rect 12897 8381 12909 8384
rect 12943 8381 12955 8415
rect 12897 8375 12955 8381
rect 13817 8415 13875 8421
rect 13817 8381 13829 8415
rect 13863 8412 13875 8415
rect 13906 8412 13912 8424
rect 13863 8384 13912 8412
rect 13863 8381 13875 8384
rect 13817 8375 13875 8381
rect 13906 8372 13912 8384
rect 13964 8372 13970 8424
rect 14090 8372 14096 8424
rect 14148 8412 14154 8424
rect 14829 8415 14887 8421
rect 14829 8412 14841 8415
rect 14148 8384 14841 8412
rect 14148 8372 14154 8384
rect 14829 8381 14841 8384
rect 14875 8381 14887 8415
rect 14829 8375 14887 8381
rect 7800 8316 9996 8344
rect 7800 8304 7806 8316
rect 10686 8304 10692 8356
rect 10744 8304 10750 8356
rect 10956 8347 11014 8353
rect 10956 8313 10968 8347
rect 11002 8313 11014 8347
rect 10956 8307 11014 8313
rect 3421 8279 3479 8285
rect 3421 8245 3433 8279
rect 3467 8245 3479 8279
rect 3421 8239 3479 8245
rect 4154 8236 4160 8288
rect 4212 8276 4218 8288
rect 4433 8279 4491 8285
rect 4433 8276 4445 8279
rect 4212 8248 4445 8276
rect 4212 8236 4218 8248
rect 4433 8245 4445 8248
rect 4479 8245 4491 8279
rect 4433 8239 4491 8245
rect 5258 8236 5264 8288
rect 5316 8236 5322 8288
rect 8938 8236 8944 8288
rect 8996 8276 9002 8288
rect 9398 8276 9404 8288
rect 8996 8248 9404 8276
rect 8996 8236 9002 8248
rect 9398 8236 9404 8248
rect 9456 8236 9462 8288
rect 10980 8276 11008 8307
rect 11698 8304 11704 8356
rect 11756 8344 11762 8356
rect 12805 8347 12863 8353
rect 12805 8344 12817 8347
rect 11756 8316 12817 8344
rect 11756 8304 11762 8316
rect 12805 8313 12817 8316
rect 12851 8313 12863 8347
rect 12805 8307 12863 8313
rect 13265 8347 13323 8353
rect 13265 8313 13277 8347
rect 13311 8344 13323 8347
rect 15028 8344 15056 8443
rect 13311 8316 15056 8344
rect 13311 8313 13323 8316
rect 13265 8307 13323 8313
rect 11054 8276 11060 8288
rect 10980 8248 11060 8276
rect 11054 8236 11060 8248
rect 11112 8236 11118 8288
rect 11882 8236 11888 8288
rect 11940 8276 11946 8288
rect 12526 8276 12532 8288
rect 11940 8248 12532 8276
rect 11940 8236 11946 8248
rect 12526 8236 12532 8248
rect 12584 8236 12590 8288
rect 13906 8276 13912 8288
rect 13867 8248 13912 8276
rect 13906 8236 13912 8248
rect 13964 8236 13970 8288
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 2133 8075 2191 8081
rect 2133 8041 2145 8075
rect 2179 8072 2191 8075
rect 2314 8072 2320 8084
rect 2179 8044 2320 8072
rect 2179 8041 2191 8044
rect 2133 8035 2191 8041
rect 2314 8032 2320 8044
rect 2372 8032 2378 8084
rect 2501 8075 2559 8081
rect 2501 8041 2513 8075
rect 2547 8072 2559 8075
rect 2958 8072 2964 8084
rect 2547 8044 2964 8072
rect 2547 8041 2559 8044
rect 2501 8035 2559 8041
rect 2958 8032 2964 8044
rect 3016 8032 3022 8084
rect 3145 8075 3203 8081
rect 3145 8041 3157 8075
rect 3191 8072 3203 8075
rect 3326 8072 3332 8084
rect 3191 8044 3332 8072
rect 3191 8041 3203 8044
rect 3145 8035 3203 8041
rect 3326 8032 3332 8044
rect 3384 8032 3390 8084
rect 4249 8075 4307 8081
rect 4249 8041 4261 8075
rect 4295 8072 4307 8075
rect 4890 8072 4896 8084
rect 4295 8044 4896 8072
rect 4295 8041 4307 8044
rect 4249 8035 4307 8041
rect 4890 8032 4896 8044
rect 4948 8032 4954 8084
rect 6365 8075 6423 8081
rect 6365 8041 6377 8075
rect 6411 8072 6423 8075
rect 6546 8072 6552 8084
rect 6411 8044 6552 8072
rect 6411 8041 6423 8044
rect 6365 8035 6423 8041
rect 6546 8032 6552 8044
rect 6604 8032 6610 8084
rect 6914 8032 6920 8084
rect 6972 8072 6978 8084
rect 7377 8075 7435 8081
rect 7377 8072 7389 8075
rect 6972 8044 7389 8072
rect 6972 8032 6978 8044
rect 7377 8041 7389 8044
rect 7423 8041 7435 8075
rect 7377 8035 7435 8041
rect 8573 8075 8631 8081
rect 8573 8041 8585 8075
rect 8619 8072 8631 8075
rect 13081 8075 13139 8081
rect 8619 8044 13032 8072
rect 8619 8041 8631 8044
rect 8573 8035 8631 8041
rect 4062 7964 4068 8016
rect 4120 8004 4126 8016
rect 4617 8007 4675 8013
rect 4617 8004 4629 8007
rect 4120 7976 4629 8004
rect 4120 7964 4126 7976
rect 4617 7973 4629 7976
rect 4663 8004 4675 8007
rect 5074 8004 5080 8016
rect 4663 7976 5080 8004
rect 4663 7973 4675 7976
rect 4617 7967 4675 7973
rect 5074 7964 5080 7976
rect 5132 7964 5138 8016
rect 5813 8007 5871 8013
rect 5813 7973 5825 8007
rect 5859 8004 5871 8007
rect 6270 8004 6276 8016
rect 5859 7976 6276 8004
rect 5859 7973 5871 7976
rect 5813 7967 5871 7973
rect 6270 7964 6276 7976
rect 6328 7964 6334 8016
rect 6733 8007 6791 8013
rect 6733 7973 6745 8007
rect 6779 8004 6791 8007
rect 8478 8004 8484 8016
rect 6779 7976 8484 8004
rect 6779 7973 6791 7976
rect 6733 7967 6791 7973
rect 8478 7964 8484 7976
rect 8536 7964 8542 8016
rect 9950 8013 9956 8016
rect 9944 7967 9956 8013
rect 10008 8004 10014 8016
rect 11974 8013 11980 8016
rect 11968 8004 11980 8013
rect 10008 7976 10044 8004
rect 11935 7976 11980 8004
rect 9950 7964 9956 7967
rect 10008 7964 10014 7976
rect 11968 7967 11980 7976
rect 11974 7964 11980 7967
rect 12032 7964 12038 8016
rect 3970 7896 3976 7948
rect 4028 7936 4034 7948
rect 5721 7939 5779 7945
rect 5721 7936 5733 7939
rect 4028 7908 5733 7936
rect 4028 7896 4034 7908
rect 5721 7905 5733 7908
rect 5767 7905 5779 7939
rect 5721 7899 5779 7905
rect 5994 7896 6000 7948
rect 6052 7936 6058 7948
rect 7745 7939 7803 7945
rect 7745 7936 7757 7939
rect 6052 7908 6960 7936
rect 6052 7896 6058 7908
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7837 2651 7871
rect 2593 7831 2651 7837
rect 2608 7800 2636 7831
rect 2682 7828 2688 7880
rect 2740 7868 2746 7880
rect 4706 7868 4712 7880
rect 2740 7840 2785 7868
rect 4667 7840 4712 7868
rect 2740 7828 2746 7840
rect 4706 7828 4712 7840
rect 4764 7828 4770 7880
rect 4890 7868 4896 7880
rect 4803 7840 4896 7868
rect 4890 7828 4896 7840
rect 4948 7868 4954 7880
rect 5905 7871 5963 7877
rect 4948 7840 5580 7868
rect 4948 7828 4954 7840
rect 5442 7800 5448 7812
rect 2608 7772 5448 7800
rect 5442 7760 5448 7772
rect 5500 7760 5506 7812
rect 5552 7800 5580 7840
rect 5905 7837 5917 7871
rect 5951 7868 5963 7871
rect 6270 7868 6276 7880
rect 5951 7840 6276 7868
rect 5951 7837 5963 7840
rect 5905 7831 5963 7837
rect 5920 7800 5948 7831
rect 6270 7828 6276 7840
rect 6328 7828 6334 7880
rect 6932 7877 6960 7908
rect 7024 7908 7757 7936
rect 7024 7880 7052 7908
rect 7745 7905 7757 7908
rect 7791 7905 7803 7939
rect 8386 7936 8392 7948
rect 7745 7899 7803 7905
rect 7852 7908 8392 7936
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7837 6883 7871
rect 6825 7831 6883 7837
rect 6917 7871 6975 7877
rect 6917 7837 6929 7871
rect 6963 7837 6975 7871
rect 6917 7831 6975 7837
rect 5552 7772 5948 7800
rect 6840 7800 6868 7831
rect 7006 7828 7012 7880
rect 7064 7828 7070 7880
rect 7098 7828 7104 7880
rect 7156 7868 7162 7880
rect 7852 7877 7880 7908
rect 8386 7896 8392 7908
rect 8444 7896 8450 7948
rect 8570 7896 8576 7948
rect 8628 7936 8634 7948
rect 8941 7939 8999 7945
rect 8941 7936 8953 7939
rect 8628 7908 8953 7936
rect 8628 7896 8634 7908
rect 8941 7905 8953 7908
rect 8987 7905 8999 7939
rect 8941 7899 8999 7905
rect 9674 7896 9680 7948
rect 9732 7936 9738 7948
rect 13004 7936 13032 8044
rect 13081 8041 13093 8075
rect 13127 8041 13139 8075
rect 13081 8035 13139 8041
rect 13096 8004 13124 8035
rect 13630 8013 13636 8016
rect 13602 8007 13636 8013
rect 13602 8004 13614 8007
rect 13096 7976 13614 8004
rect 13602 7973 13614 7976
rect 13688 8004 13694 8016
rect 13688 7976 13750 8004
rect 13602 7967 13636 7973
rect 13630 7964 13636 7967
rect 13688 7964 13694 7976
rect 17402 7936 17408 7948
rect 9732 7908 9777 7936
rect 13004 7908 17408 7936
rect 9732 7896 9738 7908
rect 17402 7896 17408 7908
rect 17460 7896 17466 7948
rect 7837 7871 7895 7877
rect 7837 7868 7849 7871
rect 7156 7840 7849 7868
rect 7156 7828 7162 7840
rect 7837 7837 7849 7840
rect 7883 7837 7895 7871
rect 8018 7868 8024 7880
rect 7979 7840 8024 7868
rect 7837 7831 7895 7837
rect 8018 7828 8024 7840
rect 8076 7828 8082 7880
rect 8662 7828 8668 7880
rect 8720 7868 8726 7880
rect 9033 7871 9091 7877
rect 9033 7868 9045 7871
rect 8720 7840 9045 7868
rect 8720 7828 8726 7840
rect 9033 7837 9045 7840
rect 9079 7837 9091 7871
rect 9214 7868 9220 7880
rect 9175 7840 9220 7868
rect 9033 7831 9091 7837
rect 9214 7828 9220 7840
rect 9272 7828 9278 7880
rect 11606 7828 11612 7880
rect 11664 7868 11670 7880
rect 11701 7871 11759 7877
rect 11701 7868 11713 7871
rect 11664 7840 11713 7868
rect 11664 7828 11670 7840
rect 11701 7837 11713 7840
rect 11747 7837 11759 7871
rect 13354 7868 13360 7880
rect 13315 7840 13360 7868
rect 11701 7831 11759 7837
rect 13354 7828 13360 7840
rect 13412 7828 13418 7880
rect 8386 7800 8392 7812
rect 6840 7772 8392 7800
rect 8386 7760 8392 7772
rect 8444 7760 8450 7812
rect 5353 7735 5411 7741
rect 5353 7701 5365 7735
rect 5399 7732 5411 7735
rect 7190 7732 7196 7744
rect 5399 7704 7196 7732
rect 5399 7701 5411 7704
rect 5353 7695 5411 7701
rect 7190 7692 7196 7704
rect 7248 7692 7254 7744
rect 9582 7692 9588 7744
rect 9640 7732 9646 7744
rect 11057 7735 11115 7741
rect 11057 7732 11069 7735
rect 9640 7704 11069 7732
rect 9640 7692 9646 7704
rect 11057 7701 11069 7704
rect 11103 7732 11115 7735
rect 13538 7732 13544 7744
rect 11103 7704 13544 7732
rect 11103 7701 11115 7704
rect 11057 7695 11115 7701
rect 13538 7692 13544 7704
rect 13596 7692 13602 7744
rect 13998 7692 14004 7744
rect 14056 7732 14062 7744
rect 14737 7735 14795 7741
rect 14737 7732 14749 7735
rect 14056 7704 14749 7732
rect 14056 7692 14062 7704
rect 14737 7701 14749 7704
rect 14783 7701 14795 7735
rect 14737 7695 14795 7701
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 5258 7528 5264 7540
rect 4632 7500 5264 7528
rect 1854 7352 1860 7404
rect 1912 7392 1918 7404
rect 2501 7395 2559 7401
rect 2501 7392 2513 7395
rect 1912 7364 2513 7392
rect 1912 7352 1918 7364
rect 2501 7361 2513 7364
rect 2547 7361 2559 7395
rect 2501 7355 2559 7361
rect 2866 7352 2872 7404
rect 2924 7392 2930 7404
rect 3513 7395 3571 7401
rect 3513 7392 3525 7395
rect 2924 7364 3525 7392
rect 2924 7352 2930 7364
rect 3513 7361 3525 7364
rect 3559 7361 3571 7395
rect 4154 7392 4160 7404
rect 4115 7364 4160 7392
rect 3513 7355 3571 7361
rect 4154 7352 4160 7364
rect 4212 7352 4218 7404
rect 4632 7401 4660 7500
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 5350 7488 5356 7540
rect 5408 7528 5414 7540
rect 6273 7531 6331 7537
rect 6273 7528 6285 7531
rect 5408 7500 6285 7528
rect 5408 7488 5414 7500
rect 6273 7497 6285 7500
rect 6319 7497 6331 7531
rect 6273 7491 6331 7497
rect 6641 7531 6699 7537
rect 6641 7497 6653 7531
rect 6687 7528 6699 7531
rect 7742 7528 7748 7540
rect 6687 7500 7748 7528
rect 6687 7497 6699 7500
rect 6641 7491 6699 7497
rect 7742 7488 7748 7500
rect 7800 7488 7806 7540
rect 8570 7528 8576 7540
rect 8531 7500 8576 7528
rect 8570 7488 8576 7500
rect 8628 7488 8634 7540
rect 14277 7531 14335 7537
rect 14277 7528 14289 7531
rect 8956 7500 14289 7528
rect 5718 7420 5724 7472
rect 5776 7460 5782 7472
rect 8018 7460 8024 7472
rect 5776 7432 8024 7460
rect 5776 7420 5782 7432
rect 8018 7420 8024 7432
rect 8076 7420 8082 7472
rect 4617 7395 4675 7401
rect 4617 7361 4629 7395
rect 4663 7361 4675 7395
rect 7377 7395 7435 7401
rect 7377 7392 7389 7395
rect 4617 7355 4675 7361
rect 5644 7364 7389 7392
rect 1394 7284 1400 7336
rect 1452 7324 1458 7336
rect 2317 7327 2375 7333
rect 2317 7324 2329 7327
rect 1452 7296 2329 7324
rect 1452 7284 1458 7296
rect 2317 7293 2329 7296
rect 2363 7293 2375 7327
rect 2317 7287 2375 7293
rect 4884 7327 4942 7333
rect 4884 7293 4896 7327
rect 4930 7324 4942 7327
rect 5166 7324 5172 7336
rect 4930 7296 5172 7324
rect 4930 7293 4942 7296
rect 4884 7287 4942 7293
rect 5166 7284 5172 7296
rect 5224 7324 5230 7336
rect 5644 7324 5672 7364
rect 7377 7361 7389 7364
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 8113 7395 8171 7401
rect 8113 7361 8125 7395
rect 8159 7392 8171 7395
rect 8956 7392 8984 7500
rect 14277 7497 14289 7500
rect 14323 7497 14335 7531
rect 14277 7491 14335 7497
rect 9950 7460 9956 7472
rect 9048 7432 9956 7460
rect 9048 7401 9076 7432
rect 9950 7420 9956 7432
rect 10008 7420 10014 7472
rect 11333 7463 11391 7469
rect 11333 7429 11345 7463
rect 11379 7429 11391 7463
rect 11333 7423 11391 7429
rect 8159 7364 8984 7392
rect 9033 7395 9091 7401
rect 8159 7361 8171 7364
rect 8113 7355 8171 7361
rect 9033 7361 9045 7395
rect 9079 7361 9091 7395
rect 9033 7355 9091 7361
rect 9217 7395 9275 7401
rect 9217 7361 9229 7395
rect 9263 7392 9275 7395
rect 9582 7392 9588 7404
rect 9263 7364 9588 7392
rect 9263 7361 9275 7364
rect 9217 7355 9275 7361
rect 9582 7352 9588 7364
rect 9640 7352 9646 7404
rect 10042 7352 10048 7404
rect 10100 7392 10106 7404
rect 10229 7395 10287 7401
rect 10100 7364 10145 7392
rect 10100 7352 10106 7364
rect 10229 7361 10241 7395
rect 10275 7392 10287 7395
rect 10502 7392 10508 7404
rect 10275 7364 10508 7392
rect 10275 7361 10287 7364
rect 10229 7355 10287 7361
rect 10502 7352 10508 7364
rect 10560 7352 10566 7404
rect 10594 7352 10600 7404
rect 10652 7392 10658 7404
rect 11241 7395 11299 7401
rect 11241 7392 11253 7395
rect 10652 7364 11253 7392
rect 10652 7352 10658 7364
rect 11241 7361 11253 7364
rect 11287 7361 11299 7395
rect 11241 7355 11299 7361
rect 5224 7296 5672 7324
rect 6457 7327 6515 7333
rect 5224 7284 5230 7296
rect 6457 7293 6469 7327
rect 6503 7324 6515 7327
rect 6641 7327 6699 7333
rect 6641 7324 6653 7327
rect 6503 7296 6653 7324
rect 6503 7293 6515 7296
rect 6457 7287 6515 7293
rect 6641 7293 6653 7296
rect 6687 7293 6699 7327
rect 7190 7324 7196 7336
rect 7151 7296 7196 7324
rect 6641 7287 6699 7293
rect 7190 7284 7196 7296
rect 7248 7284 7254 7336
rect 7282 7284 7288 7336
rect 7340 7324 7346 7336
rect 9953 7327 10011 7333
rect 9953 7324 9965 7327
rect 7340 7296 9965 7324
rect 7340 7284 7346 7296
rect 9953 7293 9965 7296
rect 9999 7293 10011 7327
rect 9953 7287 10011 7293
rect 10318 7284 10324 7336
rect 10376 7324 10382 7336
rect 10781 7327 10839 7333
rect 10781 7324 10793 7327
rect 10376 7296 10793 7324
rect 10376 7284 10382 7296
rect 10781 7293 10793 7296
rect 10827 7293 10839 7327
rect 11348 7324 11376 7423
rect 11422 7420 11428 7472
rect 11480 7460 11486 7472
rect 12526 7460 12532 7472
rect 11480 7432 12532 7460
rect 11480 7420 11486 7432
rect 12526 7420 12532 7432
rect 12584 7460 12590 7472
rect 13354 7460 13360 7472
rect 12584 7432 13360 7460
rect 12584 7420 12590 7432
rect 13354 7420 13360 7432
rect 13412 7420 13418 7472
rect 13449 7463 13507 7469
rect 13449 7429 13461 7463
rect 13495 7460 13507 7463
rect 14366 7460 14372 7472
rect 13495 7432 14372 7460
rect 13495 7429 13507 7432
rect 13449 7423 13507 7429
rect 14366 7420 14372 7432
rect 14424 7420 14430 7472
rect 11974 7392 11980 7404
rect 11935 7364 11980 7392
rect 11974 7352 11980 7364
rect 12032 7352 12038 7404
rect 12342 7352 12348 7404
rect 12400 7392 12406 7404
rect 12989 7395 13047 7401
rect 12989 7392 13001 7395
rect 12400 7364 13001 7392
rect 12400 7352 12406 7364
rect 12989 7361 13001 7364
rect 13035 7361 13047 7395
rect 12989 7355 13047 7361
rect 13630 7352 13636 7404
rect 13688 7392 13694 7404
rect 14001 7395 14059 7401
rect 14001 7392 14013 7395
rect 13688 7364 14013 7392
rect 13688 7352 13694 7364
rect 14001 7361 14013 7364
rect 14047 7361 14059 7395
rect 14001 7355 14059 7361
rect 14090 7352 14096 7404
rect 14148 7392 14154 7404
rect 14921 7395 14979 7401
rect 14921 7392 14933 7395
rect 14148 7364 14933 7392
rect 14148 7352 14154 7364
rect 14921 7361 14933 7364
rect 14967 7361 14979 7395
rect 14921 7355 14979 7361
rect 15013 7395 15071 7401
rect 15013 7361 15025 7395
rect 15059 7361 15071 7395
rect 15013 7355 15071 7361
rect 13909 7327 13967 7333
rect 13909 7324 13921 7327
rect 11348 7296 13921 7324
rect 10781 7287 10839 7293
rect 13909 7293 13921 7296
rect 13955 7293 13967 7327
rect 13909 7287 13967 7293
rect 14369 7327 14427 7333
rect 14369 7293 14381 7327
rect 14415 7324 14427 7327
rect 14829 7327 14887 7333
rect 14829 7324 14841 7327
rect 14415 7296 14841 7324
rect 14415 7293 14427 7296
rect 14369 7287 14427 7293
rect 14829 7293 14841 7296
rect 14875 7293 14887 7327
rect 14829 7287 14887 7293
rect 2409 7259 2467 7265
rect 2409 7225 2421 7259
rect 2455 7256 2467 7259
rect 2498 7256 2504 7268
rect 2455 7228 2504 7256
rect 2455 7225 2467 7228
rect 2409 7219 2467 7225
rect 2498 7216 2504 7228
rect 2556 7216 2562 7268
rect 4062 7216 4068 7268
rect 4120 7256 4126 7268
rect 13814 7256 13820 7268
rect 4120 7228 13308 7256
rect 13775 7228 13820 7256
rect 4120 7216 4126 7228
rect 1946 7188 1952 7200
rect 1907 7160 1952 7188
rect 1946 7148 1952 7160
rect 2004 7148 2010 7200
rect 2958 7188 2964 7200
rect 2919 7160 2964 7188
rect 2958 7148 2964 7160
rect 3016 7148 3022 7200
rect 3326 7188 3332 7200
rect 3287 7160 3332 7188
rect 3326 7148 3332 7160
rect 3384 7148 3390 7200
rect 3418 7148 3424 7200
rect 3476 7188 3482 7200
rect 5994 7188 6000 7200
rect 3476 7160 3521 7188
rect 5955 7160 6000 7188
rect 3476 7148 3482 7160
rect 5994 7148 6000 7160
rect 6052 7148 6058 7200
rect 6178 7148 6184 7200
rect 6236 7188 6242 7200
rect 6546 7188 6552 7200
rect 6236 7160 6552 7188
rect 6236 7148 6242 7160
rect 6546 7148 6552 7160
rect 6604 7148 6610 7200
rect 6825 7191 6883 7197
rect 6825 7157 6837 7191
rect 6871 7188 6883 7191
rect 7098 7188 7104 7200
rect 6871 7160 7104 7188
rect 6871 7157 6883 7160
rect 6825 7151 6883 7157
rect 7098 7148 7104 7160
rect 7156 7148 7162 7200
rect 7282 7188 7288 7200
rect 7243 7160 7288 7188
rect 7282 7148 7288 7160
rect 7340 7148 7346 7200
rect 8941 7191 8999 7197
rect 8941 7157 8953 7191
rect 8987 7188 8999 7191
rect 9306 7188 9312 7200
rect 8987 7160 9312 7188
rect 8987 7157 8999 7160
rect 8941 7151 8999 7157
rect 9306 7148 9312 7160
rect 9364 7148 9370 7200
rect 9585 7191 9643 7197
rect 9585 7157 9597 7191
rect 9631 7188 9643 7191
rect 10410 7188 10416 7200
rect 9631 7160 10416 7188
rect 9631 7157 9643 7160
rect 9585 7151 9643 7157
rect 10410 7148 10416 7160
rect 10468 7148 10474 7200
rect 10597 7191 10655 7197
rect 10597 7157 10609 7191
rect 10643 7188 10655 7191
rect 10686 7188 10692 7200
rect 10643 7160 10692 7188
rect 10643 7157 10655 7160
rect 10597 7151 10655 7157
rect 10686 7148 10692 7160
rect 10744 7148 10750 7200
rect 11241 7191 11299 7197
rect 11241 7157 11253 7191
rect 11287 7188 11299 7191
rect 11701 7191 11759 7197
rect 11701 7188 11713 7191
rect 11287 7160 11713 7188
rect 11287 7157 11299 7160
rect 11241 7151 11299 7157
rect 11701 7157 11713 7160
rect 11747 7157 11759 7191
rect 11701 7151 11759 7157
rect 11793 7191 11851 7197
rect 11793 7157 11805 7191
rect 11839 7188 11851 7191
rect 12437 7191 12495 7197
rect 12437 7188 12449 7191
rect 11839 7160 12449 7188
rect 11839 7157 11851 7160
rect 11793 7151 11851 7157
rect 12437 7157 12449 7160
rect 12483 7157 12495 7191
rect 12802 7188 12808 7200
rect 12763 7160 12808 7188
rect 12437 7151 12495 7157
rect 12802 7148 12808 7160
rect 12860 7148 12866 7200
rect 12897 7191 12955 7197
rect 12897 7157 12909 7191
rect 12943 7188 12955 7191
rect 13170 7188 13176 7200
rect 12943 7160 13176 7188
rect 12943 7157 12955 7160
rect 12897 7151 12955 7157
rect 13170 7148 13176 7160
rect 13228 7148 13234 7200
rect 13280 7188 13308 7228
rect 13814 7216 13820 7228
rect 13872 7216 13878 7268
rect 14274 7216 14280 7268
rect 14332 7256 14338 7268
rect 15028 7256 15056 7355
rect 14332 7228 15056 7256
rect 14332 7216 14338 7228
rect 13906 7188 13912 7200
rect 13280 7160 13912 7188
rect 13906 7148 13912 7160
rect 13964 7148 13970 7200
rect 14458 7188 14464 7200
rect 14419 7160 14464 7188
rect 14458 7148 14464 7160
rect 14516 7148 14522 7200
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 2866 6944 2872 6996
rect 2924 6984 2930 6996
rect 3053 6987 3111 6993
rect 3053 6984 3065 6987
rect 2924 6956 3065 6984
rect 2924 6944 2930 6956
rect 3053 6953 3065 6956
rect 3099 6953 3111 6987
rect 3053 6947 3111 6953
rect 5166 6944 5172 6996
rect 5224 6984 5230 6996
rect 5445 6987 5503 6993
rect 5445 6984 5457 6987
rect 5224 6956 5457 6984
rect 5224 6944 5230 6956
rect 5445 6953 5457 6956
rect 5491 6953 5503 6987
rect 5445 6947 5503 6953
rect 6822 6944 6828 6996
rect 6880 6984 6886 6996
rect 7929 6987 7987 6993
rect 7929 6984 7941 6987
rect 6880 6956 7941 6984
rect 6880 6944 6886 6956
rect 7929 6953 7941 6956
rect 7975 6953 7987 6987
rect 8570 6984 8576 6996
rect 8531 6956 8576 6984
rect 7929 6947 7987 6953
rect 8570 6944 8576 6956
rect 8628 6944 8634 6996
rect 10778 6984 10784 6996
rect 8864 6956 10784 6984
rect 4332 6919 4390 6925
rect 4332 6885 4344 6919
rect 4378 6916 4390 6919
rect 4890 6916 4896 6928
rect 4378 6888 4896 6916
rect 4378 6885 4390 6888
rect 4332 6879 4390 6885
rect 4890 6876 4896 6888
rect 4948 6876 4954 6928
rect 6914 6876 6920 6928
rect 6972 6916 6978 6928
rect 8202 6916 8208 6928
rect 6972 6888 8208 6916
rect 6972 6876 6978 6888
rect 8202 6876 8208 6888
rect 8260 6876 8266 6928
rect 8662 6876 8668 6928
rect 8720 6916 8726 6928
rect 8864 6916 8892 6956
rect 10778 6944 10784 6956
rect 10836 6944 10842 6996
rect 11054 6944 11060 6996
rect 11112 6984 11118 6996
rect 12342 6984 12348 6996
rect 11112 6956 12348 6984
rect 11112 6944 11118 6956
rect 12342 6944 12348 6956
rect 12400 6984 12406 6996
rect 12989 6987 13047 6993
rect 12989 6984 13001 6987
rect 12400 6956 13001 6984
rect 12400 6944 12406 6956
rect 12989 6953 13001 6956
rect 13035 6953 13047 6987
rect 12989 6947 13047 6953
rect 13633 6987 13691 6993
rect 13633 6953 13645 6987
rect 13679 6984 13691 6987
rect 13906 6984 13912 6996
rect 13679 6956 13912 6984
rect 13679 6953 13691 6956
rect 13633 6947 13691 6953
rect 13906 6944 13912 6956
rect 13964 6944 13970 6996
rect 14458 6944 14464 6996
rect 14516 6984 14522 6996
rect 15657 6987 15715 6993
rect 15657 6984 15669 6987
rect 14516 6956 15669 6984
rect 14516 6944 14522 6956
rect 15657 6953 15669 6956
rect 15703 6953 15715 6987
rect 15657 6947 15715 6953
rect 8720 6888 8892 6916
rect 8941 6919 8999 6925
rect 8720 6876 8726 6888
rect 8941 6885 8953 6919
rect 8987 6916 8999 6919
rect 11422 6916 11428 6928
rect 8987 6888 11428 6916
rect 8987 6885 8999 6888
rect 8941 6879 8999 6885
rect 11422 6876 11428 6888
rect 11480 6876 11486 6928
rect 13354 6876 13360 6928
rect 13412 6916 13418 6928
rect 18506 6916 18512 6928
rect 13412 6888 18512 6916
rect 13412 6876 13418 6888
rect 18506 6876 18512 6888
rect 18564 6876 18570 6928
rect 1673 6851 1731 6857
rect 1673 6817 1685 6851
rect 1719 6848 1731 6851
rect 1762 6848 1768 6860
rect 1719 6820 1768 6848
rect 1719 6817 1731 6820
rect 1673 6811 1731 6817
rect 1762 6808 1768 6820
rect 1820 6808 1826 6860
rect 1940 6851 1998 6857
rect 1940 6817 1952 6851
rect 1986 6848 1998 6851
rect 2222 6848 2228 6860
rect 1986 6820 2228 6848
rect 1986 6817 1998 6820
rect 1940 6811 1998 6817
rect 2222 6808 2228 6820
rect 2280 6808 2286 6860
rect 4065 6851 4123 6857
rect 4065 6817 4077 6851
rect 4111 6848 4123 6851
rect 4706 6848 4712 6860
rect 4111 6820 4712 6848
rect 4111 6817 4123 6820
rect 4065 6811 4123 6817
rect 4706 6808 4712 6820
rect 4764 6848 4770 6860
rect 5905 6851 5963 6857
rect 5905 6848 5917 6851
rect 4764 6820 5917 6848
rect 4764 6808 4770 6820
rect 5905 6817 5917 6820
rect 5951 6817 5963 6851
rect 5905 6811 5963 6817
rect 5994 6808 6000 6860
rect 6052 6848 6058 6860
rect 6172 6851 6230 6857
rect 6172 6848 6184 6851
rect 6052 6820 6184 6848
rect 6052 6808 6058 6820
rect 6172 6817 6184 6820
rect 6218 6848 6230 6851
rect 9582 6848 9588 6860
rect 6218 6820 6960 6848
rect 9495 6820 9588 6848
rect 6218 6817 6230 6820
rect 6172 6811 6230 6817
rect 2682 6740 2688 6792
rect 2740 6780 2746 6792
rect 3329 6783 3387 6789
rect 3329 6780 3341 6783
rect 2740 6752 3341 6780
rect 2740 6740 2746 6752
rect 3329 6749 3341 6752
rect 3375 6749 3387 6783
rect 3329 6743 3387 6749
rect 6932 6712 6960 6820
rect 9582 6808 9588 6820
rect 9640 6848 9646 6860
rect 9933 6851 9991 6857
rect 9933 6848 9945 6851
rect 9640 6820 9945 6848
rect 9640 6808 9646 6820
rect 9933 6817 9945 6820
rect 9979 6817 9991 6851
rect 11698 6848 11704 6860
rect 9933 6811 9991 6817
rect 11072 6820 11704 6848
rect 7098 6740 7104 6792
rect 7156 6780 7162 6792
rect 8021 6783 8079 6789
rect 8021 6780 8033 6783
rect 7156 6752 8033 6780
rect 7156 6740 7162 6752
rect 8021 6749 8033 6752
rect 8067 6749 8079 6783
rect 8021 6743 8079 6749
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6749 8171 6783
rect 8113 6743 8171 6749
rect 8128 6712 8156 6743
rect 8938 6740 8944 6792
rect 8996 6780 9002 6792
rect 9033 6783 9091 6789
rect 9033 6780 9045 6783
rect 8996 6752 9045 6780
rect 8996 6740 9002 6752
rect 9033 6749 9045 6752
rect 9079 6749 9091 6783
rect 9033 6743 9091 6749
rect 9217 6783 9275 6789
rect 9217 6749 9229 6783
rect 9263 6780 9275 6783
rect 9401 6783 9459 6789
rect 9401 6780 9413 6783
rect 9263 6752 9413 6780
rect 9263 6749 9275 6752
rect 9217 6743 9275 6749
rect 9401 6749 9413 6752
rect 9447 6749 9459 6783
rect 9674 6780 9680 6792
rect 9635 6752 9680 6780
rect 9401 6743 9459 6749
rect 6932 6684 8156 6712
rect 9048 6712 9076 6743
rect 9674 6740 9680 6752
rect 9732 6740 9738 6792
rect 9582 6712 9588 6724
rect 9048 6684 9588 6712
rect 9582 6672 9588 6684
rect 9640 6672 9646 6724
rect 11072 6721 11100 6820
rect 11698 6808 11704 6820
rect 11756 6808 11762 6860
rect 11882 6857 11888 6860
rect 11876 6848 11888 6857
rect 11843 6820 11888 6848
rect 11876 6811 11888 6820
rect 11882 6808 11888 6811
rect 11940 6808 11946 6860
rect 12820 6820 15884 6848
rect 11606 6780 11612 6792
rect 11567 6752 11612 6780
rect 11606 6740 11612 6752
rect 11664 6740 11670 6792
rect 11057 6715 11115 6721
rect 11057 6681 11069 6715
rect 11103 6681 11115 6715
rect 11057 6675 11115 6681
rect 7190 6604 7196 6656
rect 7248 6644 7254 6656
rect 7285 6647 7343 6653
rect 7285 6644 7297 6647
rect 7248 6616 7297 6644
rect 7248 6604 7254 6616
rect 7285 6613 7297 6616
rect 7331 6613 7343 6647
rect 7285 6607 7343 6613
rect 7374 6604 7380 6656
rect 7432 6644 7438 6656
rect 7561 6647 7619 6653
rect 7561 6644 7573 6647
rect 7432 6616 7573 6644
rect 7432 6604 7438 6616
rect 7561 6613 7573 6616
rect 7607 6613 7619 6647
rect 7561 6607 7619 6613
rect 9214 6604 9220 6656
rect 9272 6644 9278 6656
rect 11072 6644 11100 6675
rect 9272 6616 11100 6644
rect 9272 6604 9278 6616
rect 11146 6604 11152 6656
rect 11204 6644 11210 6656
rect 12820 6644 12848 6820
rect 12894 6740 12900 6792
rect 12952 6780 12958 6792
rect 13078 6780 13084 6792
rect 12952 6752 13084 6780
rect 12952 6740 12958 6752
rect 13078 6740 13084 6752
rect 13136 6780 13142 6792
rect 13725 6783 13783 6789
rect 13725 6780 13737 6783
rect 13136 6752 13737 6780
rect 13136 6740 13142 6752
rect 13725 6749 13737 6752
rect 13771 6749 13783 6783
rect 13725 6743 13783 6749
rect 13814 6740 13820 6792
rect 13872 6780 13878 6792
rect 13909 6783 13967 6789
rect 13909 6780 13921 6783
rect 13872 6752 13921 6780
rect 13872 6740 13878 6752
rect 13909 6749 13921 6752
rect 13955 6780 13967 6783
rect 14274 6780 14280 6792
rect 13955 6752 14280 6780
rect 13955 6749 13967 6752
rect 13909 6743 13967 6749
rect 14274 6740 14280 6752
rect 14332 6740 14338 6792
rect 14550 6740 14556 6792
rect 14608 6780 14614 6792
rect 15856 6789 15884 6820
rect 14737 6783 14795 6789
rect 14737 6780 14749 6783
rect 14608 6752 14749 6780
rect 14608 6740 14614 6752
rect 14737 6749 14749 6752
rect 14783 6749 14795 6783
rect 14737 6743 14795 6749
rect 15749 6783 15807 6789
rect 15749 6749 15761 6783
rect 15795 6749 15807 6783
rect 15749 6743 15807 6749
rect 15841 6783 15899 6789
rect 15841 6749 15853 6783
rect 15887 6780 15899 6783
rect 17494 6780 17500 6792
rect 15887 6752 17500 6780
rect 15887 6749 15899 6752
rect 15841 6743 15899 6749
rect 13265 6715 13323 6721
rect 13265 6681 13277 6715
rect 13311 6712 13323 6715
rect 15764 6712 15792 6743
rect 17494 6740 17500 6752
rect 17552 6740 17558 6792
rect 13311 6684 15792 6712
rect 13311 6681 13323 6684
rect 13265 6675 13323 6681
rect 15286 6644 15292 6656
rect 11204 6616 12848 6644
rect 15247 6616 15292 6644
rect 11204 6604 11210 6616
rect 15286 6604 15292 6616
rect 15344 6604 15350 6656
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 3237 6443 3295 6449
rect 3237 6409 3249 6443
rect 3283 6440 3295 6443
rect 3418 6440 3424 6452
rect 3283 6412 3424 6440
rect 3283 6409 3295 6412
rect 3237 6403 3295 6409
rect 3418 6400 3424 6412
rect 3476 6400 3482 6452
rect 5721 6443 5779 6449
rect 5721 6409 5733 6443
rect 5767 6440 5779 6443
rect 7282 6440 7288 6452
rect 5767 6412 7288 6440
rect 5767 6409 5779 6412
rect 5721 6403 5779 6409
rect 7282 6400 7288 6412
rect 7340 6400 7346 6452
rect 7650 6440 7656 6452
rect 7392 6412 7656 6440
rect 2961 6375 3019 6381
rect 2961 6341 2973 6375
rect 3007 6341 3019 6375
rect 2961 6335 3019 6341
rect 2976 6304 3004 6335
rect 3602 6332 3608 6384
rect 3660 6372 3666 6384
rect 6914 6372 6920 6384
rect 3660 6344 6920 6372
rect 3660 6332 3666 6344
rect 6914 6332 6920 6344
rect 6972 6332 6978 6384
rect 7190 6332 7196 6384
rect 7248 6372 7254 6384
rect 7392 6372 7420 6412
rect 7650 6400 7656 6412
rect 7708 6440 7714 6452
rect 10045 6443 10103 6449
rect 7708 6412 8892 6440
rect 7708 6400 7714 6412
rect 7248 6344 7420 6372
rect 7248 6332 7254 6344
rect 3789 6307 3847 6313
rect 3789 6304 3801 6307
rect 2976 6276 3801 6304
rect 1854 6245 1860 6248
rect 1581 6239 1639 6245
rect 1581 6205 1593 6239
rect 1627 6205 1639 6239
rect 1848 6236 1860 6245
rect 1767 6208 1860 6236
rect 1581 6199 1639 6205
rect 1848 6199 1860 6208
rect 1912 6236 1918 6248
rect 2866 6236 2872 6248
rect 1912 6208 2872 6236
rect 1596 6168 1624 6199
rect 1854 6196 1860 6199
rect 1912 6196 1918 6208
rect 2866 6196 2872 6208
rect 2924 6196 2930 6248
rect 1762 6168 1768 6180
rect 1596 6140 1768 6168
rect 1762 6128 1768 6140
rect 1820 6128 1826 6180
rect 2222 6060 2228 6112
rect 2280 6100 2286 6112
rect 2976 6100 3004 6276
rect 3789 6273 3801 6276
rect 3835 6273 3847 6307
rect 3789 6267 3847 6273
rect 4893 6307 4951 6313
rect 4893 6273 4905 6307
rect 4939 6304 4951 6307
rect 5258 6304 5264 6316
rect 4939 6276 5264 6304
rect 4939 6273 4951 6276
rect 4893 6267 4951 6273
rect 5258 6264 5264 6276
rect 5316 6264 5322 6316
rect 6270 6304 6276 6316
rect 5368 6276 6132 6304
rect 6231 6276 6276 6304
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6236 4767 6239
rect 5368 6236 5396 6276
rect 4755 6208 5396 6236
rect 4755 6205 4767 6208
rect 4709 6199 4767 6205
rect 5442 6196 5448 6248
rect 5500 6236 5506 6248
rect 6104 6236 6132 6276
rect 6270 6264 6276 6276
rect 6328 6264 6334 6316
rect 6638 6264 6644 6316
rect 6696 6304 6702 6316
rect 6696 6276 7236 6304
rect 6696 6264 6702 6276
rect 6914 6236 6920 6248
rect 5500 6208 5545 6236
rect 6104 6208 6920 6236
rect 5500 6196 5506 6208
rect 6914 6196 6920 6208
rect 6972 6196 6978 6248
rect 7208 6245 7236 6276
rect 7282 6264 7288 6316
rect 7340 6304 7346 6316
rect 7377 6307 7435 6313
rect 7377 6304 7389 6307
rect 7340 6276 7389 6304
rect 7340 6264 7346 6276
rect 7377 6273 7389 6276
rect 7423 6273 7435 6307
rect 8864 6304 8892 6412
rect 10045 6409 10057 6443
rect 10091 6440 10103 6443
rect 10594 6440 10600 6452
rect 10091 6412 10600 6440
rect 10091 6409 10103 6412
rect 10045 6403 10103 6409
rect 10594 6400 10600 6412
rect 10652 6400 10658 6452
rect 19150 6440 19156 6452
rect 11348 6412 19156 6440
rect 11348 6384 11376 6412
rect 19150 6400 19156 6412
rect 19208 6400 19214 6452
rect 9214 6372 9220 6384
rect 9127 6344 9220 6372
rect 9214 6332 9220 6344
rect 9272 6372 9278 6384
rect 11146 6372 11152 6384
rect 9272 6344 11152 6372
rect 9272 6332 9278 6344
rect 11146 6332 11152 6344
rect 11204 6332 11210 6384
rect 11330 6332 11336 6384
rect 11388 6332 11394 6384
rect 12710 6372 12716 6384
rect 11440 6344 12716 6372
rect 10134 6304 10140 6316
rect 8864 6276 10140 6304
rect 7377 6267 7435 6273
rect 10134 6264 10140 6276
rect 10192 6264 10198 6316
rect 10689 6307 10747 6313
rect 10689 6273 10701 6307
rect 10735 6304 10747 6307
rect 11054 6304 11060 6316
rect 10735 6276 11060 6304
rect 10735 6273 10747 6276
rect 10689 6267 10747 6273
rect 11054 6264 11060 6276
rect 11112 6264 11118 6316
rect 11241 6307 11299 6313
rect 11241 6273 11253 6307
rect 11287 6304 11299 6307
rect 11440 6304 11468 6344
rect 12710 6332 12716 6344
rect 12768 6332 12774 6384
rect 11287 6276 11468 6304
rect 11977 6307 12035 6313
rect 11287 6273 11299 6276
rect 11241 6267 11299 6273
rect 11977 6273 11989 6307
rect 12023 6304 12035 6307
rect 12250 6304 12256 6316
rect 12023 6276 12256 6304
rect 12023 6273 12035 6276
rect 11977 6267 12035 6273
rect 12250 6264 12256 6276
rect 12308 6264 12314 6316
rect 13081 6307 13139 6313
rect 13081 6273 13093 6307
rect 13127 6304 13139 6307
rect 13170 6304 13176 6316
rect 13127 6276 13176 6304
rect 13127 6273 13139 6276
rect 13081 6267 13139 6273
rect 13170 6264 13176 6276
rect 13228 6264 13234 6316
rect 13262 6264 13268 6316
rect 13320 6304 13326 6316
rect 13541 6307 13599 6313
rect 13541 6304 13553 6307
rect 13320 6276 13553 6304
rect 13320 6264 13326 6276
rect 13541 6273 13553 6276
rect 13587 6273 13599 6307
rect 13541 6267 13599 6273
rect 7193 6239 7251 6245
rect 7193 6205 7205 6239
rect 7239 6205 7251 6239
rect 7193 6199 7251 6205
rect 7466 6196 7472 6248
rect 7524 6236 7530 6248
rect 7837 6239 7895 6245
rect 7837 6236 7849 6239
rect 7524 6208 7849 6236
rect 7524 6196 7530 6208
rect 7837 6205 7849 6208
rect 7883 6205 7895 6239
rect 7837 6199 7895 6205
rect 8104 6239 8162 6245
rect 8104 6205 8116 6239
rect 8150 6236 8162 6239
rect 9122 6236 9128 6248
rect 8150 6208 9128 6236
rect 8150 6205 8162 6208
rect 8104 6199 8162 6205
rect 9122 6196 9128 6208
rect 9180 6196 9186 6248
rect 10410 6196 10416 6248
rect 10468 6236 10474 6248
rect 13446 6236 13452 6248
rect 10468 6208 13452 6236
rect 10468 6196 10474 6208
rect 13446 6196 13452 6208
rect 13504 6196 13510 6248
rect 13556 6236 13584 6267
rect 15194 6236 15200 6248
rect 13556 6208 15200 6236
rect 15194 6196 15200 6208
rect 15252 6196 15258 6248
rect 6546 6128 6552 6180
rect 6604 6168 6610 6180
rect 7285 6171 7343 6177
rect 7285 6168 7297 6171
rect 6604 6140 7297 6168
rect 6604 6128 6610 6140
rect 7285 6137 7297 6140
rect 7331 6168 7343 6171
rect 7926 6168 7932 6180
rect 7331 6140 7932 6168
rect 7331 6137 7343 6140
rect 7285 6131 7343 6137
rect 7926 6128 7932 6140
rect 7984 6128 7990 6180
rect 8018 6128 8024 6180
rect 8076 6168 8082 6180
rect 8076 6140 8147 6168
rect 8076 6128 8082 6140
rect 3602 6100 3608 6112
rect 2280 6072 3004 6100
rect 3563 6072 3608 6100
rect 2280 6060 2286 6072
rect 3602 6060 3608 6072
rect 3660 6060 3666 6112
rect 3697 6103 3755 6109
rect 3697 6069 3709 6103
rect 3743 6100 3755 6103
rect 4249 6103 4307 6109
rect 4249 6100 4261 6103
rect 3743 6072 4261 6100
rect 3743 6069 3755 6072
rect 3697 6063 3755 6069
rect 4249 6069 4261 6072
rect 4295 6069 4307 6103
rect 4614 6100 4620 6112
rect 4575 6072 4620 6100
rect 4249 6063 4307 6069
rect 4614 6060 4620 6072
rect 4672 6060 4678 6112
rect 5261 6103 5319 6109
rect 5261 6069 5273 6103
rect 5307 6100 5319 6103
rect 5350 6100 5356 6112
rect 5307 6072 5356 6100
rect 5307 6069 5319 6072
rect 5261 6063 5319 6069
rect 5350 6060 5356 6072
rect 5408 6060 5414 6112
rect 6086 6100 6092 6112
rect 6047 6072 6092 6100
rect 6086 6060 6092 6072
rect 6144 6060 6150 6112
rect 6181 6103 6239 6109
rect 6181 6069 6193 6103
rect 6227 6100 6239 6103
rect 6825 6103 6883 6109
rect 6825 6100 6837 6103
rect 6227 6072 6837 6100
rect 6227 6069 6239 6072
rect 6181 6063 6239 6069
rect 6825 6069 6837 6072
rect 6871 6069 6883 6103
rect 8119 6100 8147 6140
rect 8202 6128 8208 6180
rect 8260 6168 8266 6180
rect 11241 6171 11299 6177
rect 11241 6168 11253 6171
rect 8260 6140 11253 6168
rect 8260 6128 8266 6140
rect 11241 6137 11253 6140
rect 11287 6137 11299 6171
rect 11241 6131 11299 6137
rect 11701 6171 11759 6177
rect 11701 6137 11713 6171
rect 11747 6168 11759 6171
rect 12526 6168 12532 6180
rect 11747 6140 12532 6168
rect 11747 6137 11759 6140
rect 11701 6131 11759 6137
rect 12526 6128 12532 6140
rect 12584 6128 12590 6180
rect 12618 6128 12624 6180
rect 12676 6168 12682 6180
rect 12805 6171 12863 6177
rect 12805 6168 12817 6171
rect 12676 6140 12817 6168
rect 12676 6128 12682 6140
rect 12805 6137 12817 6140
rect 12851 6137 12863 6171
rect 12805 6131 12863 6137
rect 13808 6171 13866 6177
rect 13808 6137 13820 6171
rect 13854 6168 13866 6171
rect 13998 6168 14004 6180
rect 13854 6140 14004 6168
rect 13854 6137 13866 6140
rect 13808 6131 13866 6137
rect 13998 6128 14004 6140
rect 14056 6128 14062 6180
rect 15442 6171 15500 6177
rect 15442 6168 15454 6171
rect 15028 6140 15454 6168
rect 15028 6112 15056 6140
rect 15442 6137 15454 6140
rect 15488 6137 15500 6171
rect 15442 6131 15500 6137
rect 10226 6100 10232 6112
rect 8119 6072 10232 6100
rect 6825 6063 6883 6069
rect 10226 6060 10232 6072
rect 10284 6060 10290 6112
rect 10318 6060 10324 6112
rect 10376 6100 10382 6112
rect 10413 6103 10471 6109
rect 10413 6100 10425 6103
rect 10376 6072 10425 6100
rect 10376 6060 10382 6072
rect 10413 6069 10425 6072
rect 10459 6069 10471 6103
rect 10413 6063 10471 6069
rect 10505 6103 10563 6109
rect 10505 6069 10517 6103
rect 10551 6100 10563 6103
rect 10594 6100 10600 6112
rect 10551 6072 10600 6100
rect 10551 6069 10563 6072
rect 10505 6063 10563 6069
rect 10594 6060 10600 6072
rect 10652 6060 10658 6112
rect 10962 6060 10968 6112
rect 11020 6100 11026 6112
rect 11333 6103 11391 6109
rect 11333 6100 11345 6103
rect 11020 6072 11345 6100
rect 11020 6060 11026 6072
rect 11333 6069 11345 6072
rect 11379 6069 11391 6103
rect 11333 6063 11391 6069
rect 11793 6103 11851 6109
rect 11793 6069 11805 6103
rect 11839 6100 11851 6103
rect 12437 6103 12495 6109
rect 12437 6100 12449 6103
rect 11839 6072 12449 6100
rect 11839 6069 11851 6072
rect 11793 6063 11851 6069
rect 12437 6069 12449 6072
rect 12483 6069 12495 6103
rect 12437 6063 12495 6069
rect 12710 6060 12716 6112
rect 12768 6100 12774 6112
rect 12897 6103 12955 6109
rect 12897 6100 12909 6103
rect 12768 6072 12909 6100
rect 12768 6060 12774 6072
rect 12897 6069 12909 6072
rect 12943 6100 12955 6103
rect 13722 6100 13728 6112
rect 12943 6072 13728 6100
rect 12943 6069 12955 6072
rect 12897 6063 12955 6069
rect 13722 6060 13728 6072
rect 13780 6060 13786 6112
rect 14921 6103 14979 6109
rect 14921 6069 14933 6103
rect 14967 6100 14979 6103
rect 15010 6100 15016 6112
rect 14967 6072 15016 6100
rect 14967 6069 14979 6072
rect 14921 6063 14979 6069
rect 15010 6060 15016 6072
rect 15068 6060 15074 6112
rect 15562 6060 15568 6112
rect 15620 6100 15626 6112
rect 16577 6103 16635 6109
rect 16577 6100 16589 6103
rect 15620 6072 16589 6100
rect 15620 6060 15626 6072
rect 16577 6069 16589 6072
rect 16623 6069 16635 6103
rect 16577 6063 16635 6069
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 1946 5856 1952 5908
rect 2004 5896 2010 5908
rect 2041 5899 2099 5905
rect 2041 5896 2053 5899
rect 2004 5868 2053 5896
rect 2004 5856 2010 5868
rect 2041 5865 2053 5868
rect 2087 5865 2099 5899
rect 2041 5859 2099 5865
rect 2593 5899 2651 5905
rect 2593 5865 2605 5899
rect 2639 5896 2651 5899
rect 3602 5896 3608 5908
rect 2639 5868 3608 5896
rect 2639 5865 2651 5868
rect 2593 5859 2651 5865
rect 3602 5856 3608 5868
rect 3660 5856 3666 5908
rect 4614 5856 4620 5908
rect 4672 5896 4678 5908
rect 5442 5896 5448 5908
rect 4672 5868 5448 5896
rect 4672 5856 4678 5868
rect 5442 5856 5448 5868
rect 5500 5856 5506 5908
rect 6089 5899 6147 5905
rect 6089 5865 6101 5899
rect 6135 5896 6147 5899
rect 6270 5896 6276 5908
rect 6135 5868 6276 5896
rect 6135 5865 6147 5868
rect 6089 5859 6147 5865
rect 6270 5856 6276 5868
rect 6328 5856 6334 5908
rect 6362 5856 6368 5908
rect 6420 5896 6426 5908
rect 10318 5896 10324 5908
rect 6420 5868 10324 5896
rect 6420 5856 6426 5868
rect 9600 5840 9628 5868
rect 10318 5856 10324 5868
rect 10376 5856 10382 5908
rect 10597 5899 10655 5905
rect 10597 5865 10609 5899
rect 10643 5865 10655 5899
rect 10962 5896 10968 5908
rect 10923 5868 10968 5896
rect 10597 5859 10655 5865
rect 2774 5788 2780 5840
rect 2832 5828 2838 5840
rect 2961 5831 3019 5837
rect 2961 5828 2973 5831
rect 2832 5800 2973 5828
rect 2832 5788 2838 5800
rect 2961 5797 2973 5800
rect 3007 5797 3019 5831
rect 2961 5791 3019 5797
rect 4976 5831 5034 5837
rect 4976 5797 4988 5831
rect 5022 5828 5034 5831
rect 6914 5828 6920 5840
rect 5022 5800 6920 5828
rect 5022 5797 5034 5800
rect 4976 5791 5034 5797
rect 6914 5788 6920 5800
rect 6972 5828 6978 5840
rect 7282 5828 7288 5840
rect 6972 5800 7288 5828
rect 6972 5788 6978 5800
rect 7282 5788 7288 5800
rect 7340 5788 7346 5840
rect 7552 5831 7610 5837
rect 7552 5797 7564 5831
rect 7598 5828 7610 5831
rect 9214 5828 9220 5840
rect 7598 5800 9220 5828
rect 7598 5797 7610 5800
rect 7552 5791 7610 5797
rect 9214 5788 9220 5800
rect 9272 5788 9278 5840
rect 9582 5788 9588 5840
rect 9640 5788 9646 5840
rect 10612 5828 10640 5859
rect 10962 5856 10968 5868
rect 11020 5856 11026 5908
rect 13078 5896 13084 5908
rect 11532 5868 13084 5896
rect 11532 5828 11560 5868
rect 13078 5856 13084 5868
rect 13136 5856 13142 5908
rect 14550 5896 14556 5908
rect 14511 5868 14556 5896
rect 14550 5856 14556 5868
rect 14608 5856 14614 5908
rect 16669 5899 16727 5905
rect 16669 5896 16681 5899
rect 14660 5868 16681 5896
rect 14660 5828 14688 5868
rect 16669 5865 16681 5868
rect 16715 5865 16727 5899
rect 17402 5896 17408 5908
rect 17363 5868 17408 5896
rect 16669 5859 16727 5865
rect 17402 5856 17408 5868
rect 17460 5856 17466 5908
rect 15562 5837 15568 5840
rect 15556 5828 15568 5837
rect 10612 5800 11560 5828
rect 11624 5800 14688 5828
rect 15523 5800 15568 5828
rect 1949 5763 2007 5769
rect 1949 5729 1961 5763
rect 1995 5760 2007 5763
rect 2682 5760 2688 5772
rect 1995 5732 2688 5760
rect 1995 5729 2007 5732
rect 1949 5723 2007 5729
rect 2682 5720 2688 5732
rect 2740 5720 2746 5772
rect 2866 5720 2872 5772
rect 2924 5760 2930 5772
rect 5258 5760 5264 5772
rect 2924 5732 5264 5760
rect 2924 5720 2930 5732
rect 2222 5692 2228 5704
rect 2183 5664 2228 5692
rect 2222 5652 2228 5664
rect 2280 5652 2286 5704
rect 2958 5652 2964 5704
rect 3016 5692 3022 5704
rect 3252 5701 3280 5732
rect 5258 5720 5264 5732
rect 5316 5760 5322 5772
rect 11624 5760 11652 5800
rect 15556 5791 15568 5800
rect 15562 5788 15568 5791
rect 15620 5788 15626 5840
rect 5316 5732 11652 5760
rect 11876 5763 11934 5769
rect 5316 5720 5322 5732
rect 11876 5729 11888 5763
rect 11922 5760 11934 5763
rect 12250 5760 12256 5772
rect 11922 5732 12256 5760
rect 11922 5729 11934 5732
rect 11876 5723 11934 5729
rect 12250 5720 12256 5732
rect 12308 5760 12314 5772
rect 12618 5760 12624 5772
rect 12308 5732 12624 5760
rect 12308 5720 12314 5732
rect 12618 5720 12624 5732
rect 12676 5720 12682 5772
rect 13446 5720 13452 5772
rect 13504 5760 13510 5772
rect 14645 5763 14703 5769
rect 14645 5760 14657 5763
rect 13504 5732 14657 5760
rect 13504 5720 13510 5732
rect 14645 5729 14657 5732
rect 14691 5729 14703 5763
rect 14645 5723 14703 5729
rect 15194 5720 15200 5772
rect 15252 5760 15258 5772
rect 15289 5763 15347 5769
rect 15289 5760 15301 5763
rect 15252 5732 15301 5760
rect 15252 5720 15258 5732
rect 15289 5729 15301 5732
rect 15335 5729 15347 5763
rect 15289 5723 15347 5729
rect 15378 5720 15384 5772
rect 15436 5760 15442 5772
rect 17313 5763 17371 5769
rect 17313 5760 17325 5763
rect 15436 5732 17325 5760
rect 15436 5720 15442 5732
rect 17313 5729 17325 5732
rect 17359 5729 17371 5763
rect 17313 5723 17371 5729
rect 17954 5720 17960 5772
rect 18012 5760 18018 5772
rect 18877 5763 18935 5769
rect 18877 5760 18889 5763
rect 18012 5732 18889 5760
rect 18012 5720 18018 5732
rect 18877 5729 18889 5732
rect 18923 5729 18935 5763
rect 18877 5723 18935 5729
rect 3053 5695 3111 5701
rect 3053 5692 3065 5695
rect 3016 5664 3065 5692
rect 3016 5652 3022 5664
rect 3053 5661 3065 5664
rect 3099 5661 3111 5695
rect 3053 5655 3111 5661
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5661 3295 5695
rect 3237 5655 3295 5661
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5661 4767 5695
rect 4709 5655 4767 5661
rect 1581 5627 1639 5633
rect 1581 5593 1593 5627
rect 1627 5624 1639 5627
rect 3326 5624 3332 5636
rect 1627 5596 3332 5624
rect 1627 5593 1639 5596
rect 1581 5587 1639 5593
rect 3326 5584 3332 5596
rect 3384 5584 3390 5636
rect 4724 5568 4752 5655
rect 5810 5652 5816 5704
rect 5868 5692 5874 5704
rect 6270 5692 6276 5704
rect 5868 5664 6276 5692
rect 5868 5652 5874 5664
rect 6270 5652 6276 5664
rect 6328 5652 6334 5704
rect 6822 5652 6828 5704
rect 6880 5692 6886 5704
rect 7285 5695 7343 5701
rect 7285 5692 7297 5695
rect 6880 5664 7297 5692
rect 6880 5652 6886 5664
rect 7285 5661 7297 5664
rect 7331 5661 7343 5695
rect 11054 5692 11060 5704
rect 11015 5664 11060 5692
rect 7285 5655 7343 5661
rect 11054 5652 11060 5664
rect 11112 5652 11118 5704
rect 11241 5695 11299 5701
rect 11241 5661 11253 5695
rect 11287 5692 11299 5695
rect 11606 5692 11612 5704
rect 11287 5664 11468 5692
rect 11567 5664 11612 5692
rect 11287 5661 11299 5664
rect 11241 5655 11299 5661
rect 6638 5584 6644 5636
rect 6696 5624 6702 5636
rect 9490 5624 9496 5636
rect 6696 5596 7328 5624
rect 6696 5584 6702 5596
rect 2958 5516 2964 5568
rect 3016 5556 3022 5568
rect 3970 5556 3976 5568
rect 3016 5528 3976 5556
rect 3016 5516 3022 5528
rect 3970 5516 3976 5528
rect 4028 5516 4034 5568
rect 4706 5556 4712 5568
rect 4619 5528 4712 5556
rect 4706 5516 4712 5528
rect 4764 5556 4770 5568
rect 5350 5556 5356 5568
rect 4764 5528 5356 5556
rect 4764 5516 4770 5528
rect 5350 5516 5356 5528
rect 5408 5556 5414 5568
rect 6822 5556 6828 5568
rect 5408 5528 6828 5556
rect 5408 5516 5414 5528
rect 6822 5516 6828 5528
rect 6880 5516 6886 5568
rect 7300 5556 7328 5596
rect 8588 5596 9496 5624
rect 8588 5556 8616 5596
rect 9490 5584 9496 5596
rect 9548 5624 9554 5636
rect 11330 5624 11336 5636
rect 9548 5596 11336 5624
rect 9548 5584 9554 5596
rect 11330 5584 11336 5596
rect 11388 5584 11394 5636
rect 7300 5528 8616 5556
rect 8665 5559 8723 5565
rect 8665 5525 8677 5559
rect 8711 5556 8723 5559
rect 8846 5556 8852 5568
rect 8711 5528 8852 5556
rect 8711 5525 8723 5528
rect 8665 5519 8723 5525
rect 8846 5516 8852 5528
rect 8904 5516 8910 5568
rect 11440 5556 11468 5664
rect 11606 5652 11612 5664
rect 11664 5652 11670 5704
rect 13262 5692 13268 5704
rect 13223 5664 13268 5692
rect 13262 5652 13268 5664
rect 13320 5652 13326 5704
rect 14829 5695 14887 5701
rect 14829 5661 14841 5695
rect 14875 5692 14887 5695
rect 15010 5692 15016 5704
rect 14875 5664 15016 5692
rect 14875 5661 14887 5664
rect 14829 5655 14887 5661
rect 15010 5652 15016 5664
rect 15068 5652 15074 5704
rect 17494 5692 17500 5704
rect 17455 5664 17500 5692
rect 17494 5652 17500 5664
rect 17552 5652 17558 5704
rect 19153 5695 19211 5701
rect 19153 5661 19165 5695
rect 19199 5692 19211 5695
rect 19794 5692 19800 5704
rect 19199 5664 19800 5692
rect 19199 5661 19211 5664
rect 19153 5655 19211 5661
rect 19794 5652 19800 5664
rect 19852 5652 19858 5704
rect 11882 5556 11888 5568
rect 11440 5528 11888 5556
rect 11882 5516 11888 5528
rect 11940 5556 11946 5568
rect 12989 5559 13047 5565
rect 12989 5556 13001 5559
rect 11940 5528 13001 5556
rect 11940 5516 11946 5528
rect 12989 5525 13001 5528
rect 13035 5525 13047 5559
rect 12989 5519 13047 5525
rect 14185 5559 14243 5565
rect 14185 5525 14197 5559
rect 14231 5556 14243 5559
rect 15470 5556 15476 5568
rect 14231 5528 15476 5556
rect 14231 5525 14243 5528
rect 14185 5519 14243 5525
rect 15470 5516 15476 5528
rect 15528 5516 15534 5568
rect 16942 5556 16948 5568
rect 16903 5528 16948 5556
rect 16942 5516 16948 5528
rect 17000 5516 17006 5568
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 4062 5312 4068 5364
rect 4120 5352 4126 5364
rect 4120 5324 5580 5352
rect 4120 5312 4126 5324
rect 5552 5284 5580 5324
rect 5718 5312 5724 5364
rect 5776 5352 5782 5364
rect 5997 5355 6055 5361
rect 5997 5352 6009 5355
rect 5776 5324 6009 5352
rect 5776 5312 5782 5324
rect 5997 5321 6009 5324
rect 6043 5321 6055 5355
rect 8478 5352 8484 5364
rect 5997 5315 6055 5321
rect 6104 5324 7788 5352
rect 8439 5324 8484 5352
rect 6104 5284 6132 5324
rect 5552 5256 6132 5284
rect 7760 5284 7788 5324
rect 8478 5312 8484 5324
rect 8536 5312 8542 5364
rect 11054 5312 11060 5364
rect 11112 5352 11118 5364
rect 11333 5355 11391 5361
rect 11333 5352 11345 5355
rect 11112 5324 11345 5352
rect 11112 5312 11118 5324
rect 11333 5321 11345 5324
rect 11379 5321 11391 5355
rect 12526 5352 12532 5364
rect 12487 5324 12532 5352
rect 11333 5315 11391 5321
rect 12526 5312 12532 5324
rect 12584 5312 12590 5364
rect 13449 5355 13507 5361
rect 13449 5352 13461 5355
rect 13004 5324 13461 5352
rect 12894 5284 12900 5296
rect 7760 5256 12900 5284
rect 12894 5244 12900 5256
rect 12952 5244 12958 5296
rect 3878 5216 3884 5228
rect 3839 5188 3884 5216
rect 3878 5176 3884 5188
rect 3936 5176 3942 5228
rect 8202 5176 8208 5228
rect 8260 5216 8266 5228
rect 8941 5219 8999 5225
rect 8941 5216 8953 5219
rect 8260 5188 8953 5216
rect 8260 5176 8266 5188
rect 8941 5185 8953 5188
rect 8987 5185 8999 5219
rect 9122 5216 9128 5228
rect 9083 5188 9128 5216
rect 8941 5179 8999 5185
rect 9122 5176 9128 5188
rect 9180 5176 9186 5228
rect 10502 5216 10508 5228
rect 10463 5188 10508 5216
rect 10502 5176 10508 5188
rect 10560 5176 10566 5228
rect 11977 5219 12035 5225
rect 11977 5185 11989 5219
rect 12023 5216 12035 5219
rect 12618 5216 12624 5228
rect 12023 5188 12624 5216
rect 12023 5185 12035 5188
rect 11977 5179 12035 5185
rect 12618 5176 12624 5188
rect 12676 5176 12682 5228
rect 13004 5225 13032 5324
rect 13449 5321 13461 5324
rect 13495 5352 13507 5355
rect 13538 5352 13544 5364
rect 13495 5324 13544 5352
rect 13495 5321 13507 5324
rect 13449 5315 13507 5321
rect 13538 5312 13544 5324
rect 13596 5312 13602 5364
rect 15197 5287 15255 5293
rect 15197 5253 15209 5287
rect 15243 5284 15255 5287
rect 15243 5256 16988 5284
rect 15243 5253 15255 5256
rect 15197 5247 15255 5253
rect 12989 5219 13047 5225
rect 12989 5185 13001 5219
rect 13035 5185 13047 5219
rect 13170 5216 13176 5228
rect 13083 5188 13176 5216
rect 12989 5179 13047 5185
rect 13170 5176 13176 5188
rect 13228 5216 13234 5228
rect 13630 5216 13636 5228
rect 13228 5188 13636 5216
rect 13228 5176 13234 5188
rect 13630 5176 13636 5188
rect 13688 5176 13694 5228
rect 13998 5176 14004 5228
rect 14056 5216 14062 5228
rect 14737 5219 14795 5225
rect 14737 5216 14749 5219
rect 14056 5188 14749 5216
rect 14056 5176 14062 5188
rect 14737 5185 14749 5188
rect 14783 5185 14795 5219
rect 14737 5179 14795 5185
rect 15562 5176 15568 5228
rect 15620 5216 15626 5228
rect 15749 5219 15807 5225
rect 15749 5216 15761 5219
rect 15620 5188 15761 5216
rect 15620 5176 15626 5188
rect 15749 5185 15761 5188
rect 15795 5185 15807 5219
rect 15749 5179 15807 5185
rect 1762 5108 1768 5160
rect 1820 5148 1826 5160
rect 2041 5151 2099 5157
rect 2041 5148 2053 5151
rect 1820 5120 2053 5148
rect 1820 5108 1826 5120
rect 2041 5117 2053 5120
rect 2087 5117 2099 5151
rect 2041 5111 2099 5117
rect 2308 5151 2366 5157
rect 2308 5117 2320 5151
rect 2354 5148 2366 5151
rect 2590 5148 2596 5160
rect 2354 5120 2596 5148
rect 2354 5117 2366 5120
rect 2308 5111 2366 5117
rect 2590 5108 2596 5120
rect 2648 5108 2654 5160
rect 2866 5108 2872 5160
rect 2924 5148 2930 5160
rect 3510 5148 3516 5160
rect 2924 5120 3516 5148
rect 2924 5108 2930 5120
rect 3510 5108 3516 5120
rect 3568 5108 3574 5160
rect 3697 5151 3755 5157
rect 3697 5117 3709 5151
rect 3743 5148 3755 5151
rect 4154 5148 4160 5160
rect 3743 5120 4160 5148
rect 3743 5117 3755 5120
rect 3697 5111 3755 5117
rect 4154 5108 4160 5120
rect 4212 5108 4218 5160
rect 4617 5151 4675 5157
rect 4617 5117 4629 5151
rect 4663 5148 4675 5151
rect 4706 5148 4712 5160
rect 4663 5120 4712 5148
rect 4663 5117 4675 5120
rect 4617 5111 4675 5117
rect 4706 5108 4712 5120
rect 4764 5108 4770 5160
rect 4884 5151 4942 5157
rect 4884 5117 4896 5151
rect 4930 5148 4942 5151
rect 5902 5148 5908 5160
rect 4930 5120 5908 5148
rect 4930 5117 4942 5120
rect 4884 5111 4942 5117
rect 5902 5108 5908 5120
rect 5960 5108 5966 5160
rect 6822 5148 6828 5160
rect 6783 5120 6828 5148
rect 6822 5108 6828 5120
rect 6880 5108 6886 5160
rect 7092 5151 7150 5157
rect 7092 5117 7104 5151
rect 7138 5148 7150 5151
rect 8846 5148 8852 5160
rect 7138 5120 8852 5148
rect 7138 5117 7150 5120
rect 7092 5111 7150 5117
rect 8846 5108 8852 5120
rect 8904 5108 8910 5160
rect 9214 5108 9220 5160
rect 9272 5148 9278 5160
rect 10321 5151 10379 5157
rect 10321 5148 10333 5151
rect 9272 5120 10333 5148
rect 9272 5108 9278 5120
rect 10321 5117 10333 5120
rect 10367 5117 10379 5151
rect 10321 5111 10379 5117
rect 12897 5151 12955 5157
rect 12897 5117 12909 5151
rect 12943 5148 12955 5151
rect 13262 5148 13268 5160
rect 12943 5120 13268 5148
rect 12943 5117 12955 5120
rect 12897 5111 12955 5117
rect 13262 5108 13268 5120
rect 13320 5108 13326 5160
rect 13538 5148 13544 5160
rect 13499 5120 13544 5148
rect 13538 5108 13544 5120
rect 13596 5108 13602 5160
rect 14182 5108 14188 5160
rect 14240 5148 14246 5160
rect 14458 5148 14464 5160
rect 14240 5120 14464 5148
rect 14240 5108 14246 5120
rect 14458 5108 14464 5120
rect 14516 5148 14522 5160
rect 14553 5151 14611 5157
rect 14553 5148 14565 5151
rect 14516 5120 14565 5148
rect 14516 5108 14522 5120
rect 14553 5117 14565 5120
rect 14599 5117 14611 5151
rect 14553 5111 14611 5117
rect 14645 5151 14703 5157
rect 14645 5117 14657 5151
rect 14691 5148 14703 5151
rect 15102 5148 15108 5160
rect 14691 5120 15108 5148
rect 14691 5117 14703 5120
rect 14645 5111 14703 5117
rect 15102 5108 15108 5120
rect 15160 5148 15166 5160
rect 16850 5148 16856 5160
rect 15160 5120 16856 5148
rect 15160 5108 15166 5120
rect 16850 5108 16856 5120
rect 16908 5108 16914 5160
rect 16960 5157 16988 5256
rect 16945 5151 17003 5157
rect 16945 5117 16957 5151
rect 16991 5117 17003 5151
rect 19794 5148 19800 5160
rect 19755 5120 19800 5148
rect 16945 5111 17003 5117
rect 19794 5108 19800 5120
rect 19852 5108 19858 5160
rect 5810 5040 5816 5092
rect 5868 5080 5874 5092
rect 11146 5080 11152 5092
rect 5868 5052 8892 5080
rect 5868 5040 5874 5052
rect 3418 5012 3424 5024
rect 3379 4984 3424 5012
rect 3418 4972 3424 4984
rect 3476 4972 3482 5024
rect 4890 4972 4896 5024
rect 4948 5012 4954 5024
rect 5534 5012 5540 5024
rect 4948 4984 5540 5012
rect 4948 4972 4954 4984
rect 5534 4972 5540 4984
rect 5592 4972 5598 5024
rect 6914 4972 6920 5024
rect 6972 5012 6978 5024
rect 8864 5021 8892 5052
rect 9876 5052 11152 5080
rect 9876 5021 9904 5052
rect 11146 5040 11152 5052
rect 11204 5040 11210 5092
rect 15470 5040 15476 5092
rect 15528 5080 15534 5092
rect 15565 5083 15623 5089
rect 15565 5080 15577 5083
rect 15528 5052 15577 5080
rect 15528 5040 15534 5052
rect 15565 5049 15577 5052
rect 15611 5049 15623 5083
rect 15565 5043 15623 5049
rect 17221 5083 17279 5089
rect 17221 5049 17233 5083
rect 17267 5080 17279 5083
rect 17862 5080 17868 5092
rect 17267 5052 17868 5080
rect 17267 5049 17279 5052
rect 17221 5043 17279 5049
rect 17862 5040 17868 5052
rect 17920 5040 17926 5092
rect 8205 5015 8263 5021
rect 8205 5012 8217 5015
rect 6972 4984 8217 5012
rect 6972 4972 6978 4984
rect 8205 4981 8217 4984
rect 8251 4981 8263 5015
rect 8205 4975 8263 4981
rect 8849 5015 8907 5021
rect 8849 4981 8861 5015
rect 8895 4981 8907 5015
rect 8849 4975 8907 4981
rect 9861 5015 9919 5021
rect 9861 4981 9873 5015
rect 9907 4981 9919 5015
rect 9861 4975 9919 4981
rect 10134 4972 10140 5024
rect 10192 5012 10198 5024
rect 10229 5015 10287 5021
rect 10229 5012 10241 5015
rect 10192 4984 10241 5012
rect 10192 4972 10198 4984
rect 10229 4981 10241 4984
rect 10275 4981 10287 5015
rect 10229 4975 10287 4981
rect 11054 4972 11060 5024
rect 11112 5012 11118 5024
rect 11701 5015 11759 5021
rect 11701 5012 11713 5015
rect 11112 4984 11713 5012
rect 11112 4972 11118 4984
rect 11701 4981 11713 4984
rect 11747 4981 11759 5015
rect 11701 4975 11759 4981
rect 11790 4972 11796 5024
rect 11848 5012 11854 5024
rect 13725 5015 13783 5021
rect 11848 4984 11893 5012
rect 11848 4972 11854 4984
rect 13725 4981 13737 5015
rect 13771 5012 13783 5015
rect 13998 5012 14004 5024
rect 13771 4984 14004 5012
rect 13771 4981 13783 4984
rect 13725 4975 13783 4981
rect 13998 4972 14004 4984
rect 14056 4972 14062 5024
rect 14182 5012 14188 5024
rect 14143 4984 14188 5012
rect 14182 4972 14188 4984
rect 14240 4972 14246 5024
rect 15102 4972 15108 5024
rect 15160 5012 15166 5024
rect 15657 5015 15715 5021
rect 15657 5012 15669 5015
rect 15160 4984 15669 5012
rect 15160 4972 15166 4984
rect 15657 4981 15669 4984
rect 15703 4981 15715 5015
rect 15657 4975 15715 4981
rect 19981 5015 20039 5021
rect 19981 4981 19993 5015
rect 20027 5012 20039 5015
rect 20622 5012 20628 5024
rect 20027 4984 20628 5012
rect 20027 4981 20039 4984
rect 19981 4975 20039 4981
rect 20622 4972 20628 4984
rect 20680 4972 20686 5024
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 4614 4808 4620 4820
rect 4172 4780 4620 4808
rect 2777 4743 2835 4749
rect 2777 4709 2789 4743
rect 2823 4740 2835 4743
rect 2823 4712 3556 4740
rect 2823 4709 2835 4712
rect 2777 4703 2835 4709
rect 2222 4672 2228 4684
rect 2183 4644 2228 4672
rect 2222 4632 2228 4644
rect 2280 4632 2286 4684
rect 2314 4632 2320 4684
rect 2372 4672 2378 4684
rect 3234 4672 3240 4684
rect 2372 4644 2417 4672
rect 3195 4644 3240 4672
rect 2372 4632 2378 4644
rect 3234 4632 3240 4644
rect 3292 4632 3298 4684
rect 2406 4604 2412 4616
rect 2367 4576 2412 4604
rect 2406 4564 2412 4576
rect 2464 4564 2470 4616
rect 3326 4604 3332 4616
rect 3287 4576 3332 4604
rect 3326 4564 3332 4576
rect 3384 4564 3390 4616
rect 3421 4607 3479 4613
rect 3421 4573 3433 4607
rect 3467 4573 3479 4607
rect 3528 4604 3556 4712
rect 3970 4632 3976 4684
rect 4028 4672 4034 4684
rect 4172 4681 4200 4780
rect 4614 4768 4620 4780
rect 4672 4768 4678 4820
rect 5537 4811 5595 4817
rect 5537 4777 5549 4811
rect 5583 4808 5595 4811
rect 5902 4808 5908 4820
rect 5583 4780 5908 4808
rect 5583 4777 5595 4780
rect 5537 4771 5595 4777
rect 5902 4768 5908 4780
rect 5960 4768 5966 4820
rect 6086 4768 6092 4820
rect 6144 4808 6150 4820
rect 6181 4811 6239 4817
rect 6181 4808 6193 4811
rect 6144 4780 6193 4808
rect 6144 4768 6150 4780
rect 6181 4777 6193 4780
rect 6227 4777 6239 4811
rect 6181 4771 6239 4777
rect 7377 4811 7435 4817
rect 7377 4777 7389 4811
rect 7423 4808 7435 4811
rect 10137 4811 10195 4817
rect 10137 4808 10149 4811
rect 7423 4780 10149 4808
rect 7423 4777 7435 4780
rect 7377 4771 7435 4777
rect 10137 4777 10149 4780
rect 10183 4777 10195 4811
rect 10137 4771 10195 4777
rect 11146 4768 11152 4820
rect 11204 4808 11210 4820
rect 11204 4780 11744 4808
rect 11204 4768 11210 4780
rect 4706 4740 4712 4752
rect 4264 4712 4712 4740
rect 4157 4675 4215 4681
rect 4157 4672 4169 4675
rect 4028 4644 4169 4672
rect 4028 4632 4034 4644
rect 4157 4641 4169 4644
rect 4203 4641 4215 4675
rect 4157 4635 4215 4641
rect 4264 4604 4292 4712
rect 4706 4700 4712 4712
rect 4764 4700 4770 4752
rect 5442 4700 5448 4752
rect 5500 4740 5506 4752
rect 6549 4743 6607 4749
rect 6549 4740 6561 4743
rect 5500 4712 6561 4740
rect 5500 4700 5506 4712
rect 6549 4709 6561 4712
rect 6595 4709 6607 4743
rect 6549 4703 6607 4709
rect 7745 4743 7803 4749
rect 7745 4709 7757 4743
rect 7791 4740 7803 4743
rect 7926 4740 7932 4752
rect 7791 4712 7932 4740
rect 7791 4709 7803 4712
rect 7745 4703 7803 4709
rect 7926 4700 7932 4712
rect 7984 4700 7990 4752
rect 8754 4740 8760 4752
rect 8715 4712 8760 4740
rect 8754 4700 8760 4712
rect 8812 4700 8818 4752
rect 8846 4700 8852 4752
rect 8904 4740 8910 4752
rect 11514 4749 11520 4752
rect 11508 4740 11520 4749
rect 8904 4712 10180 4740
rect 11475 4712 11520 4740
rect 8904 4700 8910 4712
rect 4424 4675 4482 4681
rect 4424 4641 4436 4675
rect 4470 4672 4482 4675
rect 5534 4672 5540 4684
rect 4470 4644 5540 4672
rect 4470 4641 4482 4644
rect 4424 4635 4482 4641
rect 5534 4632 5540 4644
rect 5592 4632 5598 4684
rect 8297 4675 8355 4681
rect 8297 4641 8309 4675
rect 8343 4672 8355 4675
rect 8343 4644 9076 4672
rect 8343 4641 8355 4644
rect 8297 4635 8355 4641
rect 3528 4576 4292 4604
rect 6641 4607 6699 4613
rect 3421 4567 3479 4573
rect 6641 4573 6653 4607
rect 6687 4573 6699 4607
rect 6641 4567 6699 4573
rect 6825 4607 6883 4613
rect 6825 4573 6837 4607
rect 6871 4604 6883 4607
rect 6914 4604 6920 4616
rect 6871 4576 6920 4604
rect 6871 4573 6883 4576
rect 6825 4567 6883 4573
rect 2424 4536 2452 4564
rect 3436 4536 3464 4567
rect 2424 4508 3464 4536
rect 5902 4496 5908 4548
rect 5960 4536 5966 4548
rect 6656 4536 6684 4567
rect 6914 4564 6920 4576
rect 6972 4564 6978 4616
rect 7834 4604 7840 4616
rect 7795 4576 7840 4604
rect 7834 4564 7840 4576
rect 7892 4564 7898 4616
rect 8021 4607 8079 4613
rect 8021 4573 8033 4607
rect 8067 4604 8079 4607
rect 8110 4604 8116 4616
rect 8067 4576 8116 4604
rect 8067 4573 8079 4576
rect 8021 4567 8079 4573
rect 8110 4564 8116 4576
rect 8168 4564 8174 4616
rect 9048 4613 9076 4644
rect 9306 4632 9312 4684
rect 9364 4672 9370 4684
rect 10045 4675 10103 4681
rect 10045 4672 10057 4675
rect 9364 4644 10057 4672
rect 9364 4632 9370 4644
rect 10045 4641 10057 4644
rect 10091 4641 10103 4675
rect 10152 4672 10180 4712
rect 11508 4703 11520 4712
rect 11514 4700 11520 4703
rect 11572 4700 11578 4752
rect 11716 4740 11744 4780
rect 11790 4768 11796 4820
rect 11848 4808 11854 4820
rect 12897 4811 12955 4817
rect 12897 4808 12909 4811
rect 11848 4780 12909 4808
rect 11848 4768 11854 4780
rect 12897 4777 12909 4780
rect 12943 4777 12955 4811
rect 12897 4771 12955 4777
rect 14182 4768 14188 4820
rect 14240 4808 14246 4820
rect 14645 4811 14703 4817
rect 14645 4808 14657 4811
rect 14240 4780 14657 4808
rect 14240 4768 14246 4780
rect 14645 4777 14657 4780
rect 14691 4777 14703 4811
rect 14645 4771 14703 4777
rect 15286 4768 15292 4820
rect 15344 4808 15350 4820
rect 15657 4811 15715 4817
rect 15657 4808 15669 4811
rect 15344 4780 15669 4808
rect 15344 4768 15350 4780
rect 15657 4777 15669 4780
rect 15703 4777 15715 4811
rect 15657 4771 15715 4777
rect 15749 4811 15807 4817
rect 15749 4777 15761 4811
rect 15795 4808 15807 4811
rect 16942 4808 16948 4820
rect 15795 4780 16948 4808
rect 15795 4777 15807 4780
rect 15749 4771 15807 4777
rect 16942 4768 16948 4780
rect 17000 4768 17006 4820
rect 14553 4743 14611 4749
rect 14553 4740 14565 4743
rect 11716 4712 14565 4740
rect 14553 4709 14565 4712
rect 14599 4709 14611 4743
rect 14553 4703 14611 4709
rect 15013 4743 15071 4749
rect 15013 4709 15025 4743
rect 15059 4740 15071 4743
rect 15102 4740 15108 4752
rect 15059 4712 15108 4740
rect 15059 4709 15071 4712
rect 15013 4703 15071 4709
rect 15102 4700 15108 4712
rect 15160 4700 15166 4752
rect 10152 4644 13216 4672
rect 10045 4635 10103 4641
rect 8849 4607 8907 4613
rect 8849 4573 8861 4607
rect 8895 4573 8907 4607
rect 8849 4567 8907 4573
rect 9033 4607 9091 4613
rect 9033 4573 9045 4607
rect 9079 4604 9091 4607
rect 9122 4604 9128 4616
rect 9079 4576 9128 4604
rect 9079 4573 9091 4576
rect 9033 4567 9091 4573
rect 6730 4536 6736 4548
rect 5960 4508 6736 4536
rect 5960 4496 5966 4508
rect 6730 4496 6736 4508
rect 6788 4496 6794 4548
rect 7282 4496 7288 4548
rect 7340 4536 7346 4548
rect 8864 4536 8892 4567
rect 9122 4564 9128 4576
rect 9180 4564 9186 4616
rect 10226 4604 10232 4616
rect 10187 4576 10232 4604
rect 10226 4564 10232 4576
rect 10284 4564 10290 4616
rect 10778 4564 10784 4616
rect 10836 4604 10842 4616
rect 11238 4604 11244 4616
rect 10836 4576 11244 4604
rect 10836 4564 10842 4576
rect 11238 4564 11244 4576
rect 11296 4564 11302 4616
rect 12618 4536 12624 4548
rect 7340 4508 8892 4536
rect 12579 4508 12624 4536
rect 7340 4496 7346 4508
rect 12618 4496 12624 4508
rect 12676 4496 12682 4548
rect 13188 4536 13216 4644
rect 13262 4632 13268 4684
rect 13320 4672 13326 4684
rect 17862 4672 17868 4684
rect 13320 4644 15976 4672
rect 17823 4644 17868 4672
rect 13320 4632 13326 4644
rect 13354 4604 13360 4616
rect 13315 4576 13360 4604
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 13541 4607 13599 4613
rect 13541 4573 13553 4607
rect 13587 4604 13599 4607
rect 13630 4604 13636 4616
rect 13587 4576 13636 4604
rect 13587 4573 13599 4576
rect 13541 4567 13599 4573
rect 13630 4564 13636 4576
rect 13688 4564 13694 4616
rect 14829 4607 14887 4613
rect 14829 4573 14841 4607
rect 14875 4604 14887 4607
rect 15010 4604 15016 4616
rect 14875 4576 15016 4604
rect 14875 4573 14887 4576
rect 14829 4567 14887 4573
rect 15010 4564 15016 4576
rect 15068 4564 15074 4616
rect 15841 4607 15899 4613
rect 15841 4573 15853 4607
rect 15887 4573 15899 4607
rect 15948 4604 15976 4644
rect 17862 4632 17868 4644
rect 17920 4632 17926 4684
rect 19334 4604 19340 4616
rect 15948 4576 19340 4604
rect 15841 4567 15899 4573
rect 15856 4536 15884 4567
rect 19334 4564 19340 4576
rect 19392 4564 19398 4616
rect 13188 4508 15884 4536
rect 1857 4471 1915 4477
rect 1857 4437 1869 4471
rect 1903 4468 1915 4471
rect 2777 4471 2835 4477
rect 2777 4468 2789 4471
rect 1903 4440 2789 4468
rect 1903 4437 1915 4440
rect 1857 4431 1915 4437
rect 2777 4437 2789 4440
rect 2823 4437 2835 4471
rect 2777 4431 2835 4437
rect 2869 4471 2927 4477
rect 2869 4437 2881 4471
rect 2915 4468 2927 4471
rect 5074 4468 5080 4480
rect 2915 4440 5080 4468
rect 2915 4437 2927 4440
rect 2869 4431 2927 4437
rect 5074 4428 5080 4440
rect 5132 4428 5138 4480
rect 5534 4428 5540 4480
rect 5592 4468 5598 4480
rect 8205 4471 8263 4477
rect 8205 4468 8217 4471
rect 5592 4440 8217 4468
rect 5592 4428 5598 4440
rect 8205 4437 8217 4440
rect 8251 4437 8263 4471
rect 8386 4468 8392 4480
rect 8347 4440 8392 4468
rect 8205 4431 8263 4437
rect 8386 4428 8392 4440
rect 8444 4428 8450 4480
rect 9677 4471 9735 4477
rect 9677 4437 9689 4471
rect 9723 4468 9735 4471
rect 11146 4468 11152 4480
rect 9723 4440 11152 4468
rect 9723 4437 9735 4440
rect 9677 4431 9735 4437
rect 11146 4428 11152 4440
rect 11204 4428 11210 4480
rect 14185 4471 14243 4477
rect 14185 4437 14197 4471
rect 14231 4468 14243 4471
rect 15013 4471 15071 4477
rect 15013 4468 15025 4471
rect 14231 4440 15025 4468
rect 14231 4437 14243 4440
rect 14185 4431 14243 4437
rect 15013 4437 15025 4440
rect 15059 4437 15071 4471
rect 15013 4431 15071 4437
rect 15102 4428 15108 4480
rect 15160 4468 15166 4480
rect 15289 4471 15347 4477
rect 15289 4468 15301 4471
rect 15160 4440 15301 4468
rect 15160 4428 15166 4440
rect 15289 4437 15301 4440
rect 15335 4437 15347 4471
rect 15289 4431 15347 4437
rect 18049 4471 18107 4477
rect 18049 4437 18061 4471
rect 18095 4468 18107 4471
rect 18782 4468 18788 4480
rect 18095 4440 18788 4468
rect 18095 4437 18107 4440
rect 18049 4431 18107 4437
rect 18782 4428 18788 4440
rect 18840 4428 18846 4480
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 2406 4224 2412 4276
rect 2464 4264 2470 4276
rect 3145 4267 3203 4273
rect 3145 4264 3157 4267
rect 2464 4236 3157 4264
rect 2464 4224 2470 4236
rect 3145 4233 3157 4236
rect 3191 4233 3203 4267
rect 3145 4227 3203 4233
rect 5629 4267 5687 4273
rect 5629 4233 5641 4267
rect 5675 4264 5687 4267
rect 5718 4264 5724 4276
rect 5675 4236 5724 4264
rect 5675 4233 5687 4236
rect 5629 4227 5687 4233
rect 5718 4224 5724 4236
rect 5776 4224 5782 4276
rect 7101 4267 7159 4273
rect 7101 4233 7113 4267
rect 7147 4264 7159 4267
rect 7834 4264 7840 4276
rect 7147 4236 7840 4264
rect 7147 4233 7159 4236
rect 7101 4227 7159 4233
rect 7834 4224 7840 4236
rect 7892 4224 7898 4276
rect 7926 4224 7932 4276
rect 7984 4264 7990 4276
rect 8113 4267 8171 4273
rect 8113 4264 8125 4267
rect 7984 4236 8125 4264
rect 7984 4224 7990 4236
rect 8113 4233 8125 4236
rect 8159 4233 8171 4267
rect 9306 4264 9312 4276
rect 9267 4236 9312 4264
rect 8113 4227 8171 4233
rect 9306 4224 9312 4236
rect 9364 4224 9370 4276
rect 9950 4224 9956 4276
rect 10008 4264 10014 4276
rect 10962 4264 10968 4276
rect 10008 4236 10968 4264
rect 10008 4224 10014 4236
rect 10962 4224 10968 4236
rect 11020 4264 11026 4276
rect 13170 4264 13176 4276
rect 11020 4236 13176 4264
rect 11020 4224 11026 4236
rect 13170 4224 13176 4236
rect 13228 4224 13234 4276
rect 4798 4196 4804 4208
rect 4711 4168 4804 4196
rect 4798 4156 4804 4168
rect 4856 4196 4862 4208
rect 4856 4168 6316 4196
rect 4856 4156 4862 4168
rect 5718 4128 5724 4140
rect 4724 4100 5724 4128
rect 1762 4060 1768 4072
rect 1675 4032 1768 4060
rect 1762 4020 1768 4032
rect 1820 4060 1826 4072
rect 3421 4063 3479 4069
rect 3421 4060 3433 4063
rect 1820 4032 3433 4060
rect 1820 4020 1826 4032
rect 3421 4029 3433 4032
rect 3467 4060 3479 4063
rect 3970 4060 3976 4072
rect 3467 4032 3976 4060
rect 3467 4029 3479 4032
rect 3421 4023 3479 4029
rect 3970 4020 3976 4032
rect 4028 4020 4034 4072
rect 2032 3995 2090 4001
rect 2032 3961 2044 3995
rect 2078 3992 2090 3995
rect 2130 3992 2136 4004
rect 2078 3964 2136 3992
rect 2078 3961 2090 3964
rect 2032 3955 2090 3961
rect 2130 3952 2136 3964
rect 2188 3952 2194 4004
rect 3602 3952 3608 4004
rect 3660 4001 3666 4004
rect 3660 3995 3724 4001
rect 3660 3961 3678 3995
rect 3712 3961 3724 3995
rect 3660 3955 3724 3961
rect 3660 3952 3666 3955
rect 3786 3952 3792 4004
rect 3844 3992 3850 4004
rect 4724 3992 4752 4100
rect 5718 4088 5724 4100
rect 5776 4088 5782 4140
rect 6288 4137 6316 4168
rect 6914 4156 6920 4208
rect 6972 4196 6978 4208
rect 8202 4196 8208 4208
rect 6972 4168 8208 4196
rect 6972 4156 6978 4168
rect 8202 4156 8208 4168
rect 8260 4156 8266 4208
rect 11606 4196 11612 4208
rect 11532 4168 11612 4196
rect 6273 4131 6331 4137
rect 6273 4097 6285 4131
rect 6319 4128 6331 4131
rect 6362 4128 6368 4140
rect 6319 4100 6368 4128
rect 6319 4097 6331 4100
rect 6273 4091 6331 4097
rect 6362 4088 6368 4100
rect 6420 4088 6426 4140
rect 7650 4128 7656 4140
rect 7611 4100 7656 4128
rect 7650 4088 7656 4100
rect 7708 4088 7714 4140
rect 8662 4128 8668 4140
rect 8623 4100 8668 4128
rect 8662 4088 8668 4100
rect 8720 4088 8726 4140
rect 9766 4128 9772 4140
rect 9727 4100 9772 4128
rect 9766 4088 9772 4100
rect 9824 4088 9830 4140
rect 9858 4088 9864 4140
rect 9916 4088 9922 4140
rect 9953 4131 10011 4137
rect 9953 4097 9965 4131
rect 9999 4128 10011 4131
rect 10502 4128 10508 4140
rect 9999 4100 10508 4128
rect 9999 4097 10011 4100
rect 9953 4091 10011 4097
rect 10502 4088 10508 4100
rect 10560 4088 10566 4140
rect 11532 4137 11560 4168
rect 11606 4156 11612 4168
rect 11664 4156 11670 4208
rect 13722 4156 13728 4208
rect 13780 4196 13786 4208
rect 13780 4168 14688 4196
rect 13780 4156 13786 4168
rect 11517 4131 11575 4137
rect 11517 4097 11529 4131
rect 11563 4097 11575 4131
rect 11517 4091 11575 4097
rect 13906 4088 13912 4140
rect 13964 4128 13970 4140
rect 14660 4137 14688 4168
rect 14645 4131 14703 4137
rect 13964 4100 14596 4128
rect 13964 4088 13970 4100
rect 5994 4060 6000 4072
rect 3844 3964 4752 3992
rect 4816 4032 6000 4060
rect 3844 3952 3850 3964
rect 2958 3884 2964 3936
rect 3016 3924 3022 3936
rect 4816 3924 4844 4032
rect 5994 4020 6000 4032
rect 6052 4020 6058 4072
rect 6089 4063 6147 4069
rect 6089 4029 6101 4063
rect 6135 4060 6147 4063
rect 6638 4060 6644 4072
rect 6135 4032 6644 4060
rect 6135 4029 6147 4032
rect 6089 4023 6147 4029
rect 6638 4020 6644 4032
rect 6696 4060 6702 4072
rect 9876 4060 9904 4088
rect 6696 4032 9904 4060
rect 10321 4063 10379 4069
rect 6696 4020 6702 4032
rect 10321 4029 10333 4063
rect 10367 4060 10379 4063
rect 12066 4060 12072 4072
rect 10367 4032 12072 4060
rect 10367 4029 10379 4032
rect 10321 4023 10379 4029
rect 12066 4020 12072 4032
rect 12124 4020 12130 4072
rect 12342 4020 12348 4072
rect 12400 4060 12406 4072
rect 12437 4063 12495 4069
rect 12437 4060 12449 4063
rect 12400 4032 12449 4060
rect 12400 4020 12406 4032
rect 12437 4029 12449 4032
rect 12483 4029 12495 4063
rect 12437 4023 12495 4029
rect 13170 4020 13176 4072
rect 13228 4060 13234 4072
rect 14461 4063 14519 4069
rect 14461 4060 14473 4063
rect 13228 4032 14473 4060
rect 13228 4020 13234 4032
rect 14461 4029 14473 4032
rect 14507 4029 14519 4063
rect 14568 4060 14596 4100
rect 14645 4097 14657 4131
rect 14691 4097 14703 4131
rect 14645 4091 14703 4097
rect 19334 4088 19340 4140
rect 19392 4128 19398 4140
rect 22462 4128 22468 4140
rect 19392 4100 22468 4128
rect 19392 4088 19398 4100
rect 22462 4088 22468 4100
rect 22520 4088 22526 4140
rect 15105 4063 15163 4069
rect 15105 4060 15117 4063
rect 14568 4032 15117 4060
rect 14461 4023 14519 4029
rect 15105 4029 15117 4032
rect 15151 4029 15163 4063
rect 15105 4023 15163 4029
rect 4982 3952 4988 4004
rect 5040 3992 5046 4004
rect 7561 3995 7619 4001
rect 7561 3992 7573 3995
rect 5040 3964 7573 3992
rect 5040 3952 5046 3964
rect 7561 3961 7573 3964
rect 7607 3992 7619 3995
rect 10134 3992 10140 4004
rect 7607 3964 10140 3992
rect 7607 3961 7619 3964
rect 7561 3955 7619 3961
rect 10134 3952 10140 3964
rect 10192 3952 10198 4004
rect 12526 3992 12532 4004
rect 10520 3964 12532 3992
rect 5166 3924 5172 3936
rect 3016 3896 4844 3924
rect 5127 3896 5172 3924
rect 3016 3884 3022 3896
rect 5166 3884 5172 3896
rect 5224 3884 5230 3936
rect 5258 3884 5264 3936
rect 5316 3924 5322 3936
rect 5997 3927 6055 3933
rect 5997 3924 6009 3927
rect 5316 3896 6009 3924
rect 5316 3884 5322 3896
rect 5997 3893 6009 3896
rect 6043 3893 6055 3927
rect 5997 3887 6055 3893
rect 6086 3884 6092 3936
rect 6144 3924 6150 3936
rect 7469 3927 7527 3933
rect 7469 3924 7481 3927
rect 6144 3896 7481 3924
rect 6144 3884 6150 3896
rect 7469 3893 7481 3896
rect 7515 3893 7527 3927
rect 8478 3924 8484 3936
rect 8439 3896 8484 3924
rect 7469 3887 7527 3893
rect 8478 3884 8484 3896
rect 8536 3884 8542 3936
rect 8570 3884 8576 3936
rect 8628 3924 8634 3936
rect 9674 3924 9680 3936
rect 8628 3896 8673 3924
rect 9635 3896 9680 3924
rect 8628 3884 8634 3896
rect 9674 3884 9680 3896
rect 9732 3884 9738 3936
rect 10520 3933 10548 3964
rect 12526 3952 12532 3964
rect 12584 3952 12590 4004
rect 12704 3995 12762 4001
rect 12704 3961 12716 3995
rect 12750 3992 12762 3995
rect 12894 3992 12900 4004
rect 12750 3964 12900 3992
rect 12750 3961 12762 3964
rect 12704 3955 12762 3961
rect 12894 3952 12900 3964
rect 12952 3952 12958 4004
rect 14553 3995 14611 4001
rect 14553 3992 14565 3995
rect 13004 3964 14565 3992
rect 10505 3927 10563 3933
rect 10505 3893 10517 3927
rect 10551 3893 10563 3927
rect 10505 3887 10563 3893
rect 10873 3927 10931 3933
rect 10873 3893 10885 3927
rect 10919 3924 10931 3927
rect 11054 3924 11060 3936
rect 10919 3896 11060 3924
rect 10919 3893 10931 3896
rect 10873 3887 10931 3893
rect 11054 3884 11060 3896
rect 11112 3884 11118 3936
rect 11238 3924 11244 3936
rect 11199 3896 11244 3924
rect 11238 3884 11244 3896
rect 11296 3884 11302 3936
rect 11330 3884 11336 3936
rect 11388 3924 11394 3936
rect 13004 3924 13032 3964
rect 14553 3961 14565 3964
rect 14599 3961 14611 3995
rect 14553 3955 14611 3961
rect 14642 3952 14648 4004
rect 14700 3992 14706 4004
rect 14700 3964 15332 3992
rect 14700 3952 14706 3964
rect 11388 3896 13032 3924
rect 11388 3884 11394 3896
rect 13630 3884 13636 3936
rect 13688 3924 13694 3936
rect 13817 3927 13875 3933
rect 13817 3924 13829 3927
rect 13688 3896 13829 3924
rect 13688 3884 13694 3896
rect 13817 3893 13829 3896
rect 13863 3893 13875 3927
rect 14090 3924 14096 3936
rect 14051 3896 14096 3924
rect 13817 3887 13875 3893
rect 14090 3884 14096 3896
rect 14148 3884 14154 3936
rect 15304 3933 15332 3964
rect 15289 3927 15347 3933
rect 15289 3893 15301 3927
rect 15335 3893 15347 3927
rect 15289 3887 15347 3893
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 2498 3680 2504 3732
rect 2556 3720 2562 3732
rect 4614 3720 4620 3732
rect 2556 3692 4620 3720
rect 2556 3680 2562 3692
rect 4614 3680 4620 3692
rect 4672 3680 4678 3732
rect 5166 3680 5172 3732
rect 5224 3720 5230 3732
rect 6181 3723 6239 3729
rect 6181 3720 6193 3723
rect 5224 3692 6193 3720
rect 5224 3680 5230 3692
rect 6181 3689 6193 3692
rect 6227 3689 6239 3723
rect 6181 3683 6239 3689
rect 6730 3680 6736 3732
rect 6788 3720 6794 3732
rect 8938 3720 8944 3732
rect 6788 3692 8944 3720
rect 6788 3680 6794 3692
rect 8938 3680 8944 3692
rect 8996 3680 9002 3732
rect 9125 3723 9183 3729
rect 9125 3689 9137 3723
rect 9171 3720 9183 3723
rect 9674 3720 9680 3732
rect 9171 3692 9680 3720
rect 9171 3689 9183 3692
rect 9125 3683 9183 3689
rect 9674 3680 9680 3692
rect 9732 3680 9738 3732
rect 11241 3723 11299 3729
rect 10060 3692 11192 3720
rect 2032 3655 2090 3661
rect 2032 3621 2044 3655
rect 2078 3652 2090 3655
rect 2406 3652 2412 3664
rect 2078 3624 2412 3652
rect 2078 3621 2090 3624
rect 2032 3615 2090 3621
rect 2406 3612 2412 3624
rect 2464 3612 2470 3664
rect 2590 3612 2596 3664
rect 2648 3652 2654 3664
rect 3142 3652 3148 3664
rect 2648 3624 3148 3652
rect 2648 3612 2654 3624
rect 3142 3612 3148 3624
rect 3200 3612 3206 3664
rect 4424 3655 4482 3661
rect 4424 3621 4436 3655
rect 4470 3652 4482 3655
rect 4798 3652 4804 3664
rect 4470 3624 4804 3652
rect 4470 3621 4482 3624
rect 4424 3615 4482 3621
rect 4798 3612 4804 3624
rect 4856 3612 4862 3664
rect 4890 3612 4896 3664
rect 4948 3652 4954 3664
rect 8570 3652 8576 3664
rect 4948 3624 8576 3652
rect 4948 3612 4954 3624
rect 8570 3612 8576 3624
rect 8628 3652 8634 3664
rect 10060 3652 10088 3692
rect 8628 3624 10088 3652
rect 10128 3655 10186 3661
rect 8628 3612 8634 3624
rect 10128 3621 10140 3655
rect 10174 3652 10186 3655
rect 10226 3652 10232 3664
rect 10174 3624 10232 3652
rect 10174 3621 10186 3624
rect 10128 3615 10186 3621
rect 10226 3612 10232 3624
rect 10284 3612 10290 3664
rect 1578 3544 1584 3596
rect 1636 3584 1642 3596
rect 7006 3584 7012 3596
rect 1636 3556 7012 3584
rect 1636 3544 1642 3556
rect 7006 3544 7012 3556
rect 7064 3544 7070 3596
rect 7368 3587 7426 3593
rect 7368 3553 7380 3587
rect 7414 3584 7426 3587
rect 7650 3584 7656 3596
rect 7414 3556 7656 3584
rect 7414 3553 7426 3556
rect 7368 3547 7426 3553
rect 7650 3544 7656 3556
rect 7708 3584 7714 3596
rect 7926 3584 7932 3596
rect 7708 3556 7932 3584
rect 7708 3544 7714 3556
rect 7926 3544 7932 3556
rect 7984 3544 7990 3596
rect 8478 3544 8484 3596
rect 8536 3584 8542 3596
rect 11164 3584 11192 3692
rect 11241 3689 11253 3723
rect 11287 3689 11299 3723
rect 11241 3683 11299 3689
rect 11256 3652 11284 3683
rect 11514 3680 11520 3732
rect 11572 3720 11578 3732
rect 12342 3720 12348 3732
rect 11572 3692 12348 3720
rect 11572 3680 11578 3692
rect 12342 3680 12348 3692
rect 12400 3680 12406 3732
rect 12894 3720 12900 3732
rect 12855 3692 12900 3720
rect 12894 3680 12900 3692
rect 12952 3720 12958 3732
rect 13173 3723 13231 3729
rect 12952 3692 13124 3720
rect 12952 3680 12958 3692
rect 11606 3652 11612 3664
rect 11256 3624 11612 3652
rect 11606 3612 11612 3624
rect 11664 3652 11670 3664
rect 11762 3655 11820 3661
rect 11762 3652 11774 3655
rect 11664 3624 11774 3652
rect 11664 3612 11670 3624
rect 11762 3621 11774 3624
rect 11808 3621 11820 3655
rect 11762 3615 11820 3621
rect 11974 3612 11980 3664
rect 12032 3652 12038 3664
rect 13096 3652 13124 3692
rect 13173 3689 13185 3723
rect 13219 3720 13231 3723
rect 13354 3720 13360 3732
rect 13219 3692 13360 3720
rect 13219 3689 13231 3692
rect 13173 3683 13231 3689
rect 13354 3680 13360 3692
rect 13412 3680 13418 3732
rect 13630 3680 13636 3732
rect 13688 3720 13694 3732
rect 16209 3723 16267 3729
rect 16209 3720 16221 3723
rect 13688 3692 16221 3720
rect 13688 3680 13694 3692
rect 16209 3689 16221 3692
rect 16255 3689 16267 3723
rect 16209 3683 16267 3689
rect 12032 3624 13032 3652
rect 13096 3624 13676 3652
rect 12032 3612 12038 3624
rect 11238 3584 11244 3596
rect 8536 3556 11008 3584
rect 11164 3556 11244 3584
rect 8536 3544 8542 3556
rect 1762 3516 1768 3528
rect 1723 3488 1768 3516
rect 1762 3476 1768 3488
rect 1820 3476 1826 3528
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3485 3479 3519
rect 3421 3479 3479 3485
rect 3436 3448 3464 3479
rect 3970 3476 3976 3528
rect 4028 3516 4034 3528
rect 4157 3519 4215 3525
rect 4157 3516 4169 3519
rect 4028 3488 4169 3516
rect 4028 3476 4034 3488
rect 4157 3485 4169 3488
rect 4203 3485 4215 3519
rect 4157 3479 4215 3485
rect 5718 3476 5724 3528
rect 5776 3516 5782 3528
rect 6273 3519 6331 3525
rect 6273 3516 6285 3519
rect 5776 3488 6285 3516
rect 5776 3476 5782 3488
rect 6273 3485 6285 3488
rect 6319 3485 6331 3519
rect 6273 3479 6331 3485
rect 6362 3476 6368 3528
rect 6420 3516 6426 3528
rect 6420 3488 6465 3516
rect 6420 3476 6426 3488
rect 6822 3476 6828 3528
rect 6880 3516 6886 3528
rect 7101 3519 7159 3525
rect 7101 3516 7113 3519
rect 6880 3488 7113 3516
rect 6880 3476 6886 3488
rect 7101 3485 7113 3488
rect 7147 3485 7159 3519
rect 7101 3479 7159 3485
rect 8202 3476 8208 3528
rect 8260 3516 8266 3528
rect 9766 3516 9772 3528
rect 8260 3488 9772 3516
rect 8260 3476 8266 3488
rect 9766 3476 9772 3488
rect 9824 3516 9830 3528
rect 9861 3519 9919 3525
rect 9861 3516 9873 3519
rect 9824 3488 9873 3516
rect 9824 3476 9830 3488
rect 9861 3485 9873 3488
rect 9907 3485 9919 3519
rect 9861 3479 9919 3485
rect 5534 3448 5540 3460
rect 2700 3420 3464 3448
rect 5495 3420 5540 3448
rect 2038 3340 2044 3392
rect 2096 3380 2102 3392
rect 2700 3380 2728 3420
rect 5534 3408 5540 3420
rect 5592 3408 5598 3460
rect 5810 3448 5816 3460
rect 5771 3420 5816 3448
rect 5810 3408 5816 3420
rect 5868 3408 5874 3460
rect 8220 3448 8248 3476
rect 8036 3420 8248 3448
rect 10980 3448 11008 3556
rect 11238 3544 11244 3556
rect 11296 3584 11302 3596
rect 12802 3584 12808 3596
rect 11296 3556 12808 3584
rect 11296 3544 11302 3556
rect 12802 3544 12808 3556
rect 12860 3544 12866 3596
rect 13004 3584 13032 3624
rect 13081 3587 13139 3593
rect 13081 3584 13093 3587
rect 12991 3556 13093 3584
rect 13081 3553 13093 3556
rect 13127 3584 13139 3587
rect 13541 3587 13599 3593
rect 13541 3584 13553 3587
rect 13127 3556 13553 3584
rect 13127 3553 13139 3556
rect 13081 3547 13139 3553
rect 13541 3553 13553 3556
rect 13587 3553 13599 3587
rect 13648 3584 13676 3624
rect 13722 3612 13728 3664
rect 13780 3652 13786 3664
rect 13780 3624 14228 3652
rect 13780 3612 13786 3624
rect 14200 3593 14228 3624
rect 14185 3587 14243 3593
rect 13648 3556 13768 3584
rect 13541 3547 13599 3553
rect 11514 3476 11520 3528
rect 11572 3516 11578 3528
rect 11572 3488 11617 3516
rect 11572 3476 11578 3488
rect 12526 3476 12532 3528
rect 12584 3516 12590 3528
rect 13170 3516 13176 3528
rect 12584 3488 13176 3516
rect 12584 3476 12590 3488
rect 13170 3476 13176 3488
rect 13228 3476 13234 3528
rect 13354 3476 13360 3528
rect 13412 3516 13418 3528
rect 13740 3525 13768 3556
rect 14185 3553 14197 3587
rect 14231 3553 14243 3587
rect 14185 3547 14243 3553
rect 14366 3544 14372 3596
rect 14424 3584 14430 3596
rect 15289 3587 15347 3593
rect 15289 3584 15301 3587
rect 14424 3556 15301 3584
rect 14424 3544 14430 3556
rect 15289 3553 15301 3556
rect 15335 3553 15347 3587
rect 16022 3584 16028 3596
rect 15983 3556 16028 3584
rect 15289 3547 15347 3553
rect 16022 3544 16028 3556
rect 16080 3544 16086 3596
rect 13633 3519 13691 3525
rect 13633 3516 13645 3519
rect 13412 3488 13645 3516
rect 13412 3476 13418 3488
rect 13633 3485 13645 3488
rect 13679 3485 13691 3519
rect 13633 3479 13691 3485
rect 13725 3519 13783 3525
rect 13725 3485 13737 3519
rect 13771 3485 13783 3519
rect 13725 3479 13783 3485
rect 15565 3519 15623 3525
rect 15565 3485 15577 3519
rect 15611 3516 15623 3519
rect 16114 3516 16120 3528
rect 15611 3488 16120 3516
rect 15611 3485 15623 3488
rect 15565 3479 15623 3485
rect 16114 3476 16120 3488
rect 16172 3476 16178 3528
rect 11330 3448 11336 3460
rect 10980 3420 11336 3448
rect 2096 3352 2728 3380
rect 3145 3383 3203 3389
rect 2096 3340 2102 3352
rect 3145 3349 3157 3383
rect 3191 3380 3203 3383
rect 3602 3380 3608 3392
rect 3191 3352 3608 3380
rect 3191 3349 3203 3352
rect 3145 3343 3203 3349
rect 3602 3340 3608 3352
rect 3660 3380 3666 3392
rect 5258 3380 5264 3392
rect 3660 3352 5264 3380
rect 3660 3340 3666 3352
rect 5258 3340 5264 3352
rect 5316 3340 5322 3392
rect 5718 3340 5724 3392
rect 5776 3380 5782 3392
rect 6546 3380 6552 3392
rect 5776 3352 6552 3380
rect 5776 3340 5782 3352
rect 6546 3340 6552 3352
rect 6604 3340 6610 3392
rect 7466 3340 7472 3392
rect 7524 3380 7530 3392
rect 8036 3380 8064 3420
rect 11330 3408 11336 3420
rect 11388 3408 11394 3460
rect 7524 3352 8064 3380
rect 7524 3340 7530 3352
rect 8110 3340 8116 3392
rect 8168 3380 8174 3392
rect 8481 3383 8539 3389
rect 8481 3380 8493 3383
rect 8168 3352 8493 3380
rect 8168 3340 8174 3352
rect 8481 3349 8493 3352
rect 8527 3380 8539 3383
rect 10502 3380 10508 3392
rect 8527 3352 10508 3380
rect 8527 3349 8539 3352
rect 8481 3343 8539 3349
rect 10502 3340 10508 3352
rect 10560 3340 10566 3392
rect 13081 3383 13139 3389
rect 13081 3349 13093 3383
rect 13127 3380 13139 3383
rect 13906 3380 13912 3392
rect 13127 3352 13912 3380
rect 13127 3349 13139 3352
rect 13081 3343 13139 3349
rect 13906 3340 13912 3352
rect 13964 3340 13970 3392
rect 14369 3383 14427 3389
rect 14369 3349 14381 3383
rect 14415 3380 14427 3383
rect 15010 3380 15016 3392
rect 14415 3352 15016 3380
rect 14415 3349 14427 3352
rect 14369 3343 14427 3349
rect 15010 3340 15016 3352
rect 15068 3340 15074 3392
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 1673 3179 1731 3185
rect 1673 3145 1685 3179
rect 1719 3176 1731 3179
rect 2222 3176 2228 3188
rect 1719 3148 2228 3176
rect 1719 3145 1731 3148
rect 1673 3139 1731 3145
rect 2222 3136 2228 3148
rect 2280 3136 2286 3188
rect 2501 3179 2559 3185
rect 2501 3145 2513 3179
rect 2547 3176 2559 3179
rect 2590 3176 2596 3188
rect 2547 3148 2596 3176
rect 2547 3145 2559 3148
rect 2501 3139 2559 3145
rect 2590 3136 2596 3148
rect 2648 3136 2654 3188
rect 2685 3179 2743 3185
rect 2685 3145 2697 3179
rect 2731 3176 2743 3179
rect 3234 3176 3240 3188
rect 2731 3148 3240 3176
rect 2731 3145 2743 3148
rect 2685 3139 2743 3145
rect 3234 3136 3240 3148
rect 3292 3136 3298 3188
rect 3326 3136 3332 3188
rect 3384 3176 3390 3188
rect 3697 3179 3755 3185
rect 3697 3176 3709 3179
rect 3384 3148 3709 3176
rect 3384 3136 3390 3148
rect 3697 3145 3709 3148
rect 3743 3145 3755 3179
rect 3697 3139 3755 3145
rect 4154 3136 4160 3188
rect 4212 3176 4218 3188
rect 4709 3179 4767 3185
rect 4709 3176 4721 3179
rect 4212 3148 4721 3176
rect 4212 3136 4218 3148
rect 4709 3145 4721 3148
rect 4755 3145 4767 3179
rect 5350 3176 5356 3188
rect 4709 3139 4767 3145
rect 4908 3148 5356 3176
rect 4908 3108 4936 3148
rect 5350 3136 5356 3148
rect 5408 3136 5414 3188
rect 5721 3179 5779 3185
rect 5721 3145 5733 3179
rect 5767 3176 5779 3179
rect 8386 3176 8392 3188
rect 5767 3148 8392 3176
rect 5767 3145 5779 3148
rect 5721 3139 5779 3145
rect 8386 3136 8392 3148
rect 8444 3136 8450 3188
rect 8938 3136 8944 3188
rect 8996 3176 9002 3188
rect 8996 3148 9260 3176
rect 8996 3136 9002 3148
rect 6178 3108 6184 3120
rect 4264 3080 4936 3108
rect 5092 3080 6184 3108
rect 2130 3000 2136 3052
rect 2188 3040 2194 3052
rect 2317 3043 2375 3049
rect 2317 3040 2329 3043
rect 2188 3012 2329 3040
rect 2188 3000 2194 3012
rect 2317 3009 2329 3012
rect 2363 3040 2375 3043
rect 3329 3043 3387 3049
rect 3329 3040 3341 3043
rect 2363 3012 3341 3040
rect 2363 3009 2375 3012
rect 2317 3003 2375 3009
rect 3329 3009 3341 3012
rect 3375 3040 3387 3043
rect 3418 3040 3424 3052
rect 3375 3012 3424 3040
rect 3375 3009 3387 3012
rect 3329 3003 3387 3009
rect 3418 3000 3424 3012
rect 3476 3000 3482 3052
rect 4157 3043 4215 3049
rect 4157 3009 4169 3043
rect 4203 3040 4215 3043
rect 4264 3040 4292 3080
rect 4203 3012 4292 3040
rect 4203 3009 4215 3012
rect 4157 3003 4215 3009
rect 4338 3000 4344 3052
rect 4396 3040 4402 3052
rect 5092 3040 5120 3080
rect 6178 3068 6184 3080
rect 6236 3068 6242 3120
rect 7558 3068 7564 3120
rect 7616 3108 7622 3120
rect 7616 3080 8064 3108
rect 7616 3068 7622 3080
rect 5258 3040 5264 3052
rect 4396 3012 4441 3040
rect 5000 3012 5120 3040
rect 5219 3012 5264 3040
rect 4396 3000 4402 3012
rect 2038 2972 2044 2984
rect 1999 2944 2044 2972
rect 2038 2932 2044 2944
rect 2096 2932 2102 2984
rect 3145 2975 3203 2981
rect 3145 2941 3157 2975
rect 3191 2972 3203 2975
rect 5000 2972 5028 3012
rect 5258 3000 5264 3012
rect 5316 3000 5322 3052
rect 5718 3000 5724 3052
rect 5776 3040 5782 3052
rect 6270 3040 6276 3052
rect 5776 3012 6276 3040
rect 5776 3000 5782 3012
rect 6270 3000 6276 3012
rect 6328 3000 6334 3052
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3040 6423 3043
rect 7745 3043 7803 3049
rect 6411 3012 7696 3040
rect 6411 3009 6423 3012
rect 6365 3003 6423 3009
rect 3191 2944 5028 2972
rect 3191 2941 3203 2944
rect 3145 2935 3203 2941
rect 5074 2932 5080 2984
rect 5132 2972 5138 2984
rect 5169 2975 5227 2981
rect 5169 2972 5181 2975
rect 5132 2944 5181 2972
rect 5132 2932 5138 2944
rect 5169 2941 5181 2944
rect 5215 2941 5227 2975
rect 7466 2972 7472 2984
rect 7427 2944 7472 2972
rect 5169 2935 5227 2941
rect 7466 2932 7472 2944
rect 7524 2932 7530 2984
rect 198 2864 204 2916
rect 256 2904 262 2916
rect 1946 2904 1952 2916
rect 256 2876 1952 2904
rect 256 2864 262 2876
rect 1946 2864 1952 2876
rect 2004 2864 2010 2916
rect 2133 2907 2191 2913
rect 2133 2873 2145 2907
rect 2179 2904 2191 2907
rect 2501 2907 2559 2913
rect 2501 2904 2513 2907
rect 2179 2876 2513 2904
rect 2179 2873 2191 2876
rect 2133 2867 2191 2873
rect 2501 2873 2513 2876
rect 2547 2873 2559 2907
rect 2501 2867 2559 2873
rect 4065 2907 4123 2913
rect 4065 2873 4077 2907
rect 4111 2904 4123 2907
rect 4246 2904 4252 2916
rect 4111 2876 4252 2904
rect 4111 2873 4123 2876
rect 4065 2867 4123 2873
rect 4246 2864 4252 2876
rect 4304 2864 4310 2916
rect 5902 2904 5908 2916
rect 4632 2876 5908 2904
rect 2866 2796 2872 2848
rect 2924 2836 2930 2848
rect 3050 2836 3056 2848
rect 2924 2808 3056 2836
rect 2924 2796 2930 2808
rect 3050 2796 3056 2808
rect 3108 2796 3114 2848
rect 3142 2796 3148 2848
rect 3200 2836 3206 2848
rect 4632 2836 4660 2876
rect 5902 2864 5908 2876
rect 5960 2864 5966 2916
rect 6089 2907 6147 2913
rect 6089 2873 6101 2907
rect 6135 2904 6147 2907
rect 6822 2904 6828 2916
rect 6135 2876 6828 2904
rect 6135 2873 6147 2876
rect 6089 2867 6147 2873
rect 6822 2864 6828 2876
rect 6880 2864 6886 2916
rect 7668 2904 7696 3012
rect 7745 3009 7757 3043
rect 7791 3040 7803 3043
rect 7926 3040 7932 3052
rect 7791 3012 7932 3040
rect 7791 3009 7803 3012
rect 7745 3003 7803 3009
rect 7926 3000 7932 3012
rect 7984 3000 7990 3052
rect 8036 2972 8064 3080
rect 8193 3000 8199 3052
rect 8251 3049 8257 3052
rect 8251 3040 8263 3049
rect 9232 3040 9260 3148
rect 9306 3136 9312 3188
rect 9364 3176 9370 3188
rect 9585 3179 9643 3185
rect 9585 3176 9597 3179
rect 9364 3148 9597 3176
rect 9364 3136 9370 3148
rect 9585 3145 9597 3148
rect 9631 3176 9643 3179
rect 10226 3176 10232 3188
rect 9631 3148 10232 3176
rect 9631 3145 9643 3148
rect 9585 3139 9643 3145
rect 10226 3136 10232 3148
rect 10284 3136 10290 3188
rect 13265 3179 13323 3185
rect 13265 3145 13277 3179
rect 13311 3176 13323 3179
rect 14274 3176 14280 3188
rect 13311 3148 14280 3176
rect 13311 3145 13323 3148
rect 13265 3139 13323 3145
rect 14274 3136 14280 3148
rect 14332 3136 14338 3188
rect 14369 3179 14427 3185
rect 14369 3145 14381 3179
rect 14415 3176 14427 3179
rect 20162 3176 20168 3188
rect 14415 3148 20168 3176
rect 14415 3145 14427 3148
rect 14369 3139 14427 3145
rect 20162 3136 20168 3148
rect 20220 3136 20226 3188
rect 11790 3068 11796 3120
rect 11848 3108 11854 3120
rect 12710 3108 12716 3120
rect 11848 3080 12716 3108
rect 11848 3068 11854 3080
rect 12710 3068 12716 3080
rect 12768 3068 12774 3120
rect 14090 3108 14096 3120
rect 12912 3080 14096 3108
rect 10134 3040 10140 3052
rect 8251 3012 8296 3040
rect 9232 3012 10140 3040
rect 8251 3003 8263 3012
rect 8251 3000 8257 3003
rect 10134 3000 10140 3012
rect 10192 3000 10198 3052
rect 10318 3000 10324 3052
rect 10376 3040 10382 3052
rect 10413 3043 10471 3049
rect 10413 3040 10425 3043
rect 10376 3012 10425 3040
rect 10376 3000 10382 3012
rect 10413 3009 10425 3012
rect 10459 3009 10471 3043
rect 10413 3003 10471 3009
rect 10502 3000 10508 3052
rect 10560 3040 10566 3052
rect 12912 3049 12940 3080
rect 14090 3068 14096 3080
rect 14148 3068 14154 3120
rect 14921 3111 14979 3117
rect 14921 3077 14933 3111
rect 14967 3108 14979 3111
rect 16022 3108 16028 3120
rect 14967 3080 16028 3108
rect 14967 3077 14979 3080
rect 14921 3071 14979 3077
rect 16022 3068 16028 3080
rect 16080 3068 16086 3120
rect 11425 3043 11483 3049
rect 11425 3040 11437 3043
rect 10560 3012 11437 3040
rect 10560 3000 10566 3012
rect 11425 3009 11437 3012
rect 11471 3009 11483 3043
rect 11425 3003 11483 3009
rect 12897 3043 12955 3049
rect 12897 3009 12909 3043
rect 12943 3009 12955 3043
rect 12897 3003 12955 3009
rect 13081 3043 13139 3049
rect 13081 3009 13093 3043
rect 13127 3040 13139 3043
rect 13265 3043 13323 3049
rect 13265 3040 13277 3043
rect 13127 3012 13277 3040
rect 13127 3009 13139 3012
rect 13081 3003 13139 3009
rect 13265 3009 13277 3012
rect 13311 3009 13323 3043
rect 13265 3003 13323 3009
rect 13372 3012 14780 3040
rect 9950 2972 9956 2984
rect 8036 2944 9956 2972
rect 9950 2932 9956 2944
rect 10008 2932 10014 2984
rect 10152 2972 10180 3000
rect 10594 2972 10600 2984
rect 10152 2944 10600 2972
rect 10594 2932 10600 2944
rect 10652 2932 10658 2984
rect 10686 2932 10692 2984
rect 10744 2972 10750 2984
rect 13372 2972 13400 3012
rect 10744 2944 13400 2972
rect 13449 2975 13507 2981
rect 10744 2932 10750 2944
rect 13449 2941 13461 2975
rect 13495 2941 13507 2975
rect 13722 2972 13728 2984
rect 13683 2944 13728 2972
rect 13449 2935 13507 2941
rect 8110 2904 8116 2916
rect 7668 2876 8116 2904
rect 8110 2864 8116 2876
rect 8168 2904 8174 2916
rect 8450 2907 8508 2913
rect 8450 2904 8462 2907
rect 8168 2876 8462 2904
rect 8168 2864 8174 2876
rect 8450 2873 8462 2876
rect 8496 2873 8508 2907
rect 8450 2867 8508 2873
rect 8570 2864 8576 2916
rect 8628 2904 8634 2916
rect 9490 2904 9496 2916
rect 8628 2876 9496 2904
rect 8628 2864 8634 2876
rect 9490 2864 9496 2876
rect 9548 2864 9554 2916
rect 11333 2907 11391 2913
rect 11333 2904 11345 2907
rect 9876 2876 11345 2904
rect 3200 2808 4660 2836
rect 3200 2796 3206 2808
rect 4706 2796 4712 2848
rect 4764 2836 4770 2848
rect 5077 2839 5135 2845
rect 5077 2836 5089 2839
rect 4764 2808 5089 2836
rect 4764 2796 4770 2808
rect 5077 2805 5089 2808
rect 5123 2805 5135 2839
rect 5077 2799 5135 2805
rect 6181 2839 6239 2845
rect 6181 2805 6193 2839
rect 6227 2836 6239 2839
rect 7101 2839 7159 2845
rect 7101 2836 7113 2839
rect 6227 2808 7113 2836
rect 6227 2805 6239 2808
rect 6181 2799 6239 2805
rect 7101 2805 7113 2808
rect 7147 2805 7159 2839
rect 7101 2799 7159 2805
rect 7190 2796 7196 2848
rect 7248 2836 7254 2848
rect 7561 2839 7619 2845
rect 7561 2836 7573 2839
rect 7248 2808 7573 2836
rect 7248 2796 7254 2808
rect 7561 2805 7573 2808
rect 7607 2836 7619 2839
rect 9214 2836 9220 2848
rect 7607 2808 9220 2836
rect 7607 2805 7619 2808
rect 7561 2799 7619 2805
rect 9214 2796 9220 2808
rect 9272 2796 9278 2848
rect 9876 2845 9904 2876
rect 11333 2873 11345 2876
rect 11379 2873 11391 2907
rect 12802 2904 12808 2916
rect 12763 2876 12808 2904
rect 11333 2867 11391 2873
rect 12802 2864 12808 2876
rect 12860 2864 12866 2916
rect 13078 2864 13084 2916
rect 13136 2904 13142 2916
rect 13464 2904 13492 2935
rect 13722 2932 13728 2944
rect 13780 2932 13786 2984
rect 13814 2932 13820 2984
rect 13872 2972 13878 2984
rect 14752 2981 14780 3012
rect 14185 2975 14243 2981
rect 14185 2972 14197 2975
rect 13872 2944 14197 2972
rect 13872 2932 13878 2944
rect 14185 2941 14197 2944
rect 14231 2941 14243 2975
rect 14185 2935 14243 2941
rect 14737 2975 14795 2981
rect 14737 2941 14749 2975
rect 14783 2941 14795 2975
rect 14737 2935 14795 2941
rect 15289 2975 15347 2981
rect 15289 2941 15301 2975
rect 15335 2941 15347 2975
rect 16114 2972 16120 2984
rect 16075 2944 16120 2972
rect 15289 2935 15347 2941
rect 13136 2876 13492 2904
rect 13136 2864 13142 2876
rect 14458 2864 14464 2916
rect 14516 2904 14522 2916
rect 15304 2904 15332 2935
rect 16114 2932 16120 2944
rect 16172 2932 16178 2984
rect 16850 2932 16856 2984
rect 16908 2972 16914 2984
rect 17037 2975 17095 2981
rect 17037 2972 17049 2975
rect 16908 2944 17049 2972
rect 16908 2932 16914 2944
rect 17037 2941 17049 2944
rect 17083 2941 17095 2975
rect 17037 2935 17095 2941
rect 18325 2975 18383 2981
rect 18325 2941 18337 2975
rect 18371 2972 18383 2975
rect 18506 2972 18512 2984
rect 18371 2944 18512 2972
rect 18371 2941 18383 2944
rect 18325 2935 18383 2941
rect 18506 2932 18512 2944
rect 18564 2932 18570 2984
rect 19150 2972 19156 2984
rect 19111 2944 19156 2972
rect 19150 2932 19156 2944
rect 19208 2932 19214 2984
rect 22002 2904 22008 2916
rect 14516 2876 15332 2904
rect 15488 2876 22008 2904
rect 14516 2864 14522 2876
rect 9861 2839 9919 2845
rect 9861 2805 9873 2839
rect 9907 2805 9919 2839
rect 10226 2836 10232 2848
rect 10187 2808 10232 2836
rect 9861 2799 9919 2805
rect 10226 2796 10232 2808
rect 10284 2796 10290 2848
rect 10321 2839 10379 2845
rect 10321 2805 10333 2839
rect 10367 2836 10379 2839
rect 10502 2836 10508 2848
rect 10367 2808 10508 2836
rect 10367 2805 10379 2808
rect 10321 2799 10379 2805
rect 10502 2796 10508 2808
rect 10560 2796 10566 2848
rect 10594 2796 10600 2848
rect 10652 2836 10658 2848
rect 10873 2839 10931 2845
rect 10873 2836 10885 2839
rect 10652 2808 10885 2836
rect 10652 2796 10658 2808
rect 10873 2805 10885 2808
rect 10919 2805 10931 2839
rect 10873 2799 10931 2805
rect 11054 2796 11060 2848
rect 11112 2836 11118 2848
rect 11241 2839 11299 2845
rect 11241 2836 11253 2839
rect 11112 2808 11253 2836
rect 11112 2796 11118 2808
rect 11241 2805 11253 2808
rect 11287 2805 11299 2839
rect 11241 2799 11299 2805
rect 12437 2839 12495 2845
rect 12437 2805 12449 2839
rect 12483 2836 12495 2839
rect 15286 2836 15292 2848
rect 12483 2808 15292 2836
rect 12483 2805 12495 2808
rect 12437 2799 12495 2805
rect 15286 2796 15292 2808
rect 15344 2796 15350 2848
rect 15488 2845 15516 2876
rect 22002 2864 22008 2876
rect 22060 2864 22066 2916
rect 15473 2839 15531 2845
rect 15473 2805 15485 2839
rect 15519 2805 15531 2839
rect 15473 2799 15531 2805
rect 16301 2839 16359 2845
rect 16301 2805 16313 2839
rect 16347 2836 16359 2839
rect 16942 2836 16948 2848
rect 16347 2808 16948 2836
rect 16347 2805 16359 2808
rect 16301 2799 16359 2805
rect 16942 2796 16948 2808
rect 17000 2796 17006 2848
rect 17221 2839 17279 2845
rect 17221 2805 17233 2839
rect 17267 2836 17279 2839
rect 17862 2836 17868 2848
rect 17267 2808 17868 2836
rect 17267 2805 17279 2808
rect 17221 2799 17279 2805
rect 17862 2796 17868 2808
rect 17920 2796 17926 2848
rect 18509 2839 18567 2845
rect 18509 2805 18521 2839
rect 18555 2836 18567 2839
rect 19242 2836 19248 2848
rect 18555 2808 19248 2836
rect 18555 2805 18567 2808
rect 18509 2799 18567 2805
rect 19242 2796 19248 2808
rect 19300 2796 19306 2848
rect 19337 2839 19395 2845
rect 19337 2805 19349 2839
rect 19383 2836 19395 2839
rect 19702 2836 19708 2848
rect 19383 2808 19708 2836
rect 19383 2805 19395 2808
rect 19337 2799 19395 2805
rect 19702 2796 19708 2808
rect 19760 2796 19766 2848
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 2314 2632 2320 2644
rect 2275 2604 2320 2632
rect 2314 2592 2320 2604
rect 2372 2592 2378 2644
rect 2682 2632 2688 2644
rect 2643 2604 2688 2632
rect 2682 2592 2688 2604
rect 2740 2592 2746 2644
rect 5353 2635 5411 2641
rect 5353 2601 5365 2635
rect 5399 2632 5411 2635
rect 7282 2632 7288 2644
rect 5399 2604 7288 2632
rect 5399 2601 5411 2604
rect 5353 2595 5411 2601
rect 7282 2592 7288 2604
rect 7340 2592 7346 2644
rect 8386 2592 8392 2644
rect 8444 2632 8450 2644
rect 9033 2635 9091 2641
rect 9033 2632 9045 2635
rect 8444 2604 9045 2632
rect 8444 2592 8450 2604
rect 9033 2601 9045 2604
rect 9079 2601 9091 2635
rect 10134 2632 10140 2644
rect 10095 2604 10140 2632
rect 9033 2595 9091 2601
rect 10134 2592 10140 2604
rect 10192 2592 10198 2644
rect 10229 2635 10287 2641
rect 10229 2601 10241 2635
rect 10275 2632 10287 2635
rect 10962 2632 10968 2644
rect 10275 2604 10968 2632
rect 10275 2601 10287 2604
rect 10229 2595 10287 2601
rect 10962 2592 10968 2604
rect 11020 2592 11026 2644
rect 11146 2632 11152 2644
rect 11107 2604 11152 2632
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 15102 2632 15108 2644
rect 11808 2604 15108 2632
rect 4062 2524 4068 2576
rect 4120 2564 4126 2576
rect 4709 2567 4767 2573
rect 4709 2564 4721 2567
rect 4120 2536 4721 2564
rect 4120 2524 4126 2536
rect 4709 2533 4721 2536
rect 4755 2564 4767 2567
rect 5626 2564 5632 2576
rect 4755 2536 5632 2564
rect 4755 2533 4767 2536
rect 4709 2527 4767 2533
rect 5626 2524 5632 2536
rect 5684 2524 5690 2576
rect 7006 2524 7012 2576
rect 7064 2564 7070 2576
rect 8113 2567 8171 2573
rect 8113 2564 8125 2567
rect 7064 2536 8125 2564
rect 7064 2524 7070 2536
rect 8113 2533 8125 2536
rect 8159 2564 8171 2567
rect 8478 2564 8484 2576
rect 8159 2536 8484 2564
rect 8159 2533 8171 2536
rect 8113 2527 8171 2533
rect 8478 2524 8484 2536
rect 8536 2524 8542 2576
rect 9125 2567 9183 2573
rect 9125 2533 9137 2567
rect 9171 2564 9183 2567
rect 10594 2564 10600 2576
rect 9171 2536 10600 2564
rect 9171 2533 9183 2536
rect 9125 2527 9183 2533
rect 10594 2524 10600 2536
rect 10652 2524 10658 2576
rect 4816 2468 5212 2496
rect 2774 2388 2780 2440
rect 2832 2428 2838 2440
rect 2961 2431 3019 2437
rect 2832 2400 2877 2428
rect 2832 2388 2838 2400
rect 2961 2397 2973 2431
rect 3007 2428 3019 2431
rect 3418 2428 3424 2440
rect 3007 2400 3424 2428
rect 3007 2397 3019 2400
rect 2961 2391 3019 2397
rect 3418 2388 3424 2400
rect 3476 2388 3482 2440
rect 4062 2388 4068 2440
rect 4120 2428 4126 2440
rect 4816 2437 4844 2468
rect 4801 2431 4859 2437
rect 4801 2428 4813 2431
rect 4120 2400 4813 2428
rect 4120 2388 4126 2400
rect 4801 2397 4813 2400
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2397 5043 2431
rect 5184 2428 5212 2468
rect 5258 2456 5264 2508
rect 5316 2496 5322 2508
rect 5721 2499 5779 2505
rect 5721 2496 5733 2499
rect 5316 2468 5733 2496
rect 5316 2456 5322 2468
rect 5721 2465 5733 2468
rect 5767 2465 5779 2499
rect 5721 2459 5779 2465
rect 5813 2499 5871 2505
rect 5813 2465 5825 2499
rect 5859 2496 5871 2499
rect 6454 2496 6460 2508
rect 5859 2468 6460 2496
rect 5859 2465 5871 2468
rect 5813 2459 5871 2465
rect 6454 2456 6460 2468
rect 6512 2456 6518 2508
rect 6917 2499 6975 2505
rect 6917 2465 6929 2499
rect 6963 2496 6975 2499
rect 7374 2496 7380 2508
rect 6963 2468 7380 2496
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 7374 2456 7380 2468
rect 7432 2456 7438 2508
rect 8018 2496 8024 2508
rect 7979 2468 8024 2496
rect 8018 2456 8024 2468
rect 8076 2456 8082 2508
rect 11698 2496 11704 2508
rect 8128 2468 11704 2496
rect 5902 2428 5908 2440
rect 5184 2400 5908 2428
rect 4985 2391 5043 2397
rect 5000 2360 5028 2391
rect 5902 2388 5908 2400
rect 5960 2388 5966 2440
rect 5997 2431 6055 2437
rect 5997 2397 6009 2431
rect 6043 2428 6055 2431
rect 6362 2428 6368 2440
rect 6043 2400 6368 2428
rect 6043 2397 6055 2400
rect 5997 2391 6055 2397
rect 6012 2360 6040 2391
rect 6362 2388 6368 2400
rect 6420 2388 6426 2440
rect 7193 2431 7251 2437
rect 7193 2397 7205 2431
rect 7239 2428 7251 2431
rect 8128 2428 8156 2468
rect 11698 2456 11704 2468
rect 11756 2456 11762 2508
rect 11808 2505 11836 2604
rect 15102 2592 15108 2604
rect 15160 2592 15166 2644
rect 12066 2564 12072 2576
rect 12027 2536 12072 2564
rect 12066 2524 12072 2536
rect 12124 2524 12130 2576
rect 12897 2567 12955 2573
rect 12897 2533 12909 2567
rect 12943 2564 12955 2567
rect 13538 2564 13544 2576
rect 12943 2536 13544 2564
rect 12943 2533 12955 2536
rect 12897 2527 12955 2533
rect 13538 2524 13544 2536
rect 13596 2524 13602 2576
rect 13725 2567 13783 2573
rect 13725 2533 13737 2567
rect 13771 2564 13783 2567
rect 21542 2564 21548 2576
rect 13771 2536 21548 2564
rect 13771 2533 13783 2536
rect 13725 2527 13783 2533
rect 21542 2524 21548 2536
rect 21600 2524 21606 2576
rect 11793 2499 11851 2505
rect 11793 2465 11805 2499
rect 11839 2465 11851 2499
rect 11793 2459 11851 2465
rect 12631 2499 12689 2505
rect 12631 2465 12643 2499
rect 12677 2465 12689 2499
rect 12631 2459 12689 2465
rect 7239 2400 8156 2428
rect 8205 2431 8263 2437
rect 7239 2397 7251 2400
rect 7193 2391 7251 2397
rect 8205 2397 8217 2431
rect 8251 2397 8263 2431
rect 9306 2428 9312 2440
rect 9267 2400 9312 2428
rect 8205 2391 8263 2397
rect 5000 2332 6040 2360
rect 7742 2320 7748 2372
rect 7800 2360 7806 2372
rect 8220 2360 8248 2391
rect 9306 2388 9312 2400
rect 9364 2388 9370 2440
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 10318 2428 10324 2440
rect 9732 2400 10324 2428
rect 9732 2388 9738 2400
rect 10318 2388 10324 2400
rect 10376 2388 10382 2440
rect 11241 2431 11299 2437
rect 11241 2428 11253 2431
rect 10428 2400 11253 2428
rect 7800 2332 8248 2360
rect 7800 2320 7806 2332
rect 4341 2295 4399 2301
rect 4341 2261 4353 2295
rect 4387 2292 4399 2295
rect 6914 2292 6920 2304
rect 4387 2264 6920 2292
rect 4387 2261 4399 2264
rect 4341 2255 4399 2261
rect 6914 2252 6920 2264
rect 6972 2252 6978 2304
rect 7006 2252 7012 2304
rect 7064 2292 7070 2304
rect 7653 2295 7711 2301
rect 7653 2292 7665 2295
rect 7064 2264 7665 2292
rect 7064 2252 7070 2264
rect 7653 2261 7665 2264
rect 7699 2261 7711 2295
rect 8220 2292 8248 2332
rect 8665 2363 8723 2369
rect 8665 2329 8677 2363
rect 8711 2360 8723 2363
rect 10428 2360 10456 2400
rect 11241 2397 11253 2400
rect 11287 2397 11299 2431
rect 11241 2391 11299 2397
rect 11425 2431 11483 2437
rect 11425 2397 11437 2431
rect 11471 2428 11483 2431
rect 11606 2428 11612 2440
rect 11471 2400 11612 2428
rect 11471 2397 11483 2400
rect 11425 2391 11483 2397
rect 11606 2388 11612 2400
rect 11664 2388 11670 2440
rect 8711 2332 10456 2360
rect 10781 2363 10839 2369
rect 8711 2329 8723 2332
rect 8665 2323 8723 2329
rect 10781 2329 10793 2363
rect 10827 2360 10839 2363
rect 12636 2360 12664 2459
rect 12986 2456 12992 2508
rect 13044 2496 13050 2508
rect 13357 2499 13415 2505
rect 13357 2496 13369 2499
rect 13044 2468 13369 2496
rect 13044 2456 13050 2468
rect 13357 2465 13369 2468
rect 13403 2465 13415 2499
rect 13906 2496 13912 2508
rect 13867 2468 13912 2496
rect 13357 2459 13415 2465
rect 13906 2456 13912 2468
rect 13964 2456 13970 2508
rect 14182 2456 14188 2508
rect 14240 2496 14246 2508
rect 14737 2499 14795 2505
rect 14737 2496 14749 2499
rect 14240 2468 14749 2496
rect 14240 2456 14246 2468
rect 14737 2465 14749 2468
rect 14783 2465 14795 2499
rect 15654 2496 15660 2508
rect 15615 2468 15660 2496
rect 14737 2459 14795 2465
rect 15654 2456 15660 2468
rect 15712 2456 15718 2508
rect 16574 2496 16580 2508
rect 16535 2468 16580 2496
rect 16574 2456 16580 2468
rect 16632 2456 16638 2508
rect 17034 2456 17040 2508
rect 17092 2496 17098 2508
rect 17497 2499 17555 2505
rect 17497 2496 17509 2499
rect 17092 2468 17509 2496
rect 17092 2456 17098 2468
rect 17497 2465 17509 2468
rect 17543 2465 17555 2499
rect 17497 2459 17555 2465
rect 10827 2332 12664 2360
rect 13541 2363 13599 2369
rect 10827 2329 10839 2332
rect 10781 2323 10839 2329
rect 13541 2329 13553 2363
rect 13587 2360 13599 2363
rect 13725 2363 13783 2369
rect 13725 2360 13737 2363
rect 13587 2332 13737 2360
rect 13587 2329 13599 2332
rect 13541 2323 13599 2329
rect 13725 2329 13737 2332
rect 13771 2329 13783 2363
rect 13725 2323 13783 2329
rect 14093 2363 14151 2369
rect 14093 2329 14105 2363
rect 14139 2360 14151 2363
rect 21082 2360 21088 2372
rect 14139 2332 21088 2360
rect 14139 2329 14151 2332
rect 14093 2323 14151 2329
rect 21082 2320 21088 2332
rect 21140 2320 21146 2372
rect 8754 2292 8760 2304
rect 8220 2264 8760 2292
rect 7653 2255 7711 2261
rect 8754 2252 8760 2264
rect 8812 2292 8818 2304
rect 9674 2292 9680 2304
rect 8812 2264 9680 2292
rect 8812 2252 8818 2264
rect 9674 2252 9680 2264
rect 9732 2252 9738 2304
rect 9769 2295 9827 2301
rect 9769 2261 9781 2295
rect 9815 2292 9827 2295
rect 11054 2292 11060 2304
rect 9815 2264 11060 2292
rect 9815 2261 9827 2264
rect 9769 2255 9827 2261
rect 11054 2252 11060 2264
rect 11112 2252 11118 2304
rect 14921 2295 14979 2301
rect 14921 2261 14933 2295
rect 14967 2292 14979 2295
rect 15562 2292 15568 2304
rect 14967 2264 15568 2292
rect 14967 2261 14979 2264
rect 14921 2255 14979 2261
rect 15562 2252 15568 2264
rect 15620 2252 15626 2304
rect 15841 2295 15899 2301
rect 15841 2261 15853 2295
rect 15887 2292 15899 2295
rect 16482 2292 16488 2304
rect 15887 2264 16488 2292
rect 15887 2261 15899 2264
rect 15841 2255 15899 2261
rect 16482 2252 16488 2264
rect 16540 2252 16546 2304
rect 16761 2295 16819 2301
rect 16761 2261 16773 2295
rect 16807 2292 16819 2295
rect 17402 2292 17408 2304
rect 16807 2264 17408 2292
rect 16807 2261 16819 2264
rect 16761 2255 16819 2261
rect 17402 2252 17408 2264
rect 17460 2252 17466 2304
rect 17681 2295 17739 2301
rect 17681 2261 17693 2295
rect 17727 2292 17739 2295
rect 17954 2292 17960 2304
rect 17727 2264 17960 2292
rect 17727 2261 17739 2264
rect 17681 2255 17739 2261
rect 17954 2252 17960 2264
rect 18012 2252 18018 2304
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 6454 2048 6460 2100
rect 6512 2088 6518 2100
rect 13354 2088 13360 2100
rect 6512 2060 13360 2088
rect 6512 2048 6518 2060
rect 13354 2048 13360 2060
rect 13412 2088 13418 2100
rect 15654 2088 15660 2100
rect 13412 2060 15660 2088
rect 13412 2048 13418 2060
rect 15654 2048 15660 2060
rect 15712 2048 15718 2100
rect 2038 1980 2044 2032
rect 2096 2020 2102 2032
rect 8018 2020 8024 2032
rect 2096 1992 8024 2020
rect 2096 1980 2102 1992
rect 8018 1980 8024 1992
rect 8076 2020 8082 2032
rect 9582 2020 9588 2032
rect 8076 1992 9588 2020
rect 8076 1980 8082 1992
rect 9582 1980 9588 1992
rect 9640 1980 9646 2032
rect 658 1912 664 1964
rect 716 1952 722 1964
rect 7190 1952 7196 1964
rect 716 1924 7196 1952
rect 716 1912 722 1924
rect 7190 1912 7196 1924
rect 7248 1912 7254 1964
rect 1118 1844 1124 1896
rect 1176 1884 1182 1896
rect 5442 1884 5448 1896
rect 1176 1856 5448 1884
rect 1176 1844 1182 1856
rect 5442 1844 5448 1856
rect 5500 1884 5506 1896
rect 7466 1884 7472 1896
rect 5500 1856 7472 1884
rect 5500 1844 5506 1856
rect 7466 1844 7472 1856
rect 7524 1844 7530 1896
rect 11330 1368 11336 1420
rect 11388 1408 11394 1420
rect 12158 1408 12164 1420
rect 11388 1380 12164 1408
rect 11388 1368 11394 1380
rect 12158 1368 12164 1380
rect 12216 1368 12222 1420
rect 3510 1300 3516 1352
rect 3568 1340 3574 1352
rect 5166 1340 5172 1352
rect 3568 1312 5172 1340
rect 3568 1300 3574 1312
rect 5166 1300 5172 1312
rect 5224 1300 5230 1352
<< via1 >>
rect 3700 20816 3752 20868
rect 6920 20816 6972 20868
rect 4068 20272 4120 20324
rect 6368 20272 6420 20324
rect 3700 20204 3752 20256
rect 6736 20204 6788 20256
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 5172 20000 5224 20052
rect 5540 20000 5592 20052
rect 6920 20000 6972 20052
rect 10876 20000 10928 20052
rect 12900 20000 12952 20052
rect 13360 20043 13412 20052
rect 13360 20009 13369 20043
rect 13369 20009 13403 20043
rect 13403 20009 13412 20043
rect 13360 20000 13412 20009
rect 14556 20000 14608 20052
rect 15200 20000 15252 20052
rect 15660 20043 15712 20052
rect 15660 20009 15669 20043
rect 15669 20009 15703 20043
rect 15703 20009 15712 20043
rect 15660 20000 15712 20009
rect 16580 20000 16632 20052
rect 17960 20000 18012 20052
rect 2872 19864 2924 19916
rect 3056 19907 3108 19916
rect 3056 19873 3065 19907
rect 3065 19873 3099 19907
rect 3099 19873 3108 19907
rect 3056 19864 3108 19873
rect 5264 19864 5316 19916
rect 6460 19864 6512 19916
rect 8852 19864 8904 19916
rect 12440 19932 12492 19984
rect 9864 19864 9916 19916
rect 3240 19839 3292 19848
rect 3240 19805 3249 19839
rect 3249 19805 3283 19839
rect 3283 19805 3292 19839
rect 3240 19796 3292 19805
rect 3516 19728 3568 19780
rect 4896 19796 4948 19848
rect 5080 19796 5132 19848
rect 7380 19839 7432 19848
rect 1860 19703 1912 19712
rect 1860 19669 1869 19703
rect 1869 19669 1903 19703
rect 1903 19669 1912 19703
rect 1860 19660 1912 19669
rect 4068 19703 4120 19712
rect 4068 19669 4077 19703
rect 4077 19669 4111 19703
rect 4111 19669 4120 19703
rect 4068 19660 4120 19669
rect 4988 19728 5040 19780
rect 7380 19805 7389 19839
rect 7389 19805 7423 19839
rect 7423 19805 7432 19839
rect 7380 19796 7432 19805
rect 10968 19839 11020 19848
rect 10968 19805 10977 19839
rect 10977 19805 11011 19839
rect 11011 19805 11020 19839
rect 10968 19796 11020 19805
rect 13912 19864 13964 19916
rect 14188 19907 14240 19916
rect 14188 19873 14197 19907
rect 14197 19873 14231 19907
rect 14231 19873 14240 19907
rect 14188 19864 14240 19873
rect 14464 19864 14516 19916
rect 15476 19907 15528 19916
rect 15476 19873 15485 19907
rect 15485 19873 15519 19907
rect 15519 19873 15528 19907
rect 15476 19864 15528 19873
rect 15568 19864 15620 19916
rect 17040 19907 17092 19916
rect 17040 19873 17049 19907
rect 17049 19873 17083 19907
rect 17083 19873 17092 19907
rect 17040 19864 17092 19873
rect 11704 19796 11756 19848
rect 12072 19839 12124 19848
rect 12072 19805 12081 19839
rect 12081 19805 12115 19839
rect 12115 19805 12124 19839
rect 12072 19796 12124 19805
rect 19800 19728 19852 19780
rect 6920 19660 6972 19712
rect 11796 19660 11848 19712
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 3240 19456 3292 19508
rect 5816 19456 5868 19508
rect 6460 19499 6512 19508
rect 6460 19465 6469 19499
rect 6469 19465 6503 19499
rect 6503 19465 6512 19499
rect 6460 19456 6512 19465
rect 7380 19456 7432 19508
rect 10968 19456 11020 19508
rect 3976 19320 4028 19372
rect 2136 19295 2188 19304
rect 2136 19261 2145 19295
rect 2145 19261 2179 19295
rect 2179 19261 2188 19295
rect 2136 19252 2188 19261
rect 2228 19184 2280 19236
rect 2596 19184 2648 19236
rect 1768 19159 1820 19168
rect 1768 19125 1777 19159
rect 1777 19125 1811 19159
rect 1811 19125 1820 19159
rect 1768 19116 1820 19125
rect 4896 19252 4948 19304
rect 5080 19295 5132 19304
rect 5080 19261 5089 19295
rect 5089 19261 5123 19295
rect 5123 19261 5132 19295
rect 5080 19252 5132 19261
rect 4252 19184 4304 19236
rect 5724 19184 5776 19236
rect 5816 19184 5868 19236
rect 6920 19184 6972 19236
rect 7104 19252 7156 19304
rect 8760 19252 8812 19304
rect 10324 19252 10376 19304
rect 12072 19252 12124 19304
rect 12164 19252 12216 19304
rect 14096 19295 14148 19304
rect 14096 19261 14105 19295
rect 14105 19261 14139 19295
rect 14139 19261 14148 19295
rect 14096 19252 14148 19261
rect 3240 19116 3292 19168
rect 3332 19116 3384 19168
rect 3516 19116 3568 19168
rect 3608 19116 3660 19168
rect 4436 19116 4488 19168
rect 6644 19116 6696 19168
rect 7012 19116 7064 19168
rect 8392 19116 8444 19168
rect 9036 19116 9088 19168
rect 9404 19159 9456 19168
rect 9404 19125 9413 19159
rect 9413 19125 9447 19159
rect 9447 19125 9456 19159
rect 9404 19116 9456 19125
rect 10968 19184 11020 19236
rect 11796 19227 11848 19236
rect 11796 19193 11805 19227
rect 11805 19193 11839 19227
rect 11839 19193 11848 19227
rect 11796 19184 11848 19193
rect 12716 19227 12768 19236
rect 12716 19193 12750 19227
rect 12750 19193 12768 19227
rect 12716 19184 12768 19193
rect 13728 19184 13780 19236
rect 16580 19295 16632 19304
rect 16580 19261 16589 19295
rect 16589 19261 16623 19295
rect 16623 19261 16632 19295
rect 16580 19252 16632 19261
rect 17132 19295 17184 19304
rect 17132 19261 17141 19295
rect 17141 19261 17175 19295
rect 17175 19261 17184 19295
rect 17132 19252 17184 19261
rect 17224 19252 17276 19304
rect 18604 19295 18656 19304
rect 18604 19261 18613 19295
rect 18613 19261 18647 19295
rect 18647 19261 18656 19295
rect 18604 19252 18656 19261
rect 18788 19252 18840 19304
rect 22100 19184 22152 19236
rect 11428 19116 11480 19168
rect 14280 19159 14332 19168
rect 14280 19125 14289 19159
rect 14289 19125 14323 19159
rect 14323 19125 14332 19159
rect 14280 19116 14332 19125
rect 15108 19116 15160 19168
rect 16120 19116 16172 19168
rect 16948 19116 17000 19168
rect 17500 19116 17552 19168
rect 18512 19116 18564 19168
rect 18880 19116 18932 19168
rect 20260 19116 20312 19168
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 1492 18912 1544 18964
rect 2504 18912 2556 18964
rect 2872 18912 2924 18964
rect 3332 18955 3384 18964
rect 3332 18921 3341 18955
rect 3341 18921 3375 18955
rect 3375 18921 3384 18955
rect 3332 18912 3384 18921
rect 4068 18912 4120 18964
rect 4344 18912 4396 18964
rect 5172 18912 5224 18964
rect 3976 18844 4028 18896
rect 4528 18887 4580 18896
rect 4528 18853 4537 18887
rect 4537 18853 4571 18887
rect 4571 18853 4580 18887
rect 4528 18844 4580 18853
rect 5540 18912 5592 18964
rect 5724 18912 5776 18964
rect 6736 18912 6788 18964
rect 8852 18955 8904 18964
rect 8852 18921 8861 18955
rect 8861 18921 8895 18955
rect 8895 18921 8904 18955
rect 8852 18912 8904 18921
rect 9312 18912 9364 18964
rect 1400 18819 1452 18828
rect 1400 18785 1409 18819
rect 1409 18785 1443 18819
rect 1443 18785 1452 18819
rect 1400 18776 1452 18785
rect 3332 18776 3384 18828
rect 204 18708 256 18760
rect 1584 18683 1636 18692
rect 1584 18649 1593 18683
rect 1593 18649 1627 18683
rect 1627 18649 1636 18683
rect 1584 18640 1636 18649
rect 4344 18776 4396 18828
rect 3608 18751 3660 18760
rect 3608 18717 3617 18751
rect 3617 18717 3651 18751
rect 3651 18717 3660 18751
rect 3608 18708 3660 18717
rect 7380 18844 7432 18896
rect 9404 18844 9456 18896
rect 11888 18912 11940 18964
rect 12716 18912 12768 18964
rect 19340 18912 19392 18964
rect 21180 18912 21232 18964
rect 2780 18640 2832 18692
rect 3056 18640 3108 18692
rect 4160 18572 4212 18624
rect 4804 18708 4856 18760
rect 5080 18708 5132 18760
rect 5816 18776 5868 18828
rect 6000 18776 6052 18828
rect 7380 18708 7432 18760
rect 8392 18572 8444 18624
rect 11336 18819 11388 18828
rect 10140 18751 10192 18760
rect 10140 18717 10149 18751
rect 10149 18717 10183 18751
rect 10183 18717 10192 18751
rect 10140 18708 10192 18717
rect 11336 18785 11345 18819
rect 11345 18785 11379 18819
rect 11379 18785 11388 18819
rect 11336 18776 11388 18785
rect 11796 18776 11848 18828
rect 12348 18844 12400 18896
rect 13912 18887 13964 18896
rect 12072 18776 12124 18828
rect 12992 18776 13044 18828
rect 13912 18853 13921 18887
rect 13921 18853 13955 18887
rect 13955 18853 13964 18887
rect 13912 18844 13964 18853
rect 14188 18844 14240 18896
rect 15568 18887 15620 18896
rect 15568 18853 15577 18887
rect 15577 18853 15611 18887
rect 15611 18853 15620 18887
rect 15568 18844 15620 18853
rect 18788 18887 18840 18896
rect 18788 18853 18797 18887
rect 18797 18853 18831 18887
rect 18831 18853 18840 18887
rect 18788 18844 18840 18853
rect 15200 18776 15252 18828
rect 18512 18819 18564 18828
rect 18512 18785 18521 18819
rect 18521 18785 18555 18819
rect 18555 18785 18564 18819
rect 18512 18776 18564 18785
rect 15568 18708 15620 18760
rect 10692 18572 10744 18624
rect 10968 18615 11020 18624
rect 10968 18581 10977 18615
rect 10977 18581 11011 18615
rect 11011 18581 11020 18615
rect 10968 18572 11020 18581
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 1032 18368 1084 18420
rect 2596 18368 2648 18420
rect 2780 18368 2832 18420
rect 3056 18368 3108 18420
rect 10968 18368 11020 18420
rect 11796 18368 11848 18420
rect 13452 18411 13504 18420
rect 13452 18377 13461 18411
rect 13461 18377 13495 18411
rect 13495 18377 13504 18411
rect 13452 18368 13504 18377
rect 21640 18368 21692 18420
rect 1676 18343 1728 18352
rect 1676 18309 1685 18343
rect 1685 18309 1719 18343
rect 1719 18309 1728 18343
rect 1676 18300 1728 18309
rect 4896 18343 4948 18352
rect 4896 18309 4905 18343
rect 4905 18309 4939 18343
rect 4939 18309 4948 18343
rect 4896 18300 4948 18309
rect 5724 18275 5776 18284
rect 2228 18164 2280 18216
rect 572 18028 624 18080
rect 2688 18028 2740 18080
rect 5724 18241 5733 18275
rect 5733 18241 5767 18275
rect 5767 18241 5776 18275
rect 5724 18232 5776 18241
rect 8116 18232 8168 18284
rect 8392 18275 8444 18284
rect 8392 18241 8401 18275
rect 8401 18241 8435 18275
rect 8435 18241 8444 18275
rect 8392 18232 8444 18241
rect 8852 18232 8904 18284
rect 10048 18300 10100 18352
rect 11612 18300 11664 18352
rect 13084 18300 13136 18352
rect 4068 18164 4120 18216
rect 4160 18164 4212 18216
rect 11152 18232 11204 18284
rect 11796 18232 11848 18284
rect 12992 18275 13044 18284
rect 12992 18241 13001 18275
rect 13001 18241 13035 18275
rect 13035 18241 13044 18275
rect 12992 18232 13044 18241
rect 13912 18232 13964 18284
rect 4804 18096 4856 18148
rect 4896 18096 4948 18148
rect 9128 18096 9180 18148
rect 9680 18096 9732 18148
rect 13176 18164 13228 18216
rect 6368 18071 6420 18080
rect 6368 18037 6377 18071
rect 6377 18037 6411 18071
rect 6411 18037 6420 18071
rect 6368 18028 6420 18037
rect 6460 18028 6512 18080
rect 7196 18071 7248 18080
rect 7196 18037 7205 18071
rect 7205 18037 7239 18071
rect 7239 18037 7248 18071
rect 7196 18028 7248 18037
rect 7288 18071 7340 18080
rect 7288 18037 7297 18071
rect 7297 18037 7331 18071
rect 7331 18037 7340 18071
rect 7288 18028 7340 18037
rect 7472 18028 7524 18080
rect 8300 18071 8352 18080
rect 8300 18037 8309 18071
rect 8309 18037 8343 18071
rect 8343 18037 8352 18071
rect 8300 18028 8352 18037
rect 9956 18028 10008 18080
rect 10876 18071 10928 18080
rect 10876 18037 10885 18071
rect 10885 18037 10919 18071
rect 10919 18037 10928 18071
rect 10876 18028 10928 18037
rect 11060 18028 11112 18080
rect 12440 18028 12492 18080
rect 12900 18071 12952 18080
rect 12900 18037 12909 18071
rect 12909 18037 12943 18071
rect 12943 18037 12952 18071
rect 12900 18028 12952 18037
rect 13544 18028 13596 18080
rect 14004 18028 14056 18080
rect 19524 18028 19576 18080
rect 22560 18028 22612 18080
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 4252 17824 4304 17876
rect 7196 17824 7248 17876
rect 9128 17867 9180 17876
rect 9128 17833 9137 17867
rect 9137 17833 9171 17867
rect 9171 17833 9180 17867
rect 9128 17824 9180 17833
rect 9680 17867 9732 17876
rect 9680 17833 9689 17867
rect 9689 17833 9723 17867
rect 9723 17833 9732 17867
rect 9680 17824 9732 17833
rect 13912 17867 13964 17876
rect 6000 17799 6052 17808
rect 6000 17765 6009 17799
rect 6009 17765 6043 17799
rect 6043 17765 6052 17799
rect 6000 17756 6052 17765
rect 1400 17620 1452 17672
rect 3240 17688 3292 17740
rect 4068 17731 4120 17740
rect 4068 17697 4077 17731
rect 4077 17697 4111 17731
rect 4111 17697 4120 17731
rect 4068 17688 4120 17697
rect 4712 17688 4764 17740
rect 7472 17756 7524 17808
rect 7104 17688 7156 17740
rect 12164 17756 12216 17808
rect 13912 17833 13921 17867
rect 13921 17833 13955 17867
rect 13955 17833 13964 17867
rect 13912 17824 13964 17833
rect 20628 17824 20680 17876
rect 3424 17663 3476 17672
rect 3424 17629 3433 17663
rect 3433 17629 3467 17663
rect 3467 17629 3476 17663
rect 3424 17620 3476 17629
rect 3976 17484 4028 17536
rect 5816 17620 5868 17672
rect 6736 17620 6788 17672
rect 7012 17663 7064 17672
rect 7012 17629 7021 17663
rect 7021 17629 7055 17663
rect 7055 17629 7064 17663
rect 7012 17620 7064 17629
rect 8208 17688 8260 17740
rect 9496 17688 9548 17740
rect 10140 17731 10192 17740
rect 10140 17697 10149 17731
rect 10149 17697 10183 17731
rect 10183 17697 10192 17731
rect 10140 17688 10192 17697
rect 10416 17688 10468 17740
rect 11704 17688 11756 17740
rect 11980 17688 12032 17740
rect 7472 17663 7524 17672
rect 7472 17629 7481 17663
rect 7481 17629 7515 17663
rect 7515 17629 7524 17663
rect 7472 17620 7524 17629
rect 8484 17620 8536 17672
rect 9864 17620 9916 17672
rect 9680 17552 9732 17604
rect 10508 17620 10560 17672
rect 12072 17620 12124 17672
rect 12532 17663 12584 17672
rect 12532 17629 12541 17663
rect 12541 17629 12575 17663
rect 12575 17629 12584 17663
rect 12532 17620 12584 17629
rect 10876 17484 10928 17536
rect 11796 17484 11848 17536
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 1768 17323 1820 17332
rect 1768 17289 1777 17323
rect 1777 17289 1811 17323
rect 1811 17289 1820 17323
rect 1768 17280 1820 17289
rect 3424 17280 3476 17332
rect 5632 17280 5684 17332
rect 6276 17280 6328 17332
rect 8208 17323 8260 17332
rect 4712 17212 4764 17264
rect 3240 17187 3292 17196
rect 1584 17119 1636 17128
rect 1584 17085 1593 17119
rect 1593 17085 1627 17119
rect 1627 17085 1636 17119
rect 1584 17076 1636 17085
rect 2320 17008 2372 17060
rect 3240 17153 3249 17187
rect 3249 17153 3283 17187
rect 3283 17153 3292 17187
rect 3240 17144 3292 17153
rect 5172 17144 5224 17196
rect 5540 17212 5592 17264
rect 8208 17289 8217 17323
rect 8217 17289 8251 17323
rect 8251 17289 8260 17323
rect 8208 17280 8260 17289
rect 10048 17323 10100 17332
rect 10048 17289 10057 17323
rect 10057 17289 10091 17323
rect 10091 17289 10100 17323
rect 10048 17280 10100 17289
rect 11704 17323 11756 17332
rect 11704 17289 11713 17323
rect 11713 17289 11747 17323
rect 11747 17289 11756 17323
rect 11704 17280 11756 17289
rect 12440 17323 12492 17332
rect 12440 17289 12449 17323
rect 12449 17289 12483 17323
rect 12483 17289 12492 17323
rect 12440 17280 12492 17289
rect 13820 17280 13872 17332
rect 19340 17280 19392 17332
rect 11428 17212 11480 17264
rect 6460 17144 6512 17196
rect 10048 17144 10100 17196
rect 5908 17119 5960 17128
rect 5908 17085 5917 17119
rect 5917 17085 5951 17119
rect 5951 17085 5960 17119
rect 5908 17076 5960 17085
rect 6736 17076 6788 17128
rect 6828 17119 6880 17128
rect 6828 17085 6837 17119
rect 6837 17085 6871 17119
rect 6871 17085 6880 17119
rect 6828 17076 6880 17085
rect 7472 17076 7524 17128
rect 8668 17119 8720 17128
rect 8668 17085 8677 17119
rect 8677 17085 8711 17119
rect 8711 17085 8720 17119
rect 8668 17076 8720 17085
rect 9680 17076 9732 17128
rect 10324 17119 10376 17128
rect 10324 17085 10333 17119
rect 10333 17085 10367 17119
rect 10367 17085 10376 17119
rect 10324 17076 10376 17085
rect 11704 17144 11756 17196
rect 10876 17076 10928 17128
rect 11980 17076 12032 17128
rect 12164 17119 12216 17128
rect 12164 17085 12173 17119
rect 12173 17085 12207 17119
rect 12207 17085 12216 17119
rect 12164 17076 12216 17085
rect 12808 17076 12860 17128
rect 3608 17008 3660 17060
rect 3792 17008 3844 17060
rect 4804 17008 4856 17060
rect 1676 16940 1728 16992
rect 5264 16983 5316 16992
rect 5264 16949 5273 16983
rect 5273 16949 5307 16983
rect 5307 16949 5316 16983
rect 5264 16940 5316 16949
rect 6828 16940 6880 16992
rect 7380 17008 7432 17060
rect 12256 17008 12308 17060
rect 14556 17008 14608 17060
rect 8208 16940 8260 16992
rect 9680 16940 9732 16992
rect 10324 16940 10376 16992
rect 12072 16940 12124 16992
rect 12808 16983 12860 16992
rect 12808 16949 12817 16983
rect 12817 16949 12851 16983
rect 12851 16949 12860 16983
rect 12808 16940 12860 16949
rect 13084 16940 13136 16992
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 1860 16779 1912 16788
rect 1860 16745 1869 16779
rect 1869 16745 1903 16779
rect 1903 16745 1912 16779
rect 1860 16736 1912 16745
rect 2964 16736 3016 16788
rect 3424 16779 3476 16788
rect 3424 16745 3433 16779
rect 3433 16745 3467 16779
rect 3467 16745 3476 16779
rect 3424 16736 3476 16745
rect 3976 16736 4028 16788
rect 6184 16736 6236 16788
rect 7288 16736 7340 16788
rect 8300 16736 8352 16788
rect 9956 16779 10008 16788
rect 9956 16745 9965 16779
rect 9965 16745 9999 16779
rect 9999 16745 10008 16779
rect 9956 16736 10008 16745
rect 10876 16736 10928 16788
rect 11060 16736 11112 16788
rect 1584 16668 1636 16720
rect 3148 16668 3200 16720
rect 3516 16668 3568 16720
rect 1676 16643 1728 16652
rect 1676 16609 1685 16643
rect 1685 16609 1719 16643
rect 1719 16609 1728 16643
rect 1676 16600 1728 16609
rect 4252 16600 4304 16652
rect 5816 16600 5868 16652
rect 6828 16668 6880 16720
rect 7196 16668 7248 16720
rect 6552 16643 6604 16652
rect 6552 16609 6586 16643
rect 6586 16609 6604 16643
rect 6552 16600 6604 16609
rect 7012 16600 7064 16652
rect 7380 16600 7432 16652
rect 8484 16643 8536 16652
rect 2688 16532 2740 16584
rect 3240 16532 3292 16584
rect 3792 16532 3844 16584
rect 3424 16464 3476 16516
rect 3700 16464 3752 16516
rect 8484 16609 8493 16643
rect 8493 16609 8527 16643
rect 8527 16609 8536 16643
rect 8484 16600 8536 16609
rect 9956 16600 10008 16652
rect 10140 16668 10192 16720
rect 12072 16668 12124 16720
rect 9680 16532 9732 16584
rect 8852 16464 8904 16516
rect 9772 16464 9824 16516
rect 11152 16600 11204 16652
rect 11796 16600 11848 16652
rect 10508 16575 10560 16584
rect 10508 16541 10517 16575
rect 10517 16541 10551 16575
rect 10551 16541 10560 16575
rect 10508 16532 10560 16541
rect 11428 16575 11480 16584
rect 11428 16541 11437 16575
rect 11437 16541 11471 16575
rect 11471 16541 11480 16575
rect 11428 16532 11480 16541
rect 11704 16532 11756 16584
rect 12532 16600 12584 16652
rect 12900 16643 12952 16652
rect 12900 16609 12934 16643
rect 12934 16609 12952 16643
rect 12900 16600 12952 16609
rect 14556 16711 14608 16720
rect 14556 16677 14565 16711
rect 14565 16677 14599 16711
rect 14599 16677 14608 16711
rect 14556 16668 14608 16677
rect 19432 16600 19484 16652
rect 2964 16439 3016 16448
rect 2964 16405 2973 16439
rect 2973 16405 3007 16439
rect 3007 16405 3016 16439
rect 2964 16396 3016 16405
rect 3332 16396 3384 16448
rect 5264 16396 5316 16448
rect 6000 16439 6052 16448
rect 6000 16405 6009 16439
rect 6009 16405 6043 16439
rect 6043 16405 6052 16439
rect 6000 16396 6052 16405
rect 6460 16396 6512 16448
rect 9956 16396 10008 16448
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 1952 16235 2004 16244
rect 1952 16201 1961 16235
rect 1961 16201 1995 16235
rect 1995 16201 2004 16235
rect 1952 16192 2004 16201
rect 2780 16192 2832 16244
rect 3056 16192 3108 16244
rect 3516 16192 3568 16244
rect 3700 16192 3752 16244
rect 6460 16192 6512 16244
rect 10140 16235 10192 16244
rect 10140 16201 10149 16235
rect 10149 16201 10183 16235
rect 10183 16201 10192 16235
rect 10140 16192 10192 16201
rect 6828 16124 6880 16176
rect 3792 16056 3844 16108
rect 4068 16056 4120 16108
rect 4528 16056 4580 16108
rect 5356 16056 5408 16108
rect 5816 16099 5868 16108
rect 5816 16065 5825 16099
rect 5825 16065 5859 16099
rect 5859 16065 5868 16099
rect 5816 16056 5868 16065
rect 8208 16056 8260 16108
rect 9312 16056 9364 16108
rect 10968 16056 11020 16108
rect 1768 16031 1820 16040
rect 1768 15997 1777 16031
rect 1777 15997 1811 16031
rect 1811 15997 1820 16031
rect 1768 15988 1820 15997
rect 2320 16031 2372 16040
rect 2320 15997 2329 16031
rect 2329 15997 2363 16031
rect 2363 15997 2372 16031
rect 2320 15988 2372 15997
rect 2596 15920 2648 15972
rect 4988 15988 5040 16040
rect 5264 15988 5316 16040
rect 6460 15988 6512 16040
rect 7196 16031 7248 16040
rect 7196 15997 7205 16031
rect 7205 15997 7239 16031
rect 7239 15997 7248 16031
rect 7196 15988 7248 15997
rect 9772 15988 9824 16040
rect 9956 15988 10008 16040
rect 3516 15920 3568 15972
rect 4068 15920 4120 15972
rect 5816 15920 5868 15972
rect 2504 15852 2556 15904
rect 3608 15852 3660 15904
rect 4252 15852 4304 15904
rect 4436 15895 4488 15904
rect 4436 15861 4445 15895
rect 4445 15861 4479 15895
rect 4479 15861 4488 15895
rect 4436 15852 4488 15861
rect 5264 15852 5316 15904
rect 5540 15895 5592 15904
rect 5540 15861 5549 15895
rect 5549 15861 5583 15895
rect 5583 15861 5592 15895
rect 5540 15852 5592 15861
rect 5724 15852 5776 15904
rect 6184 15852 6236 15904
rect 6828 15895 6880 15904
rect 6828 15861 6837 15895
rect 6837 15861 6871 15895
rect 6871 15861 6880 15895
rect 6828 15852 6880 15861
rect 8852 15852 8904 15904
rect 10048 15852 10100 15904
rect 10876 15988 10928 16040
rect 12072 16056 12124 16108
rect 12440 16056 12492 16108
rect 14188 16124 14240 16176
rect 13820 16099 13872 16108
rect 13820 16065 13829 16099
rect 13829 16065 13863 16099
rect 13863 16065 13872 16099
rect 13820 16056 13872 16065
rect 11520 16031 11572 16040
rect 11520 15997 11529 16031
rect 11529 15997 11563 16031
rect 11563 15997 11572 16031
rect 11520 15988 11572 15997
rect 11612 15988 11664 16040
rect 10692 15920 10744 15972
rect 11980 15852 12032 15904
rect 12992 15895 13044 15904
rect 12992 15861 13001 15895
rect 13001 15861 13035 15895
rect 13035 15861 13044 15895
rect 12992 15852 13044 15861
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 1584 15691 1636 15700
rect 1584 15657 1593 15691
rect 1593 15657 1627 15691
rect 1627 15657 1636 15691
rect 1584 15648 1636 15657
rect 2964 15648 3016 15700
rect 4436 15648 4488 15700
rect 4528 15691 4580 15700
rect 4528 15657 4537 15691
rect 4537 15657 4571 15691
rect 4571 15657 4580 15691
rect 4528 15648 4580 15657
rect 3424 15580 3476 15632
rect 5264 15648 5316 15700
rect 6828 15648 6880 15700
rect 7104 15691 7156 15700
rect 7104 15657 7113 15691
rect 7113 15657 7147 15691
rect 7147 15657 7156 15691
rect 7104 15648 7156 15657
rect 6184 15580 6236 15632
rect 6368 15580 6420 15632
rect 6552 15623 6604 15632
rect 6552 15589 6561 15623
rect 6561 15589 6595 15623
rect 6595 15589 6604 15623
rect 11152 15648 11204 15700
rect 11428 15648 11480 15700
rect 11612 15691 11664 15700
rect 11612 15657 11621 15691
rect 11621 15657 11655 15691
rect 11655 15657 11664 15691
rect 11612 15648 11664 15657
rect 11980 15691 12032 15700
rect 11980 15657 11989 15691
rect 11989 15657 12023 15691
rect 12023 15657 12032 15691
rect 11980 15648 12032 15657
rect 12992 15648 13044 15700
rect 6552 15580 6604 15589
rect 1676 15512 1728 15564
rect 2412 15555 2464 15564
rect 2412 15521 2421 15555
rect 2421 15521 2455 15555
rect 2455 15521 2464 15555
rect 2412 15512 2464 15521
rect 3240 15512 3292 15564
rect 3792 15512 3844 15564
rect 4988 15512 5040 15564
rect 9220 15580 9272 15632
rect 9312 15580 9364 15632
rect 10232 15580 10284 15632
rect 11704 15580 11756 15632
rect 14004 15580 14056 15632
rect 8024 15512 8076 15564
rect 2596 15487 2648 15496
rect 2596 15453 2605 15487
rect 2605 15453 2639 15487
rect 2639 15453 2648 15487
rect 2596 15444 2648 15453
rect 3516 15444 3568 15496
rect 3976 15444 4028 15496
rect 4712 15487 4764 15496
rect 4712 15453 4721 15487
rect 4721 15453 4755 15487
rect 4755 15453 4764 15487
rect 4712 15444 4764 15453
rect 3700 15308 3752 15360
rect 6000 15444 6052 15496
rect 7380 15444 7432 15496
rect 5724 15308 5776 15360
rect 5816 15308 5868 15360
rect 6552 15308 6604 15360
rect 6736 15308 6788 15360
rect 8668 15308 8720 15360
rect 10324 15512 10376 15564
rect 12532 15512 12584 15564
rect 14188 15512 14240 15564
rect 12256 15487 12308 15496
rect 12256 15453 12265 15487
rect 12265 15453 12299 15487
rect 12299 15453 12308 15487
rect 12256 15444 12308 15453
rect 9312 15419 9364 15428
rect 9312 15385 9321 15419
rect 9321 15385 9355 15419
rect 9355 15385 9364 15419
rect 9312 15376 9364 15385
rect 13636 15376 13688 15428
rect 10876 15308 10928 15360
rect 10968 15308 11020 15360
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 3424 15147 3476 15156
rect 3424 15113 3433 15147
rect 3433 15113 3467 15147
rect 3467 15113 3476 15147
rect 3424 15104 3476 15113
rect 8760 15104 8812 15156
rect 1676 15011 1728 15020
rect 1676 14977 1685 15011
rect 1685 14977 1719 15011
rect 1719 14977 1728 15011
rect 1676 14968 1728 14977
rect 1768 14832 1820 14884
rect 8024 15036 8076 15088
rect 3516 14968 3568 15020
rect 4988 14968 5040 15020
rect 13728 15104 13780 15156
rect 14004 15147 14056 15156
rect 14004 15113 14013 15147
rect 14013 15113 14047 15147
rect 14047 15113 14056 15147
rect 14004 15104 14056 15113
rect 14188 15104 14240 15156
rect 15016 15147 15068 15156
rect 3240 14943 3292 14952
rect 3240 14909 3249 14943
rect 3249 14909 3283 14943
rect 3283 14909 3292 14943
rect 3240 14900 3292 14909
rect 3700 14900 3752 14952
rect 3884 14900 3936 14952
rect 4712 14900 4764 14952
rect 5908 14900 5960 14952
rect 9312 15036 9364 15088
rect 10232 15036 10284 15088
rect 11612 15036 11664 15088
rect 9496 15011 9548 15020
rect 9496 14977 9505 15011
rect 9505 14977 9539 15011
rect 9539 14977 9548 15011
rect 10324 15011 10376 15020
rect 9496 14968 9548 14977
rect 10324 14977 10333 15011
rect 10333 14977 10367 15011
rect 10367 14977 10376 15011
rect 10324 14968 10376 14977
rect 12440 15011 12492 15020
rect 12440 14977 12449 15011
rect 12449 14977 12483 15011
rect 12483 14977 12492 15011
rect 12440 14968 12492 14977
rect 9588 14900 9640 14952
rect 10968 14900 11020 14952
rect 11060 14900 11112 14952
rect 12164 14900 12216 14952
rect 5448 14832 5500 14884
rect 6368 14832 6420 14884
rect 7104 14875 7156 14884
rect 7104 14841 7138 14875
rect 7138 14841 7156 14875
rect 7104 14832 7156 14841
rect 7196 14832 7248 14884
rect 7380 14832 7432 14884
rect 2228 14807 2280 14816
rect 2228 14773 2237 14807
rect 2237 14773 2271 14807
rect 2271 14773 2280 14807
rect 2228 14764 2280 14773
rect 2688 14807 2740 14816
rect 2688 14773 2697 14807
rect 2697 14773 2731 14807
rect 2731 14773 2740 14807
rect 2688 14764 2740 14773
rect 3056 14764 3108 14816
rect 3332 14764 3384 14816
rect 5356 14807 5408 14816
rect 5356 14773 5365 14807
rect 5365 14773 5399 14807
rect 5399 14773 5408 14807
rect 5356 14764 5408 14773
rect 8484 14807 8536 14816
rect 8484 14773 8493 14807
rect 8493 14773 8527 14807
rect 8527 14773 8536 14807
rect 8484 14764 8536 14773
rect 8944 14764 8996 14816
rect 12716 14832 12768 14884
rect 11060 14764 11112 14816
rect 11428 14764 11480 14816
rect 11888 14764 11940 14816
rect 13820 14968 13872 15020
rect 15016 15113 15025 15147
rect 15025 15113 15059 15147
rect 15059 15113 15068 15147
rect 15016 15104 15068 15113
rect 15844 14968 15896 15020
rect 14372 14943 14424 14952
rect 14372 14909 14381 14943
rect 14381 14909 14415 14943
rect 14415 14909 14424 14943
rect 14372 14900 14424 14909
rect 12992 14764 13044 14816
rect 18604 14832 18656 14884
rect 15384 14807 15436 14816
rect 15384 14773 15393 14807
rect 15393 14773 15427 14807
rect 15427 14773 15436 14807
rect 15384 14764 15436 14773
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 1676 14603 1728 14612
rect 1676 14569 1685 14603
rect 1685 14569 1719 14603
rect 1719 14569 1728 14603
rect 1676 14560 1728 14569
rect 2228 14560 2280 14612
rect 5264 14560 5316 14612
rect 9220 14560 9272 14612
rect 9496 14560 9548 14612
rect 14004 14560 14056 14612
rect 14188 14603 14240 14612
rect 14188 14569 14197 14603
rect 14197 14569 14231 14603
rect 14231 14569 14240 14603
rect 14188 14560 14240 14569
rect 1492 14467 1544 14476
rect 1492 14433 1501 14467
rect 1501 14433 1535 14467
rect 1535 14433 1544 14467
rect 1492 14424 1544 14433
rect 2136 14424 2188 14476
rect 2320 14467 2372 14476
rect 2320 14433 2343 14467
rect 2343 14433 2372 14467
rect 2320 14424 2372 14433
rect 2596 14492 2648 14544
rect 2780 14424 2832 14476
rect 5356 14492 5408 14544
rect 8484 14492 8536 14544
rect 8760 14492 8812 14544
rect 5816 14424 5868 14476
rect 6552 14424 6604 14476
rect 6736 14467 6788 14476
rect 6736 14433 6745 14467
rect 6745 14433 6779 14467
rect 6779 14433 6788 14467
rect 6736 14424 6788 14433
rect 7840 14467 7892 14476
rect 7840 14433 7849 14467
rect 7849 14433 7883 14467
rect 7883 14433 7892 14467
rect 7840 14424 7892 14433
rect 5724 14356 5776 14408
rect 3792 14288 3844 14340
rect 7472 14356 7524 14408
rect 3516 14220 3568 14272
rect 5080 14263 5132 14272
rect 5080 14229 5089 14263
rect 5089 14229 5123 14263
rect 5123 14229 5132 14263
rect 5080 14220 5132 14229
rect 5908 14263 5960 14272
rect 5908 14229 5917 14263
rect 5917 14229 5951 14263
rect 5951 14229 5960 14263
rect 5908 14220 5960 14229
rect 6368 14263 6420 14272
rect 6368 14229 6377 14263
rect 6377 14229 6411 14263
rect 6411 14229 6420 14263
rect 6368 14220 6420 14229
rect 7104 14288 7156 14340
rect 8208 14356 8260 14408
rect 8760 14399 8812 14408
rect 8760 14365 8769 14399
rect 8769 14365 8803 14399
rect 8803 14365 8812 14399
rect 8760 14356 8812 14365
rect 9404 14424 9456 14476
rect 10416 14424 10468 14476
rect 11428 14467 11480 14476
rect 11428 14433 11462 14467
rect 11462 14433 11480 14467
rect 11428 14424 11480 14433
rect 11888 14492 11940 14544
rect 15476 14560 15528 14612
rect 15660 14603 15712 14612
rect 15660 14569 15669 14603
rect 15669 14569 15703 14603
rect 15703 14569 15712 14603
rect 15660 14560 15712 14569
rect 12900 14424 12952 14476
rect 13820 14424 13872 14476
rect 19524 14560 19576 14612
rect 9680 14356 9732 14408
rect 10508 14356 10560 14408
rect 10692 14399 10744 14408
rect 10692 14365 10701 14399
rect 10701 14365 10735 14399
rect 10735 14365 10744 14399
rect 10692 14356 10744 14365
rect 12256 14356 12308 14408
rect 7012 14220 7064 14272
rect 7840 14220 7892 14272
rect 9312 14220 9364 14272
rect 9496 14220 9548 14272
rect 12348 14220 12400 14272
rect 12532 14263 12584 14272
rect 12532 14229 12541 14263
rect 12541 14229 12575 14263
rect 12575 14229 12584 14263
rect 12532 14220 12584 14229
rect 13728 14220 13780 14272
rect 15844 14399 15896 14408
rect 15844 14365 15853 14399
rect 15853 14365 15887 14399
rect 15887 14365 15896 14399
rect 15844 14356 15896 14365
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 1768 14016 1820 14068
rect 2136 13923 2188 13932
rect 2136 13889 2145 13923
rect 2145 13889 2179 13923
rect 2179 13889 2188 13923
rect 2136 13880 2188 13889
rect 2780 14016 2832 14068
rect 3700 14016 3752 14068
rect 4160 14016 4212 14068
rect 5448 14016 5500 14068
rect 8760 14016 8812 14068
rect 9496 14016 9548 14068
rect 10048 14016 10100 14068
rect 12440 14016 12492 14068
rect 12716 14016 12768 14068
rect 13820 14059 13872 14068
rect 3516 13880 3568 13932
rect 5816 13948 5868 14000
rect 5448 13923 5500 13932
rect 5448 13889 5457 13923
rect 5457 13889 5491 13923
rect 5491 13889 5500 13923
rect 5448 13880 5500 13889
rect 6920 13880 6972 13932
rect 8116 13923 8168 13932
rect 8116 13889 8125 13923
rect 8125 13889 8159 13923
rect 8159 13889 8168 13923
rect 8116 13880 8168 13889
rect 8944 13880 8996 13932
rect 9864 13880 9916 13932
rect 9956 13923 10008 13932
rect 9956 13889 9965 13923
rect 9965 13889 9999 13923
rect 9999 13889 10008 13923
rect 9956 13880 10008 13889
rect 10232 13880 10284 13932
rect 11888 13948 11940 14000
rect 12256 13948 12308 14000
rect 13820 14025 13829 14059
rect 13829 14025 13863 14059
rect 13863 14025 13872 14059
rect 13820 14016 13872 14025
rect 10876 13923 10928 13932
rect 10876 13889 10885 13923
rect 10885 13889 10919 13923
rect 10919 13889 10928 13923
rect 10876 13880 10928 13889
rect 11060 13880 11112 13932
rect 1400 13812 1452 13864
rect 4252 13812 4304 13864
rect 3424 13744 3476 13796
rect 5080 13812 5132 13864
rect 5264 13855 5316 13864
rect 5264 13821 5273 13855
rect 5273 13821 5307 13855
rect 5307 13821 5316 13855
rect 5264 13812 5316 13821
rect 6184 13855 6236 13864
rect 6184 13821 6193 13855
rect 6193 13821 6227 13855
rect 6227 13821 6236 13855
rect 6184 13812 6236 13821
rect 6368 13812 6420 13864
rect 5540 13744 5592 13796
rect 7288 13744 7340 13796
rect 8208 13744 8260 13796
rect 9680 13744 9732 13796
rect 11152 13812 11204 13864
rect 11612 13812 11664 13864
rect 12164 13812 12216 13864
rect 12348 13812 12400 13864
rect 13544 13812 13596 13864
rect 14188 13812 14240 13864
rect 13820 13744 13872 13796
rect 3516 13676 3568 13728
rect 4712 13676 4764 13728
rect 5724 13719 5776 13728
rect 5724 13685 5733 13719
rect 5733 13685 5767 13719
rect 5767 13685 5776 13719
rect 5724 13676 5776 13685
rect 6000 13676 6052 13728
rect 7656 13676 7708 13728
rect 8760 13676 8812 13728
rect 9128 13676 9180 13728
rect 11152 13676 11204 13728
rect 11704 13676 11756 13728
rect 18696 13812 18748 13864
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 2688 13472 2740 13524
rect 3332 13515 3384 13524
rect 3332 13481 3341 13515
rect 3341 13481 3375 13515
rect 3375 13481 3384 13515
rect 3332 13472 3384 13481
rect 3608 13472 3660 13524
rect 6368 13472 6420 13524
rect 7104 13515 7156 13524
rect 7104 13481 7113 13515
rect 7113 13481 7147 13515
rect 7147 13481 7156 13515
rect 7104 13472 7156 13481
rect 8760 13472 8812 13524
rect 1492 13404 1544 13456
rect 2504 13379 2556 13388
rect 2504 13345 2513 13379
rect 2513 13345 2547 13379
rect 2547 13345 2556 13379
rect 2504 13336 2556 13345
rect 2872 13336 2924 13388
rect 3884 13336 3936 13388
rect 4160 13404 4212 13456
rect 5448 13404 5500 13456
rect 6920 13404 6972 13456
rect 8300 13404 8352 13456
rect 9772 13472 9824 13524
rect 10692 13472 10744 13524
rect 10784 13472 10836 13524
rect 11152 13472 11204 13524
rect 12440 13472 12492 13524
rect 13820 13472 13872 13524
rect 6552 13336 6604 13388
rect 7012 13336 7064 13388
rect 8208 13336 8260 13388
rect 9680 13336 9732 13388
rect 10416 13336 10468 13388
rect 2136 13268 2188 13320
rect 3700 13268 3752 13320
rect 5724 13311 5776 13320
rect 5724 13277 5733 13311
rect 5733 13277 5767 13311
rect 5767 13277 5776 13311
rect 5724 13268 5776 13277
rect 7380 13311 7432 13320
rect 7380 13277 7389 13311
rect 7389 13277 7423 13311
rect 7423 13277 7432 13311
rect 7380 13268 7432 13277
rect 8484 13268 8536 13320
rect 9772 13268 9824 13320
rect 10876 13268 10928 13320
rect 11336 13336 11388 13388
rect 11060 13268 11112 13320
rect 11152 13311 11204 13320
rect 11152 13277 11161 13311
rect 11161 13277 11195 13311
rect 11195 13277 11204 13311
rect 12256 13311 12308 13320
rect 11152 13268 11204 13277
rect 12256 13277 12265 13311
rect 12265 13277 12299 13311
rect 12299 13277 12308 13311
rect 12256 13268 12308 13277
rect 9956 13200 10008 13252
rect 12992 13336 13044 13388
rect 13728 13336 13780 13388
rect 14280 13379 14332 13388
rect 14280 13345 14289 13379
rect 14289 13345 14323 13379
rect 14323 13345 14332 13379
rect 14280 13336 14332 13345
rect 14832 13336 14884 13388
rect 15108 13336 15160 13388
rect 15292 13336 15344 13388
rect 15752 13379 15804 13388
rect 15752 13345 15761 13379
rect 15761 13345 15795 13379
rect 15795 13345 15804 13379
rect 15752 13336 15804 13345
rect 12532 13268 12584 13320
rect 14648 13268 14700 13320
rect 15844 13311 15896 13320
rect 3424 13132 3476 13184
rect 4068 13132 4120 13184
rect 5724 13132 5776 13184
rect 5908 13132 5960 13184
rect 15016 13200 15068 13252
rect 15844 13277 15853 13311
rect 15853 13277 15887 13311
rect 15887 13277 15896 13311
rect 15844 13268 15896 13277
rect 16764 13311 16816 13320
rect 16764 13277 16773 13311
rect 16773 13277 16807 13311
rect 16807 13277 16816 13311
rect 16764 13268 16816 13277
rect 10324 13132 10376 13184
rect 13544 13132 13596 13184
rect 14924 13132 14976 13184
rect 15844 13132 15896 13184
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 3148 12928 3200 12980
rect 6000 12928 6052 12980
rect 6184 12928 6236 12980
rect 7288 12928 7340 12980
rect 7656 12928 7708 12980
rect 9680 12971 9732 12980
rect 9680 12937 9689 12971
rect 9689 12937 9723 12971
rect 9723 12937 9732 12971
rect 9680 12928 9732 12937
rect 4160 12860 4212 12912
rect 9312 12860 9364 12912
rect 9864 12860 9916 12912
rect 2412 12835 2464 12844
rect 2412 12801 2421 12835
rect 2421 12801 2455 12835
rect 2455 12801 2464 12835
rect 2412 12792 2464 12801
rect 3424 12835 3476 12844
rect 3424 12801 3433 12835
rect 3433 12801 3467 12835
rect 3467 12801 3476 12835
rect 3424 12792 3476 12801
rect 3700 12792 3752 12844
rect 3332 12724 3384 12776
rect 3516 12724 3568 12776
rect 3792 12767 3844 12776
rect 3792 12733 3801 12767
rect 3801 12733 3835 12767
rect 3835 12733 3844 12767
rect 3792 12724 3844 12733
rect 3976 12792 4028 12844
rect 2964 12656 3016 12708
rect 1584 12588 1636 12640
rect 2136 12631 2188 12640
rect 2136 12597 2145 12631
rect 2145 12597 2179 12631
rect 2179 12597 2188 12631
rect 2136 12588 2188 12597
rect 2780 12631 2832 12640
rect 2780 12597 2789 12631
rect 2789 12597 2823 12631
rect 2823 12597 2832 12631
rect 3148 12631 3200 12640
rect 2780 12588 2832 12597
rect 3148 12597 3157 12631
rect 3157 12597 3191 12631
rect 3191 12597 3200 12631
rect 3148 12588 3200 12597
rect 5724 12792 5776 12844
rect 5816 12724 5868 12776
rect 9036 12792 9088 12844
rect 9496 12792 9548 12844
rect 12164 12928 12216 12980
rect 14280 12928 14332 12980
rect 15568 12971 15620 12980
rect 15568 12937 15577 12971
rect 15577 12937 15611 12971
rect 15611 12937 15620 12971
rect 15568 12928 15620 12937
rect 12348 12860 12400 12912
rect 12440 12835 12492 12844
rect 12440 12801 12449 12835
rect 12449 12801 12483 12835
rect 12483 12801 12492 12835
rect 12440 12792 12492 12801
rect 15108 12835 15160 12844
rect 15108 12801 15117 12835
rect 15117 12801 15151 12835
rect 15151 12801 15160 12835
rect 15108 12792 15160 12801
rect 5908 12656 5960 12708
rect 7012 12724 7064 12776
rect 5540 12588 5592 12640
rect 7380 12656 7432 12708
rect 9956 12724 10008 12776
rect 10416 12724 10468 12776
rect 10324 12656 10376 12708
rect 12716 12724 12768 12776
rect 11152 12656 11204 12708
rect 11612 12656 11664 12708
rect 11704 12656 11756 12708
rect 12440 12656 12492 12708
rect 13820 12656 13872 12708
rect 6184 12588 6236 12640
rect 6368 12588 6420 12640
rect 9128 12588 9180 12640
rect 9496 12588 9548 12640
rect 11888 12588 11940 12640
rect 12072 12588 12124 12640
rect 14648 12724 14700 12776
rect 14924 12767 14976 12776
rect 14924 12733 14933 12767
rect 14933 12733 14967 12767
rect 14967 12733 14976 12767
rect 14924 12724 14976 12733
rect 15016 12767 15068 12776
rect 15016 12733 15025 12767
rect 15025 12733 15059 12767
rect 15059 12733 15068 12767
rect 15016 12724 15068 12733
rect 14280 12631 14332 12640
rect 14280 12597 14289 12631
rect 14289 12597 14323 12631
rect 14323 12597 14332 12631
rect 14280 12588 14332 12597
rect 15936 12631 15988 12640
rect 15936 12597 15945 12631
rect 15945 12597 15979 12631
rect 15979 12597 15988 12631
rect 15936 12588 15988 12597
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 2136 12384 2188 12436
rect 3056 12384 3108 12436
rect 4804 12384 4856 12436
rect 9864 12384 9916 12436
rect 4436 12359 4488 12368
rect 4436 12325 4445 12359
rect 4445 12325 4479 12359
rect 4479 12325 4488 12359
rect 4436 12316 4488 12325
rect 4988 12316 5040 12368
rect 8760 12316 8812 12368
rect 10784 12384 10836 12436
rect 10968 12384 11020 12436
rect 11612 12427 11664 12436
rect 2780 12248 2832 12300
rect 3516 12248 3568 12300
rect 3424 12223 3476 12232
rect 1676 12112 1728 12164
rect 3424 12189 3433 12223
rect 3433 12189 3467 12223
rect 3467 12189 3476 12223
rect 3424 12180 3476 12189
rect 3976 12180 4028 12232
rect 5540 12248 5592 12300
rect 6184 12291 6236 12300
rect 6184 12257 6218 12291
rect 6218 12257 6236 12291
rect 6184 12248 6236 12257
rect 7104 12248 7156 12300
rect 7564 12248 7616 12300
rect 9220 12248 9272 12300
rect 4804 12180 4856 12232
rect 5172 12180 5224 12232
rect 8576 12223 8628 12232
rect 8576 12189 8585 12223
rect 8585 12189 8619 12223
rect 8619 12189 8628 12223
rect 8576 12180 8628 12189
rect 9864 12180 9916 12232
rect 10416 12316 10468 12368
rect 10692 12316 10744 12368
rect 11612 12393 11621 12427
rect 11621 12393 11655 12427
rect 11655 12393 11664 12427
rect 11612 12384 11664 12393
rect 11888 12427 11940 12436
rect 11888 12393 11897 12427
rect 11897 12393 11931 12427
rect 11931 12393 11940 12427
rect 11888 12384 11940 12393
rect 13820 12384 13872 12436
rect 15108 12384 15160 12436
rect 11060 12248 11112 12300
rect 14280 12316 14332 12368
rect 14556 12248 14608 12300
rect 12348 12223 12400 12232
rect 12348 12189 12357 12223
rect 12357 12189 12391 12223
rect 12391 12189 12400 12223
rect 12348 12180 12400 12189
rect 3700 12112 3752 12164
rect 4252 12112 4304 12164
rect 7196 12112 7248 12164
rect 7564 12112 7616 12164
rect 7288 12087 7340 12096
rect 7288 12053 7297 12087
rect 7297 12053 7331 12087
rect 7331 12053 7340 12087
rect 7288 12044 7340 12053
rect 7380 12044 7432 12096
rect 11612 12112 11664 12164
rect 12532 12180 12584 12232
rect 11704 12044 11756 12096
rect 14464 12044 14516 12096
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 3976 11840 4028 11892
rect 4160 11840 4212 11892
rect 6736 11840 6788 11892
rect 7012 11840 7064 11892
rect 7472 11840 7524 11892
rect 10048 11840 10100 11892
rect 10600 11840 10652 11892
rect 10692 11840 10744 11892
rect 12348 11840 12400 11892
rect 3424 11772 3476 11824
rect 3700 11815 3752 11824
rect 3700 11781 3709 11815
rect 3709 11781 3743 11815
rect 3743 11781 3752 11815
rect 3700 11772 3752 11781
rect 1584 11679 1636 11688
rect 1584 11645 1593 11679
rect 1593 11645 1627 11679
rect 1627 11645 1636 11679
rect 1584 11636 1636 11645
rect 2228 11636 2280 11688
rect 4804 11704 4856 11756
rect 5172 11704 5224 11756
rect 7104 11772 7156 11824
rect 7748 11772 7800 11824
rect 13636 11840 13688 11892
rect 13820 11883 13872 11892
rect 13820 11849 13829 11883
rect 13829 11849 13863 11883
rect 13863 11849 13872 11883
rect 13820 11840 13872 11849
rect 15936 11840 15988 11892
rect 6920 11704 6972 11756
rect 3700 11636 3752 11688
rect 5908 11636 5960 11688
rect 6000 11568 6052 11620
rect 8484 11704 8536 11756
rect 9588 11704 9640 11756
rect 10324 11704 10376 11756
rect 11060 11704 11112 11756
rect 12440 11747 12492 11756
rect 12440 11713 12449 11747
rect 12449 11713 12483 11747
rect 12483 11713 12492 11747
rect 12440 11704 12492 11713
rect 13820 11704 13872 11756
rect 17224 11704 17276 11756
rect 12348 11636 12400 11688
rect 8484 11568 8536 11620
rect 5448 11500 5500 11552
rect 6460 11500 6512 11552
rect 7472 11500 7524 11552
rect 9312 11500 9364 11552
rect 9404 11500 9456 11552
rect 10324 11500 10376 11552
rect 12624 11568 12676 11620
rect 13360 11568 13412 11620
rect 14096 11636 14148 11688
rect 17040 11568 17092 11620
rect 13912 11500 13964 11552
rect 14280 11500 14332 11552
rect 15108 11500 15160 11552
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 2412 11296 2464 11348
rect 4068 11339 4120 11348
rect 4068 11305 4077 11339
rect 4077 11305 4111 11339
rect 4111 11305 4120 11339
rect 4068 11296 4120 11305
rect 5356 11296 5408 11348
rect 7380 11296 7432 11348
rect 1676 11271 1728 11280
rect 1676 11237 1710 11271
rect 1710 11237 1728 11271
rect 1676 11228 1728 11237
rect 3792 11228 3844 11280
rect 2228 11160 2280 11212
rect 3056 11203 3108 11212
rect 3056 11169 3065 11203
rect 3065 11169 3099 11203
rect 3099 11169 3108 11203
rect 3056 11160 3108 11169
rect 3608 11160 3660 11212
rect 7472 11228 7524 11280
rect 5816 11160 5868 11212
rect 4252 11092 4304 11144
rect 9588 11296 9640 11348
rect 9680 11296 9732 11348
rect 11060 11339 11112 11348
rect 11060 11305 11069 11339
rect 11069 11305 11103 11339
rect 11103 11305 11112 11339
rect 11060 11296 11112 11305
rect 11704 11296 11756 11348
rect 12716 11296 12768 11348
rect 12900 11296 12952 11348
rect 14096 11339 14148 11348
rect 14096 11305 14105 11339
rect 14105 11305 14139 11339
rect 14139 11305 14148 11339
rect 14096 11296 14148 11305
rect 8576 11228 8628 11280
rect 6184 11067 6236 11076
rect 6184 11033 6193 11067
rect 6193 11033 6227 11067
rect 6227 11033 6236 11067
rect 6184 11024 6236 11033
rect 3976 10956 4028 11008
rect 7012 10956 7064 11008
rect 7748 11024 7800 11076
rect 8760 11160 8812 11212
rect 9588 11160 9640 11212
rect 11704 11203 11756 11212
rect 11704 11169 11738 11203
rect 11738 11169 11756 11203
rect 11704 11160 11756 11169
rect 12440 11160 12492 11212
rect 13176 11160 13228 11212
rect 11060 11092 11112 11144
rect 13636 11135 13688 11144
rect 13636 11101 13645 11135
rect 13645 11101 13679 11135
rect 13679 11101 13688 11135
rect 13636 11092 13688 11101
rect 13820 11160 13872 11212
rect 12716 11024 12768 11076
rect 14004 11092 14056 11144
rect 14648 11135 14700 11144
rect 14648 11101 14657 11135
rect 14657 11101 14691 11135
rect 14691 11101 14700 11135
rect 14648 11092 14700 11101
rect 17132 11024 17184 11076
rect 8668 10956 8720 11008
rect 10876 10956 10928 11008
rect 11612 10956 11664 11008
rect 16764 10956 16816 11008
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 4068 10752 4120 10804
rect 5816 10727 5868 10736
rect 5816 10693 5825 10727
rect 5825 10693 5859 10727
rect 5859 10693 5868 10727
rect 5816 10684 5868 10693
rect 6920 10684 6972 10736
rect 7196 10684 7248 10736
rect 8576 10752 8628 10804
rect 8760 10752 8812 10804
rect 10876 10752 10928 10804
rect 12992 10752 13044 10804
rect 3148 10616 3200 10668
rect 12808 10684 12860 10736
rect 13084 10684 13136 10736
rect 2136 10548 2188 10600
rect 4252 10548 4304 10600
rect 6368 10548 6420 10600
rect 8668 10616 8720 10668
rect 9220 10659 9272 10668
rect 8576 10548 8628 10600
rect 9220 10625 9229 10659
rect 9229 10625 9263 10659
rect 9263 10625 9272 10659
rect 9220 10616 9272 10625
rect 11244 10616 11296 10668
rect 12992 10616 13044 10668
rect 9680 10591 9732 10600
rect 9680 10557 9689 10591
rect 9689 10557 9723 10591
rect 9723 10557 9732 10591
rect 9680 10548 9732 10557
rect 9956 10591 10008 10600
rect 9956 10557 9990 10591
rect 9990 10557 10008 10591
rect 9956 10548 10008 10557
rect 10232 10548 10284 10600
rect 14280 10752 14332 10804
rect 13360 10616 13412 10668
rect 14004 10659 14056 10668
rect 14004 10625 14013 10659
rect 14013 10625 14047 10659
rect 14047 10625 14056 10659
rect 14004 10616 14056 10625
rect 13452 10548 13504 10600
rect 2412 10480 2464 10532
rect 5724 10480 5776 10532
rect 7656 10480 7708 10532
rect 8668 10480 8720 10532
rect 4988 10412 5040 10464
rect 7196 10412 7248 10464
rect 7288 10412 7340 10464
rect 8208 10412 8260 10464
rect 8852 10412 8904 10464
rect 9220 10412 9272 10464
rect 9772 10412 9824 10464
rect 9956 10412 10008 10464
rect 11152 10455 11204 10464
rect 11152 10421 11161 10455
rect 11161 10421 11195 10455
rect 11195 10421 11204 10455
rect 11152 10412 11204 10421
rect 11520 10455 11572 10464
rect 11520 10421 11529 10455
rect 11529 10421 11563 10455
rect 11563 10421 11572 10455
rect 11520 10412 11572 10421
rect 11980 10455 12032 10464
rect 11980 10421 11989 10455
rect 11989 10421 12023 10455
rect 12023 10421 12032 10455
rect 11980 10412 12032 10421
rect 12900 10412 12952 10464
rect 16580 10412 16632 10464
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 3240 10140 3292 10192
rect 3424 10208 3476 10260
rect 4712 10208 4764 10260
rect 7472 10208 7524 10260
rect 8668 10208 8720 10260
rect 9680 10208 9732 10260
rect 7380 10140 7432 10192
rect 8208 10140 8260 10192
rect 10508 10140 10560 10192
rect 11060 10208 11112 10260
rect 11704 10208 11756 10260
rect 12900 10251 12952 10260
rect 11244 10140 11296 10192
rect 11520 10140 11572 10192
rect 12900 10217 12909 10251
rect 12909 10217 12943 10251
rect 12943 10217 12952 10251
rect 12900 10208 12952 10217
rect 15108 10208 15160 10260
rect 12532 10140 12584 10192
rect 2872 10072 2924 10124
rect 3424 10072 3476 10124
rect 3700 10072 3752 10124
rect 4804 10072 4856 10124
rect 5080 10072 5132 10124
rect 6368 10115 6420 10124
rect 6368 10081 6377 10115
rect 6377 10081 6411 10115
rect 6411 10081 6420 10115
rect 6368 10072 6420 10081
rect 6460 10072 6512 10124
rect 8852 10072 8904 10124
rect 10324 10072 10376 10124
rect 10600 10115 10652 10124
rect 10600 10081 10609 10115
rect 10609 10081 10643 10115
rect 10643 10081 10652 10115
rect 10600 10072 10652 10081
rect 10692 10072 10744 10124
rect 2228 10004 2280 10056
rect 4988 10004 5040 10056
rect 5724 10047 5776 10056
rect 5724 10013 5733 10047
rect 5733 10013 5767 10047
rect 5767 10013 5776 10047
rect 5724 10004 5776 10013
rect 8300 10004 8352 10056
rect 8760 10047 8812 10056
rect 8760 10013 8769 10047
rect 8769 10013 8803 10047
rect 8803 10013 8812 10047
rect 8760 10004 8812 10013
rect 10508 10004 10560 10056
rect 12624 10072 12676 10124
rect 14464 10072 14516 10124
rect 13728 10047 13780 10056
rect 13728 10013 13737 10047
rect 13737 10013 13771 10047
rect 13771 10013 13780 10047
rect 13728 10004 13780 10013
rect 14004 10004 14056 10056
rect 5816 9936 5868 9988
rect 3792 9868 3844 9920
rect 7748 9868 7800 9920
rect 12072 9936 12124 9988
rect 12256 9936 12308 9988
rect 13084 9868 13136 9920
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 4344 9596 4396 9648
rect 5264 9664 5316 9716
rect 6368 9664 6420 9716
rect 6460 9639 6512 9648
rect 2596 9571 2648 9580
rect 2596 9537 2605 9571
rect 2605 9537 2639 9571
rect 2639 9537 2648 9571
rect 2596 9528 2648 9537
rect 2688 9528 2740 9580
rect 4988 9528 5040 9580
rect 6460 9605 6469 9639
rect 6469 9605 6503 9639
rect 6503 9605 6512 9639
rect 6460 9596 6512 9605
rect 3700 9460 3752 9512
rect 4896 9460 4948 9512
rect 8300 9596 8352 9648
rect 7196 9503 7248 9512
rect 3056 9392 3108 9444
rect 4160 9392 4212 9444
rect 7196 9469 7205 9503
rect 7205 9469 7239 9503
rect 7239 9469 7248 9503
rect 7196 9460 7248 9469
rect 8208 9528 8260 9580
rect 8668 9571 8720 9580
rect 8668 9537 8677 9571
rect 8677 9537 8711 9571
rect 8711 9537 8720 9571
rect 8668 9528 8720 9537
rect 9772 9528 9824 9580
rect 10692 9528 10744 9580
rect 11244 9528 11296 9580
rect 7472 9460 7524 9512
rect 9404 9460 9456 9512
rect 9588 9460 9640 9512
rect 10508 9460 10560 9512
rect 6460 9392 6512 9444
rect 2320 9367 2372 9376
rect 2320 9333 2329 9367
rect 2329 9333 2363 9367
rect 2363 9333 2372 9367
rect 2320 9324 2372 9333
rect 2412 9367 2464 9376
rect 2412 9333 2421 9367
rect 2421 9333 2455 9367
rect 2455 9333 2464 9367
rect 2964 9367 3016 9376
rect 2412 9324 2464 9333
rect 2964 9333 2973 9367
rect 2973 9333 3007 9367
rect 3007 9333 3016 9367
rect 2964 9324 3016 9333
rect 3332 9367 3384 9376
rect 3332 9333 3341 9367
rect 3341 9333 3375 9367
rect 3375 9333 3384 9367
rect 3332 9324 3384 9333
rect 3516 9324 3568 9376
rect 4252 9324 4304 9376
rect 6276 9324 6328 9376
rect 9496 9392 9548 9444
rect 7012 9324 7064 9376
rect 7196 9324 7248 9376
rect 7748 9324 7800 9376
rect 8300 9324 8352 9376
rect 8576 9367 8628 9376
rect 8576 9333 8585 9367
rect 8585 9333 8619 9367
rect 8619 9333 8628 9367
rect 8576 9324 8628 9333
rect 9404 9324 9456 9376
rect 9680 9324 9732 9376
rect 10048 9324 10100 9376
rect 11428 9367 11480 9376
rect 11428 9333 11437 9367
rect 11437 9333 11471 9367
rect 11471 9333 11480 9367
rect 11428 9324 11480 9333
rect 11704 9528 11756 9580
rect 12992 9571 13044 9580
rect 12992 9537 13001 9571
rect 13001 9537 13035 9571
rect 13035 9537 13044 9571
rect 12992 9528 13044 9537
rect 13084 9528 13136 9580
rect 13176 9460 13228 9512
rect 13820 9392 13872 9444
rect 14280 9392 14332 9444
rect 13636 9367 13688 9376
rect 13636 9333 13645 9367
rect 13645 9333 13679 9367
rect 13679 9333 13688 9367
rect 13636 9324 13688 9333
rect 14096 9367 14148 9376
rect 14096 9333 14105 9367
rect 14105 9333 14139 9367
rect 14139 9333 14148 9367
rect 14096 9324 14148 9333
rect 14556 9367 14608 9376
rect 14556 9333 14565 9367
rect 14565 9333 14599 9367
rect 14599 9333 14608 9367
rect 14556 9324 14608 9333
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 2228 9120 2280 9172
rect 4344 9120 4396 9172
rect 6828 9120 6880 9172
rect 7472 9163 7524 9172
rect 7472 9129 7481 9163
rect 7481 9129 7515 9163
rect 7515 9129 7524 9163
rect 7472 9120 7524 9129
rect 1492 8984 1544 9036
rect 2688 9052 2740 9104
rect 3056 9052 3108 9104
rect 3424 9052 3476 9104
rect 4068 8984 4120 9036
rect 5632 8984 5684 9036
rect 6736 8984 6788 9036
rect 7472 8984 7524 9036
rect 7656 8984 7708 9036
rect 7932 9027 7984 9036
rect 7932 8993 7941 9027
rect 7941 8993 7975 9027
rect 7975 8993 7984 9027
rect 7932 8984 7984 8993
rect 9496 9120 9548 9172
rect 11704 9163 11756 9172
rect 11704 9129 11713 9163
rect 11713 9129 11747 9163
rect 11747 9129 11756 9163
rect 11704 9120 11756 9129
rect 8392 9052 8444 9104
rect 11520 9052 11572 9104
rect 12256 9052 12308 9104
rect 8116 8984 8168 9036
rect 8208 8984 8260 9036
rect 4896 8959 4948 8968
rect 4896 8925 4905 8959
rect 4905 8925 4939 8959
rect 4939 8925 4948 8959
rect 4896 8916 4948 8925
rect 5172 8916 5224 8968
rect 6000 8959 6052 8968
rect 6000 8925 6009 8959
rect 6009 8925 6043 8959
rect 6043 8925 6052 8959
rect 6000 8916 6052 8925
rect 6920 8959 6972 8968
rect 6920 8925 6929 8959
rect 6929 8925 6963 8959
rect 6963 8925 6972 8959
rect 6920 8916 6972 8925
rect 9312 8984 9364 9036
rect 10048 9027 10100 9036
rect 10048 8993 10057 9027
rect 10057 8993 10091 9027
rect 10091 8993 10100 9027
rect 10048 8984 10100 8993
rect 11612 8984 11664 9036
rect 11980 8984 12032 9036
rect 12348 8984 12400 9036
rect 13084 9027 13136 9036
rect 13084 8993 13093 9027
rect 13093 8993 13127 9027
rect 13127 8993 13136 9027
rect 13084 8984 13136 8993
rect 5356 8848 5408 8900
rect 9680 8916 9732 8968
rect 10232 8959 10284 8968
rect 10232 8925 10241 8959
rect 10241 8925 10275 8959
rect 10275 8925 10284 8959
rect 10232 8916 10284 8925
rect 10784 8848 10836 8900
rect 11244 8959 11296 8968
rect 11244 8925 11253 8959
rect 11253 8925 11287 8959
rect 11287 8925 11296 8959
rect 11244 8916 11296 8925
rect 13636 9052 13688 9104
rect 13820 9052 13872 9104
rect 15108 9052 15160 9104
rect 13544 8984 13596 9036
rect 3424 8823 3476 8832
rect 3424 8789 3433 8823
rect 3433 8789 3467 8823
rect 3467 8789 3476 8823
rect 3424 8780 3476 8789
rect 5448 8823 5500 8832
rect 5448 8789 5457 8823
rect 5457 8789 5491 8823
rect 5491 8789 5500 8823
rect 5448 8780 5500 8789
rect 6368 8780 6420 8832
rect 7380 8780 7432 8832
rect 8760 8780 8812 8832
rect 9588 8780 9640 8832
rect 10048 8780 10100 8832
rect 10692 8823 10744 8832
rect 10692 8789 10701 8823
rect 10701 8789 10735 8823
rect 10735 8789 10744 8823
rect 10692 8780 10744 8789
rect 14280 8959 14332 8968
rect 13268 8848 13320 8900
rect 14280 8925 14289 8959
rect 14289 8925 14323 8959
rect 14323 8925 14332 8959
rect 14280 8916 14332 8925
rect 15292 8848 15344 8900
rect 14924 8780 14976 8832
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 2412 8576 2464 8628
rect 4068 8619 4120 8628
rect 4068 8585 4077 8619
rect 4077 8585 4111 8619
rect 4111 8585 4120 8619
rect 4068 8576 4120 8585
rect 6460 8619 6512 8628
rect 2596 8508 2648 8560
rect 3976 8508 4028 8560
rect 6460 8585 6469 8619
rect 6469 8585 6503 8619
rect 6503 8585 6512 8619
rect 6460 8576 6512 8585
rect 9680 8576 9732 8628
rect 9956 8576 10008 8628
rect 14556 8576 14608 8628
rect 10324 8551 10376 8560
rect 3516 8483 3568 8492
rect 3516 8449 3525 8483
rect 3525 8449 3559 8483
rect 3559 8449 3568 8483
rect 3516 8440 3568 8449
rect 1492 8372 1544 8424
rect 2688 8372 2740 8424
rect 3424 8372 3476 8424
rect 4160 8440 4212 8492
rect 4804 8440 4856 8492
rect 10324 8517 10333 8551
rect 10333 8517 10367 8551
rect 10367 8517 10376 8551
rect 10324 8508 10376 8517
rect 3792 8304 3844 8356
rect 8668 8415 8720 8424
rect 8668 8381 8677 8415
rect 8677 8381 8711 8415
rect 8711 8381 8720 8415
rect 8668 8372 8720 8381
rect 9772 8440 9824 8492
rect 10600 8440 10652 8492
rect 11980 8440 12032 8492
rect 13820 8508 13872 8560
rect 18512 8508 18564 8560
rect 13268 8440 13320 8492
rect 14924 8483 14976 8492
rect 14924 8449 14933 8483
rect 14933 8449 14967 8483
rect 14967 8449 14976 8483
rect 14924 8440 14976 8449
rect 9680 8372 9732 8424
rect 5724 8304 5776 8356
rect 7288 8347 7340 8356
rect 7288 8313 7322 8347
rect 7322 8313 7340 8347
rect 7288 8304 7340 8313
rect 7748 8304 7800 8356
rect 13912 8372 13964 8424
rect 14096 8372 14148 8424
rect 10692 8304 10744 8356
rect 4160 8236 4212 8288
rect 5264 8236 5316 8288
rect 8944 8236 8996 8288
rect 9404 8236 9456 8288
rect 11704 8304 11756 8356
rect 11060 8236 11112 8288
rect 11888 8236 11940 8288
rect 12532 8236 12584 8288
rect 13912 8279 13964 8288
rect 13912 8245 13921 8279
rect 13921 8245 13955 8279
rect 13955 8245 13964 8279
rect 13912 8236 13964 8245
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 2320 8032 2372 8084
rect 2964 8032 3016 8084
rect 3332 8032 3384 8084
rect 4896 8032 4948 8084
rect 6552 8032 6604 8084
rect 6920 8032 6972 8084
rect 4068 7964 4120 8016
rect 5080 7964 5132 8016
rect 6276 7964 6328 8016
rect 8484 7964 8536 8016
rect 9956 8007 10008 8016
rect 9956 7973 9990 8007
rect 9990 7973 10008 8007
rect 11980 8007 12032 8016
rect 9956 7964 10008 7973
rect 11980 7973 12014 8007
rect 12014 7973 12032 8007
rect 11980 7964 12032 7973
rect 3976 7896 4028 7948
rect 6000 7896 6052 7948
rect 2688 7871 2740 7880
rect 2688 7837 2697 7871
rect 2697 7837 2731 7871
rect 2731 7837 2740 7871
rect 4712 7871 4764 7880
rect 2688 7828 2740 7837
rect 4712 7837 4721 7871
rect 4721 7837 4755 7871
rect 4755 7837 4764 7871
rect 4712 7828 4764 7837
rect 4896 7871 4948 7880
rect 4896 7837 4905 7871
rect 4905 7837 4939 7871
rect 4939 7837 4948 7871
rect 4896 7828 4948 7837
rect 5448 7760 5500 7812
rect 6276 7828 6328 7880
rect 7012 7828 7064 7880
rect 7104 7828 7156 7880
rect 8392 7896 8444 7948
rect 8576 7896 8628 7948
rect 9680 7939 9732 7948
rect 9680 7905 9689 7939
rect 9689 7905 9723 7939
rect 9723 7905 9732 7939
rect 13636 8007 13688 8016
rect 13636 7973 13648 8007
rect 13648 7973 13688 8007
rect 13636 7964 13688 7973
rect 9680 7896 9732 7905
rect 17408 7896 17460 7948
rect 8024 7871 8076 7880
rect 8024 7837 8033 7871
rect 8033 7837 8067 7871
rect 8067 7837 8076 7871
rect 8024 7828 8076 7837
rect 8668 7828 8720 7880
rect 9220 7871 9272 7880
rect 9220 7837 9229 7871
rect 9229 7837 9263 7871
rect 9263 7837 9272 7871
rect 9220 7828 9272 7837
rect 11612 7828 11664 7880
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 8392 7760 8444 7812
rect 7196 7692 7248 7744
rect 9588 7692 9640 7744
rect 13544 7692 13596 7744
rect 14004 7692 14056 7744
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 1860 7352 1912 7404
rect 2872 7352 2924 7404
rect 4160 7395 4212 7404
rect 4160 7361 4169 7395
rect 4169 7361 4203 7395
rect 4203 7361 4212 7395
rect 4160 7352 4212 7361
rect 5264 7488 5316 7540
rect 5356 7488 5408 7540
rect 7748 7488 7800 7540
rect 8576 7531 8628 7540
rect 8576 7497 8585 7531
rect 8585 7497 8619 7531
rect 8619 7497 8628 7531
rect 8576 7488 8628 7497
rect 5724 7420 5776 7472
rect 8024 7420 8076 7472
rect 1400 7284 1452 7336
rect 5172 7284 5224 7336
rect 9956 7420 10008 7472
rect 9588 7352 9640 7404
rect 10048 7395 10100 7404
rect 10048 7361 10057 7395
rect 10057 7361 10091 7395
rect 10091 7361 10100 7395
rect 10048 7352 10100 7361
rect 10508 7352 10560 7404
rect 10600 7352 10652 7404
rect 7196 7327 7248 7336
rect 7196 7293 7205 7327
rect 7205 7293 7239 7327
rect 7239 7293 7248 7327
rect 7196 7284 7248 7293
rect 7288 7284 7340 7336
rect 10324 7284 10376 7336
rect 11428 7420 11480 7472
rect 12532 7420 12584 7472
rect 13360 7420 13412 7472
rect 14372 7420 14424 7472
rect 11980 7395 12032 7404
rect 11980 7361 11989 7395
rect 11989 7361 12023 7395
rect 12023 7361 12032 7395
rect 11980 7352 12032 7361
rect 12348 7352 12400 7404
rect 13636 7352 13688 7404
rect 14096 7352 14148 7404
rect 2504 7216 2556 7268
rect 4068 7216 4120 7268
rect 13820 7259 13872 7268
rect 1952 7191 2004 7200
rect 1952 7157 1961 7191
rect 1961 7157 1995 7191
rect 1995 7157 2004 7191
rect 1952 7148 2004 7157
rect 2964 7191 3016 7200
rect 2964 7157 2973 7191
rect 2973 7157 3007 7191
rect 3007 7157 3016 7191
rect 2964 7148 3016 7157
rect 3332 7191 3384 7200
rect 3332 7157 3341 7191
rect 3341 7157 3375 7191
rect 3375 7157 3384 7191
rect 3332 7148 3384 7157
rect 3424 7191 3476 7200
rect 3424 7157 3433 7191
rect 3433 7157 3467 7191
rect 3467 7157 3476 7191
rect 6000 7191 6052 7200
rect 3424 7148 3476 7157
rect 6000 7157 6009 7191
rect 6009 7157 6043 7191
rect 6043 7157 6052 7191
rect 6000 7148 6052 7157
rect 6184 7148 6236 7200
rect 6552 7148 6604 7200
rect 7104 7148 7156 7200
rect 7288 7191 7340 7200
rect 7288 7157 7297 7191
rect 7297 7157 7331 7191
rect 7331 7157 7340 7191
rect 7288 7148 7340 7157
rect 9312 7148 9364 7200
rect 10416 7148 10468 7200
rect 10692 7148 10744 7200
rect 12808 7191 12860 7200
rect 12808 7157 12817 7191
rect 12817 7157 12851 7191
rect 12851 7157 12860 7191
rect 12808 7148 12860 7157
rect 13176 7148 13228 7200
rect 13820 7225 13829 7259
rect 13829 7225 13863 7259
rect 13863 7225 13872 7259
rect 13820 7216 13872 7225
rect 14280 7216 14332 7268
rect 13912 7148 13964 7200
rect 14464 7191 14516 7200
rect 14464 7157 14473 7191
rect 14473 7157 14507 7191
rect 14507 7157 14516 7191
rect 14464 7148 14516 7157
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 2872 6944 2924 6996
rect 5172 6944 5224 6996
rect 6828 6944 6880 6996
rect 8576 6987 8628 6996
rect 8576 6953 8585 6987
rect 8585 6953 8619 6987
rect 8619 6953 8628 6987
rect 8576 6944 8628 6953
rect 4896 6876 4948 6928
rect 6920 6876 6972 6928
rect 8208 6876 8260 6928
rect 8668 6876 8720 6928
rect 10784 6944 10836 6996
rect 11060 6944 11112 6996
rect 12348 6944 12400 6996
rect 13912 6944 13964 6996
rect 14464 6944 14516 6996
rect 11428 6876 11480 6928
rect 13360 6876 13412 6928
rect 18512 6876 18564 6928
rect 1768 6808 1820 6860
rect 2228 6808 2280 6860
rect 4712 6808 4764 6860
rect 6000 6808 6052 6860
rect 9588 6851 9640 6860
rect 2688 6740 2740 6792
rect 9588 6817 9597 6851
rect 9597 6817 9631 6851
rect 9631 6817 9640 6851
rect 9588 6808 9640 6817
rect 7104 6740 7156 6792
rect 8944 6740 8996 6792
rect 9680 6783 9732 6792
rect 9680 6749 9689 6783
rect 9689 6749 9723 6783
rect 9723 6749 9732 6783
rect 9680 6740 9732 6749
rect 9588 6672 9640 6724
rect 11704 6808 11756 6860
rect 11888 6851 11940 6860
rect 11888 6817 11922 6851
rect 11922 6817 11940 6851
rect 11888 6808 11940 6817
rect 11612 6783 11664 6792
rect 11612 6749 11621 6783
rect 11621 6749 11655 6783
rect 11655 6749 11664 6783
rect 11612 6740 11664 6749
rect 7196 6604 7248 6656
rect 7380 6604 7432 6656
rect 9220 6604 9272 6656
rect 11152 6604 11204 6656
rect 12900 6740 12952 6792
rect 13084 6740 13136 6792
rect 13820 6740 13872 6792
rect 14280 6740 14332 6792
rect 14556 6740 14608 6792
rect 17500 6740 17552 6792
rect 15292 6647 15344 6656
rect 15292 6613 15301 6647
rect 15301 6613 15335 6647
rect 15335 6613 15344 6647
rect 15292 6604 15344 6613
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 3424 6400 3476 6452
rect 7288 6400 7340 6452
rect 3608 6332 3660 6384
rect 6920 6332 6972 6384
rect 7196 6332 7248 6384
rect 7656 6400 7708 6452
rect 1860 6239 1912 6248
rect 1860 6205 1894 6239
rect 1894 6205 1912 6239
rect 1860 6196 1912 6205
rect 2872 6196 2924 6248
rect 1768 6128 1820 6180
rect 2228 6060 2280 6112
rect 5264 6264 5316 6316
rect 6276 6307 6328 6316
rect 5448 6239 5500 6248
rect 5448 6205 5457 6239
rect 5457 6205 5491 6239
rect 5491 6205 5500 6239
rect 6276 6273 6285 6307
rect 6285 6273 6319 6307
rect 6319 6273 6328 6307
rect 6276 6264 6328 6273
rect 6644 6264 6696 6316
rect 5448 6196 5500 6205
rect 6920 6196 6972 6248
rect 7288 6264 7340 6316
rect 10600 6400 10652 6452
rect 19156 6400 19208 6452
rect 9220 6375 9272 6384
rect 9220 6341 9229 6375
rect 9229 6341 9263 6375
rect 9263 6341 9272 6375
rect 9220 6332 9272 6341
rect 11152 6332 11204 6384
rect 11336 6332 11388 6384
rect 10140 6264 10192 6316
rect 11060 6264 11112 6316
rect 12716 6332 12768 6384
rect 12256 6264 12308 6316
rect 13176 6264 13228 6316
rect 13268 6264 13320 6316
rect 7472 6196 7524 6248
rect 9128 6196 9180 6248
rect 10416 6196 10468 6248
rect 13452 6196 13504 6248
rect 15200 6239 15252 6248
rect 15200 6205 15209 6239
rect 15209 6205 15243 6239
rect 15243 6205 15252 6239
rect 15200 6196 15252 6205
rect 6552 6128 6604 6180
rect 7932 6128 7984 6180
rect 8024 6128 8076 6180
rect 3608 6103 3660 6112
rect 3608 6069 3617 6103
rect 3617 6069 3651 6103
rect 3651 6069 3660 6103
rect 3608 6060 3660 6069
rect 4620 6103 4672 6112
rect 4620 6069 4629 6103
rect 4629 6069 4663 6103
rect 4663 6069 4672 6103
rect 4620 6060 4672 6069
rect 5356 6060 5408 6112
rect 6092 6103 6144 6112
rect 6092 6069 6101 6103
rect 6101 6069 6135 6103
rect 6135 6069 6144 6103
rect 6092 6060 6144 6069
rect 8208 6128 8260 6180
rect 12532 6128 12584 6180
rect 12624 6128 12676 6180
rect 14004 6128 14056 6180
rect 10232 6060 10284 6112
rect 10324 6060 10376 6112
rect 10600 6060 10652 6112
rect 10968 6060 11020 6112
rect 12716 6060 12768 6112
rect 13728 6060 13780 6112
rect 15016 6060 15068 6112
rect 15568 6060 15620 6112
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 1952 5856 2004 5908
rect 3608 5856 3660 5908
rect 4620 5856 4672 5908
rect 5448 5856 5500 5908
rect 6276 5856 6328 5908
rect 6368 5856 6420 5908
rect 10324 5856 10376 5908
rect 10968 5899 11020 5908
rect 2780 5788 2832 5840
rect 6920 5788 6972 5840
rect 7288 5788 7340 5840
rect 9220 5788 9272 5840
rect 9588 5788 9640 5840
rect 10968 5865 10977 5899
rect 10977 5865 11011 5899
rect 11011 5865 11020 5899
rect 10968 5856 11020 5865
rect 13084 5856 13136 5908
rect 14556 5899 14608 5908
rect 14556 5865 14565 5899
rect 14565 5865 14599 5899
rect 14599 5865 14608 5899
rect 14556 5856 14608 5865
rect 17408 5899 17460 5908
rect 17408 5865 17417 5899
rect 17417 5865 17451 5899
rect 17451 5865 17460 5899
rect 17408 5856 17460 5865
rect 15568 5831 15620 5840
rect 2688 5720 2740 5772
rect 2872 5720 2924 5772
rect 2228 5695 2280 5704
rect 2228 5661 2237 5695
rect 2237 5661 2271 5695
rect 2271 5661 2280 5695
rect 2228 5652 2280 5661
rect 2964 5652 3016 5704
rect 5264 5720 5316 5772
rect 15568 5797 15602 5831
rect 15602 5797 15620 5831
rect 15568 5788 15620 5797
rect 12256 5720 12308 5772
rect 12624 5720 12676 5772
rect 13452 5720 13504 5772
rect 15200 5720 15252 5772
rect 15384 5720 15436 5772
rect 17960 5720 18012 5772
rect 3332 5584 3384 5636
rect 5816 5652 5868 5704
rect 6276 5652 6328 5704
rect 6828 5652 6880 5704
rect 11060 5695 11112 5704
rect 11060 5661 11069 5695
rect 11069 5661 11103 5695
rect 11103 5661 11112 5695
rect 11060 5652 11112 5661
rect 11612 5695 11664 5704
rect 6644 5584 6696 5636
rect 2964 5516 3016 5568
rect 3976 5516 4028 5568
rect 4712 5516 4764 5568
rect 5356 5516 5408 5568
rect 6828 5516 6880 5568
rect 9496 5584 9548 5636
rect 11336 5584 11388 5636
rect 8852 5516 8904 5568
rect 11612 5661 11621 5695
rect 11621 5661 11655 5695
rect 11655 5661 11664 5695
rect 11612 5652 11664 5661
rect 13268 5695 13320 5704
rect 13268 5661 13277 5695
rect 13277 5661 13311 5695
rect 13311 5661 13320 5695
rect 13268 5652 13320 5661
rect 15016 5652 15068 5704
rect 17500 5695 17552 5704
rect 17500 5661 17509 5695
rect 17509 5661 17543 5695
rect 17543 5661 17552 5695
rect 17500 5652 17552 5661
rect 19800 5652 19852 5704
rect 11888 5516 11940 5568
rect 15476 5516 15528 5568
rect 16948 5559 17000 5568
rect 16948 5525 16957 5559
rect 16957 5525 16991 5559
rect 16991 5525 17000 5559
rect 16948 5516 17000 5525
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 4068 5312 4120 5364
rect 5724 5312 5776 5364
rect 8484 5355 8536 5364
rect 8484 5321 8493 5355
rect 8493 5321 8527 5355
rect 8527 5321 8536 5355
rect 8484 5312 8536 5321
rect 11060 5312 11112 5364
rect 12532 5355 12584 5364
rect 12532 5321 12541 5355
rect 12541 5321 12575 5355
rect 12575 5321 12584 5355
rect 12532 5312 12584 5321
rect 12900 5244 12952 5296
rect 3884 5219 3936 5228
rect 3884 5185 3893 5219
rect 3893 5185 3927 5219
rect 3927 5185 3936 5219
rect 3884 5176 3936 5185
rect 8208 5176 8260 5228
rect 9128 5219 9180 5228
rect 9128 5185 9137 5219
rect 9137 5185 9171 5219
rect 9171 5185 9180 5219
rect 9128 5176 9180 5185
rect 10508 5219 10560 5228
rect 10508 5185 10517 5219
rect 10517 5185 10551 5219
rect 10551 5185 10560 5219
rect 10508 5176 10560 5185
rect 12624 5176 12676 5228
rect 13544 5312 13596 5364
rect 13176 5219 13228 5228
rect 13176 5185 13185 5219
rect 13185 5185 13219 5219
rect 13219 5185 13228 5219
rect 13176 5176 13228 5185
rect 13636 5176 13688 5228
rect 14004 5176 14056 5228
rect 15568 5176 15620 5228
rect 1768 5108 1820 5160
rect 2596 5108 2648 5160
rect 2872 5108 2924 5160
rect 3516 5108 3568 5160
rect 4160 5108 4212 5160
rect 4712 5108 4764 5160
rect 5908 5108 5960 5160
rect 6828 5151 6880 5160
rect 6828 5117 6837 5151
rect 6837 5117 6871 5151
rect 6871 5117 6880 5151
rect 6828 5108 6880 5117
rect 8852 5108 8904 5160
rect 9220 5108 9272 5160
rect 13268 5108 13320 5160
rect 13544 5151 13596 5160
rect 13544 5117 13553 5151
rect 13553 5117 13587 5151
rect 13587 5117 13596 5151
rect 13544 5108 13596 5117
rect 14188 5108 14240 5160
rect 14464 5108 14516 5160
rect 15108 5108 15160 5160
rect 16856 5108 16908 5160
rect 19800 5151 19852 5160
rect 19800 5117 19809 5151
rect 19809 5117 19843 5151
rect 19843 5117 19852 5151
rect 19800 5108 19852 5117
rect 5816 5040 5868 5092
rect 3424 5015 3476 5024
rect 3424 4981 3433 5015
rect 3433 4981 3467 5015
rect 3467 4981 3476 5015
rect 3424 4972 3476 4981
rect 4896 4972 4948 5024
rect 5540 4972 5592 5024
rect 6920 4972 6972 5024
rect 11152 5040 11204 5092
rect 15476 5040 15528 5092
rect 17868 5040 17920 5092
rect 10140 4972 10192 5024
rect 11060 4972 11112 5024
rect 11796 5015 11848 5024
rect 11796 4981 11805 5015
rect 11805 4981 11839 5015
rect 11839 4981 11848 5015
rect 11796 4972 11848 4981
rect 14004 4972 14056 5024
rect 14188 5015 14240 5024
rect 14188 4981 14197 5015
rect 14197 4981 14231 5015
rect 14231 4981 14240 5015
rect 14188 4972 14240 4981
rect 15108 4972 15160 5024
rect 20628 4972 20680 5024
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 2228 4675 2280 4684
rect 2228 4641 2237 4675
rect 2237 4641 2271 4675
rect 2271 4641 2280 4675
rect 2228 4632 2280 4641
rect 2320 4675 2372 4684
rect 2320 4641 2329 4675
rect 2329 4641 2363 4675
rect 2363 4641 2372 4675
rect 3240 4675 3292 4684
rect 2320 4632 2372 4641
rect 3240 4641 3249 4675
rect 3249 4641 3283 4675
rect 3283 4641 3292 4675
rect 3240 4632 3292 4641
rect 2412 4607 2464 4616
rect 2412 4573 2421 4607
rect 2421 4573 2455 4607
rect 2455 4573 2464 4607
rect 2412 4564 2464 4573
rect 3332 4607 3384 4616
rect 3332 4573 3341 4607
rect 3341 4573 3375 4607
rect 3375 4573 3384 4607
rect 3332 4564 3384 4573
rect 3976 4632 4028 4684
rect 4620 4768 4672 4820
rect 5908 4768 5960 4820
rect 6092 4768 6144 4820
rect 11152 4768 11204 4820
rect 4712 4700 4764 4752
rect 5448 4700 5500 4752
rect 7932 4700 7984 4752
rect 8760 4743 8812 4752
rect 8760 4709 8769 4743
rect 8769 4709 8803 4743
rect 8803 4709 8812 4743
rect 8760 4700 8812 4709
rect 8852 4700 8904 4752
rect 11520 4743 11572 4752
rect 5540 4632 5592 4684
rect 5908 4496 5960 4548
rect 6920 4564 6972 4616
rect 7840 4607 7892 4616
rect 7840 4573 7849 4607
rect 7849 4573 7883 4607
rect 7883 4573 7892 4607
rect 7840 4564 7892 4573
rect 8116 4564 8168 4616
rect 9312 4632 9364 4684
rect 11520 4709 11554 4743
rect 11554 4709 11572 4743
rect 11520 4700 11572 4709
rect 11796 4768 11848 4820
rect 14188 4768 14240 4820
rect 15292 4768 15344 4820
rect 16948 4768 17000 4820
rect 15108 4700 15160 4752
rect 6736 4496 6788 4548
rect 7288 4496 7340 4548
rect 9128 4564 9180 4616
rect 10232 4607 10284 4616
rect 10232 4573 10241 4607
rect 10241 4573 10275 4607
rect 10275 4573 10284 4607
rect 10232 4564 10284 4573
rect 10784 4564 10836 4616
rect 11244 4607 11296 4616
rect 11244 4573 11253 4607
rect 11253 4573 11287 4607
rect 11287 4573 11296 4607
rect 11244 4564 11296 4573
rect 12624 4539 12676 4548
rect 12624 4505 12633 4539
rect 12633 4505 12667 4539
rect 12667 4505 12676 4539
rect 12624 4496 12676 4505
rect 13268 4675 13320 4684
rect 13268 4641 13277 4675
rect 13277 4641 13311 4675
rect 13311 4641 13320 4675
rect 17868 4675 17920 4684
rect 13268 4632 13320 4641
rect 13360 4607 13412 4616
rect 13360 4573 13369 4607
rect 13369 4573 13403 4607
rect 13403 4573 13412 4607
rect 13360 4564 13412 4573
rect 13636 4564 13688 4616
rect 15016 4564 15068 4616
rect 17868 4641 17877 4675
rect 17877 4641 17911 4675
rect 17911 4641 17920 4675
rect 17868 4632 17920 4641
rect 19340 4564 19392 4616
rect 5080 4428 5132 4480
rect 5540 4428 5592 4480
rect 8392 4471 8444 4480
rect 8392 4437 8401 4471
rect 8401 4437 8435 4471
rect 8435 4437 8444 4471
rect 8392 4428 8444 4437
rect 11152 4428 11204 4480
rect 15108 4428 15160 4480
rect 18788 4428 18840 4480
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 2412 4224 2464 4276
rect 5724 4224 5776 4276
rect 7840 4224 7892 4276
rect 7932 4224 7984 4276
rect 9312 4267 9364 4276
rect 9312 4233 9321 4267
rect 9321 4233 9355 4267
rect 9355 4233 9364 4267
rect 9312 4224 9364 4233
rect 9956 4224 10008 4276
rect 10968 4224 11020 4276
rect 13176 4224 13228 4276
rect 4804 4199 4856 4208
rect 4804 4165 4813 4199
rect 4813 4165 4847 4199
rect 4847 4165 4856 4199
rect 4804 4156 4856 4165
rect 1768 4063 1820 4072
rect 1768 4029 1777 4063
rect 1777 4029 1811 4063
rect 1811 4029 1820 4063
rect 1768 4020 1820 4029
rect 3976 4020 4028 4072
rect 2136 3952 2188 4004
rect 3608 3952 3660 4004
rect 3792 3952 3844 4004
rect 5724 4088 5776 4140
rect 6920 4156 6972 4208
rect 8208 4156 8260 4208
rect 6368 4088 6420 4140
rect 7656 4131 7708 4140
rect 7656 4097 7665 4131
rect 7665 4097 7699 4131
rect 7699 4097 7708 4131
rect 7656 4088 7708 4097
rect 8668 4131 8720 4140
rect 8668 4097 8677 4131
rect 8677 4097 8711 4131
rect 8711 4097 8720 4131
rect 8668 4088 8720 4097
rect 9772 4131 9824 4140
rect 9772 4097 9781 4131
rect 9781 4097 9815 4131
rect 9815 4097 9824 4131
rect 9772 4088 9824 4097
rect 9864 4088 9916 4140
rect 10508 4088 10560 4140
rect 11612 4156 11664 4208
rect 13728 4156 13780 4208
rect 13912 4088 13964 4140
rect 2964 3884 3016 3936
rect 6000 4020 6052 4072
rect 6644 4020 6696 4072
rect 12072 4020 12124 4072
rect 12348 4020 12400 4072
rect 13176 4020 13228 4072
rect 19340 4088 19392 4140
rect 22468 4088 22520 4140
rect 4988 3952 5040 4004
rect 10140 3952 10192 4004
rect 5172 3927 5224 3936
rect 5172 3893 5181 3927
rect 5181 3893 5215 3927
rect 5215 3893 5224 3927
rect 5172 3884 5224 3893
rect 5264 3884 5316 3936
rect 6092 3884 6144 3936
rect 8484 3927 8536 3936
rect 8484 3893 8493 3927
rect 8493 3893 8527 3927
rect 8527 3893 8536 3927
rect 8484 3884 8536 3893
rect 8576 3927 8628 3936
rect 8576 3893 8585 3927
rect 8585 3893 8619 3927
rect 8619 3893 8628 3927
rect 9680 3927 9732 3936
rect 8576 3884 8628 3893
rect 9680 3893 9689 3927
rect 9689 3893 9723 3927
rect 9723 3893 9732 3927
rect 9680 3884 9732 3893
rect 12532 3952 12584 4004
rect 12900 3952 12952 4004
rect 11060 3884 11112 3936
rect 11244 3927 11296 3936
rect 11244 3893 11253 3927
rect 11253 3893 11287 3927
rect 11287 3893 11296 3927
rect 11244 3884 11296 3893
rect 11336 3927 11388 3936
rect 11336 3893 11345 3927
rect 11345 3893 11379 3927
rect 11379 3893 11388 3927
rect 14648 3952 14700 4004
rect 11336 3884 11388 3893
rect 13636 3884 13688 3936
rect 14096 3927 14148 3936
rect 14096 3893 14105 3927
rect 14105 3893 14139 3927
rect 14139 3893 14148 3927
rect 14096 3884 14148 3893
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 2504 3680 2556 3732
rect 4620 3680 4672 3732
rect 5172 3680 5224 3732
rect 6736 3680 6788 3732
rect 8944 3680 8996 3732
rect 9680 3680 9732 3732
rect 2412 3612 2464 3664
rect 2596 3612 2648 3664
rect 3148 3612 3200 3664
rect 4804 3612 4856 3664
rect 4896 3612 4948 3664
rect 8576 3612 8628 3664
rect 10232 3612 10284 3664
rect 1584 3544 1636 3596
rect 7012 3544 7064 3596
rect 7656 3544 7708 3596
rect 7932 3544 7984 3596
rect 8484 3544 8536 3596
rect 11520 3680 11572 3732
rect 12348 3680 12400 3732
rect 12900 3723 12952 3732
rect 12900 3689 12909 3723
rect 12909 3689 12943 3723
rect 12943 3689 12952 3723
rect 12900 3680 12952 3689
rect 11612 3612 11664 3664
rect 11980 3612 12032 3664
rect 13360 3680 13412 3732
rect 13636 3680 13688 3732
rect 1768 3519 1820 3528
rect 1768 3485 1777 3519
rect 1777 3485 1811 3519
rect 1811 3485 1820 3519
rect 1768 3476 1820 3485
rect 3976 3476 4028 3528
rect 5724 3476 5776 3528
rect 6368 3519 6420 3528
rect 6368 3485 6377 3519
rect 6377 3485 6411 3519
rect 6411 3485 6420 3519
rect 6368 3476 6420 3485
rect 6828 3476 6880 3528
rect 8208 3476 8260 3528
rect 9772 3476 9824 3528
rect 5540 3451 5592 3460
rect 2044 3340 2096 3392
rect 5540 3417 5549 3451
rect 5549 3417 5583 3451
rect 5583 3417 5592 3451
rect 5540 3408 5592 3417
rect 5816 3451 5868 3460
rect 5816 3417 5825 3451
rect 5825 3417 5859 3451
rect 5859 3417 5868 3451
rect 5816 3408 5868 3417
rect 11244 3544 11296 3596
rect 12808 3544 12860 3596
rect 13728 3612 13780 3664
rect 11520 3519 11572 3528
rect 11520 3485 11529 3519
rect 11529 3485 11563 3519
rect 11563 3485 11572 3519
rect 11520 3476 11572 3485
rect 12532 3476 12584 3528
rect 13176 3476 13228 3528
rect 13360 3476 13412 3528
rect 14372 3544 14424 3596
rect 16028 3587 16080 3596
rect 16028 3553 16037 3587
rect 16037 3553 16071 3587
rect 16071 3553 16080 3587
rect 16028 3544 16080 3553
rect 16120 3476 16172 3528
rect 3608 3340 3660 3392
rect 5264 3340 5316 3392
rect 5724 3340 5776 3392
rect 6552 3340 6604 3392
rect 7472 3340 7524 3392
rect 11336 3408 11388 3460
rect 8116 3340 8168 3392
rect 10508 3340 10560 3392
rect 13912 3340 13964 3392
rect 15016 3340 15068 3392
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 2228 3136 2280 3188
rect 2596 3136 2648 3188
rect 3240 3136 3292 3188
rect 3332 3136 3384 3188
rect 4160 3136 4212 3188
rect 5356 3136 5408 3188
rect 8392 3136 8444 3188
rect 8944 3136 8996 3188
rect 2136 3000 2188 3052
rect 3424 3000 3476 3052
rect 4344 3043 4396 3052
rect 4344 3009 4353 3043
rect 4353 3009 4387 3043
rect 4387 3009 4396 3043
rect 6184 3068 6236 3120
rect 7564 3068 7616 3120
rect 5264 3043 5316 3052
rect 4344 3000 4396 3009
rect 2044 2975 2096 2984
rect 2044 2941 2053 2975
rect 2053 2941 2087 2975
rect 2087 2941 2096 2975
rect 2044 2932 2096 2941
rect 5264 3009 5273 3043
rect 5273 3009 5307 3043
rect 5307 3009 5316 3043
rect 5264 3000 5316 3009
rect 5724 3000 5776 3052
rect 6276 3000 6328 3052
rect 5080 2932 5132 2984
rect 7472 2975 7524 2984
rect 7472 2941 7481 2975
rect 7481 2941 7515 2975
rect 7515 2941 7524 2975
rect 7472 2932 7524 2941
rect 204 2864 256 2916
rect 1952 2864 2004 2916
rect 4252 2864 4304 2916
rect 2872 2796 2924 2848
rect 3056 2839 3108 2848
rect 3056 2805 3065 2839
rect 3065 2805 3099 2839
rect 3099 2805 3108 2839
rect 3056 2796 3108 2805
rect 3148 2796 3200 2848
rect 5908 2864 5960 2916
rect 6828 2864 6880 2916
rect 7932 3000 7984 3052
rect 8199 3043 8251 3052
rect 8199 3009 8217 3043
rect 8217 3009 8251 3043
rect 9312 3136 9364 3188
rect 10232 3136 10284 3188
rect 14280 3136 14332 3188
rect 20168 3136 20220 3188
rect 11796 3068 11848 3120
rect 12716 3068 12768 3120
rect 8199 3000 8251 3009
rect 10140 3000 10192 3052
rect 10324 3000 10376 3052
rect 10508 3000 10560 3052
rect 14096 3068 14148 3120
rect 16028 3068 16080 3120
rect 9956 2932 10008 2984
rect 10600 2932 10652 2984
rect 10692 2932 10744 2984
rect 13728 2975 13780 2984
rect 8116 2864 8168 2916
rect 8576 2864 8628 2916
rect 9496 2864 9548 2916
rect 4712 2796 4764 2848
rect 7196 2796 7248 2848
rect 9220 2796 9272 2848
rect 12808 2907 12860 2916
rect 12808 2873 12817 2907
rect 12817 2873 12851 2907
rect 12851 2873 12860 2907
rect 12808 2864 12860 2873
rect 13084 2864 13136 2916
rect 13728 2941 13737 2975
rect 13737 2941 13771 2975
rect 13771 2941 13780 2975
rect 13728 2932 13780 2941
rect 13820 2932 13872 2984
rect 16120 2975 16172 2984
rect 14464 2864 14516 2916
rect 16120 2941 16129 2975
rect 16129 2941 16163 2975
rect 16163 2941 16172 2975
rect 16120 2932 16172 2941
rect 16856 2932 16908 2984
rect 18512 2932 18564 2984
rect 19156 2975 19208 2984
rect 19156 2941 19165 2975
rect 19165 2941 19199 2975
rect 19199 2941 19208 2975
rect 19156 2932 19208 2941
rect 10232 2839 10284 2848
rect 10232 2805 10241 2839
rect 10241 2805 10275 2839
rect 10275 2805 10284 2839
rect 10232 2796 10284 2805
rect 10508 2796 10560 2848
rect 10600 2796 10652 2848
rect 11060 2796 11112 2848
rect 15292 2796 15344 2848
rect 22008 2864 22060 2916
rect 16948 2796 17000 2848
rect 17868 2796 17920 2848
rect 19248 2796 19300 2848
rect 19708 2796 19760 2848
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 2320 2635 2372 2644
rect 2320 2601 2329 2635
rect 2329 2601 2363 2635
rect 2363 2601 2372 2635
rect 2320 2592 2372 2601
rect 2688 2635 2740 2644
rect 2688 2601 2697 2635
rect 2697 2601 2731 2635
rect 2731 2601 2740 2635
rect 2688 2592 2740 2601
rect 7288 2592 7340 2644
rect 8392 2592 8444 2644
rect 10140 2635 10192 2644
rect 10140 2601 10149 2635
rect 10149 2601 10183 2635
rect 10183 2601 10192 2635
rect 10140 2592 10192 2601
rect 10968 2592 11020 2644
rect 11152 2635 11204 2644
rect 11152 2601 11161 2635
rect 11161 2601 11195 2635
rect 11195 2601 11204 2635
rect 11152 2592 11204 2601
rect 4068 2524 4120 2576
rect 5632 2524 5684 2576
rect 7012 2524 7064 2576
rect 8484 2524 8536 2576
rect 10600 2524 10652 2576
rect 2780 2431 2832 2440
rect 2780 2397 2789 2431
rect 2789 2397 2823 2431
rect 2823 2397 2832 2431
rect 2780 2388 2832 2397
rect 3424 2388 3476 2440
rect 4068 2388 4120 2440
rect 5264 2456 5316 2508
rect 6460 2456 6512 2508
rect 7380 2456 7432 2508
rect 8024 2499 8076 2508
rect 8024 2465 8033 2499
rect 8033 2465 8067 2499
rect 8067 2465 8076 2499
rect 8024 2456 8076 2465
rect 5908 2388 5960 2440
rect 6368 2388 6420 2440
rect 11704 2456 11756 2508
rect 15108 2592 15160 2644
rect 12072 2567 12124 2576
rect 12072 2533 12081 2567
rect 12081 2533 12115 2567
rect 12115 2533 12124 2567
rect 12072 2524 12124 2533
rect 13544 2524 13596 2576
rect 21548 2524 21600 2576
rect 9312 2431 9364 2440
rect 7748 2320 7800 2372
rect 9312 2397 9321 2431
rect 9321 2397 9355 2431
rect 9355 2397 9364 2431
rect 9312 2388 9364 2397
rect 9680 2388 9732 2440
rect 10324 2431 10376 2440
rect 10324 2397 10333 2431
rect 10333 2397 10367 2431
rect 10367 2397 10376 2431
rect 10324 2388 10376 2397
rect 6920 2252 6972 2304
rect 7012 2252 7064 2304
rect 11612 2388 11664 2440
rect 12992 2456 13044 2508
rect 13912 2499 13964 2508
rect 13912 2465 13921 2499
rect 13921 2465 13955 2499
rect 13955 2465 13964 2499
rect 13912 2456 13964 2465
rect 14188 2456 14240 2508
rect 15660 2499 15712 2508
rect 15660 2465 15669 2499
rect 15669 2465 15703 2499
rect 15703 2465 15712 2499
rect 15660 2456 15712 2465
rect 16580 2499 16632 2508
rect 16580 2465 16589 2499
rect 16589 2465 16623 2499
rect 16623 2465 16632 2499
rect 16580 2456 16632 2465
rect 17040 2456 17092 2508
rect 21088 2320 21140 2372
rect 8760 2252 8812 2304
rect 9680 2252 9732 2304
rect 11060 2252 11112 2304
rect 15568 2252 15620 2304
rect 16488 2252 16540 2304
rect 17408 2252 17460 2304
rect 17960 2252 18012 2304
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 6460 2048 6512 2100
rect 13360 2048 13412 2100
rect 15660 2048 15712 2100
rect 2044 1980 2096 2032
rect 8024 1980 8076 2032
rect 9588 1980 9640 2032
rect 664 1912 716 1964
rect 7196 1912 7248 1964
rect 1124 1844 1176 1896
rect 5448 1844 5500 1896
rect 7472 1844 7524 1896
rect 11336 1368 11388 1420
rect 12164 1368 12216 1420
rect 3516 1300 3568 1352
rect 5172 1300 5224 1352
<< metal2 >>
rect 202 22320 258 22800
rect 570 22320 626 22800
rect 1030 22320 1086 22800
rect 1490 22320 1546 22800
rect 1950 22320 2006 22800
rect 2410 22320 2466 22800
rect 2778 22536 2834 22545
rect 2778 22471 2834 22480
rect 216 18766 244 22320
rect 204 18760 256 18766
rect 204 18702 256 18708
rect 584 18086 612 22320
rect 1044 18426 1072 22320
rect 1504 18970 1532 22320
rect 1860 19712 1912 19718
rect 1858 19680 1860 19689
rect 1912 19680 1914 19689
rect 1858 19615 1914 19624
rect 1766 19272 1822 19281
rect 1766 19207 1822 19216
rect 1780 19174 1808 19207
rect 1768 19168 1820 19174
rect 1768 19110 1820 19116
rect 1492 18964 1544 18970
rect 1492 18906 1544 18912
rect 1400 18828 1452 18834
rect 1400 18770 1452 18776
rect 1032 18420 1084 18426
rect 1032 18362 1084 18368
rect 572 18080 624 18086
rect 572 18022 624 18028
rect 1412 17678 1440 18770
rect 1582 18728 1638 18737
rect 1582 18663 1584 18672
rect 1636 18663 1638 18672
rect 1584 18634 1636 18640
rect 1676 18352 1728 18358
rect 1674 18320 1676 18329
rect 1728 18320 1730 18329
rect 1674 18255 1730 18264
rect 1400 17672 1452 17678
rect 1400 17614 1452 17620
rect 1766 17368 1822 17377
rect 1766 17303 1768 17312
rect 1820 17303 1822 17312
rect 1768 17274 1820 17280
rect 1584 17128 1636 17134
rect 1964 17105 1992 22320
rect 2136 19304 2188 19310
rect 2136 19246 2188 19252
rect 2148 18193 2176 19246
rect 2228 19236 2280 19242
rect 2228 19178 2280 19184
rect 2240 18222 2268 19178
rect 2228 18216 2280 18222
rect 2134 18184 2190 18193
rect 2228 18158 2280 18164
rect 2134 18119 2190 18128
rect 1584 17070 1636 17076
rect 1950 17096 2006 17105
rect 1596 16726 1624 17070
rect 1950 17031 2006 17040
rect 2320 17060 2372 17066
rect 2320 17002 2372 17008
rect 1676 16992 1728 16998
rect 1676 16934 1728 16940
rect 1584 16720 1636 16726
rect 1584 16662 1636 16668
rect 1688 16658 1716 16934
rect 1858 16824 1914 16833
rect 1858 16759 1860 16768
rect 1912 16759 1914 16768
rect 1860 16730 1912 16736
rect 1676 16652 1728 16658
rect 1676 16594 1728 16600
rect 1950 16416 2006 16425
rect 1950 16351 2006 16360
rect 1964 16250 1992 16351
rect 1952 16244 2004 16250
rect 1952 16186 2004 16192
rect 2332 16046 2360 17002
rect 1768 16040 1820 16046
rect 1766 16008 1768 16017
rect 2320 16040 2372 16046
rect 1820 16008 1822 16017
rect 2320 15982 2372 15988
rect 1766 15943 1822 15952
rect 1582 15872 1638 15881
rect 1582 15807 1638 15816
rect 1596 15706 1624 15807
rect 1584 15700 1636 15706
rect 2424 15688 2452 22320
rect 2596 19236 2648 19242
rect 2596 19178 2648 19184
rect 2504 18964 2556 18970
rect 2504 18906 2556 18912
rect 2516 15910 2544 18906
rect 2608 18601 2636 19178
rect 2792 18816 2820 22471
rect 2870 22320 2926 22800
rect 3330 22320 3386 22800
rect 3790 22320 3846 22800
rect 4250 22320 4306 22800
rect 4710 22320 4766 22800
rect 5170 22320 5226 22800
rect 5630 22320 5686 22800
rect 6090 22320 6146 22800
rect 6550 22320 6606 22800
rect 7010 22320 7066 22800
rect 7470 22320 7526 22800
rect 7930 22320 7986 22800
rect 8390 22320 8446 22800
rect 8850 22320 8906 22800
rect 9310 22320 9366 22800
rect 9770 22320 9826 22800
rect 10230 22320 10286 22800
rect 10690 22320 10746 22800
rect 11150 22320 11206 22800
rect 11610 22320 11666 22800
rect 11978 22320 12034 22800
rect 12438 22320 12494 22800
rect 12898 22320 12954 22800
rect 13358 22320 13414 22800
rect 13818 22320 13874 22800
rect 14278 22320 14334 22800
rect 14738 22320 14794 22800
rect 15198 22320 15254 22800
rect 15658 22320 15714 22800
rect 16118 22320 16174 22800
rect 16578 22320 16634 22800
rect 17038 22320 17094 22800
rect 17498 22320 17554 22800
rect 17958 22320 18014 22800
rect 18418 22320 18474 22800
rect 18878 22320 18934 22800
rect 19338 22320 19394 22800
rect 19798 22320 19854 22800
rect 20258 22320 20314 22800
rect 20718 22320 20774 22800
rect 21178 22320 21234 22800
rect 21638 22320 21694 22800
rect 22098 22320 22154 22800
rect 22558 22320 22614 22800
rect 2884 20074 2912 22320
rect 3146 21584 3202 21593
rect 3146 21519 3202 21528
rect 2884 20046 3004 20074
rect 2872 19916 2924 19922
rect 2872 19858 2924 19864
rect 2884 18970 2912 19858
rect 2872 18964 2924 18970
rect 2872 18906 2924 18912
rect 2792 18788 2912 18816
rect 2780 18692 2832 18698
rect 2780 18634 2832 18640
rect 2594 18592 2650 18601
rect 2594 18527 2650 18536
rect 2792 18426 2820 18634
rect 2596 18420 2648 18426
rect 2596 18362 2648 18368
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 2608 15978 2636 18362
rect 2688 18080 2740 18086
rect 2688 18022 2740 18028
rect 2700 16590 2728 18022
rect 2778 17776 2834 17785
rect 2778 17711 2834 17720
rect 2688 16584 2740 16590
rect 2688 16526 2740 16532
rect 2792 16250 2820 17711
rect 2780 16244 2832 16250
rect 2780 16186 2832 16192
rect 2596 15972 2648 15978
rect 2596 15914 2648 15920
rect 2504 15904 2556 15910
rect 2884 15881 2912 18788
rect 2976 16794 3004 20046
rect 3056 19916 3108 19922
rect 3056 19858 3108 19864
rect 3068 18698 3096 19858
rect 3056 18692 3108 18698
rect 3056 18634 3108 18640
rect 3056 18420 3108 18426
rect 3056 18362 3108 18368
rect 2964 16788 3016 16794
rect 2964 16730 3016 16736
rect 2964 16448 3016 16454
rect 2964 16390 3016 16396
rect 2504 15846 2556 15852
rect 2870 15872 2926 15881
rect 2870 15807 2926 15816
rect 2976 15706 3004 16390
rect 3068 16250 3096 18362
rect 3160 18329 3188 21519
rect 3240 19848 3292 19854
rect 3240 19790 3292 19796
rect 3252 19514 3280 19790
rect 3240 19508 3292 19514
rect 3240 19450 3292 19456
rect 3344 19394 3372 22320
rect 3698 22128 3754 22137
rect 3698 22063 3754 22072
rect 3606 21176 3662 21185
rect 3606 21111 3662 21120
rect 3620 20074 3648 21111
rect 3712 20874 3740 22063
rect 3700 20868 3752 20874
rect 3700 20810 3752 20816
rect 3698 20632 3754 20641
rect 3698 20567 3754 20576
rect 3712 20262 3740 20567
rect 3700 20256 3752 20262
rect 3700 20198 3752 20204
rect 3620 20046 3740 20074
rect 3516 19780 3568 19786
rect 3516 19722 3568 19728
rect 3344 19366 3464 19394
rect 3240 19168 3292 19174
rect 3240 19110 3292 19116
rect 3332 19168 3384 19174
rect 3332 19110 3384 19116
rect 3146 18320 3202 18329
rect 3146 18255 3202 18264
rect 3252 17746 3280 19110
rect 3344 18970 3372 19110
rect 3332 18964 3384 18970
rect 3332 18906 3384 18912
rect 3332 18828 3384 18834
rect 3332 18770 3384 18776
rect 3240 17740 3292 17746
rect 3240 17682 3292 17688
rect 3146 17640 3202 17649
rect 3146 17575 3202 17584
rect 3160 16726 3188 17575
rect 3252 17202 3280 17682
rect 3240 17196 3292 17202
rect 3240 17138 3292 17144
rect 3148 16720 3200 16726
rect 3148 16662 3200 16668
rect 3056 16244 3108 16250
rect 3056 16186 3108 16192
rect 2964 15700 3016 15706
rect 2424 15660 2544 15688
rect 1584 15642 1636 15648
rect 2410 15600 2466 15609
rect 1676 15564 1728 15570
rect 2410 15535 2412 15544
rect 1676 15506 1728 15512
rect 2464 15535 2466 15544
rect 2412 15506 2464 15512
rect 1688 15026 1716 15506
rect 1676 15020 1728 15026
rect 1676 14962 1728 14968
rect 1674 14920 1730 14929
rect 1674 14855 1730 14864
rect 1768 14884 1820 14890
rect 1688 14618 1716 14855
rect 1768 14826 1820 14832
rect 1676 14612 1728 14618
rect 1676 14554 1728 14560
rect 1492 14476 1544 14482
rect 1492 14418 1544 14424
rect 1400 13864 1452 13870
rect 1400 13806 1452 13812
rect 1412 10713 1440 13806
rect 1504 13462 1532 14418
rect 1780 14074 1808 14826
rect 2228 14816 2280 14822
rect 2228 14758 2280 14764
rect 2240 14618 2268 14758
rect 2516 14657 2544 15660
rect 2964 15642 3016 15648
rect 2596 15496 2648 15502
rect 2596 15438 2648 15444
rect 2608 15337 2636 15438
rect 2594 15328 2650 15337
rect 2594 15263 2650 15272
rect 2688 14816 2740 14822
rect 2688 14758 2740 14764
rect 3056 14816 3108 14822
rect 3056 14758 3108 14764
rect 2502 14648 2558 14657
rect 2228 14612 2280 14618
rect 2502 14583 2558 14592
rect 2228 14554 2280 14560
rect 2596 14544 2648 14550
rect 2596 14486 2648 14492
rect 2136 14476 2188 14482
rect 2136 14418 2188 14424
rect 2320 14476 2372 14482
rect 2372 14436 2452 14464
rect 2320 14418 2372 14424
rect 1768 14068 1820 14074
rect 1768 14010 1820 14016
rect 2148 13938 2176 14418
rect 2424 14362 2452 14436
rect 2608 14362 2636 14486
rect 2424 14334 2636 14362
rect 2136 13932 2188 13938
rect 2136 13874 2188 13880
rect 1492 13456 1544 13462
rect 1492 13398 1544 13404
rect 2148 13326 2176 13874
rect 2700 13530 2728 14758
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2792 14074 2820 14418
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 2962 13968 3018 13977
rect 2962 13903 3018 13912
rect 2688 13524 2740 13530
rect 2688 13466 2740 13472
rect 2504 13388 2556 13394
rect 2504 13330 2556 13336
rect 2872 13388 2924 13394
rect 2872 13330 2924 13336
rect 2136 13320 2188 13326
rect 2136 13262 2188 13268
rect 2412 12844 2464 12850
rect 2412 12786 2464 12792
rect 1584 12640 1636 12646
rect 1584 12582 1636 12588
rect 2136 12640 2188 12646
rect 2136 12582 2188 12588
rect 1596 11694 1624 12582
rect 2148 12442 2176 12582
rect 2136 12436 2188 12442
rect 2136 12378 2188 12384
rect 1676 12164 1728 12170
rect 1676 12106 1728 12112
rect 1584 11688 1636 11694
rect 1584 11630 1636 11636
rect 1688 11286 1716 12106
rect 2228 11688 2280 11694
rect 2228 11630 2280 11636
rect 1676 11280 1728 11286
rect 1676 11222 1728 11228
rect 2240 11218 2268 11630
rect 2424 11354 2452 12786
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2228 11212 2280 11218
rect 2228 11154 2280 11160
rect 1398 10704 1454 10713
rect 1398 10639 1454 10648
rect 1412 7342 1440 10639
rect 2136 10600 2188 10606
rect 2240 10554 2268 11154
rect 2188 10548 2268 10554
rect 2136 10542 2268 10548
rect 2148 10526 2268 10542
rect 2424 10538 2452 11290
rect 2240 10062 2268 10526
rect 2412 10532 2464 10538
rect 2412 10474 2464 10480
rect 2228 10056 2280 10062
rect 2228 9998 2280 10004
rect 2240 9178 2268 9998
rect 2320 9376 2372 9382
rect 2320 9318 2372 9324
rect 2412 9376 2464 9382
rect 2412 9318 2464 9324
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 1492 9036 1544 9042
rect 1492 8978 1544 8984
rect 1504 8430 1532 8978
rect 1492 8424 1544 8430
rect 1492 8366 1544 8372
rect 2332 8090 2360 9318
rect 2424 8634 2452 9318
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2320 8084 2372 8090
rect 2320 8026 2372 8032
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 1400 7336 1452 7342
rect 1400 7278 1452 7284
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1780 6186 1808 6802
rect 1872 6254 1900 7346
rect 2516 7313 2544 13330
rect 2780 12640 2832 12646
rect 2780 12582 2832 12588
rect 2792 12306 2820 12582
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2884 10282 2912 13330
rect 2976 12714 3004 13903
rect 2964 12708 3016 12714
rect 2964 12650 3016 12656
rect 3068 12442 3096 14758
rect 3160 12986 3188 16662
rect 3240 16584 3292 16590
rect 3240 16526 3292 16532
rect 3252 15570 3280 16526
rect 3344 16454 3372 18770
rect 3436 17785 3464 19366
rect 3528 19174 3556 19722
rect 3516 19168 3568 19174
rect 3516 19110 3568 19116
rect 3608 19168 3660 19174
rect 3608 19110 3660 19116
rect 3620 18766 3648 19110
rect 3608 18760 3660 18766
rect 3608 18702 3660 18708
rect 3514 18592 3570 18601
rect 3514 18527 3570 18536
rect 3422 17776 3478 17785
rect 3422 17711 3478 17720
rect 3424 17672 3476 17678
rect 3424 17614 3476 17620
rect 3436 17338 3464 17614
rect 3424 17332 3476 17338
rect 3424 17274 3476 17280
rect 3424 16788 3476 16794
rect 3424 16730 3476 16736
rect 3436 16697 3464 16730
rect 3528 16726 3556 18527
rect 3620 17066 3648 18702
rect 3608 17060 3660 17066
rect 3608 17002 3660 17008
rect 3516 16720 3568 16726
rect 3422 16688 3478 16697
rect 3516 16662 3568 16668
rect 3422 16623 3478 16632
rect 3712 16522 3740 20046
rect 3804 17066 3832 22320
rect 4068 20324 4120 20330
rect 4068 20266 4120 20272
rect 4080 20233 4108 20266
rect 4066 20224 4122 20233
rect 4066 20159 4122 20168
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 3976 19372 4028 19378
rect 3976 19314 4028 19320
rect 3988 18902 4016 19314
rect 4080 18970 4108 19654
rect 4264 19394 4292 22320
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 4264 19366 4384 19394
rect 4252 19236 4304 19242
rect 4252 19178 4304 19184
rect 4068 18964 4120 18970
rect 4068 18906 4120 18912
rect 3976 18896 4028 18902
rect 3976 18838 4028 18844
rect 4160 18624 4212 18630
rect 4160 18566 4212 18572
rect 4172 18222 4200 18566
rect 4068 18216 4120 18222
rect 4068 18158 4120 18164
rect 4160 18216 4212 18222
rect 4160 18158 4212 18164
rect 4080 17785 4108 18158
rect 4264 17882 4292 19178
rect 4356 18970 4384 19366
rect 4436 19168 4488 19174
rect 4436 19110 4488 19116
rect 4526 19136 4582 19145
rect 4344 18964 4396 18970
rect 4344 18906 4396 18912
rect 4448 18850 4476 19110
rect 4526 19071 4582 19080
rect 4540 18902 4568 19071
rect 4356 18834 4476 18850
rect 4528 18896 4580 18902
rect 4528 18838 4580 18844
rect 4344 18828 4476 18834
rect 4396 18822 4476 18828
rect 4344 18770 4396 18776
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4252 17876 4304 17882
rect 4724 17864 4752 22320
rect 5184 20058 5212 22320
rect 5172 20052 5224 20058
rect 5172 19994 5224 20000
rect 5540 20052 5592 20058
rect 5540 19994 5592 20000
rect 5264 19916 5316 19922
rect 5264 19858 5316 19864
rect 4896 19848 4948 19854
rect 4896 19790 4948 19796
rect 5080 19848 5132 19854
rect 5080 19790 5132 19796
rect 5276 19802 5304 19858
rect 4908 19310 4936 19790
rect 4988 19780 5040 19786
rect 4988 19722 5040 19728
rect 4896 19304 4948 19310
rect 4896 19246 4948 19252
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 4816 18154 4844 18702
rect 4908 18358 4936 19246
rect 4896 18352 4948 18358
rect 4896 18294 4948 18300
rect 4894 18184 4950 18193
rect 4804 18148 4856 18154
rect 4894 18119 4896 18128
rect 4804 18090 4856 18096
rect 4948 18119 4950 18128
rect 4896 18090 4948 18096
rect 4724 17836 4936 17864
rect 4252 17818 4304 17824
rect 4066 17776 4122 17785
rect 4066 17711 4068 17720
rect 4120 17711 4122 17720
rect 4712 17740 4764 17746
rect 4068 17682 4120 17688
rect 4712 17682 4764 17688
rect 3976 17536 4028 17542
rect 3976 17478 4028 17484
rect 3792 17060 3844 17066
rect 3792 17002 3844 17008
rect 3988 16794 4016 17478
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 4724 17270 4752 17682
rect 4712 17264 4764 17270
rect 4712 17206 4764 17212
rect 4804 17060 4856 17066
rect 4804 17002 4856 17008
rect 3976 16788 4028 16794
rect 3976 16730 4028 16736
rect 4252 16652 4304 16658
rect 4252 16594 4304 16600
rect 3792 16584 3844 16590
rect 3792 16526 3844 16532
rect 3424 16516 3476 16522
rect 3424 16458 3476 16464
rect 3700 16516 3752 16522
rect 3700 16458 3752 16464
rect 3332 16448 3384 16454
rect 3332 16390 3384 16396
rect 3240 15564 3292 15570
rect 3240 15506 3292 15512
rect 3240 14952 3292 14958
rect 3240 14894 3292 14900
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 3148 12640 3200 12646
rect 3148 12582 3200 12588
rect 3056 12436 3108 12442
rect 2792 10254 2912 10282
rect 2976 12396 3056 12424
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 2608 8566 2636 9522
rect 2700 9110 2728 9522
rect 2688 9104 2740 9110
rect 2688 9046 2740 9052
rect 2596 8560 2648 8566
rect 2596 8502 2648 8508
rect 2502 7304 2558 7313
rect 2502 7239 2504 7248
rect 2556 7239 2558 7248
rect 2504 7210 2556 7216
rect 1952 7200 2004 7206
rect 2516 7179 2544 7210
rect 1952 7142 2004 7148
rect 1860 6248 1912 6254
rect 1860 6190 1912 6196
rect 1768 6180 1820 6186
rect 1768 6122 1820 6128
rect 1780 5166 1808 6122
rect 1964 5914 1992 7142
rect 2228 6860 2280 6866
rect 2228 6802 2280 6808
rect 2240 6118 2268 6802
rect 2228 6112 2280 6118
rect 2228 6054 2280 6060
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 2240 5710 2268 6054
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 2608 5166 2636 8502
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 2700 7886 2728 8366
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2688 6792 2740 6798
rect 2688 6734 2740 6740
rect 2700 5778 2728 6734
rect 2792 5846 2820 10254
rect 2872 10124 2924 10130
rect 2872 10066 2924 10072
rect 2884 7410 2912 10066
rect 2976 9489 3004 12396
rect 3056 12378 3108 12384
rect 3056 11212 3108 11218
rect 3056 11154 3108 11160
rect 2962 9480 3018 9489
rect 3068 9450 3096 11154
rect 3160 10674 3188 12582
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3252 10198 3280 14894
rect 3344 14822 3372 16390
rect 3436 15638 3464 16458
rect 3516 16244 3568 16250
rect 3516 16186 3568 16192
rect 3700 16244 3752 16250
rect 3700 16186 3752 16192
rect 3528 15978 3556 16186
rect 3516 15972 3568 15978
rect 3516 15914 3568 15920
rect 3424 15632 3476 15638
rect 3424 15574 3476 15580
rect 3528 15502 3556 15914
rect 3608 15904 3660 15910
rect 3608 15846 3660 15852
rect 3516 15496 3568 15502
rect 3422 15464 3478 15473
rect 3516 15438 3568 15444
rect 3422 15399 3478 15408
rect 3436 15162 3464 15399
rect 3424 15156 3476 15162
rect 3424 15098 3476 15104
rect 3516 15020 3568 15026
rect 3516 14962 3568 14968
rect 3332 14816 3384 14822
rect 3332 14758 3384 14764
rect 3330 14512 3386 14521
rect 3330 14447 3386 14456
rect 3344 13530 3372 14447
rect 3528 14278 3556 14962
rect 3516 14272 3568 14278
rect 3516 14214 3568 14220
rect 3528 13938 3556 14214
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 3424 13796 3476 13802
rect 3424 13738 3476 13744
rect 3332 13524 3384 13530
rect 3332 13466 3384 13472
rect 3436 13190 3464 13738
rect 3516 13728 3568 13734
rect 3516 13670 3568 13676
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 3332 12776 3384 12782
rect 3332 12718 3384 12724
rect 3240 10192 3292 10198
rect 3240 10134 3292 10140
rect 3344 9466 3372 12718
rect 3436 12238 3464 12786
rect 3528 12782 3556 13670
rect 3620 13530 3648 15846
rect 3712 15366 3740 16186
rect 3804 16114 3832 16526
rect 4264 16402 4292 16594
rect 3896 16374 4292 16402
rect 3792 16108 3844 16114
rect 3792 16050 3844 16056
rect 3804 15745 3832 16050
rect 3790 15736 3846 15745
rect 3790 15671 3846 15680
rect 3792 15564 3844 15570
rect 3792 15506 3844 15512
rect 3700 15360 3752 15366
rect 3700 15302 3752 15308
rect 3700 14952 3752 14958
rect 3700 14894 3752 14900
rect 3712 14074 3740 14894
rect 3804 14346 3832 15506
rect 3896 14958 3924 16374
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4068 16108 4120 16114
rect 4068 16050 4120 16056
rect 4528 16108 4580 16114
rect 4528 16050 4580 16056
rect 4080 15978 4108 16050
rect 4068 15972 4120 15978
rect 4068 15914 4120 15920
rect 4252 15904 4304 15910
rect 4252 15846 4304 15852
rect 4436 15904 4488 15910
rect 4436 15846 4488 15852
rect 4066 15736 4122 15745
rect 4066 15671 4122 15680
rect 3976 15496 4028 15502
rect 4080 15484 4108 15671
rect 4028 15456 4108 15484
rect 3976 15438 4028 15444
rect 3884 14952 3936 14958
rect 3988 14929 4016 15438
rect 3884 14894 3936 14900
rect 3974 14920 4030 14929
rect 3974 14855 4030 14864
rect 3792 14340 3844 14346
rect 3792 14282 3844 14288
rect 3700 14068 3752 14074
rect 3700 14010 3752 14016
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 3608 13524 3660 13530
rect 3608 13466 3660 13472
rect 3712 13326 3740 14010
rect 4066 13560 4122 13569
rect 4066 13495 4122 13504
rect 3884 13388 3936 13394
rect 3884 13330 3936 13336
rect 3700 13320 3752 13326
rect 3700 13262 3752 13268
rect 3712 12850 3740 13262
rect 3700 12844 3752 12850
rect 3700 12786 3752 12792
rect 3516 12776 3568 12782
rect 3516 12718 3568 12724
rect 3792 12776 3844 12782
rect 3792 12718 3844 12724
rect 3516 12300 3568 12306
rect 3516 12242 3568 12248
rect 3424 12232 3476 12238
rect 3528 12209 3556 12242
rect 3424 12174 3476 12180
rect 3514 12200 3570 12209
rect 3436 11830 3464 12174
rect 3514 12135 3570 12144
rect 3700 12164 3752 12170
rect 3424 11824 3476 11830
rect 3424 11766 3476 11772
rect 3436 10266 3464 11766
rect 3528 11098 3556 12135
rect 3700 12106 3752 12112
rect 3606 12064 3662 12073
rect 3606 11999 3662 12008
rect 3620 11218 3648 11999
rect 3712 11830 3740 12106
rect 3700 11824 3752 11830
rect 3700 11766 3752 11772
rect 3700 11688 3752 11694
rect 3700 11630 3752 11636
rect 3608 11212 3660 11218
rect 3608 11154 3660 11160
rect 3528 11070 3648 11098
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3424 10124 3476 10130
rect 3424 10066 3476 10072
rect 2962 9415 3018 9424
rect 3056 9444 3108 9450
rect 3056 9386 3108 9392
rect 3160 9438 3372 9466
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2976 8090 3004 9318
rect 3056 9104 3108 9110
rect 3056 9046 3108 9052
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 2884 7002 2912 7346
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2872 6996 2924 7002
rect 2872 6938 2924 6944
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 2780 5840 2832 5846
rect 2780 5782 2832 5788
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 1768 5160 1820 5166
rect 1768 5102 1820 5108
rect 2596 5160 2648 5166
rect 2596 5102 2648 5108
rect 1780 4078 1808 5102
rect 2228 4684 2280 4690
rect 2228 4626 2280 4632
rect 2320 4684 2372 4690
rect 2320 4626 2372 4632
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 1584 3596 1636 3602
rect 1584 3538 1636 3544
rect 204 2916 256 2922
rect 204 2858 256 2864
rect 216 480 244 2858
rect 664 1964 716 1970
rect 664 1906 716 1912
rect 676 480 704 1906
rect 1124 1896 1176 1902
rect 1124 1838 1176 1844
rect 1136 480 1164 1838
rect 1596 480 1624 3538
rect 1780 3534 1808 4014
rect 2136 4004 2188 4010
rect 2136 3946 2188 3952
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 2044 3392 2096 3398
rect 2044 3334 2096 3340
rect 2056 2990 2084 3334
rect 2148 3058 2176 3946
rect 2240 3194 2268 4626
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 1952 2916 2004 2922
rect 1952 2858 2004 2864
rect 1964 2825 1992 2858
rect 1950 2816 2006 2825
rect 1950 2751 2006 2760
rect 2332 2650 2360 4626
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 2424 4282 2452 4558
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 2424 3670 2452 4218
rect 2792 4049 2820 5782
rect 2884 5778 2912 6190
rect 2976 5817 3004 7142
rect 2962 5808 3018 5817
rect 2872 5772 2924 5778
rect 2962 5743 3018 5752
rect 2872 5714 2924 5720
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 2976 5574 3004 5646
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2778 4040 2834 4049
rect 2778 3975 2834 3984
rect 2884 3890 2912 5102
rect 2976 3942 3004 5510
rect 2792 3862 2912 3890
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2412 3664 2464 3670
rect 2412 3606 2464 3612
rect 2320 2644 2372 2650
rect 2320 2586 2372 2592
rect 2044 2032 2096 2038
rect 2044 1974 2096 1980
rect 2056 480 2084 1974
rect 2516 480 2544 3674
rect 2596 3664 2648 3670
rect 2596 3606 2648 3612
rect 2608 3194 2636 3606
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 2608 3097 2636 3130
rect 2594 3088 2650 3097
rect 2594 3023 2650 3032
rect 2686 2680 2742 2689
rect 2686 2615 2688 2624
rect 2740 2615 2742 2624
rect 2688 2586 2740 2592
rect 2700 2145 2728 2586
rect 2792 2446 2820 3862
rect 2872 2848 2924 2854
rect 2872 2790 2924 2796
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 2686 2136 2742 2145
rect 2686 2071 2742 2080
rect 2792 1193 2820 2382
rect 2778 1184 2834 1193
rect 2778 1119 2834 1128
rect 202 0 258 480
rect 662 0 718 480
rect 1122 0 1178 480
rect 1582 0 1638 480
rect 2042 0 2098 480
rect 2502 0 2558 480
rect 2884 241 2912 2790
rect 2976 480 3004 3878
rect 3068 2854 3096 9046
rect 3160 3670 3188 9438
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 3344 8090 3372 9318
rect 3436 9110 3464 10066
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3424 9104 3476 9110
rect 3424 9046 3476 9052
rect 3436 8945 3464 9046
rect 3422 8936 3478 8945
rect 3422 8871 3478 8880
rect 3424 8832 3476 8838
rect 3424 8774 3476 8780
rect 3436 8430 3464 8774
rect 3528 8498 3556 9318
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3424 8424 3476 8430
rect 3620 8378 3648 11070
rect 3712 10130 3740 11630
rect 3804 11286 3832 12718
rect 3792 11280 3844 11286
rect 3792 11222 3844 11228
rect 3700 10124 3752 10130
rect 3700 10066 3752 10072
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3700 9512 3752 9518
rect 3700 9454 3752 9460
rect 3424 8366 3476 8372
rect 3528 8350 3648 8378
rect 3332 8084 3384 8090
rect 3332 8026 3384 8032
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3344 5642 3372 7142
rect 3436 6458 3464 7142
rect 3424 6452 3476 6458
rect 3424 6394 3476 6400
rect 3332 5636 3384 5642
rect 3332 5578 3384 5584
rect 3528 5166 3556 8350
rect 3606 6896 3662 6905
rect 3606 6831 3662 6840
rect 3620 6390 3648 6831
rect 3608 6384 3660 6390
rect 3608 6326 3660 6332
rect 3608 6112 3660 6118
rect 3608 6054 3660 6060
rect 3620 5914 3648 6054
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3516 5160 3568 5166
rect 3516 5102 3568 5108
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 3240 4684 3292 4690
rect 3240 4626 3292 4632
rect 3148 3664 3200 3670
rect 3148 3606 3200 3612
rect 3252 3194 3280 4626
rect 3332 4616 3384 4622
rect 3332 4558 3384 4564
rect 3344 3194 3372 4558
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3436 3097 3464 4966
rect 3608 4004 3660 4010
rect 3608 3946 3660 3952
rect 3712 3992 3740 9454
rect 3804 8362 3832 9862
rect 3792 8356 3844 8362
rect 3792 8298 3844 8304
rect 3896 5234 3924 13330
rect 4080 13308 4108 13495
rect 4172 13462 4200 14010
rect 4264 13870 4292 15846
rect 4448 15706 4476 15846
rect 4540 15706 4568 16050
rect 4436 15700 4488 15706
rect 4436 15642 4488 15648
rect 4528 15700 4580 15706
rect 4528 15642 4580 15648
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 4618 15056 4674 15065
rect 4618 14991 4674 15000
rect 4632 14260 4660 14991
rect 4724 14958 4752 15438
rect 4712 14952 4764 14958
rect 4712 14894 4764 14900
rect 4632 14232 4752 14260
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4252 13864 4304 13870
rect 4252 13806 4304 13812
rect 4724 13734 4752 14232
rect 4712 13728 4764 13734
rect 4712 13670 4764 13676
rect 4160 13456 4212 13462
rect 4160 13398 4212 13404
rect 4080 13280 4292 13308
rect 4068 13184 4120 13190
rect 4068 13126 4120 13132
rect 3976 12844 4028 12850
rect 3976 12786 4028 12792
rect 3988 12617 4016 12786
rect 3974 12608 4030 12617
rect 3974 12543 4030 12552
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 3988 11898 4016 12174
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 4080 11354 4108 13126
rect 4160 12912 4212 12918
rect 4160 12854 4212 12860
rect 4172 11898 4200 12854
rect 4264 12170 4292 13280
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4816 12442 4844 17002
rect 4908 12617 4936 17836
rect 5000 17490 5028 19722
rect 5092 19310 5120 19790
rect 5276 19774 5396 19802
rect 5080 19304 5132 19310
rect 5080 19246 5132 19252
rect 5092 18766 5120 19246
rect 5172 18964 5224 18970
rect 5172 18906 5224 18912
rect 5080 18760 5132 18766
rect 5080 18702 5132 18708
rect 5092 17785 5120 18702
rect 5078 17776 5134 17785
rect 5078 17711 5134 17720
rect 5000 17462 5120 17490
rect 4988 16040 5040 16046
rect 4988 15982 5040 15988
rect 5000 15570 5028 15982
rect 4988 15564 5040 15570
rect 4988 15506 5040 15512
rect 5000 15026 5028 15506
rect 4988 15020 5040 15026
rect 4988 14962 5040 14968
rect 5092 14362 5120 17462
rect 5184 17202 5212 18906
rect 5368 17785 5396 19774
rect 5552 18970 5580 19994
rect 5540 18964 5592 18970
rect 5540 18906 5592 18912
rect 5538 18320 5594 18329
rect 5538 18255 5594 18264
rect 5354 17776 5410 17785
rect 5410 17734 5488 17762
rect 5354 17711 5410 17720
rect 5172 17196 5224 17202
rect 5172 17138 5224 17144
rect 5264 16992 5316 16998
rect 5000 14334 5120 14362
rect 5184 16952 5264 16980
rect 4894 12608 4950 12617
rect 4894 12543 4950 12552
rect 4804 12436 4856 12442
rect 4804 12378 4856 12384
rect 5000 12374 5028 14334
rect 5080 14272 5132 14278
rect 5080 14214 5132 14220
rect 5092 13870 5120 14214
rect 5080 13864 5132 13870
rect 5080 13806 5132 13812
rect 5184 13716 5212 16952
rect 5264 16934 5316 16940
rect 5264 16448 5316 16454
rect 5264 16390 5316 16396
rect 5276 16046 5304 16390
rect 5460 16266 5488 17734
rect 5552 17270 5580 18255
rect 5644 17338 5672 22320
rect 5816 19508 5868 19514
rect 5816 19450 5868 19456
rect 5828 19394 5856 19450
rect 5828 19366 5948 19394
rect 5724 19236 5776 19242
rect 5724 19178 5776 19184
rect 5816 19236 5868 19242
rect 5816 19178 5868 19184
rect 5736 18970 5764 19178
rect 5724 18964 5776 18970
rect 5724 18906 5776 18912
rect 5736 18290 5764 18906
rect 5828 18834 5856 19178
rect 5816 18828 5868 18834
rect 5816 18770 5868 18776
rect 5724 18284 5776 18290
rect 5724 18226 5776 18232
rect 5816 17672 5868 17678
rect 5816 17614 5868 17620
rect 5632 17332 5684 17338
rect 5632 17274 5684 17280
rect 5540 17264 5592 17270
rect 5828 17218 5856 17614
rect 5540 17206 5592 17212
rect 5644 17190 5856 17218
rect 5460 16238 5580 16266
rect 5356 16108 5408 16114
rect 5356 16050 5408 16056
rect 5264 16040 5316 16046
rect 5264 15982 5316 15988
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 5276 15706 5304 15846
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5368 14822 5396 16050
rect 5552 15994 5580 16238
rect 5460 15966 5580 15994
rect 5460 15065 5488 15966
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5446 15056 5502 15065
rect 5446 14991 5502 15000
rect 5448 14884 5500 14890
rect 5448 14826 5500 14832
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5276 13870 5304 14554
rect 5368 14550 5396 14758
rect 5356 14544 5408 14550
rect 5356 14486 5408 14492
rect 5460 14362 5488 14826
rect 5368 14334 5488 14362
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 5092 13688 5212 13716
rect 4436 12368 4488 12374
rect 4434 12336 4436 12345
rect 4988 12368 5040 12374
rect 4488 12336 4490 12345
rect 4988 12310 5040 12316
rect 4434 12271 4490 12280
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4252 12164 4304 12170
rect 4252 12106 4304 12112
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 4816 11762 4844 12174
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 4158 11656 4214 11665
rect 4158 11591 4214 11600
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 3988 10169 4016 10950
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 3974 10160 4030 10169
rect 3974 10095 4030 10104
rect 4080 9761 4108 10746
rect 4066 9752 4122 9761
rect 4066 9687 4122 9696
rect 4172 9450 4200 11591
rect 5000 11370 5028 12310
rect 4816 11342 5028 11370
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4264 10606 4292 11086
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 4344 9648 4396 9654
rect 4344 9590 4396 9596
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 3974 8800 4030 8809
rect 3974 8735 4030 8744
rect 3988 8566 4016 8735
rect 4080 8634 4108 8978
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 3976 8560 4028 8566
rect 3976 8502 4028 8508
rect 4172 8498 4200 9386
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 4160 8288 4212 8294
rect 4066 8256 4122 8265
rect 4160 8230 4212 8236
rect 4066 8191 4122 8200
rect 4080 8022 4108 8191
rect 4068 8016 4120 8022
rect 4068 7958 4120 7964
rect 3976 7948 4028 7954
rect 3976 7890 4028 7896
rect 3988 5574 4016 7890
rect 4066 7848 4122 7857
rect 4066 7783 4122 7792
rect 4080 7274 4108 7783
rect 4172 7410 4200 8230
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4068 7268 4120 7274
rect 4068 7210 4120 7216
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 3976 4684 4028 4690
rect 3976 4626 4028 4632
rect 3988 4078 4016 4626
rect 4080 4457 4108 5306
rect 4160 5160 4212 5166
rect 4160 5102 4212 5108
rect 4066 4448 4122 4457
rect 4066 4383 4122 4392
rect 3976 4072 4028 4078
rect 3976 4014 4028 4020
rect 3792 4004 3844 4010
rect 3712 3964 3792 3992
rect 3620 3398 3648 3946
rect 3712 3505 3740 3964
rect 3792 3946 3844 3952
rect 3790 3632 3846 3641
rect 3790 3567 3846 3576
rect 3698 3496 3754 3505
rect 3698 3431 3754 3440
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 3422 3088 3478 3097
rect 3422 3023 3424 3032
rect 3476 3023 3478 3032
rect 3424 2994 3476 3000
rect 3056 2848 3108 2854
rect 3148 2848 3200 2854
rect 3056 2790 3108 2796
rect 3146 2816 3148 2825
rect 3200 2816 3202 2825
rect 3146 2751 3202 2760
rect 3436 2446 3464 2994
rect 3424 2440 3476 2446
rect 3424 2382 3476 2388
rect 3804 1442 3832 3567
rect 3988 3534 4016 4014
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 4172 3194 4200 5102
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 4264 3074 4292 9318
rect 4356 9178 4384 9590
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 4724 7886 4752 10202
rect 4816 10130 4844 11342
rect 5092 11268 5120 13688
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 5184 11762 5212 12174
rect 5172 11756 5224 11762
rect 5172 11698 5224 11704
rect 5368 11354 5396 14334
rect 5446 14104 5502 14113
rect 5446 14039 5448 14048
rect 5500 14039 5502 14048
rect 5448 14010 5500 14016
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5460 13462 5488 13874
rect 5552 13802 5580 15846
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5448 13456 5500 13462
rect 5448 13398 5500 13404
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5552 12306 5580 12582
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5356 11348 5408 11354
rect 5356 11290 5408 11296
rect 4908 11240 5120 11268
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4816 9364 4844 10066
rect 4908 9518 4936 11240
rect 4988 10464 5040 10470
rect 4988 10406 5040 10412
rect 5000 10062 5028 10406
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 5000 9586 5028 9998
rect 4988 9580 5040 9586
rect 4988 9522 5040 9528
rect 4896 9512 4948 9518
rect 5000 9489 5028 9522
rect 4896 9454 4948 9460
rect 4986 9480 5042 9489
rect 4986 9415 5042 9424
rect 4816 9336 5028 9364
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4712 7880 4764 7886
rect 4816 7868 4844 8434
rect 4908 8090 4936 8910
rect 4896 8084 4948 8090
rect 4896 8026 4948 8032
rect 4896 7880 4948 7886
rect 4816 7840 4896 7868
rect 4712 7822 4764 7828
rect 4896 7822 4948 7828
rect 4724 7698 4752 7822
rect 4724 7670 4844 7698
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4632 5914 4660 6054
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4724 5574 4752 6802
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4724 5166 4752 5510
rect 4712 5160 4764 5166
rect 4632 5120 4712 5148
rect 4632 4826 4660 5120
rect 4712 5102 4764 5108
rect 4816 5001 4844 7670
rect 4908 6934 4936 7822
rect 4896 6928 4948 6934
rect 4896 6870 4948 6876
rect 5000 5658 5028 9336
rect 5092 8022 5120 10066
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 5172 8968 5224 8974
rect 5172 8910 5224 8916
rect 5080 8016 5132 8022
rect 5080 7958 5132 7964
rect 5184 7342 5212 8910
rect 5276 8294 5304 9658
rect 5460 8922 5488 11494
rect 5644 9042 5672 17190
rect 5920 17134 5948 19366
rect 6000 18828 6052 18834
rect 6000 18770 6052 18776
rect 6012 17814 6040 18770
rect 6000 17808 6052 17814
rect 6000 17750 6052 17756
rect 5908 17128 5960 17134
rect 5908 17070 5960 17076
rect 5998 16824 6054 16833
rect 5998 16759 6054 16768
rect 5816 16652 5868 16658
rect 5816 16594 5868 16600
rect 5828 16114 5856 16594
rect 6012 16454 6040 16759
rect 6000 16448 6052 16454
rect 6000 16390 6052 16396
rect 5816 16108 5868 16114
rect 5816 16050 5868 16056
rect 5816 15972 5868 15978
rect 5816 15914 5868 15920
rect 5724 15904 5776 15910
rect 5724 15846 5776 15852
rect 5736 15366 5764 15846
rect 5828 15366 5856 15914
rect 6012 15502 6040 16390
rect 6000 15496 6052 15502
rect 6000 15438 6052 15444
rect 5724 15360 5776 15366
rect 5724 15302 5776 15308
rect 5816 15360 5868 15366
rect 5816 15302 5868 15308
rect 5908 14952 5960 14958
rect 5908 14894 5960 14900
rect 5816 14476 5868 14482
rect 5816 14418 5868 14424
rect 5724 14408 5776 14414
rect 5724 14350 5776 14356
rect 5736 13734 5764 14350
rect 5828 14006 5856 14418
rect 5920 14278 5948 14894
rect 5998 14648 6054 14657
rect 5998 14583 6054 14592
rect 5908 14272 5960 14278
rect 5908 14214 5960 14220
rect 5816 14000 5868 14006
rect 5816 13942 5868 13948
rect 5724 13728 5776 13734
rect 5724 13670 5776 13676
rect 5724 13320 5776 13326
rect 5920 13308 5948 14214
rect 6012 13841 6040 14583
rect 5998 13832 6054 13841
rect 5998 13767 6054 13776
rect 6012 13734 6040 13767
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 5776 13280 5948 13308
rect 5724 13262 5776 13268
rect 5724 13184 5776 13190
rect 5724 13126 5776 13132
rect 5736 12850 5764 13126
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5828 12782 5856 13280
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 5816 12776 5868 12782
rect 5816 12718 5868 12724
rect 5920 12714 5948 13126
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 5908 12708 5960 12714
rect 5908 12650 5960 12656
rect 5908 11688 5960 11694
rect 5908 11630 5960 11636
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5828 10742 5856 11154
rect 5816 10736 5868 10742
rect 5816 10678 5868 10684
rect 5920 10588 5948 11630
rect 6012 11626 6040 12922
rect 6000 11620 6052 11626
rect 6000 11562 6052 11568
rect 5828 10560 5948 10588
rect 5724 10532 5776 10538
rect 5724 10474 5776 10480
rect 5736 10062 5764 10474
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5828 9994 5856 10560
rect 5816 9988 5868 9994
rect 5816 9930 5868 9936
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 5356 8900 5408 8906
rect 5460 8894 5580 8922
rect 5356 8842 5408 8848
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5276 7546 5304 8230
rect 5368 7546 5396 8842
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 5460 7818 5488 8774
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 5184 7002 5212 7278
rect 5172 6996 5224 7002
rect 5172 6938 5224 6944
rect 5368 6610 5396 7482
rect 5368 6582 5488 6610
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5276 5778 5304 6258
rect 5460 6254 5488 6582
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 5264 5772 5316 5778
rect 5264 5714 5316 5720
rect 5000 5630 5304 5658
rect 4896 5024 4948 5030
rect 4802 4992 4858 5001
rect 4896 4966 4948 4972
rect 4802 4927 4858 4936
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4712 4752 4764 4758
rect 4712 4694 4764 4700
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 4618 3904 4674 3913
rect 4618 3839 4674 3848
rect 4632 3738 4660 3839
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 3436 1414 3832 1442
rect 3896 3046 4292 3074
rect 4342 3088 4398 3097
rect 3436 480 3464 1414
rect 3516 1352 3568 1358
rect 3516 1294 3568 1300
rect 3528 649 3556 1294
rect 3514 640 3570 649
rect 3514 575 3570 584
rect 3896 480 3924 3046
rect 4342 3023 4344 3032
rect 4396 3023 4398 3032
rect 4344 2994 4396 3000
rect 4252 2916 4304 2922
rect 4252 2858 4304 2864
rect 4068 2576 4120 2582
rect 4066 2544 4068 2553
rect 4120 2544 4122 2553
rect 4066 2479 4122 2488
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 4080 1601 4108 2382
rect 4066 1592 4122 1601
rect 4066 1527 4122 1536
rect 4264 1442 4292 2858
rect 4724 2854 4752 4694
rect 4804 4208 4856 4214
rect 4804 4150 4856 4156
rect 4816 3670 4844 4150
rect 4908 3754 4936 4966
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 4988 4004 5040 4010
rect 4988 3946 5040 3952
rect 5000 3913 5028 3946
rect 4986 3904 5042 3913
rect 4986 3839 5042 3848
rect 4908 3726 5028 3754
rect 4804 3664 4856 3670
rect 4896 3664 4948 3670
rect 4804 3606 4856 3612
rect 4894 3632 4896 3641
rect 4948 3632 4950 3641
rect 4894 3567 4950 3576
rect 5000 3516 5028 3726
rect 4816 3488 5028 3516
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4264 1414 4384 1442
rect 4356 480 4384 1414
rect 4816 480 4844 3488
rect 5092 2990 5120 4422
rect 5276 3942 5304 5630
rect 5368 5574 5396 6054
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5460 4758 5488 5850
rect 5552 5030 5580 8894
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5448 4752 5500 4758
rect 5448 4694 5500 4700
rect 5354 4040 5410 4049
rect 5354 3975 5410 3984
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 5184 3738 5212 3878
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5276 3618 5304 3878
rect 5184 3590 5304 3618
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 5184 1358 5212 3590
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 5276 3058 5304 3334
rect 5368 3194 5396 3975
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 5264 2508 5316 2514
rect 5264 2450 5316 2456
rect 5172 1352 5224 1358
rect 5172 1294 5224 1300
rect 5276 480 5304 2450
rect 5460 1902 5488 4694
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5552 4486 5580 4626
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5552 3466 5580 4422
rect 5540 3460 5592 3466
rect 5540 3402 5592 3408
rect 5644 2582 5672 8978
rect 5724 8356 5776 8362
rect 5724 8298 5776 8304
rect 5736 7478 5764 8298
rect 5724 7472 5776 7478
rect 5724 7414 5776 7420
rect 5736 5370 5764 7414
rect 5828 5710 5856 9930
rect 5998 9480 6054 9489
rect 5998 9415 6054 9424
rect 6012 8974 6040 9415
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 6012 7290 6040 7890
rect 5920 7262 6040 7290
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 5724 5364 5776 5370
rect 5724 5306 5776 5312
rect 5920 5166 5948 7262
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 6012 6866 6040 7142
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 6104 6202 6132 22320
rect 6368 20324 6420 20330
rect 6368 20266 6420 20272
rect 6380 18086 6408 20266
rect 6460 19916 6512 19922
rect 6460 19858 6512 19864
rect 6472 19514 6500 19858
rect 6460 19508 6512 19514
rect 6460 19450 6512 19456
rect 6368 18080 6420 18086
rect 6368 18022 6420 18028
rect 6460 18080 6512 18086
rect 6460 18022 6512 18028
rect 6276 17332 6328 17338
rect 6276 17274 6328 17280
rect 6184 16788 6236 16794
rect 6184 16730 6236 16736
rect 6196 16153 6224 16730
rect 6182 16144 6238 16153
rect 6182 16079 6238 16088
rect 6184 15904 6236 15910
rect 6182 15872 6184 15881
rect 6236 15872 6238 15881
rect 6182 15807 6238 15816
rect 6184 15632 6236 15638
rect 6184 15574 6236 15580
rect 6196 14521 6224 15574
rect 6182 14512 6238 14521
rect 6182 14447 6238 14456
rect 6184 13864 6236 13870
rect 6184 13806 6236 13812
rect 6196 12986 6224 13806
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 6184 12640 6236 12646
rect 6182 12608 6184 12617
rect 6236 12608 6238 12617
rect 6182 12543 6238 12552
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 6196 11082 6224 12242
rect 6184 11076 6236 11082
rect 6184 11018 6236 11024
rect 6288 9382 6316 17274
rect 6472 17202 6500 18022
rect 6460 17196 6512 17202
rect 6460 17138 6512 17144
rect 6458 17096 6514 17105
rect 6564 17082 6592 22320
rect 6920 20868 6972 20874
rect 6920 20810 6972 20816
rect 6736 20256 6788 20262
rect 6736 20198 6788 20204
rect 6644 19168 6696 19174
rect 6642 19136 6644 19145
rect 6696 19136 6698 19145
rect 6642 19071 6698 19080
rect 6748 18970 6776 20198
rect 6932 20058 6960 20810
rect 6920 20052 6972 20058
rect 6920 19994 6972 20000
rect 6920 19712 6972 19718
rect 6920 19654 6972 19660
rect 6932 19242 6960 19654
rect 7024 19292 7052 22320
rect 7380 19848 7432 19854
rect 7380 19790 7432 19796
rect 7392 19514 7420 19790
rect 7380 19508 7432 19514
rect 7380 19450 7432 19456
rect 7104 19304 7156 19310
rect 7024 19264 7104 19292
rect 7104 19246 7156 19252
rect 6920 19236 6972 19242
rect 6920 19178 6972 19184
rect 7012 19168 7064 19174
rect 6840 19116 7012 19122
rect 6840 19110 7064 19116
rect 6840 19094 7052 19110
rect 6736 18964 6788 18970
rect 6736 18906 6788 18912
rect 6736 17672 6788 17678
rect 6840 17660 6868 19094
rect 7392 18902 7420 19450
rect 7380 18896 7432 18902
rect 7380 18838 7432 18844
rect 7392 18766 7420 18838
rect 7380 18760 7432 18766
rect 7380 18702 7432 18708
rect 7196 18080 7248 18086
rect 7196 18022 7248 18028
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7208 17882 7236 18022
rect 7196 17876 7248 17882
rect 7196 17818 7248 17824
rect 7104 17740 7156 17746
rect 7104 17682 7156 17688
rect 6788 17632 6868 17660
rect 7012 17672 7064 17678
rect 6736 17614 6788 17620
rect 7012 17614 7064 17620
rect 6736 17128 6788 17134
rect 6564 17054 6684 17082
rect 6736 17070 6788 17076
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 6458 17031 6514 17040
rect 6366 16688 6422 16697
rect 6366 16623 6422 16632
rect 6380 15638 6408 16623
rect 6472 16538 6500 17031
rect 6550 16824 6606 16833
rect 6550 16759 6606 16768
rect 6564 16658 6592 16759
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6472 16510 6592 16538
rect 6460 16448 6512 16454
rect 6460 16390 6512 16396
rect 6472 16250 6500 16390
rect 6460 16244 6512 16250
rect 6460 16186 6512 16192
rect 6458 16144 6514 16153
rect 6458 16079 6514 16088
rect 6472 16046 6500 16079
rect 6460 16040 6512 16046
rect 6460 15982 6512 15988
rect 6564 15638 6592 16510
rect 6368 15632 6420 15638
rect 6368 15574 6420 15580
rect 6552 15632 6604 15638
rect 6552 15574 6604 15580
rect 6380 14890 6408 15574
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 6458 15056 6514 15065
rect 6458 14991 6514 15000
rect 6368 14884 6420 14890
rect 6368 14826 6420 14832
rect 6368 14272 6420 14278
rect 6368 14214 6420 14220
rect 6380 13870 6408 14214
rect 6368 13864 6420 13870
rect 6368 13806 6420 13812
rect 6368 13524 6420 13530
rect 6368 13466 6420 13472
rect 6380 12646 6408 13466
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6472 11558 6500 14991
rect 6564 14482 6592 15302
rect 6552 14476 6604 14482
rect 6552 14418 6604 14424
rect 6552 13388 6604 13394
rect 6552 13330 6604 13336
rect 6460 11552 6512 11558
rect 6460 11494 6512 11500
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6380 10130 6408 10542
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 6380 9722 6408 10066
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6472 9654 6500 10066
rect 6460 9648 6512 9654
rect 6460 9590 6512 9596
rect 6460 9444 6512 9450
rect 6460 9386 6512 9392
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6288 8106 6316 9318
rect 6368 8832 6420 8838
rect 6472 8820 6500 9386
rect 6420 8792 6500 8820
rect 6368 8774 6420 8780
rect 6472 8634 6500 8792
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 6196 8078 6316 8106
rect 6564 8090 6592 13330
rect 6552 8084 6604 8090
rect 6196 7206 6224 8078
rect 6552 8026 6604 8032
rect 6276 8016 6328 8022
rect 6328 7976 6408 8004
rect 6276 7958 6328 7964
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6184 7200 6236 7206
rect 6184 7142 6236 7148
rect 6288 6322 6316 7822
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 6012 6174 6132 6202
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5816 5092 5868 5098
rect 5816 5034 5868 5040
rect 5722 4312 5778 4321
rect 5722 4247 5724 4256
rect 5776 4247 5778 4256
rect 5724 4218 5776 4224
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 5736 3534 5764 4082
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5828 3466 5856 5034
rect 5920 4826 5948 5102
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 5908 4548 5960 4554
rect 5908 4490 5960 4496
rect 5816 3460 5868 3466
rect 5816 3402 5868 3408
rect 5724 3392 5776 3398
rect 5776 3340 5856 3346
rect 5724 3334 5856 3340
rect 5736 3318 5856 3334
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5632 2576 5684 2582
rect 5632 2518 5684 2524
rect 5448 1896 5500 1902
rect 5448 1838 5500 1844
rect 5736 480 5764 2994
rect 5828 2530 5856 3318
rect 5920 2922 5948 4490
rect 6012 4185 6040 6174
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 6104 4826 6132 6054
rect 6288 5914 6316 6258
rect 6380 5914 6408 7976
rect 6656 7562 6684 17054
rect 6748 15366 6776 17070
rect 6840 16998 6868 17070
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6840 16726 6868 16934
rect 6828 16720 6880 16726
rect 6828 16662 6880 16668
rect 7024 16658 7052 17614
rect 7012 16652 7064 16658
rect 7012 16594 7064 16600
rect 6828 16176 6880 16182
rect 6826 16144 6828 16153
rect 6880 16144 6882 16153
rect 6826 16079 6882 16088
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6840 15706 6868 15846
rect 7116 15706 7144 17682
rect 7300 16794 7328 18022
rect 7392 17660 7420 18702
rect 7484 18408 7512 22320
rect 7944 20346 7972 22320
rect 7944 20318 8248 20346
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 7484 18380 7788 18408
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 7484 17814 7512 18022
rect 7472 17808 7524 17814
rect 7472 17750 7524 17756
rect 7472 17672 7524 17678
rect 7392 17632 7472 17660
rect 7472 17614 7524 17620
rect 7484 17134 7512 17614
rect 7472 17128 7524 17134
rect 7472 17070 7524 17076
rect 7380 17060 7432 17066
rect 7380 17002 7432 17008
rect 7288 16788 7340 16794
rect 7288 16730 7340 16736
rect 7196 16720 7248 16726
rect 7196 16662 7248 16668
rect 7208 16046 7236 16662
rect 7392 16658 7420 17002
rect 7380 16652 7432 16658
rect 7380 16594 7432 16600
rect 7196 16040 7248 16046
rect 7248 16000 7328 16028
rect 7196 15982 7248 15988
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 7104 15700 7156 15706
rect 7104 15642 7156 15648
rect 6736 15360 6788 15366
rect 6736 15302 6788 15308
rect 7102 14920 7158 14929
rect 7102 14855 7104 14864
rect 7156 14855 7158 14864
rect 7196 14884 7248 14890
rect 7104 14826 7156 14832
rect 7196 14826 7248 14832
rect 6736 14476 6788 14482
rect 6736 14418 6788 14424
rect 6748 11898 6776 14418
rect 7104 14340 7156 14346
rect 7104 14282 7156 14288
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 6932 13462 6960 13874
rect 6920 13456 6972 13462
rect 6920 13398 6972 13404
rect 6932 12617 6960 13398
rect 7024 13394 7052 14214
rect 7116 13530 7144 14282
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 7024 12782 7052 13330
rect 7012 12776 7064 12782
rect 7012 12718 7064 12724
rect 6918 12608 6974 12617
rect 6918 12543 6974 12552
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 6932 11762 6960 12543
rect 7104 12300 7156 12306
rect 7104 12242 7156 12248
rect 7116 12050 7144 12242
rect 7208 12170 7236 14826
rect 7300 13802 7328 16000
rect 7380 15496 7432 15502
rect 7380 15438 7432 15444
rect 7392 14890 7420 15438
rect 7380 14884 7432 14890
rect 7380 14826 7432 14832
rect 7472 14408 7524 14414
rect 7472 14350 7524 14356
rect 7288 13796 7340 13802
rect 7288 13738 7340 13744
rect 7300 12986 7328 13738
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 7392 12714 7420 13262
rect 7380 12708 7432 12714
rect 7380 12650 7432 12656
rect 7196 12164 7248 12170
rect 7196 12106 7248 12112
rect 7288 12096 7340 12102
rect 7116 12022 7236 12050
rect 7288 12038 7340 12044
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 7024 11014 7052 11834
rect 7104 11824 7156 11830
rect 7104 11766 7156 11772
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 6734 9480 6790 9489
rect 6734 9415 6790 9424
rect 6748 9042 6776 9415
rect 6932 9194 6960 10678
rect 7024 9382 7052 10950
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 6828 9172 6880 9178
rect 6932 9166 7052 9194
rect 6828 9114 6880 9120
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 6472 7534 6684 7562
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6368 5908 6420 5914
rect 6368 5850 6420 5856
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 5998 4176 6054 4185
rect 5998 4111 6054 4120
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 6012 3924 6040 4014
rect 6092 3936 6144 3942
rect 6012 3896 6092 3924
rect 6092 3878 6144 3884
rect 6182 3632 6238 3641
rect 6182 3567 6238 3576
rect 6196 3126 6224 3567
rect 6184 3120 6236 3126
rect 6184 3062 6236 3068
rect 5908 2916 5960 2922
rect 5908 2858 5960 2864
rect 5828 2502 5948 2530
rect 5920 2446 5948 2502
rect 5908 2440 5960 2446
rect 5908 2382 5960 2388
rect 6196 480 6224 3062
rect 6288 3058 6316 5646
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6380 3534 6408 4082
rect 6368 3528 6420 3534
rect 6368 3470 6420 3476
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 6380 2446 6408 3470
rect 6472 2514 6500 7534
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6564 6186 6592 7142
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6552 6180 6604 6186
rect 6552 6122 6604 6128
rect 6656 5642 6684 6258
rect 6644 5636 6696 5642
rect 6644 5578 6696 5584
rect 6748 5114 6776 8978
rect 6840 7002 6868 9114
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6932 8090 6960 8910
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 7024 7970 7052 9166
rect 6932 7942 7052 7970
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6932 6934 6960 7942
rect 7116 7886 7144 11766
rect 7208 10742 7236 12022
rect 7196 10736 7248 10742
rect 7196 10678 7248 10684
rect 7300 10470 7328 12038
rect 7392 11354 7420 12038
rect 7484 11898 7512 14350
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7668 13138 7696 13670
rect 7576 13110 7696 13138
rect 7576 12306 7604 13110
rect 7656 12980 7708 12986
rect 7656 12922 7708 12928
rect 7564 12300 7616 12306
rect 7564 12242 7616 12248
rect 7564 12164 7616 12170
rect 7564 12106 7616 12112
rect 7472 11892 7524 11898
rect 7472 11834 7524 11840
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7484 11286 7512 11494
rect 7472 11280 7524 11286
rect 7472 11222 7524 11228
rect 7576 10826 7604 12106
rect 7484 10798 7604 10826
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 7208 9518 7236 10406
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7208 8242 7236 9318
rect 7300 8362 7328 10406
rect 7484 10266 7512 10798
rect 7668 10690 7696 12922
rect 7760 11830 7788 18380
rect 8116 18284 8168 18290
rect 8116 18226 8168 18232
rect 8128 18068 8156 18226
rect 8220 18170 8248 20318
rect 8404 19174 8432 22320
rect 8864 20074 8892 22320
rect 8772 20046 8892 20074
rect 8772 19310 8800 20046
rect 8852 19916 8904 19922
rect 8852 19858 8904 19864
rect 8760 19304 8812 19310
rect 8760 19246 8812 19252
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 8864 18970 8892 19858
rect 9036 19168 9088 19174
rect 9036 19110 9088 19116
rect 8852 18964 8904 18970
rect 8852 18906 8904 18912
rect 8392 18624 8444 18630
rect 8392 18566 8444 18572
rect 8404 18290 8432 18566
rect 8864 18290 8892 18906
rect 8392 18284 8444 18290
rect 8392 18226 8444 18232
rect 8852 18284 8904 18290
rect 8852 18226 8904 18232
rect 8220 18142 8432 18170
rect 8300 18080 8352 18086
rect 8128 18040 8248 18068
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 8220 17746 8248 18040
rect 8300 18022 8352 18028
rect 8208 17740 8260 17746
rect 8208 17682 8260 17688
rect 8220 17338 8248 17682
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 8208 16992 8260 16998
rect 8208 16934 8260 16940
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 8220 16114 8248 16934
rect 8312 16794 8340 18022
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 8298 16008 8354 16017
rect 8298 15943 8354 15952
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 8024 15564 8076 15570
rect 8024 15506 8076 15512
rect 8036 15473 8064 15506
rect 8022 15464 8078 15473
rect 8022 15399 8078 15408
rect 8036 15094 8064 15399
rect 8024 15088 8076 15094
rect 8024 15030 8076 15036
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 7840 14476 7892 14482
rect 7840 14418 7892 14424
rect 7852 14278 7880 14418
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 8220 13954 8248 14350
rect 8128 13938 8248 13954
rect 8116 13932 8248 13938
rect 8168 13926 8248 13932
rect 8116 13874 8168 13880
rect 8208 13796 8260 13802
rect 8208 13738 8260 13744
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 8220 13394 8248 13738
rect 8312 13462 8340 15943
rect 8300 13456 8352 13462
rect 8300 13398 8352 13404
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 7748 11824 7800 11830
rect 7748 11766 7800 11772
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 7748 11076 7800 11082
rect 7748 11018 7800 11024
rect 7576 10662 7696 10690
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7380 10192 7432 10198
rect 7380 10134 7432 10140
rect 7392 8838 7420 10134
rect 7484 9518 7512 10202
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7470 9208 7526 9217
rect 7470 9143 7472 9152
rect 7524 9143 7526 9152
rect 7472 9114 7524 9120
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7484 8945 7512 8978
rect 7470 8936 7526 8945
rect 7470 8871 7526 8880
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7288 8356 7340 8362
rect 7288 8298 7340 8304
rect 7208 8214 7328 8242
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 6920 6928 6972 6934
rect 6920 6870 6972 6876
rect 6932 6390 6960 6870
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 6920 6248 6972 6254
rect 6918 6216 6920 6225
rect 6972 6216 6974 6225
rect 6918 6151 6974 6160
rect 6920 5840 6972 5846
rect 6920 5782 6972 5788
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6840 5574 6868 5646
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6840 5166 6868 5510
rect 6564 5086 6776 5114
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6564 3398 6592 5086
rect 6736 4548 6788 4554
rect 6736 4490 6788 4496
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 6460 2508 6512 2514
rect 6460 2450 6512 2456
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 6472 2106 6500 2450
rect 6460 2100 6512 2106
rect 6460 2042 6512 2048
rect 6656 480 6684 4014
rect 6748 3738 6776 4490
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6840 3534 6868 5102
rect 6932 5030 6960 5782
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6932 4622 6960 4966
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6920 4208 6972 4214
rect 6920 4150 6972 4156
rect 7024 4162 7052 7822
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 7208 7342 7236 7686
rect 7300 7342 7328 8214
rect 7196 7336 7248 7342
rect 7196 7278 7248 7284
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 7116 6798 7144 7142
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7208 6390 7236 6598
rect 7300 6458 7328 7142
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7196 6384 7248 6390
rect 7196 6326 7248 6332
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7300 5846 7328 6258
rect 7288 5840 7340 5846
rect 7288 5782 7340 5788
rect 7288 4548 7340 4554
rect 7288 4490 7340 4496
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 6828 2916 6880 2922
rect 6828 2858 6880 2864
rect 6840 2122 6868 2858
rect 6932 2310 6960 4150
rect 7024 4134 7144 4162
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 7024 2582 7052 3538
rect 7012 2576 7064 2582
rect 7012 2518 7064 2524
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 7024 2122 7052 2246
rect 6840 2094 7052 2122
rect 7116 480 7144 4134
rect 7196 2848 7248 2854
rect 7196 2790 7248 2796
rect 7208 1970 7236 2790
rect 7300 2650 7328 4490
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 7392 2514 7420 6598
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7484 3398 7512 6190
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7576 3126 7604 10662
rect 7656 10532 7708 10538
rect 7656 10474 7708 10480
rect 7668 9042 7696 10474
rect 7760 9926 7788 11018
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 8220 10198 8248 10406
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 8312 9654 8340 9998
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7760 8362 7788 9318
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 8220 9042 8248 9522
rect 8300 9376 8352 9382
rect 8404 9364 8432 18142
rect 8484 17672 8536 17678
rect 8484 17614 8536 17620
rect 8496 16658 8524 17614
rect 8668 17128 8720 17134
rect 8668 17070 8720 17076
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8680 15366 8708 17070
rect 8852 16516 8904 16522
rect 8852 16458 8904 16464
rect 8864 15910 8892 16458
rect 8852 15904 8904 15910
rect 8852 15846 8904 15852
rect 8668 15360 8720 15366
rect 8668 15302 8720 15308
rect 8760 15156 8812 15162
rect 8760 15098 8812 15104
rect 8484 14816 8536 14822
rect 8484 14758 8536 14764
rect 8496 14550 8524 14758
rect 8772 14550 8800 15098
rect 8484 14544 8536 14550
rect 8484 14486 8536 14492
rect 8760 14544 8812 14550
rect 8760 14486 8812 14492
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 8772 14074 8800 14350
rect 8760 14068 8812 14074
rect 8760 14010 8812 14016
rect 8758 13832 8814 13841
rect 8758 13767 8814 13776
rect 8772 13734 8800 13767
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8772 13530 8800 13670
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 8496 11762 8524 13262
rect 8760 12368 8812 12374
rect 8760 12310 8812 12316
rect 8576 12232 8628 12238
rect 8772 12209 8800 12310
rect 8576 12174 8628 12180
rect 8758 12200 8814 12209
rect 8484 11756 8536 11762
rect 8484 11698 8536 11704
rect 8484 11620 8536 11626
rect 8484 11562 8536 11568
rect 8496 11121 8524 11562
rect 8588 11286 8616 12174
rect 8758 12135 8814 12144
rect 8758 11384 8814 11393
rect 8758 11319 8814 11328
rect 8576 11280 8628 11286
rect 8576 11222 8628 11228
rect 8482 11112 8538 11121
rect 8482 11047 8538 11056
rect 8588 10810 8616 11222
rect 8772 11218 8800 11319
rect 8760 11212 8812 11218
rect 8760 11154 8812 11160
rect 8668 11008 8720 11014
rect 8668 10950 8720 10956
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 8680 10674 8708 10950
rect 8760 10804 8812 10810
rect 8760 10746 8812 10752
rect 8668 10668 8720 10674
rect 8668 10610 8720 10616
rect 8576 10600 8628 10606
rect 8574 10568 8576 10577
rect 8628 10568 8630 10577
rect 8574 10503 8630 10512
rect 8668 10532 8720 10538
rect 8668 10474 8720 10480
rect 8680 10266 8708 10474
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8680 9586 8708 10202
rect 8772 10062 8800 10746
rect 8864 10470 8892 15846
rect 8942 15056 8998 15065
rect 8942 14991 8998 15000
rect 9048 15008 9076 19110
rect 9324 18970 9352 22320
rect 9404 19168 9456 19174
rect 9404 19110 9456 19116
rect 9312 18964 9364 18970
rect 9312 18906 9364 18912
rect 9416 18902 9444 19110
rect 9404 18896 9456 18902
rect 9404 18838 9456 18844
rect 9128 18148 9180 18154
rect 9128 18090 9180 18096
rect 9680 18148 9732 18154
rect 9680 18090 9732 18096
rect 9140 17882 9168 18090
rect 9692 17882 9720 18090
rect 9128 17876 9180 17882
rect 9128 17818 9180 17824
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9496 17740 9548 17746
rect 9496 17682 9548 17688
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 9324 15638 9352 16050
rect 9220 15632 9272 15638
rect 9220 15574 9272 15580
rect 9312 15632 9364 15638
rect 9312 15574 9364 15580
rect 8956 14822 8984 14991
rect 9048 14980 9168 15008
rect 9034 14920 9090 14929
rect 9034 14855 9090 14864
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 8942 14376 8998 14385
rect 8942 14311 8998 14320
rect 8956 13938 8984 14311
rect 8944 13932 8996 13938
rect 8944 13874 8996 13880
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8852 10124 8904 10130
rect 8852 10066 8904 10072
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8576 9376 8628 9382
rect 8404 9336 8576 9364
rect 8300 9318 8352 9324
rect 8576 9318 8628 9324
rect 8312 9217 8340 9318
rect 8298 9208 8354 9217
rect 8298 9143 8354 9152
rect 7932 9036 7984 9042
rect 7932 8978 7984 8984
rect 8116 9036 8168 9042
rect 8116 8978 8168 8984
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 7944 8809 7972 8978
rect 7930 8800 7986 8809
rect 7930 8735 7986 8744
rect 8128 8673 8156 8978
rect 8114 8664 8170 8673
rect 8114 8599 8170 8608
rect 7748 8356 7800 8362
rect 7748 8298 7800 8304
rect 7760 7546 7788 8298
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 8036 7478 8064 7822
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 8206 7440 8262 7449
rect 8206 7375 8262 7384
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 8220 6934 8248 7375
rect 8208 6928 8260 6934
rect 8208 6870 8260 6876
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 7668 4146 7696 6394
rect 7932 6180 7984 6186
rect 8024 6180 8076 6186
rect 7984 6140 8024 6168
rect 7932 6122 7984 6128
rect 8024 6122 8076 6128
rect 8208 6180 8260 6186
rect 8208 6122 8260 6128
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 8220 5681 8248 6122
rect 8206 5672 8262 5681
rect 8206 5607 8262 5616
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 7932 4752 7984 4758
rect 7932 4694 7984 4700
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 7852 4282 7880 4558
rect 7944 4282 7972 4694
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 7840 4276 7892 4282
rect 7840 4218 7892 4224
rect 7932 4276 7984 4282
rect 7932 4218 7984 4224
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 7668 3602 7696 4082
rect 8128 4060 8156 4558
rect 8220 4214 8248 5170
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 8128 4032 8248 4060
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 8220 3720 8248 4032
rect 8128 3692 8248 3720
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7932 3596 7984 3602
rect 7932 3538 7984 3544
rect 7564 3120 7616 3126
rect 7564 3062 7616 3068
rect 7668 3040 7696 3538
rect 7944 3058 7972 3538
rect 8128 3398 8156 3692
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 7932 3052 7984 3058
rect 7668 3012 7788 3040
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 7562 2952 7618 2961
rect 7380 2508 7432 2514
rect 7380 2450 7432 2456
rect 7196 1964 7248 1970
rect 7196 1906 7248 1912
rect 7484 1902 7512 2926
rect 7562 2887 7618 2896
rect 7472 1896 7524 1902
rect 7472 1838 7524 1844
rect 7576 480 7604 2887
rect 7760 2378 7788 3012
rect 7932 2994 7984 3000
rect 8128 2922 8156 3334
rect 8220 3058 8248 3470
rect 8199 3052 8251 3058
rect 8199 2994 8251 3000
rect 8116 2916 8168 2922
rect 8116 2858 8168 2864
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 8312 2632 8340 9143
rect 8392 9104 8444 9110
rect 8390 9072 8392 9081
rect 8444 9072 8446 9081
rect 8390 9007 8446 9016
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8680 8265 8708 8366
rect 8666 8256 8722 8265
rect 8666 8191 8722 8200
rect 8484 8016 8536 8022
rect 8390 7984 8446 7993
rect 8484 7958 8536 7964
rect 8390 7919 8392 7928
rect 8444 7919 8446 7928
rect 8392 7890 8444 7896
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 8404 4486 8432 7754
rect 8496 5370 8524 7958
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 8588 7546 8616 7890
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8680 7256 8708 7822
rect 8588 7228 8708 7256
rect 8588 7002 8616 7228
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 8668 6928 8720 6934
rect 8668 6870 8720 6876
rect 8680 6361 8708 6870
rect 8666 6352 8722 6361
rect 8666 6287 8722 6296
rect 8484 5364 8536 5370
rect 8484 5306 8536 5312
rect 8772 5273 8800 8774
rect 8864 6474 8892 10066
rect 8956 8294 8984 13874
rect 9048 12850 9076 14855
rect 9140 13818 9168 14980
rect 9232 14618 9260 15574
rect 9324 15434 9352 15574
rect 9312 15428 9364 15434
rect 9312 15370 9364 15376
rect 9312 15088 9364 15094
rect 9312 15030 9364 15036
rect 9220 14612 9272 14618
rect 9220 14554 9272 14560
rect 9324 14362 9352 15030
rect 9508 15026 9536 17682
rect 9680 17604 9732 17610
rect 9680 17546 9732 17552
rect 9692 17134 9720 17546
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9692 16590 9720 16934
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9784 16522 9812 22320
rect 9864 19916 9916 19922
rect 9864 19858 9916 19864
rect 9876 17678 9904 19858
rect 10138 18864 10194 18873
rect 10138 18799 10194 18808
rect 10152 18766 10180 18799
rect 10140 18760 10192 18766
rect 10140 18702 10192 18708
rect 10048 18352 10100 18358
rect 10048 18294 10100 18300
rect 9956 18080 10008 18086
rect 9956 18022 10008 18028
rect 9864 17672 9916 17678
rect 9864 17614 9916 17620
rect 9772 16516 9824 16522
rect 9772 16458 9824 16464
rect 9772 16040 9824 16046
rect 9772 15982 9824 15988
rect 9496 15020 9548 15026
rect 9496 14962 9548 14968
rect 9588 14952 9640 14958
rect 9508 14900 9588 14906
rect 9508 14894 9640 14900
rect 9508 14878 9628 14894
rect 9508 14618 9536 14878
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 9404 14476 9456 14482
rect 9404 14418 9456 14424
rect 9232 14334 9352 14362
rect 9232 14113 9260 14334
rect 9312 14272 9364 14278
rect 9312 14214 9364 14220
rect 9218 14104 9274 14113
rect 9218 14039 9274 14048
rect 9140 13790 9260 13818
rect 9128 13728 9180 13734
rect 9128 13670 9180 13676
rect 9036 12844 9088 12850
rect 9036 12786 9088 12792
rect 9140 12646 9168 13670
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 9232 12424 9260 13790
rect 9324 12918 9352 14214
rect 9312 12912 9364 12918
rect 9312 12854 9364 12860
rect 9232 12396 9352 12424
rect 9034 12336 9090 12345
rect 9034 12271 9090 12280
rect 9220 12300 9272 12306
rect 8944 8288 8996 8294
rect 8944 8230 8996 8236
rect 9048 8106 9076 12271
rect 9220 12242 9272 12248
rect 9126 11792 9182 11801
rect 9126 11727 9182 11736
rect 8956 8078 9076 8106
rect 8956 6798 8984 8078
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 9140 6633 9168 11727
rect 9232 10674 9260 12242
rect 9324 11801 9352 12396
rect 9310 11792 9366 11801
rect 9310 11727 9366 11736
rect 9416 11558 9444 14418
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9508 14074 9536 14214
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9692 13802 9720 14350
rect 9680 13796 9732 13802
rect 9680 13738 9732 13744
rect 9784 13530 9812 15982
rect 9876 14113 9904 17614
rect 9968 16794 9996 18022
rect 10060 17338 10088 18294
rect 10138 17776 10194 17785
rect 10138 17711 10140 17720
rect 10192 17711 10194 17720
rect 10140 17682 10192 17688
rect 10048 17332 10100 17338
rect 10048 17274 10100 17280
rect 10060 17202 10088 17274
rect 10048 17196 10100 17202
rect 10048 17138 10100 17144
rect 10244 16810 10272 22320
rect 10324 19304 10376 19310
rect 10324 19246 10376 19252
rect 10336 17728 10364 19246
rect 10704 18873 10732 22320
rect 10876 20052 10928 20058
rect 10796 20012 10876 20040
rect 10690 18864 10746 18873
rect 10690 18799 10746 18808
rect 10692 18624 10744 18630
rect 10692 18566 10744 18572
rect 10416 17740 10468 17746
rect 10336 17700 10416 17728
rect 10336 17134 10364 17700
rect 10416 17682 10468 17688
rect 10508 17672 10560 17678
rect 10508 17614 10560 17620
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 10336 16998 10364 17070
rect 10324 16992 10376 16998
rect 10324 16934 10376 16940
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 10060 16782 10272 16810
rect 9956 16652 10008 16658
rect 10060 16640 10088 16782
rect 10140 16720 10192 16726
rect 10140 16662 10192 16668
rect 10008 16612 10088 16640
rect 9956 16594 10008 16600
rect 9968 16561 9996 16594
rect 9954 16552 10010 16561
rect 9954 16487 10010 16496
rect 9956 16448 10008 16454
rect 9956 16390 10008 16396
rect 9968 16046 9996 16390
rect 10152 16250 10180 16662
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 9956 16040 10008 16046
rect 9956 15982 10008 15988
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 9862 14104 9918 14113
rect 10060 14074 10088 15846
rect 10232 15632 10284 15638
rect 10232 15574 10284 15580
rect 10244 15094 10272 15574
rect 10336 15570 10364 16934
rect 10520 16590 10548 17614
rect 10508 16584 10560 16590
rect 10508 16526 10560 16532
rect 10704 15978 10732 18566
rect 10692 15972 10744 15978
rect 10612 15932 10692 15960
rect 10324 15564 10376 15570
rect 10324 15506 10376 15512
rect 10232 15088 10284 15094
rect 10232 15030 10284 15036
rect 10336 15026 10364 15506
rect 10324 15020 10376 15026
rect 10324 14962 10376 14968
rect 10336 14464 10364 14962
rect 10416 14476 10468 14482
rect 10336 14436 10416 14464
rect 10416 14418 10468 14424
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 9862 14039 9918 14048
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9770 13424 9826 13433
rect 9680 13388 9732 13394
rect 9770 13359 9826 13368
rect 9680 13330 9732 13336
rect 9692 12986 9720 13330
rect 9784 13326 9812 13359
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9876 13002 9904 13874
rect 9968 13258 9996 13874
rect 10138 13832 10194 13841
rect 10138 13767 10194 13776
rect 10152 13433 10180 13767
rect 10138 13424 10194 13433
rect 10138 13359 10194 13368
rect 9956 13252 10008 13258
rect 9956 13194 10008 13200
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9784 12974 9904 13002
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 9508 12646 9536 12786
rect 9678 12744 9734 12753
rect 9678 12679 9734 12688
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9692 11880 9720 12679
rect 9508 11852 9720 11880
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9220 10668 9272 10674
rect 9220 10610 9272 10616
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 9232 8922 9260 10406
rect 9324 9042 9352 11494
rect 9416 9518 9444 11494
rect 9508 9897 9536 11852
rect 9586 11758 9642 11767
rect 9586 11693 9642 11702
rect 9588 11348 9640 11354
rect 9680 11348 9732 11354
rect 9640 11308 9680 11336
rect 9588 11290 9640 11296
rect 9680 11290 9732 11296
rect 9784 11257 9812 12974
rect 9864 12912 9916 12918
rect 9864 12854 9916 12860
rect 9876 12442 9904 12854
rect 9968 12782 9996 13194
rect 9956 12776 10008 12782
rect 9956 12718 10008 12724
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 9876 11801 9904 12174
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 9862 11792 9918 11801
rect 9862 11727 9918 11736
rect 9770 11248 9826 11257
rect 9588 11212 9640 11218
rect 9770 11183 9826 11192
rect 9588 11154 9640 11160
rect 9600 11098 9628 11154
rect 9876 11098 9904 11727
rect 9600 11070 9904 11098
rect 9954 11112 10010 11121
rect 9954 11047 10010 11056
rect 9862 10840 9918 10849
rect 9862 10775 9918 10784
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9692 10266 9720 10542
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9494 9888 9550 9897
rect 9494 9823 9550 9832
rect 9784 9586 9812 10406
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9588 9512 9640 9518
rect 9588 9454 9640 9460
rect 9496 9444 9548 9450
rect 9496 9386 9548 9392
rect 9404 9376 9456 9382
rect 9402 9344 9404 9353
rect 9456 9344 9458 9353
rect 9402 9279 9458 9288
rect 9508 9178 9536 9386
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9312 9036 9364 9042
rect 9312 8978 9364 8984
rect 9232 8894 9536 8922
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9232 6662 9260 7822
rect 9312 7200 9364 7206
rect 9312 7142 9364 7148
rect 9220 6656 9272 6662
rect 9126 6624 9182 6633
rect 9220 6598 9272 6604
rect 9126 6559 9182 6568
rect 9232 6474 9260 6598
rect 8864 6446 9076 6474
rect 8852 5568 8904 5574
rect 8852 5510 8904 5516
rect 8482 5264 8538 5273
rect 8482 5199 8538 5208
rect 8758 5264 8814 5273
rect 8758 5199 8814 5208
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8496 3942 8524 5199
rect 8864 5166 8892 5510
rect 8852 5160 8904 5166
rect 8852 5102 8904 5108
rect 8864 4758 8892 5102
rect 8760 4752 8812 4758
rect 8760 4694 8812 4700
rect 8852 4752 8904 4758
rect 8852 4694 8904 4700
rect 8772 4321 8800 4694
rect 8758 4312 8814 4321
rect 8758 4247 8814 4256
rect 8668 4140 8720 4146
rect 8668 4082 8720 4088
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8588 3670 8616 3878
rect 8576 3664 8628 3670
rect 8576 3606 8628 3612
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8404 2650 8432 3130
rect 8128 2604 8340 2632
rect 8392 2644 8444 2650
rect 8024 2508 8076 2514
rect 8024 2450 8076 2456
rect 7748 2372 7800 2378
rect 7748 2314 7800 2320
rect 8036 2038 8064 2450
rect 8024 2032 8076 2038
rect 8024 1974 8076 1980
rect 8128 480 8156 2604
rect 8392 2586 8444 2592
rect 8496 2582 8524 3538
rect 8576 2916 8628 2922
rect 8576 2858 8628 2864
rect 8484 2576 8536 2582
rect 8484 2518 8536 2524
rect 8588 480 8616 2858
rect 8680 2258 8708 4082
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 8956 3194 8984 3674
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 8760 2304 8812 2310
rect 8680 2252 8760 2258
rect 8680 2246 8812 2252
rect 8680 2230 8800 2246
rect 9048 480 9076 6446
rect 9140 6446 9260 6474
rect 9140 6254 9168 6446
rect 9220 6384 9272 6390
rect 9220 6326 9272 6332
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 9232 5846 9260 6326
rect 9220 5840 9272 5846
rect 9220 5782 9272 5788
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9140 4622 9168 5170
rect 9220 5160 9272 5166
rect 9324 5148 9352 7142
rect 9272 5120 9352 5148
rect 9220 5102 9272 5108
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 9232 2854 9260 5102
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 9324 4282 9352 4626
rect 9312 4276 9364 4282
rect 9312 4218 9364 4224
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9220 2848 9272 2854
rect 9220 2790 9272 2796
rect 9324 2446 9352 3130
rect 9416 2802 9444 8230
rect 9508 5642 9536 8894
rect 9600 8838 9628 9454
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9692 8974 9720 9318
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9692 8634 9720 8910
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9678 8528 9734 8537
rect 9678 8463 9734 8472
rect 9772 8492 9824 8498
rect 9692 8430 9720 8463
rect 9772 8434 9824 8440
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9784 8265 9812 8434
rect 9770 8256 9826 8265
rect 9770 8191 9826 8200
rect 9680 7948 9732 7954
rect 9784 7936 9812 8191
rect 9732 7908 9812 7936
rect 9680 7890 9732 7896
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9600 7410 9628 7686
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 9600 6866 9628 7346
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9692 6798 9720 7890
rect 9876 7721 9904 10775
rect 9968 10606 9996 11047
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 9968 10470 9996 10542
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 10060 9489 10088 11834
rect 10046 9480 10102 9489
rect 10046 9415 10102 9424
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 10060 9042 10088 9318
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 10048 8832 10100 8838
rect 10048 8774 10100 8780
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 9968 8022 9996 8570
rect 9956 8016 10008 8022
rect 9956 7958 10008 7964
rect 9862 7712 9918 7721
rect 9862 7647 9918 7656
rect 10060 7562 10088 8774
rect 9784 7534 10088 7562
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9588 6724 9640 6730
rect 9588 6666 9640 6672
rect 9600 5953 9628 6666
rect 9586 5944 9642 5953
rect 9586 5879 9642 5888
rect 9588 5840 9640 5846
rect 9588 5782 9640 5788
rect 9496 5636 9548 5642
rect 9496 5578 9548 5584
rect 9494 3224 9550 3233
rect 9494 3159 9550 3168
rect 9508 2922 9536 3159
rect 9496 2916 9548 2922
rect 9496 2858 9548 2864
rect 9416 2774 9536 2802
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 9508 480 9536 2774
rect 9600 2038 9628 5782
rect 9784 4146 9812 7534
rect 9956 7472 10008 7478
rect 9956 7414 10008 7420
rect 10046 7440 10102 7449
rect 9862 7304 9918 7313
rect 9862 7239 9918 7248
rect 9876 4146 9904 7239
rect 9968 4282 9996 7414
rect 10046 7375 10048 7384
rect 10100 7375 10102 7384
rect 10048 7346 10100 7352
rect 10152 7290 10180 13359
rect 10244 10606 10272 13874
rect 10414 13832 10470 13841
rect 10414 13767 10470 13776
rect 10428 13394 10456 13767
rect 10416 13388 10468 13394
rect 10416 13330 10468 13336
rect 10324 13184 10376 13190
rect 10324 13126 10376 13132
rect 10336 12714 10364 13126
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 10324 12708 10376 12714
rect 10324 12650 10376 12656
rect 10428 12374 10456 12718
rect 10416 12368 10468 12374
rect 10416 12310 10468 12316
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10336 11558 10364 11698
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10232 10600 10284 10606
rect 10520 10577 10548 14350
rect 10612 11898 10640 15932
rect 10692 15914 10744 15920
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10704 13530 10732 14350
rect 10796 13530 10824 20012
rect 10876 19994 10928 20000
rect 10968 19848 11020 19854
rect 10968 19790 11020 19796
rect 10980 19514 11008 19790
rect 10968 19508 11020 19514
rect 10968 19450 11020 19456
rect 10980 19242 11008 19450
rect 11164 19258 11192 22320
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 10968 19236 11020 19242
rect 10968 19178 11020 19184
rect 11072 19230 11192 19258
rect 10968 18624 11020 18630
rect 10968 18566 11020 18572
rect 10980 18426 11008 18566
rect 10968 18420 11020 18426
rect 10968 18362 11020 18368
rect 11072 18170 11100 19230
rect 11428 19168 11480 19174
rect 11428 19110 11480 19116
rect 11440 18952 11468 19110
rect 11164 18924 11468 18952
rect 11164 18290 11192 18924
rect 11336 18828 11388 18834
rect 11336 18770 11388 18776
rect 11348 18737 11376 18770
rect 11334 18728 11390 18737
rect 11334 18663 11390 18672
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 11624 18358 11652 22320
rect 11704 19848 11756 19854
rect 11704 19790 11756 19796
rect 11612 18352 11664 18358
rect 11612 18294 11664 18300
rect 11152 18284 11204 18290
rect 11152 18226 11204 18232
rect 11072 18142 11192 18170
rect 10876 18080 10928 18086
rect 10876 18022 10928 18028
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 10888 17542 10916 18022
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10888 16794 10916 17070
rect 11072 16794 11100 18022
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 11164 16658 11192 18142
rect 11716 17898 11744 19790
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11808 19242 11836 19654
rect 11796 19236 11848 19242
rect 11796 19178 11848 19184
rect 11888 18964 11940 18970
rect 11888 18906 11940 18912
rect 11796 18828 11848 18834
rect 11796 18770 11848 18776
rect 11808 18426 11836 18770
rect 11796 18420 11848 18426
rect 11796 18362 11848 18368
rect 11796 18284 11848 18290
rect 11796 18226 11848 18232
rect 11624 17870 11744 17898
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 11428 17264 11480 17270
rect 11428 17206 11480 17212
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 11440 16590 11468 17206
rect 11428 16584 11480 16590
rect 11428 16526 11480 16532
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11518 16144 11574 16153
rect 10968 16108 11020 16114
rect 11624 16130 11652 17870
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11716 17338 11744 17682
rect 11808 17542 11836 18226
rect 11796 17536 11848 17542
rect 11796 17478 11848 17484
rect 11704 17332 11756 17338
rect 11704 17274 11756 17280
rect 11716 17202 11744 17274
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11716 16590 11744 17138
rect 11796 16652 11848 16658
rect 11796 16594 11848 16600
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11624 16102 11744 16130
rect 11518 16079 11574 16088
rect 10968 16050 11020 16056
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10888 15366 10916 15982
rect 10980 15366 11008 16050
rect 11532 16046 11560 16079
rect 11520 16040 11572 16046
rect 11520 15982 11572 15988
rect 11612 16040 11664 16046
rect 11612 15982 11664 15988
rect 11624 15706 11652 15982
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11428 15700 11480 15706
rect 11428 15642 11480 15648
rect 11612 15700 11664 15706
rect 11612 15642 11664 15648
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 10968 15360 11020 15366
rect 10968 15302 11020 15308
rect 10888 13938 10916 15302
rect 10980 14958 11008 15302
rect 10968 14952 11020 14958
rect 10968 14894 11020 14900
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 11072 14822 11100 14894
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 11058 14512 11114 14521
rect 11058 14447 11114 14456
rect 11072 13938 11100 14447
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10784 13524 10836 13530
rect 10784 13466 10836 13472
rect 10796 12442 10824 13466
rect 10888 13326 10916 13874
rect 11164 13870 11192 15642
rect 11440 15450 11468 15642
rect 11716 15638 11744 16102
rect 11704 15632 11756 15638
rect 11704 15574 11756 15580
rect 11440 15422 11652 15450
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11624 15094 11652 15422
rect 11612 15088 11664 15094
rect 11612 15030 11664 15036
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 11440 14482 11468 14758
rect 11428 14476 11480 14482
rect 11480 14436 11652 14464
rect 11428 14418 11480 14424
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11624 13870 11652 14436
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 11612 13864 11664 13870
rect 11612 13806 11664 13812
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11164 13530 11192 13670
rect 11334 13560 11390 13569
rect 11152 13524 11204 13530
rect 11334 13495 11390 13504
rect 11152 13466 11204 13472
rect 11348 13394 11376 13495
rect 11336 13388 11388 13394
rect 11336 13330 11388 13336
rect 10876 13320 10928 13326
rect 11060 13320 11112 13326
rect 10876 13262 10928 13268
rect 11058 13288 11060 13297
rect 11152 13320 11204 13326
rect 11112 13288 11114 13297
rect 11152 13262 11204 13268
rect 11058 13223 11114 13232
rect 11164 12714 11192 13262
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11716 12714 11744 13670
rect 11152 12708 11204 12714
rect 11152 12650 11204 12656
rect 11612 12708 11664 12714
rect 11612 12650 11664 12656
rect 11704 12708 11756 12714
rect 11704 12650 11756 12656
rect 11624 12442 11652 12650
rect 10784 12436 10836 12442
rect 10784 12378 10836 12384
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 10692 12368 10744 12374
rect 10692 12310 10744 12316
rect 10704 11898 10732 12310
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10876 11008 10928 11014
rect 10876 10950 10928 10956
rect 10888 10810 10916 10950
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10232 10542 10284 10548
rect 10506 10568 10562 10577
rect 10506 10503 10562 10512
rect 10508 10192 10560 10198
rect 10506 10160 10508 10169
rect 10560 10160 10562 10169
rect 10324 10124 10376 10130
rect 10506 10095 10562 10104
rect 10600 10124 10652 10130
rect 10324 10066 10376 10072
rect 10600 10066 10652 10072
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10060 7262 10180 7290
rect 10060 5794 10088 7262
rect 10244 6474 10272 8910
rect 10336 8566 10364 10066
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 10520 9518 10548 9998
rect 10508 9512 10560 9518
rect 10508 9454 10560 9460
rect 10324 8560 10376 8566
rect 10324 8502 10376 8508
rect 10336 7342 10364 8502
rect 10612 8498 10640 10066
rect 10704 9586 10732 10066
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10784 8900 10836 8906
rect 10784 8842 10836 8848
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 10704 8362 10732 8774
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10324 7336 10376 7342
rect 10324 7278 10376 7284
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10152 6446 10272 6474
rect 10152 6322 10180 6446
rect 10230 6352 10286 6361
rect 10140 6316 10192 6322
rect 10230 6287 10286 6296
rect 10140 6258 10192 6264
rect 10244 6118 10272 6287
rect 10428 6254 10456 7142
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10336 5914 10364 6054
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10060 5766 10456 5794
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 10152 4049 10180 4966
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 9862 4040 9918 4049
rect 9862 3975 9918 3984
rect 10138 4040 10194 4049
rect 10138 3975 10140 3984
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9692 3738 9720 3878
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9772 3528 9824 3534
rect 9770 3496 9772 3505
rect 9824 3496 9826 3505
rect 9770 3431 9826 3440
rect 9876 2961 9904 3975
rect 10192 3975 10194 3984
rect 10140 3946 10192 3952
rect 10244 3670 10272 4558
rect 10232 3664 10284 3670
rect 10232 3606 10284 3612
rect 10244 3194 10272 3606
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10230 3088 10286 3097
rect 10140 3052 10192 3058
rect 10230 3023 10286 3032
rect 10324 3052 10376 3058
rect 10140 2994 10192 3000
rect 9956 2984 10008 2990
rect 9862 2952 9918 2961
rect 9956 2926 10008 2932
rect 9862 2887 9918 2896
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9692 2310 9720 2382
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 9588 2032 9640 2038
rect 9588 1974 9640 1980
rect 9968 480 9996 2926
rect 10152 2650 10180 2994
rect 10244 2854 10272 3023
rect 10324 2994 10376 3000
rect 10232 2848 10284 2854
rect 10232 2790 10284 2796
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 10336 2446 10364 2994
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10428 480 10456 5766
rect 10520 5273 10548 7346
rect 10612 6458 10640 7346
rect 10692 7200 10744 7206
rect 10690 7168 10692 7177
rect 10744 7168 10746 7177
rect 10690 7103 10746 7112
rect 10690 7032 10746 7041
rect 10796 7002 10824 8842
rect 10690 6967 10746 6976
rect 10784 6996 10836 7002
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 10600 6112 10652 6118
rect 10600 6054 10652 6060
rect 10506 5264 10562 5273
rect 10506 5199 10508 5208
rect 10560 5199 10562 5208
rect 10508 5170 10560 5176
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10520 3398 10548 4082
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 10520 3058 10548 3334
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10612 2990 10640 6054
rect 10704 3233 10732 6967
rect 10784 6938 10836 6944
rect 10980 6236 11008 12378
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 11072 11762 11100 12242
rect 11624 12170 11652 12378
rect 11612 12164 11664 12170
rect 11612 12106 11664 12112
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11060 11756 11112 11762
rect 11060 11698 11112 11704
rect 11072 11354 11100 11698
rect 11716 11354 11744 12038
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 11072 10266 11100 11086
rect 11612 11008 11664 11014
rect 11612 10950 11664 10956
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 11164 9568 11192 10406
rect 11256 10198 11284 10610
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11532 10198 11560 10406
rect 11244 10192 11296 10198
rect 11244 10134 11296 10140
rect 11520 10192 11572 10198
rect 11520 10134 11572 10140
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11244 9580 11296 9586
rect 11164 9540 11244 9568
rect 11244 9522 11296 9528
rect 11426 9480 11482 9489
rect 11426 9415 11482 9424
rect 11440 9382 11468 9415
rect 11428 9376 11480 9382
rect 11428 9318 11480 9324
rect 11520 9104 11572 9110
rect 11518 9072 11520 9081
rect 11572 9072 11574 9081
rect 11624 9042 11652 10950
rect 11716 10266 11744 11154
rect 11704 10260 11756 10266
rect 11704 10202 11756 10208
rect 11716 9586 11744 10202
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11518 9007 11574 9016
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11244 8968 11296 8974
rect 11072 8928 11244 8956
rect 11072 8294 11100 8928
rect 11244 8910 11296 8916
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11716 8362 11744 9114
rect 11704 8356 11756 8362
rect 11704 8298 11756 8304
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 11072 7002 11100 8230
rect 11612 7880 11664 7886
rect 11610 7848 11612 7857
rect 11664 7848 11666 7857
rect 11610 7783 11666 7792
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 11428 7472 11480 7478
rect 11428 7414 11480 7420
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 11072 6322 11100 6938
rect 11440 6934 11468 7414
rect 11624 7177 11652 7783
rect 11610 7168 11666 7177
rect 11808 7154 11836 16594
rect 11900 14822 11928 18906
rect 11992 18193 12020 22320
rect 12452 19990 12480 22320
rect 12912 20058 12940 22320
rect 13372 20058 13400 22320
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 13360 20052 13412 20058
rect 13360 19994 13412 20000
rect 12440 19984 12492 19990
rect 12440 19926 12492 19932
rect 12072 19848 12124 19854
rect 12072 19790 12124 19796
rect 12084 19310 12112 19790
rect 12072 19304 12124 19310
rect 12072 19246 12124 19252
rect 12164 19304 12216 19310
rect 12164 19246 12216 19252
rect 12072 18828 12124 18834
rect 12176 18816 12204 19246
rect 12716 19236 12768 19242
rect 12716 19178 12768 19184
rect 13728 19236 13780 19242
rect 13728 19178 13780 19184
rect 12728 18970 12756 19178
rect 12716 18964 12768 18970
rect 12716 18906 12768 18912
rect 12348 18896 12400 18902
rect 12348 18838 12400 18844
rect 12124 18788 12204 18816
rect 12072 18770 12124 18776
rect 11978 18184 12034 18193
rect 11978 18119 12034 18128
rect 11980 17740 12032 17746
rect 11980 17682 12032 17688
rect 11992 17134 12020 17682
rect 12084 17678 12112 18770
rect 12164 17808 12216 17814
rect 12164 17750 12216 17756
rect 12072 17672 12124 17678
rect 12072 17614 12124 17620
rect 11980 17128 12032 17134
rect 11980 17070 12032 17076
rect 11992 15994 12020 17070
rect 12084 16998 12112 17614
rect 12176 17241 12204 17750
rect 12162 17232 12218 17241
rect 12162 17167 12218 17176
rect 12164 17128 12216 17134
rect 12164 17070 12216 17076
rect 12254 17096 12310 17105
rect 12072 16992 12124 16998
rect 12072 16934 12124 16940
rect 12072 16720 12124 16726
rect 12072 16662 12124 16668
rect 12084 16114 12112 16662
rect 12072 16108 12124 16114
rect 12072 16050 12124 16056
rect 11992 15966 12112 15994
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 11992 15706 12020 15846
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 11888 14816 11940 14822
rect 11940 14776 12020 14804
rect 11888 14758 11940 14764
rect 11888 14544 11940 14550
rect 11888 14486 11940 14492
rect 11900 14006 11928 14486
rect 11888 14000 11940 14006
rect 11888 13942 11940 13948
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 11900 12442 11928 12582
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 11992 10554 12020 14776
rect 12084 13002 12112 15966
rect 12176 14958 12204 17070
rect 12254 17031 12256 17040
rect 12308 17031 12310 17040
rect 12256 17002 12308 17008
rect 12256 15496 12308 15502
rect 12254 15464 12256 15473
rect 12308 15464 12310 15473
rect 12254 15399 12310 15408
rect 12164 14952 12216 14958
rect 12164 14894 12216 14900
rect 12176 13870 12204 14894
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 12268 14006 12296 14350
rect 12360 14278 12388 18838
rect 12992 18828 13044 18834
rect 12992 18770 13044 18776
rect 13004 18290 13032 18770
rect 13450 18728 13506 18737
rect 13450 18663 13506 18672
rect 13464 18426 13492 18663
rect 13452 18420 13504 18426
rect 13452 18362 13504 18368
rect 13084 18352 13136 18358
rect 13084 18294 13136 18300
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 12898 18184 12954 18193
rect 12898 18119 12954 18128
rect 12912 18086 12940 18119
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12900 18080 12952 18086
rect 12900 18022 12952 18028
rect 12452 17338 12480 18022
rect 12532 17672 12584 17678
rect 12532 17614 12584 17620
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12544 16658 12572 17614
rect 12808 17128 12860 17134
rect 12808 17070 12860 17076
rect 12820 16998 12848 17070
rect 13096 16998 13124 18294
rect 13176 18216 13228 18222
rect 13176 18158 13228 18164
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 13084 16992 13136 16998
rect 13084 16934 13136 16940
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 12452 15026 12480 16050
rect 12544 15570 12572 16594
rect 12532 15564 12584 15570
rect 12532 15506 12584 15512
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12716 14884 12768 14890
rect 12716 14826 12768 14832
rect 12348 14272 12400 14278
rect 12348 14214 12400 14220
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12256 14000 12308 14006
rect 12256 13942 12308 13948
rect 12164 13864 12216 13870
rect 12164 13806 12216 13812
rect 12348 13864 12400 13870
rect 12348 13806 12400 13812
rect 12256 13320 12308 13326
rect 12256 13262 12308 13268
rect 12084 12986 12204 13002
rect 12084 12980 12216 12986
rect 12084 12974 12164 12980
rect 12164 12922 12216 12928
rect 12070 12880 12126 12889
rect 12070 12815 12126 12824
rect 12084 12646 12112 12815
rect 12072 12640 12124 12646
rect 12072 12582 12124 12588
rect 11900 10526 12020 10554
rect 11900 8294 11928 10526
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11992 9042 12020 10406
rect 12084 9994 12112 12582
rect 12072 9988 12124 9994
rect 12072 9930 12124 9936
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11992 8022 12020 8434
rect 11980 8016 12032 8022
rect 11980 7958 12032 7964
rect 11992 7410 12020 7958
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 11808 7126 12112 7154
rect 11610 7103 11666 7112
rect 11428 6928 11480 6934
rect 11428 6870 11480 6876
rect 11624 6798 11652 7103
rect 11702 6896 11758 6905
rect 11702 6831 11704 6840
rect 11756 6831 11758 6840
rect 11888 6860 11940 6866
rect 11704 6802 11756 6808
rect 11888 6802 11940 6808
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11164 6390 11192 6598
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11152 6384 11204 6390
rect 11152 6326 11204 6332
rect 11336 6384 11388 6390
rect 11336 6326 11388 6332
rect 11060 6316 11112 6322
rect 11060 6258 11112 6264
rect 10888 6208 11008 6236
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 10796 3505 10824 4558
rect 10782 3496 10838 3505
rect 10782 3431 10838 3440
rect 10690 3224 10746 3233
rect 10690 3159 10746 3168
rect 10600 2984 10652 2990
rect 10506 2952 10562 2961
rect 10692 2984 10744 2990
rect 10600 2926 10652 2932
rect 10690 2952 10692 2961
rect 10744 2952 10746 2961
rect 10506 2887 10562 2896
rect 10690 2887 10746 2896
rect 10520 2854 10548 2887
rect 10508 2848 10560 2854
rect 10508 2790 10560 2796
rect 10600 2848 10652 2854
rect 10600 2790 10652 2796
rect 10612 2582 10640 2790
rect 10600 2576 10652 2582
rect 10600 2518 10652 2524
rect 10888 480 10916 6208
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10980 5914 11008 6054
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 11072 5370 11100 5646
rect 11348 5642 11376 6326
rect 11624 5710 11652 6734
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 11336 5636 11388 5642
rect 11336 5578 11388 5584
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11060 5364 11112 5370
rect 11624 5352 11652 5646
rect 11900 5574 11928 6802
rect 11888 5568 11940 5574
rect 11888 5510 11940 5516
rect 11060 5306 11112 5312
rect 11256 5324 11652 5352
rect 11152 5092 11204 5098
rect 11152 5034 11204 5040
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 10980 2650 11008 4218
rect 11072 3942 11100 4966
rect 11164 4826 11192 5034
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 11256 4622 11284 5324
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11518 4856 11574 4865
rect 11808 4826 11836 4966
rect 11518 4791 11574 4800
rect 11796 4820 11848 4826
rect 11532 4758 11560 4791
rect 11796 4762 11848 4768
rect 11520 4752 11572 4758
rect 11572 4712 11652 4740
rect 11520 4694 11572 4700
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 11072 2310 11100 2790
rect 11164 2650 11192 4422
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 11624 4214 11652 4712
rect 11612 4208 11664 4214
rect 12084 4162 12112 7126
rect 11612 4150 11664 4156
rect 11992 4134 12112 4162
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11256 3602 11284 3878
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 11348 3466 11376 3878
rect 11520 3732 11572 3738
rect 11520 3674 11572 3680
rect 11532 3534 11560 3674
rect 11992 3670 12020 4134
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 11612 3664 11664 3670
rect 11612 3606 11664 3612
rect 11980 3664 12032 3670
rect 11980 3606 12032 3612
rect 11520 3528 11572 3534
rect 11518 3496 11520 3505
rect 11572 3496 11574 3505
rect 11336 3460 11388 3466
rect 11518 3431 11574 3440
rect 11336 3402 11388 3408
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11624 2446 11652 3606
rect 11702 3224 11758 3233
rect 11702 3159 11758 3168
rect 11716 2514 11744 3159
rect 11796 3120 11848 3126
rect 11796 3062 11848 3068
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11336 1420 11388 1426
rect 11336 1362 11388 1368
rect 11348 480 11376 1362
rect 11808 480 11836 3062
rect 12084 2582 12112 4014
rect 12072 2576 12124 2582
rect 12072 2518 12124 2524
rect 12176 1426 12204 12922
rect 12268 10169 12296 13262
rect 12360 12918 12388 13806
rect 12452 13530 12480 14010
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12544 13326 12572 14214
rect 12728 14074 12756 14826
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12532 13320 12584 13326
rect 12438 13288 12494 13297
rect 12584 13280 12664 13308
rect 12532 13262 12584 13268
rect 12438 13223 12494 13232
rect 12348 12912 12400 12918
rect 12348 12854 12400 12860
rect 12452 12850 12480 13223
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 12440 12708 12492 12714
rect 12440 12650 12492 12656
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 12452 12220 12480 12650
rect 12532 12232 12584 12238
rect 12452 12192 12532 12220
rect 12360 11898 12388 12174
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 12452 11801 12480 12192
rect 12532 12174 12584 12180
rect 12438 11792 12494 11801
rect 12438 11727 12440 11736
rect 12492 11727 12494 11736
rect 12440 11698 12492 11704
rect 12348 11688 12400 11694
rect 12348 11630 12400 11636
rect 12254 10160 12310 10169
rect 12254 10095 12310 10104
rect 12256 9988 12308 9994
rect 12256 9930 12308 9936
rect 12268 9110 12296 9930
rect 12256 9104 12308 9110
rect 12256 9046 12308 9052
rect 12360 9042 12388 11630
rect 12636 11626 12664 13280
rect 12714 12880 12770 12889
rect 12714 12815 12770 12824
rect 12728 12782 12756 12815
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 12624 11620 12676 11626
rect 12624 11562 12676 11568
rect 12714 11384 12770 11393
rect 12714 11319 12716 11328
rect 12768 11319 12770 11328
rect 12716 11290 12768 11296
rect 12820 11234 12848 16934
rect 12900 16652 12952 16658
rect 12900 16594 12952 16600
rect 12912 15473 12940 16594
rect 12992 15904 13044 15910
rect 12992 15846 13044 15852
rect 13004 15706 13032 15846
rect 12992 15700 13044 15706
rect 12992 15642 13044 15648
rect 12898 15464 12954 15473
rect 12898 15399 12954 15408
rect 12992 14816 13044 14822
rect 12992 14758 13044 14764
rect 12900 14476 12952 14482
rect 12900 14418 12952 14424
rect 12912 11354 12940 14418
rect 13004 14385 13032 14758
rect 12990 14376 13046 14385
rect 12990 14311 13046 14320
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12544 11206 12848 11234
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 12360 7562 12388 8978
rect 12268 7534 12388 7562
rect 12268 7041 12296 7534
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12254 7032 12310 7041
rect 12360 7002 12388 7346
rect 12254 6967 12310 6976
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12256 6316 12308 6322
rect 12256 6258 12308 6264
rect 12268 5778 12296 6258
rect 12256 5772 12308 5778
rect 12256 5714 12308 5720
rect 12348 4072 12400 4078
rect 12348 4014 12400 4020
rect 12360 3738 12388 4014
rect 12348 3732 12400 3738
rect 12348 3674 12400 3680
rect 12452 3210 12480 11154
rect 12544 10554 12572 11206
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 12544 10526 12664 10554
rect 12532 10192 12584 10198
rect 12532 10134 12584 10140
rect 12544 9081 12572 10134
rect 12636 10130 12664 10526
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 12530 9072 12586 9081
rect 12636 9058 12664 10066
rect 12728 9217 12756 11018
rect 13004 10810 13032 13330
rect 12992 10804 13044 10810
rect 12992 10746 13044 10752
rect 13096 10742 13124 16934
rect 13188 11218 13216 18158
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 13556 13870 13584 18022
rect 13634 15464 13690 15473
rect 13634 15399 13636 15408
rect 13688 15399 13690 15408
rect 13636 15370 13688 15376
rect 13740 15314 13768 19178
rect 13832 17338 13860 22320
rect 13912 19916 13964 19922
rect 13912 19858 13964 19864
rect 14188 19916 14240 19922
rect 14188 19858 14240 19864
rect 13924 18902 13952 19858
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 13912 18896 13964 18902
rect 13912 18838 13964 18844
rect 13912 18284 13964 18290
rect 13912 18226 13964 18232
rect 13924 17882 13952 18226
rect 14004 18080 14056 18086
rect 14004 18022 14056 18028
rect 13912 17876 13964 17882
rect 13912 17818 13964 17824
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 13818 17096 13874 17105
rect 13818 17031 13874 17040
rect 13832 16114 13860 17031
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 14016 15722 14044 18022
rect 13648 15286 13768 15314
rect 13924 15694 14044 15722
rect 13544 13864 13596 13870
rect 13544 13806 13596 13812
rect 13544 13184 13596 13190
rect 13544 13126 13596 13132
rect 13360 11620 13412 11626
rect 13360 11562 13412 11568
rect 13176 11212 13228 11218
rect 13176 11154 13228 11160
rect 12808 10736 12860 10742
rect 12808 10678 12860 10684
rect 13084 10736 13136 10742
rect 13084 10678 13136 10684
rect 12714 9208 12770 9217
rect 12714 9143 12770 9152
rect 12636 9030 12756 9058
rect 12530 9007 12586 9016
rect 12622 8936 12678 8945
rect 12622 8871 12678 8880
rect 12532 8288 12584 8294
rect 12532 8230 12584 8236
rect 12544 7478 12572 8230
rect 12532 7472 12584 7478
rect 12532 7414 12584 7420
rect 12636 6186 12664 8871
rect 12728 7018 12756 9030
rect 12820 7206 12848 10678
rect 13372 10674 13400 11562
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 12912 10266 12940 10406
rect 12900 10260 12952 10266
rect 12900 10202 12952 10208
rect 12912 9625 12940 10202
rect 12898 9616 12954 9625
rect 13004 9586 13032 10610
rect 13452 10600 13504 10606
rect 13174 10568 13230 10577
rect 13452 10542 13504 10548
rect 13174 10503 13230 10512
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 13096 9586 13124 9862
rect 12898 9551 12954 9560
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 13188 9518 13216 10503
rect 13266 10160 13322 10169
rect 13266 10095 13322 10104
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 12808 7200 12860 7206
rect 12860 7148 13032 7154
rect 12808 7142 13032 7148
rect 12820 7126 13032 7142
rect 12728 6990 12848 7018
rect 12716 6384 12768 6390
rect 12716 6326 12768 6332
rect 12532 6180 12584 6186
rect 12532 6122 12584 6128
rect 12624 6180 12676 6186
rect 12624 6122 12676 6128
rect 12544 5370 12572 6122
rect 12728 6118 12756 6326
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 12820 5930 12848 6990
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 12728 5902 12848 5930
rect 12624 5772 12676 5778
rect 12624 5714 12676 5720
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 12636 5234 12664 5714
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12636 4554 12664 5170
rect 12624 4548 12676 4554
rect 12624 4490 12676 4496
rect 12532 4004 12584 4010
rect 12532 3946 12584 3952
rect 12544 3534 12572 3946
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 12268 3182 12480 3210
rect 12164 1420 12216 1426
rect 12164 1362 12216 1368
rect 12268 480 12296 3182
rect 12728 3126 12756 5902
rect 12912 5302 12940 6734
rect 12900 5296 12952 5302
rect 12900 5238 12952 5244
rect 12900 4004 12952 4010
rect 12900 3946 12952 3952
rect 12912 3738 12940 3946
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 12716 3120 12768 3126
rect 12716 3062 12768 3068
rect 12714 2952 12770 2961
rect 12820 2922 12848 3538
rect 12714 2887 12770 2896
rect 12808 2916 12860 2922
rect 12728 480 12756 2887
rect 12808 2858 12860 2864
rect 13004 2514 13032 7126
rect 13096 6798 13124 8978
rect 13280 8906 13308 10095
rect 13268 8900 13320 8906
rect 13268 8842 13320 8848
rect 13280 8498 13308 8842
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 13174 7984 13230 7993
rect 13174 7919 13230 7928
rect 13188 7206 13216 7919
rect 13360 7880 13412 7886
rect 13358 7848 13360 7857
rect 13412 7848 13414 7857
rect 13280 7806 13358 7834
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13084 6792 13136 6798
rect 13188 6769 13216 7142
rect 13084 6734 13136 6740
rect 13174 6760 13230 6769
rect 13174 6695 13230 6704
rect 13280 6322 13308 7806
rect 13358 7783 13414 7792
rect 13360 7472 13412 7478
rect 13360 7414 13412 7420
rect 13372 6934 13400 7414
rect 13360 6928 13412 6934
rect 13360 6870 13412 6876
rect 13464 6338 13492 10542
rect 13556 9042 13584 13126
rect 13648 11898 13676 15286
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13740 14278 13768 15098
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13832 14482 13860 14962
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13740 13394 13768 14214
rect 13832 14074 13860 14418
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13820 13796 13872 13802
rect 13820 13738 13872 13744
rect 13832 13530 13860 13738
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 13924 12753 13952 15694
rect 14004 15632 14056 15638
rect 14004 15574 14056 15580
rect 14016 15162 14044 15574
rect 14004 15156 14056 15162
rect 14004 15098 14056 15104
rect 14108 15065 14136 19246
rect 14200 18902 14228 19858
rect 14292 19174 14320 22320
rect 14752 20754 14780 22320
rect 14568 20726 14780 20754
rect 14568 20058 14596 20726
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 15212 20058 15240 22320
rect 15672 20058 15700 22320
rect 14556 20052 14608 20058
rect 14556 19994 14608 20000
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 15660 20052 15712 20058
rect 15660 19994 15712 20000
rect 14464 19916 14516 19922
rect 14464 19858 14516 19864
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 15568 19916 15620 19922
rect 15568 19858 15620 19864
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 14188 18896 14240 18902
rect 14188 18838 14240 18844
rect 14188 16176 14240 16182
rect 14188 16118 14240 16124
rect 14200 15570 14228 16118
rect 14188 15564 14240 15570
rect 14188 15506 14240 15512
rect 14200 15162 14228 15506
rect 14476 15416 14504 19858
rect 15108 19168 15160 19174
rect 15108 19110 15160 19116
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 14556 17060 14608 17066
rect 14556 17002 14608 17008
rect 14568 16726 14596 17002
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 14556 16720 14608 16726
rect 14556 16662 14608 16668
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 15014 15600 15070 15609
rect 15014 15535 15070 15544
rect 14476 15388 14596 15416
rect 14188 15156 14240 15162
rect 14188 15098 14240 15104
rect 14094 15056 14150 15065
rect 14094 14991 14150 15000
rect 14200 14618 14228 15098
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 13910 12744 13966 12753
rect 13820 12708 13872 12714
rect 13910 12679 13966 12688
rect 13820 12650 13872 12656
rect 13832 12442 13860 12650
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13832 11898 13860 12378
rect 13636 11892 13688 11898
rect 13636 11834 13688 11840
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13832 11762 13860 11834
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 13634 11384 13690 11393
rect 13634 11319 13690 11328
rect 13648 11150 13676 11319
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 13636 11144 13688 11150
rect 13636 11086 13688 11092
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13648 9110 13676 9318
rect 13636 9104 13688 9110
rect 13636 9046 13688 9052
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13636 8016 13688 8022
rect 13636 7958 13688 7964
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13556 7290 13584 7686
rect 13648 7410 13676 7958
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13556 7262 13676 7290
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 13268 6316 13320 6322
rect 13464 6310 13584 6338
rect 13268 6258 13320 6264
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 13096 2922 13124 5850
rect 13188 5234 13216 6258
rect 13452 6248 13504 6254
rect 13452 6190 13504 6196
rect 13464 5778 13492 6190
rect 13452 5772 13504 5778
rect 13452 5714 13504 5720
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 13188 4865 13216 5170
rect 13280 5166 13308 5646
rect 13556 5370 13584 6310
rect 13648 5930 13676 7262
rect 13740 6118 13768 9998
rect 13832 9450 13860 11154
rect 13820 9444 13872 9450
rect 13820 9386 13872 9392
rect 13818 9344 13874 9353
rect 13818 9279 13874 9288
rect 13832 9110 13860 9279
rect 13820 9104 13872 9110
rect 13820 9046 13872 9052
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 13832 7274 13860 8502
rect 13924 8430 13952 11494
rect 14016 11150 14044 14554
rect 14188 13864 14240 13870
rect 14188 13806 14240 13812
rect 14096 11688 14148 11694
rect 14096 11630 14148 11636
rect 14108 11354 14136 11630
rect 14096 11348 14148 11354
rect 14096 11290 14148 11296
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 14016 10062 14044 10610
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 14108 8430 14136 9318
rect 13912 8424 13964 8430
rect 14096 8424 14148 8430
rect 13964 8372 14044 8378
rect 13912 8366 14044 8372
rect 14096 8366 14148 8372
rect 13924 8350 14044 8366
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 13924 7206 13952 8230
rect 14016 7834 14044 8350
rect 14016 7806 14136 7834
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 13912 7200 13964 7206
rect 13912 7142 13964 7148
rect 13924 7002 13952 7142
rect 13912 6996 13964 7002
rect 13912 6938 13964 6944
rect 13818 6896 13874 6905
rect 13818 6831 13874 6840
rect 13832 6798 13860 6831
rect 13820 6792 13872 6798
rect 13820 6734 13872 6740
rect 14016 6186 14044 7686
rect 14108 7410 14136 7806
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 14094 6352 14150 6361
rect 14094 6287 14150 6296
rect 14004 6180 14056 6186
rect 14004 6122 14056 6128
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13910 5944 13966 5953
rect 13648 5902 13768 5930
rect 13544 5364 13596 5370
rect 13544 5306 13596 5312
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 13268 5160 13320 5166
rect 13268 5102 13320 5108
rect 13544 5160 13596 5166
rect 13544 5102 13596 5108
rect 13174 4856 13230 4865
rect 13174 4791 13230 4800
rect 13268 4684 13320 4690
rect 13188 4644 13268 4672
rect 13188 4282 13216 4644
rect 13268 4626 13320 4632
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13176 4276 13228 4282
rect 13176 4218 13228 4224
rect 13176 4072 13228 4078
rect 13174 4040 13176 4049
rect 13228 4040 13230 4049
rect 13174 3975 13230 3984
rect 13372 3738 13400 4558
rect 13360 3732 13412 3738
rect 13360 3674 13412 3680
rect 13176 3528 13228 3534
rect 13176 3470 13228 3476
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13084 2916 13136 2922
rect 13084 2858 13136 2864
rect 12992 2508 13044 2514
rect 12992 2450 13044 2456
rect 13188 480 13216 3470
rect 13372 2106 13400 3470
rect 13556 2582 13584 5102
rect 13648 4622 13676 5170
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 13648 3942 13676 4558
rect 13740 4214 13768 5902
rect 13910 5879 13966 5888
rect 13728 4208 13780 4214
rect 13728 4150 13780 4156
rect 13924 4146 13952 5879
rect 14016 5273 14044 6122
rect 14002 5264 14058 5273
rect 14002 5199 14004 5208
rect 14056 5199 14058 5208
rect 14004 5170 14056 5176
rect 14016 5139 14044 5170
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 13544 2576 13596 2582
rect 13544 2518 13596 2524
rect 13360 2100 13412 2106
rect 13360 2042 13412 2048
rect 13648 480 13676 3674
rect 13728 3664 13780 3670
rect 13728 3606 13780 3612
rect 13740 2990 13768 3606
rect 13912 3392 13964 3398
rect 13912 3334 13964 3340
rect 13818 3088 13874 3097
rect 13818 3023 13874 3032
rect 13832 2990 13860 3023
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 13924 2514 13952 3334
rect 13912 2508 13964 2514
rect 13912 2450 13964 2456
rect 14016 626 14044 4966
rect 14108 4706 14136 6287
rect 14200 5166 14228 13806
rect 14280 13388 14332 13394
rect 14280 13330 14332 13336
rect 14292 12986 14320 13330
rect 14280 12980 14332 12986
rect 14280 12922 14332 12928
rect 14280 12640 14332 12646
rect 14280 12582 14332 12588
rect 14292 12374 14320 12582
rect 14280 12368 14332 12374
rect 14280 12310 14332 12316
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14292 10810 14320 11494
rect 14280 10804 14332 10810
rect 14280 10746 14332 10752
rect 14280 9444 14332 9450
rect 14280 9386 14332 9392
rect 14292 8974 14320 9386
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14292 8537 14320 8910
rect 14278 8528 14334 8537
rect 14278 8463 14334 8472
rect 14384 7585 14412 14894
rect 14568 12306 14596 15388
rect 15028 15162 15056 15535
rect 15016 15156 15068 15162
rect 15016 15098 15068 15104
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 15120 13394 15148 19110
rect 15200 18828 15252 18834
rect 15200 18770 15252 18776
rect 14832 13388 14884 13394
rect 14832 13330 14884 13336
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 14648 13320 14700 13326
rect 14648 13262 14700 13268
rect 14660 12782 14688 13262
rect 14648 12776 14700 12782
rect 14648 12718 14700 12724
rect 14844 12628 14872 13330
rect 15016 13252 15068 13258
rect 15016 13194 15068 13200
rect 14924 13184 14976 13190
rect 14924 13126 14976 13132
rect 14936 12782 14964 13126
rect 15028 12782 15056 13194
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 14924 12776 14976 12782
rect 14924 12718 14976 12724
rect 15016 12776 15068 12782
rect 15016 12718 15068 12724
rect 14844 12600 15056 12628
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 14556 12300 14608 12306
rect 14556 12242 14608 12248
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14476 10130 14504 12038
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 14646 11248 14702 11257
rect 14646 11183 14702 11192
rect 14660 11150 14688 11183
rect 14648 11144 14700 11150
rect 14648 11086 14700 11092
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 14464 10124 14516 10130
rect 14464 10066 14516 10072
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 14568 8634 14596 9318
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 14924 8832 14976 8838
rect 14924 8774 14976 8780
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14936 8498 14964 8774
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 14370 7576 14426 7585
rect 14370 7511 14426 7520
rect 14372 7472 14424 7478
rect 14372 7414 14424 7420
rect 14280 7268 14332 7274
rect 14280 7210 14332 7216
rect 14292 6798 14320 7210
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14200 4826 14228 4966
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 14108 4678 14228 4706
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 14108 3126 14136 3878
rect 14096 3120 14148 3126
rect 14096 3062 14148 3068
rect 14200 2514 14228 4678
rect 14292 3194 14320 6734
rect 14384 3602 14412 7414
rect 15028 7313 15056 12600
rect 15120 12442 15148 12786
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 15120 10266 15148 11494
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 15212 9489 15240 18770
rect 15384 14816 15436 14822
rect 15384 14758 15436 14764
rect 15396 13841 15424 14758
rect 15488 14618 15516 19858
rect 15580 18902 15608 19858
rect 16132 19174 16160 22320
rect 16592 20058 16620 22320
rect 17052 20074 17080 22320
rect 16580 20052 16632 20058
rect 16580 19994 16632 20000
rect 16960 20046 17080 20074
rect 16580 19304 16632 19310
rect 16580 19246 16632 19252
rect 16120 19168 16172 19174
rect 16120 19110 16172 19116
rect 15568 18896 15620 18902
rect 15568 18838 15620 18844
rect 15568 18760 15620 18766
rect 15568 18702 15620 18708
rect 15476 14612 15528 14618
rect 15476 14554 15528 14560
rect 15382 13832 15438 13841
rect 15382 13767 15438 13776
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15198 9480 15254 9489
rect 15198 9415 15254 9424
rect 15108 9104 15160 9110
rect 15108 9046 15160 9052
rect 15014 7304 15070 7313
rect 15014 7239 15070 7248
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 14476 7002 14504 7142
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 14556 6792 14608 6798
rect 14556 6734 14608 6740
rect 14568 5914 14596 6734
rect 15016 6112 15068 6118
rect 15016 6054 15068 6060
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 14556 5908 14608 5914
rect 14556 5850 14608 5856
rect 15028 5710 15056 6054
rect 15016 5704 15068 5710
rect 15016 5646 15068 5652
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 14372 3596 14424 3602
rect 14372 3538 14424 3544
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14476 2922 14504 5102
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 15028 4622 15056 5646
rect 15120 5166 15148 9046
rect 15304 8906 15332 13330
rect 15580 12986 15608 18702
rect 15844 15020 15896 15026
rect 15844 14962 15896 14968
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 15568 12980 15620 12986
rect 15568 12922 15620 12928
rect 15292 8900 15344 8906
rect 15292 8842 15344 8848
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15200 6248 15252 6254
rect 15200 6190 15252 6196
rect 15212 5778 15240 6190
rect 15200 5772 15252 5778
rect 15200 5714 15252 5720
rect 15108 5160 15160 5166
rect 15108 5102 15160 5108
rect 15108 5024 15160 5030
rect 15108 4966 15160 4972
rect 15120 4758 15148 4966
rect 15304 4826 15332 6598
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15580 5846 15608 6054
rect 15568 5840 15620 5846
rect 15568 5782 15620 5788
rect 15384 5772 15436 5778
rect 15384 5714 15436 5720
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 15108 4752 15160 4758
rect 15108 4694 15160 4700
rect 15016 4616 15068 4622
rect 15016 4558 15068 4564
rect 15108 4480 15160 4486
rect 15108 4422 15160 4428
rect 14568 4010 14688 4026
rect 14568 4004 14700 4010
rect 14568 3998 14648 4004
rect 14464 2916 14516 2922
rect 14464 2858 14516 2864
rect 14188 2508 14240 2514
rect 14188 2450 14240 2456
rect 14016 598 14136 626
rect 14108 480 14136 598
rect 14568 480 14596 3998
rect 14648 3946 14700 3952
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 15016 3392 15068 3398
rect 15016 3334 15068 3340
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 15028 480 15056 3334
rect 15120 2650 15148 4422
rect 15396 3720 15424 5714
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 15488 5098 15516 5510
rect 15580 5234 15608 5782
rect 15568 5228 15620 5234
rect 15568 5170 15620 5176
rect 15476 5092 15528 5098
rect 15476 5034 15528 5040
rect 15304 3692 15424 3720
rect 15304 2854 15332 3692
rect 15672 3641 15700 14554
rect 15856 14414 15884 14962
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 15750 13424 15806 13433
rect 15750 13359 15752 13368
rect 15804 13359 15806 13368
rect 15752 13330 15804 13336
rect 15856 13326 15884 14350
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 15856 13190 15884 13262
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15856 12889 15884 13126
rect 15842 12880 15898 12889
rect 15842 12815 15898 12824
rect 15936 12640 15988 12646
rect 15936 12582 15988 12588
rect 15948 11898 15976 12582
rect 15936 11892 15988 11898
rect 15936 11834 15988 11840
rect 16592 10470 16620 19246
rect 16960 19174 16988 20046
rect 17040 19916 17092 19922
rect 17040 19858 17092 19864
rect 16948 19168 17000 19174
rect 16948 19110 17000 19116
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16776 11014 16804 13262
rect 17052 11626 17080 19858
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 17224 19304 17276 19310
rect 17224 19246 17276 19252
rect 17040 11620 17092 11626
rect 17040 11562 17092 11568
rect 17144 11082 17172 19246
rect 17236 11762 17264 19246
rect 17512 19174 17540 22320
rect 17972 20058 18000 22320
rect 17960 20052 18012 20058
rect 17960 19994 18012 20000
rect 18432 19802 18460 22320
rect 18432 19774 18552 19802
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 18524 19174 18552 19774
rect 18604 19304 18656 19310
rect 18604 19246 18656 19252
rect 18788 19304 18840 19310
rect 18788 19246 18840 19252
rect 17500 19168 17552 19174
rect 17500 19110 17552 19116
rect 18512 19168 18564 19174
rect 18512 19110 18564 19116
rect 18512 18828 18564 18834
rect 18512 18770 18564 18776
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 17224 11756 17276 11762
rect 17224 11698 17276 11704
rect 17132 11076 17184 11082
rect 17132 11018 17184 11024
rect 16764 11008 16816 11014
rect 16764 10950 16816 10956
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 18524 8566 18552 18770
rect 18616 14890 18644 19246
rect 18800 18902 18828 19246
rect 18892 19174 18920 22320
rect 18880 19168 18932 19174
rect 18880 19110 18932 19116
rect 19352 19122 19380 22320
rect 19812 19786 19840 22320
rect 19800 19780 19852 19786
rect 19800 19722 19852 19728
rect 20272 19174 20300 22320
rect 20260 19168 20312 19174
rect 19352 19094 19472 19122
rect 20260 19110 20312 19116
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 18788 18896 18840 18902
rect 18788 18838 18840 18844
rect 19352 17338 19380 18906
rect 19340 17332 19392 17338
rect 19340 17274 19392 17280
rect 19444 16658 19472 19094
rect 19524 18080 19576 18086
rect 20732 18034 20760 22320
rect 21192 18970 21220 22320
rect 21180 18964 21232 18970
rect 21180 18906 21232 18912
rect 21652 18426 21680 22320
rect 22112 19242 22140 22320
rect 22100 19236 22152 19242
rect 22100 19178 22152 19184
rect 21640 18420 21692 18426
rect 21640 18362 21692 18368
rect 22572 18086 22600 22320
rect 19524 18022 19576 18028
rect 19432 16652 19484 16658
rect 19432 16594 19484 16600
rect 18604 14884 18656 14890
rect 18604 14826 18656 14832
rect 19536 14618 19564 18022
rect 20640 18006 20760 18034
rect 22560 18080 22612 18086
rect 22560 18022 22612 18028
rect 20640 17882 20668 18006
rect 20628 17876 20680 17882
rect 20628 17818 20680 17824
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 18696 13864 18748 13870
rect 18696 13806 18748 13812
rect 18512 8560 18564 8566
rect 18512 8502 18564 8508
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 16578 6760 16634 6769
rect 16578 6695 16634 6704
rect 15658 3632 15714 3641
rect 15658 3567 15714 3576
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 16040 3233 16068 3538
rect 16120 3528 16172 3534
rect 16120 3470 16172 3476
rect 16026 3224 16082 3233
rect 16026 3159 16082 3168
rect 16028 3120 16080 3126
rect 16028 3062 16080 3068
rect 15292 2848 15344 2854
rect 15292 2790 15344 2796
rect 15108 2644 15160 2650
rect 15108 2586 15160 2592
rect 15660 2508 15712 2514
rect 15660 2450 15712 2456
rect 15568 2304 15620 2310
rect 15568 2246 15620 2252
rect 15580 480 15608 2246
rect 15672 2106 15700 2450
rect 15660 2100 15712 2106
rect 15660 2042 15712 2048
rect 16040 480 16068 3062
rect 16132 2990 16160 3470
rect 16120 2984 16172 2990
rect 16120 2926 16172 2932
rect 16592 2514 16620 6695
rect 17038 6216 17094 6225
rect 17038 6151 17094 6160
rect 16948 5568 17000 5574
rect 16948 5510 17000 5516
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 16868 2990 16896 5102
rect 16960 4826 16988 5510
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 16856 2984 16908 2990
rect 16856 2926 16908 2932
rect 16948 2848 17000 2854
rect 16948 2790 17000 2796
rect 16580 2508 16632 2514
rect 16580 2450 16632 2456
rect 16488 2304 16540 2310
rect 16488 2246 16540 2252
rect 16500 480 16528 2246
rect 16960 480 16988 2790
rect 17052 2514 17080 6151
rect 17420 5914 17448 7890
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 18512 6928 18564 6934
rect 18512 6870 18564 6876
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17512 5710 17540 6734
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 17958 5808 18014 5817
rect 17958 5743 17960 5752
rect 18012 5743 18014 5752
rect 17960 5714 18012 5720
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 17868 5092 17920 5098
rect 17868 5034 17920 5040
rect 17880 4690 17908 5034
rect 17868 4684 17920 4690
rect 17868 4626 17920 4632
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 18524 2990 18552 6870
rect 18708 5817 18736 13806
rect 19156 6452 19208 6458
rect 19156 6394 19208 6400
rect 18694 5808 18750 5817
rect 18694 5743 18750 5752
rect 18788 4480 18840 4486
rect 18788 4422 18840 4428
rect 18512 2984 18564 2990
rect 18512 2926 18564 2932
rect 17868 2848 17920 2854
rect 17868 2790 17920 2796
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 17420 480 17448 2246
rect 17880 480 17908 2790
rect 17960 2304 18012 2310
rect 17960 2246 18012 2252
rect 17972 1170 18000 2246
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 17972 1142 18368 1170
rect 18340 480 18368 1142
rect 18800 480 18828 4422
rect 19168 2990 19196 6394
rect 19800 5704 19852 5710
rect 19800 5646 19852 5652
rect 19812 5166 19840 5646
rect 19800 5160 19852 5166
rect 19800 5102 19852 5108
rect 20628 5024 20680 5030
rect 20628 4966 20680 4972
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 19352 4146 19380 4558
rect 19340 4140 19392 4146
rect 19340 4082 19392 4088
rect 20168 3188 20220 3194
rect 20168 3130 20220 3136
rect 19156 2984 19208 2990
rect 19156 2926 19208 2932
rect 19248 2848 19300 2854
rect 19248 2790 19300 2796
rect 19708 2848 19760 2854
rect 19708 2790 19760 2796
rect 19260 480 19288 2790
rect 19720 480 19748 2790
rect 20180 480 20208 3130
rect 20640 480 20668 4966
rect 22468 4140 22520 4146
rect 22468 4082 22520 4088
rect 22008 2916 22060 2922
rect 22008 2858 22060 2864
rect 21548 2576 21600 2582
rect 21548 2518 21600 2524
rect 21088 2372 21140 2378
rect 21088 2314 21140 2320
rect 21100 480 21128 2314
rect 21560 480 21588 2518
rect 22020 480 22048 2858
rect 22480 480 22508 4082
rect 2870 232 2926 241
rect 2870 167 2926 176
rect 2962 0 3018 480
rect 3422 0 3478 480
rect 3882 0 3938 480
rect 4342 0 4398 480
rect 4802 0 4858 480
rect 5262 0 5318 480
rect 5722 0 5778 480
rect 6182 0 6238 480
rect 6642 0 6698 480
rect 7102 0 7158 480
rect 7562 0 7618 480
rect 8114 0 8170 480
rect 8574 0 8630 480
rect 9034 0 9090 480
rect 9494 0 9550 480
rect 9954 0 10010 480
rect 10414 0 10470 480
rect 10874 0 10930 480
rect 11334 0 11390 480
rect 11794 0 11850 480
rect 12254 0 12310 480
rect 12714 0 12770 480
rect 13174 0 13230 480
rect 13634 0 13690 480
rect 14094 0 14150 480
rect 14554 0 14610 480
rect 15014 0 15070 480
rect 15566 0 15622 480
rect 16026 0 16082 480
rect 16486 0 16542 480
rect 16946 0 17002 480
rect 17406 0 17462 480
rect 17866 0 17922 480
rect 18326 0 18382 480
rect 18786 0 18842 480
rect 19246 0 19302 480
rect 19706 0 19762 480
rect 20166 0 20222 480
rect 20626 0 20682 480
rect 21086 0 21142 480
rect 21546 0 21602 480
rect 22006 0 22062 480
rect 22466 0 22522 480
<< via2 >>
rect 2778 22480 2834 22536
rect 1858 19660 1860 19680
rect 1860 19660 1912 19680
rect 1912 19660 1914 19680
rect 1858 19624 1914 19660
rect 1766 19216 1822 19272
rect 1582 18692 1638 18728
rect 1582 18672 1584 18692
rect 1584 18672 1636 18692
rect 1636 18672 1638 18692
rect 1674 18300 1676 18320
rect 1676 18300 1728 18320
rect 1728 18300 1730 18320
rect 1674 18264 1730 18300
rect 1766 17332 1822 17368
rect 1766 17312 1768 17332
rect 1768 17312 1820 17332
rect 1820 17312 1822 17332
rect 2134 18128 2190 18184
rect 1950 17040 2006 17096
rect 1858 16788 1914 16824
rect 1858 16768 1860 16788
rect 1860 16768 1912 16788
rect 1912 16768 1914 16788
rect 1950 16360 2006 16416
rect 1766 15988 1768 16008
rect 1768 15988 1820 16008
rect 1820 15988 1822 16008
rect 1766 15952 1822 15988
rect 1582 15816 1638 15872
rect 3146 21528 3202 21584
rect 2594 18536 2650 18592
rect 2778 17720 2834 17776
rect 2870 15816 2926 15872
rect 3698 22072 3754 22128
rect 3606 21120 3662 21176
rect 3698 20576 3754 20632
rect 3146 18264 3202 18320
rect 3146 17584 3202 17640
rect 2410 15564 2466 15600
rect 2410 15544 2412 15564
rect 2412 15544 2464 15564
rect 2464 15544 2466 15564
rect 1674 14864 1730 14920
rect 2594 15272 2650 15328
rect 2502 14592 2558 14648
rect 2962 13912 3018 13968
rect 1398 10648 1454 10704
rect 3514 18536 3570 18592
rect 3422 17720 3478 17776
rect 3422 16632 3478 16688
rect 4066 20168 4122 20224
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 4526 19080 4582 19136
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4894 18148 4950 18184
rect 4894 18128 4896 18148
rect 4896 18128 4948 18148
rect 4948 18128 4950 18148
rect 4066 17740 4122 17776
rect 4066 17720 4068 17740
rect 4068 17720 4120 17740
rect 4120 17720 4122 17740
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 2502 7268 2558 7304
rect 2502 7248 2504 7268
rect 2504 7248 2556 7268
rect 2556 7248 2558 7268
rect 2962 9424 3018 9480
rect 3422 15408 3478 15464
rect 3330 14456 3386 14512
rect 3790 15680 3846 15736
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 4066 15680 4122 15736
rect 3974 14864 4030 14920
rect 4066 13504 4122 13560
rect 3514 12144 3570 12200
rect 3606 12008 3662 12064
rect 1950 2760 2006 2816
rect 2962 5752 3018 5808
rect 2778 3984 2834 4040
rect 2594 3032 2650 3088
rect 2686 2644 2742 2680
rect 2686 2624 2688 2644
rect 2688 2624 2740 2644
rect 2740 2624 2742 2644
rect 2686 2080 2742 2136
rect 2778 1128 2834 1184
rect 3422 8880 3478 8936
rect 3606 6840 3662 6896
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 4618 15000 4674 15056
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 3974 12552 4030 12608
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 5078 17720 5134 17776
rect 5538 18264 5594 18320
rect 5354 17720 5410 17776
rect 4894 12552 4950 12608
rect 5446 15000 5502 15056
rect 4434 12316 4436 12336
rect 4436 12316 4488 12336
rect 4488 12316 4490 12336
rect 4434 12280 4490 12316
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4158 11600 4214 11656
rect 3974 10104 4030 10160
rect 4066 9696 4122 9752
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 3974 8744 4030 8800
rect 4066 8200 4122 8256
rect 4066 7792 4122 7848
rect 4066 4392 4122 4448
rect 3790 3576 3846 3632
rect 3698 3440 3754 3496
rect 3422 3052 3478 3088
rect 3422 3032 3424 3052
rect 3424 3032 3476 3052
rect 3476 3032 3478 3052
rect 3146 2796 3148 2816
rect 3148 2796 3200 2816
rect 3200 2796 3202 2816
rect 3146 2760 3202 2796
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 5446 14068 5502 14104
rect 5446 14048 5448 14068
rect 5448 14048 5500 14068
rect 5500 14048 5502 14068
rect 4986 9424 5042 9480
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 5998 16768 6054 16824
rect 5998 14592 6054 14648
rect 5998 13776 6054 13832
rect 4802 4936 4858 4992
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4618 3848 4674 3904
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 4342 3052 4398 3088
rect 3514 584 3570 640
rect 4342 3032 4344 3052
rect 4344 3032 4396 3052
rect 4396 3032 4398 3052
rect 4066 2524 4068 2544
rect 4068 2524 4120 2544
rect 4120 2524 4122 2544
rect 4066 2488 4122 2524
rect 4066 1536 4122 1592
rect 4986 3848 5042 3904
rect 4894 3612 4896 3632
rect 4896 3612 4948 3632
rect 4948 3612 4950 3632
rect 4894 3576 4950 3612
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 5354 3984 5410 4040
rect 5998 9424 6054 9480
rect 6182 16088 6238 16144
rect 6182 15852 6184 15872
rect 6184 15852 6236 15872
rect 6236 15852 6238 15872
rect 6182 15816 6238 15852
rect 6182 14456 6238 14512
rect 6182 12588 6184 12608
rect 6184 12588 6236 12608
rect 6236 12588 6238 12608
rect 6182 12552 6238 12588
rect 6458 17040 6514 17096
rect 6642 19116 6644 19136
rect 6644 19116 6696 19136
rect 6696 19116 6698 19136
rect 6642 19080 6698 19116
rect 6366 16632 6422 16688
rect 6550 16768 6606 16824
rect 6458 16088 6514 16144
rect 6458 15000 6514 15056
rect 5722 4276 5778 4312
rect 5722 4256 5724 4276
rect 5724 4256 5776 4276
rect 5776 4256 5778 4276
rect 6826 16124 6828 16144
rect 6828 16124 6880 16144
rect 6880 16124 6882 16144
rect 6826 16088 6882 16124
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 7102 14884 7158 14920
rect 7102 14864 7104 14884
rect 7104 14864 7156 14884
rect 7156 14864 7158 14884
rect 6918 12552 6974 12608
rect 6734 9424 6790 9480
rect 5998 4120 6054 4176
rect 6182 3576 6238 3632
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 8298 15952 8354 16008
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 8022 15408 8078 15464
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 7470 9172 7526 9208
rect 7470 9152 7472 9172
rect 7472 9152 7524 9172
rect 7524 9152 7526 9172
rect 7470 8880 7526 8936
rect 6918 6196 6920 6216
rect 6920 6196 6972 6216
rect 6972 6196 6974 6216
rect 6918 6160 6974 6196
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 8758 13776 8814 13832
rect 8758 12144 8814 12200
rect 8758 11328 8814 11384
rect 8482 11056 8538 11112
rect 8574 10548 8576 10568
rect 8576 10548 8628 10568
rect 8628 10548 8630 10568
rect 8574 10512 8630 10548
rect 8942 15000 8998 15056
rect 9034 14864 9090 14920
rect 8942 14320 8998 14376
rect 8298 9152 8354 9208
rect 7930 8744 7986 8800
rect 8114 8608 8170 8664
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 8206 7384 8262 7440
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 8206 5616 8262 5672
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 7562 2896 7618 2952
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 8390 9052 8392 9072
rect 8392 9052 8444 9072
rect 8444 9052 8446 9072
rect 8390 9016 8446 9052
rect 8666 8200 8722 8256
rect 8390 7948 8446 7984
rect 8390 7928 8392 7948
rect 8392 7928 8444 7948
rect 8444 7928 8446 7948
rect 8666 6296 8722 6352
rect 10138 18808 10194 18864
rect 9218 14048 9274 14104
rect 9034 12280 9090 12336
rect 9126 11736 9182 11792
rect 9310 11736 9366 11792
rect 10138 17740 10194 17776
rect 10138 17720 10140 17740
rect 10140 17720 10192 17740
rect 10192 17720 10194 17740
rect 10690 18808 10746 18864
rect 9954 16496 10010 16552
rect 9862 14048 9918 14104
rect 9770 13368 9826 13424
rect 10138 13776 10194 13832
rect 10138 13368 10194 13424
rect 9678 12688 9734 12744
rect 9586 11756 9642 11758
rect 9586 11704 9588 11756
rect 9588 11704 9640 11756
rect 9640 11704 9642 11756
rect 9586 11702 9642 11704
rect 9862 11736 9918 11792
rect 9770 11192 9826 11248
rect 9954 11056 10010 11112
rect 9862 10784 9918 10840
rect 9494 9832 9550 9888
rect 9402 9324 9404 9344
rect 9404 9324 9456 9344
rect 9456 9324 9458 9344
rect 9402 9288 9458 9324
rect 9126 6568 9182 6624
rect 8482 5208 8538 5264
rect 8758 5208 8814 5264
rect 8758 4256 8814 4312
rect 9678 8472 9734 8528
rect 9770 8200 9826 8256
rect 10046 9424 10102 9480
rect 9862 7656 9918 7712
rect 9586 5888 9642 5944
rect 9494 3168 9550 3224
rect 9862 7248 9918 7304
rect 10046 7404 10102 7440
rect 10046 7384 10048 7404
rect 10048 7384 10100 7404
rect 10100 7384 10102 7404
rect 10414 13776 10470 13832
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 11334 18672 11390 18728
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 11518 16088 11574 16144
rect 11058 14456 11114 14512
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11334 13504 11390 13560
rect 11058 13268 11060 13288
rect 11060 13268 11112 13288
rect 11112 13268 11114 13288
rect 11058 13232 11114 13268
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 10506 10512 10562 10568
rect 10506 10140 10508 10160
rect 10508 10140 10560 10160
rect 10560 10140 10562 10160
rect 10506 10104 10562 10140
rect 10230 6296 10286 6352
rect 9862 3984 9918 4040
rect 10138 4004 10194 4040
rect 10138 3984 10140 4004
rect 10140 3984 10192 4004
rect 10192 3984 10194 4004
rect 9770 3476 9772 3496
rect 9772 3476 9824 3496
rect 9824 3476 9826 3496
rect 9770 3440 9826 3476
rect 10230 3032 10286 3088
rect 9862 2896 9918 2952
rect 10690 7148 10692 7168
rect 10692 7148 10744 7168
rect 10744 7148 10746 7168
rect 10690 7112 10746 7148
rect 10690 6976 10746 7032
rect 10506 5228 10562 5264
rect 10506 5208 10508 5228
rect 10508 5208 10560 5228
rect 10560 5208 10562 5228
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11426 9424 11482 9480
rect 11518 9052 11520 9072
rect 11520 9052 11572 9072
rect 11572 9052 11574 9072
rect 11518 9016 11574 9052
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11610 7828 11612 7848
rect 11612 7828 11664 7848
rect 11664 7828 11666 7848
rect 11610 7792 11666 7828
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11610 7112 11666 7168
rect 11978 18128 12034 18184
rect 12162 17176 12218 17232
rect 12254 17060 12310 17096
rect 12254 17040 12256 17060
rect 12256 17040 12308 17060
rect 12308 17040 12310 17060
rect 12254 15444 12256 15464
rect 12256 15444 12308 15464
rect 12308 15444 12310 15464
rect 12254 15408 12310 15444
rect 13450 18672 13506 18728
rect 12898 18128 12954 18184
rect 12070 12824 12126 12880
rect 11702 6860 11758 6896
rect 11702 6840 11704 6860
rect 11704 6840 11756 6860
rect 11756 6840 11758 6860
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 10782 3440 10838 3496
rect 10690 3168 10746 3224
rect 10506 2896 10562 2952
rect 10690 2932 10692 2952
rect 10692 2932 10744 2952
rect 10744 2932 10746 2952
rect 10690 2896 10746 2932
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 11518 4800 11574 4856
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 11518 3476 11520 3496
rect 11520 3476 11572 3496
rect 11572 3476 11574 3496
rect 11518 3440 11574 3476
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 11702 3168 11758 3224
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 12438 13232 12494 13288
rect 12438 11756 12494 11792
rect 12438 11736 12440 11756
rect 12440 11736 12492 11756
rect 12492 11736 12494 11756
rect 12254 10104 12310 10160
rect 12714 12824 12770 12880
rect 12714 11348 12770 11384
rect 12714 11328 12716 11348
rect 12716 11328 12768 11348
rect 12768 11328 12770 11348
rect 12898 15408 12954 15464
rect 12990 14320 13046 14376
rect 12254 6976 12310 7032
rect 12530 9016 12586 9072
rect 13634 15428 13690 15464
rect 13634 15408 13636 15428
rect 13636 15408 13688 15428
rect 13688 15408 13690 15428
rect 13818 17040 13874 17096
rect 12714 9152 12770 9208
rect 12622 8880 12678 8936
rect 12898 9560 12954 9616
rect 13174 10512 13230 10568
rect 13266 10104 13322 10160
rect 12714 2896 12770 2952
rect 13174 7928 13230 7984
rect 13358 7828 13360 7848
rect 13360 7828 13412 7848
rect 13412 7828 13414 7848
rect 13174 6704 13230 6760
rect 13358 7792 13414 7828
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 15014 15544 15070 15600
rect 14094 15000 14150 15056
rect 13910 12688 13966 12744
rect 13634 11328 13690 11384
rect 13818 9288 13874 9344
rect 13818 6840 13874 6896
rect 14094 6296 14150 6352
rect 13174 4800 13230 4856
rect 13174 4020 13176 4040
rect 13176 4020 13228 4040
rect 13228 4020 13230 4040
rect 13174 3984 13230 4020
rect 13910 5888 13966 5944
rect 14002 5228 14058 5264
rect 14002 5208 14004 5228
rect 14004 5208 14056 5228
rect 14056 5208 14058 5228
rect 13818 3032 13874 3088
rect 14278 8472 14334 8528
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 14646 11192 14702 11248
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 14370 7520 14426 7576
rect 15382 13776 15438 13832
rect 15198 9424 15254 9480
rect 15014 7248 15070 7304
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 15750 13388 15806 13424
rect 15750 13368 15752 13388
rect 15752 13368 15804 13388
rect 15804 13368 15806 13388
rect 15842 12824 15898 12880
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 16578 6704 16634 6760
rect 15658 3576 15714 3632
rect 16026 3168 16082 3224
rect 17038 6160 17094 6216
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 17958 5772 18014 5808
rect 17958 5752 17960 5772
rect 17960 5752 18012 5772
rect 18012 5752 18014 5772
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 18694 5752 18750 5808
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 2870 176 2926 232
<< metal3 >>
rect 0 22538 480 22568
rect 2773 22538 2839 22541
rect 0 22536 2839 22538
rect 0 22480 2778 22536
rect 2834 22480 2839 22536
rect 0 22478 2839 22480
rect 0 22448 480 22478
rect 2773 22475 2839 22478
rect 0 22130 480 22160
rect 3693 22130 3759 22133
rect 0 22128 3759 22130
rect 0 22072 3698 22128
rect 3754 22072 3759 22128
rect 0 22070 3759 22072
rect 0 22040 480 22070
rect 3693 22067 3759 22070
rect 0 21586 480 21616
rect 3141 21586 3207 21589
rect 0 21584 3207 21586
rect 0 21528 3146 21584
rect 3202 21528 3207 21584
rect 0 21526 3207 21528
rect 0 21496 480 21526
rect 3141 21523 3207 21526
rect 0 21178 480 21208
rect 3601 21178 3667 21181
rect 0 21176 3667 21178
rect 0 21120 3606 21176
rect 3662 21120 3667 21176
rect 0 21118 3667 21120
rect 0 21088 480 21118
rect 3601 21115 3667 21118
rect 0 20634 480 20664
rect 3693 20634 3759 20637
rect 0 20632 3759 20634
rect 0 20576 3698 20632
rect 3754 20576 3759 20632
rect 0 20574 3759 20576
rect 0 20544 480 20574
rect 3693 20571 3759 20574
rect 0 20226 480 20256
rect 4061 20226 4127 20229
rect 0 20224 4127 20226
rect 0 20168 4066 20224
rect 4122 20168 4127 20224
rect 0 20166 4127 20168
rect 0 20136 480 20166
rect 4061 20163 4127 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 20095 14992 20096
rect 0 19682 480 19712
rect 1853 19682 1919 19685
rect 0 19680 1919 19682
rect 0 19624 1858 19680
rect 1914 19624 1919 19680
rect 0 19622 1919 19624
rect 0 19592 480 19622
rect 1853 19619 1919 19622
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 0 19274 480 19304
rect 1761 19274 1827 19277
rect 0 19272 1827 19274
rect 0 19216 1766 19272
rect 1822 19216 1827 19272
rect 0 19214 1827 19216
rect 0 19184 480 19214
rect 1761 19211 1827 19214
rect 4521 19138 4587 19141
rect 6637 19138 6703 19141
rect 4521 19136 6703 19138
rect 4521 19080 4526 19136
rect 4582 19080 6642 19136
rect 6698 19080 6703 19136
rect 4521 19078 6703 19080
rect 4521 19075 4587 19078
rect 6637 19075 6703 19078
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 10133 18866 10199 18869
rect 10685 18866 10751 18869
rect 10133 18864 10751 18866
rect 10133 18808 10138 18864
rect 10194 18808 10690 18864
rect 10746 18808 10751 18864
rect 10133 18806 10751 18808
rect 10133 18803 10199 18806
rect 10685 18803 10751 18806
rect 0 18730 480 18760
rect 1577 18730 1643 18733
rect 0 18728 1643 18730
rect 0 18672 1582 18728
rect 1638 18672 1643 18728
rect 0 18670 1643 18672
rect 0 18640 480 18670
rect 1577 18667 1643 18670
rect 11329 18730 11395 18733
rect 13445 18730 13511 18733
rect 11329 18728 13511 18730
rect 11329 18672 11334 18728
rect 11390 18672 13450 18728
rect 13506 18672 13511 18728
rect 11329 18670 13511 18672
rect 11329 18667 11395 18670
rect 13445 18667 13511 18670
rect 2589 18594 2655 18597
rect 3509 18594 3575 18597
rect 2589 18592 3575 18594
rect 2589 18536 2594 18592
rect 2650 18536 3514 18592
rect 3570 18536 3575 18592
rect 2589 18534 3575 18536
rect 2589 18531 2655 18534
rect 3509 18531 3575 18534
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 0 18322 480 18352
rect 1669 18322 1735 18325
rect 0 18320 1735 18322
rect 0 18264 1674 18320
rect 1730 18264 1735 18320
rect 0 18262 1735 18264
rect 0 18232 480 18262
rect 1669 18259 1735 18262
rect 3141 18322 3207 18325
rect 5533 18322 5599 18325
rect 3141 18320 5599 18322
rect 3141 18264 3146 18320
rect 3202 18264 5538 18320
rect 5594 18264 5599 18320
rect 3141 18262 5599 18264
rect 3141 18259 3207 18262
rect 5533 18259 5599 18262
rect 2129 18186 2195 18189
rect 4889 18186 4955 18189
rect 2129 18184 4955 18186
rect 2129 18128 2134 18184
rect 2190 18128 4894 18184
rect 4950 18128 4955 18184
rect 2129 18126 4955 18128
rect 2129 18123 2195 18126
rect 4889 18123 4955 18126
rect 11973 18186 12039 18189
rect 12893 18186 12959 18189
rect 11973 18184 12959 18186
rect 11973 18128 11978 18184
rect 12034 18128 12898 18184
rect 12954 18128 12959 18184
rect 11973 18126 12959 18128
rect 11973 18123 12039 18126
rect 12893 18123 12959 18126
rect 7808 17984 8128 17985
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 0 17778 480 17808
rect 2773 17778 2839 17781
rect 0 17776 2839 17778
rect 0 17720 2778 17776
rect 2834 17720 2839 17776
rect 0 17718 2839 17720
rect 0 17688 480 17718
rect 2773 17715 2839 17718
rect 3417 17776 3483 17781
rect 3417 17720 3422 17776
rect 3478 17720 3483 17776
rect 3417 17715 3483 17720
rect 4061 17778 4127 17781
rect 5073 17778 5139 17781
rect 4061 17776 5139 17778
rect 4061 17720 4066 17776
rect 4122 17720 5078 17776
rect 5134 17720 5139 17776
rect 4061 17718 5139 17720
rect 4061 17715 4127 17718
rect 5073 17715 5139 17718
rect 5349 17778 5415 17781
rect 10133 17778 10199 17781
rect 5349 17776 10199 17778
rect 5349 17720 5354 17776
rect 5410 17720 10138 17776
rect 10194 17720 10199 17776
rect 5349 17718 10199 17720
rect 5349 17715 5415 17718
rect 10133 17715 10199 17718
rect 3141 17642 3207 17645
rect 3420 17642 3480 17715
rect 3141 17640 3480 17642
rect 3141 17584 3146 17640
rect 3202 17584 3480 17640
rect 3141 17582 3480 17584
rect 3141 17579 3207 17582
rect 4376 17440 4696 17441
rect 0 17370 480 17400
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 1761 17370 1827 17373
rect 0 17368 1827 17370
rect 0 17312 1766 17368
rect 1822 17312 1827 17368
rect 0 17310 1827 17312
rect 0 17280 480 17310
rect 1761 17307 1827 17310
rect 12157 17234 12223 17237
rect 22320 17234 22800 17264
rect 12157 17232 22800 17234
rect 12157 17176 12162 17232
rect 12218 17176 22800 17232
rect 12157 17174 22800 17176
rect 12157 17171 12223 17174
rect 22320 17144 22800 17174
rect 1945 17098 2011 17101
rect 6453 17098 6519 17101
rect 1945 17096 6519 17098
rect 1945 17040 1950 17096
rect 2006 17040 6458 17096
rect 6514 17040 6519 17096
rect 1945 17038 6519 17040
rect 1945 17035 2011 17038
rect 6453 17035 6519 17038
rect 12249 17098 12315 17101
rect 13813 17098 13879 17101
rect 12249 17096 13879 17098
rect 12249 17040 12254 17096
rect 12310 17040 13818 17096
rect 13874 17040 13879 17096
rect 12249 17038 13879 17040
rect 12249 17035 12315 17038
rect 13813 17035 13879 17038
rect 7808 16896 8128 16897
rect 0 16826 480 16856
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 16831 14992 16832
rect 1853 16826 1919 16829
rect 0 16824 1919 16826
rect 0 16768 1858 16824
rect 1914 16768 1919 16824
rect 0 16766 1919 16768
rect 0 16736 480 16766
rect 1853 16763 1919 16766
rect 5993 16826 6059 16829
rect 6545 16826 6611 16829
rect 5993 16824 6611 16826
rect 5993 16768 5998 16824
rect 6054 16768 6550 16824
rect 6606 16768 6611 16824
rect 5993 16766 6611 16768
rect 5993 16763 6059 16766
rect 6545 16763 6611 16766
rect 3417 16690 3483 16693
rect 6361 16690 6427 16693
rect 3417 16688 6427 16690
rect 3417 16632 3422 16688
rect 3478 16632 6366 16688
rect 6422 16632 6427 16688
rect 3417 16630 6427 16632
rect 3417 16627 3483 16630
rect 6361 16627 6427 16630
rect 9949 16556 10015 16557
rect 9949 16554 9996 16556
rect 9904 16552 9996 16554
rect 9904 16496 9954 16552
rect 9904 16494 9996 16496
rect 9949 16492 9996 16494
rect 10060 16492 10066 16556
rect 9949 16491 10015 16492
rect 0 16418 480 16448
rect 1945 16418 2011 16421
rect 0 16416 2011 16418
rect 0 16360 1950 16416
rect 2006 16360 2011 16416
rect 0 16358 2011 16360
rect 0 16328 480 16358
rect 1945 16355 2011 16358
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 6177 16146 6243 16149
rect 6453 16146 6519 16149
rect 6177 16144 6519 16146
rect 6177 16088 6182 16144
rect 6238 16088 6458 16144
rect 6514 16088 6519 16144
rect 6177 16086 6519 16088
rect 6177 16083 6243 16086
rect 6453 16083 6519 16086
rect 6821 16146 6887 16149
rect 11513 16146 11579 16149
rect 6821 16144 11579 16146
rect 6821 16088 6826 16144
rect 6882 16088 11518 16144
rect 11574 16088 11579 16144
rect 6821 16086 11579 16088
rect 6821 16083 6887 16086
rect 11513 16083 11579 16086
rect 1761 16010 1827 16013
rect 8293 16010 8359 16013
rect 1761 16008 8359 16010
rect 1761 15952 1766 16008
rect 1822 15952 8298 16008
rect 8354 15952 8359 16008
rect 1761 15950 8359 15952
rect 1761 15947 1827 15950
rect 8293 15947 8359 15950
rect 0 15874 480 15904
rect 1577 15874 1643 15877
rect 0 15872 1643 15874
rect 0 15816 1582 15872
rect 1638 15816 1643 15872
rect 0 15814 1643 15816
rect 0 15784 480 15814
rect 1577 15811 1643 15814
rect 2865 15874 2931 15877
rect 6177 15874 6243 15877
rect 2865 15872 6243 15874
rect 2865 15816 2870 15872
rect 2926 15816 6182 15872
rect 6238 15816 6243 15872
rect 2865 15814 6243 15816
rect 2865 15811 2931 15814
rect 6177 15811 6243 15814
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 3785 15738 3851 15741
rect 4061 15738 4127 15741
rect 3785 15736 4127 15738
rect 3785 15680 3790 15736
rect 3846 15680 4066 15736
rect 4122 15680 4127 15736
rect 3785 15678 4127 15680
rect 3785 15675 3851 15678
rect 4061 15675 4127 15678
rect 2405 15602 2471 15605
rect 15009 15602 15075 15605
rect 2405 15600 15075 15602
rect 2405 15544 2410 15600
rect 2466 15544 15014 15600
rect 15070 15544 15075 15600
rect 2405 15542 15075 15544
rect 2405 15539 2471 15542
rect 15009 15539 15075 15542
rect 0 15466 480 15496
rect 3417 15466 3483 15469
rect 8017 15466 8083 15469
rect 0 15464 3483 15466
rect 0 15408 3422 15464
rect 3478 15408 3483 15464
rect 0 15406 3483 15408
rect 0 15376 480 15406
rect 3417 15403 3483 15406
rect 4156 15464 8083 15466
rect 4156 15408 8022 15464
rect 8078 15408 8083 15464
rect 4156 15406 8083 15408
rect 2589 15330 2655 15333
rect 4156 15330 4216 15406
rect 8017 15403 8083 15406
rect 12249 15466 12315 15469
rect 12893 15466 12959 15469
rect 13629 15466 13695 15469
rect 12249 15464 13695 15466
rect 12249 15408 12254 15464
rect 12310 15408 12898 15464
rect 12954 15408 13634 15464
rect 13690 15408 13695 15464
rect 12249 15406 13695 15408
rect 12249 15403 12315 15406
rect 12893 15403 12959 15406
rect 13629 15403 13695 15406
rect 2589 15328 4216 15330
rect 2589 15272 2594 15328
rect 2650 15272 4216 15328
rect 2589 15270 4216 15272
rect 2589 15267 2655 15270
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 4613 15058 4679 15061
rect 5441 15058 5507 15061
rect 4613 15056 5507 15058
rect 4613 15000 4618 15056
rect 4674 15000 5446 15056
rect 5502 15000 5507 15056
rect 4613 14998 5507 15000
rect 4613 14995 4679 14998
rect 5441 14995 5507 14998
rect 6453 15058 6519 15061
rect 8937 15058 9003 15061
rect 14089 15058 14155 15061
rect 6453 15056 14155 15058
rect 6453 15000 6458 15056
rect 6514 15000 8942 15056
rect 8998 15000 14094 15056
rect 14150 15000 14155 15056
rect 6453 14998 14155 15000
rect 6453 14995 6519 14998
rect 8937 14995 9003 14998
rect 14089 14995 14155 14998
rect 0 14922 480 14952
rect 1669 14922 1735 14925
rect 0 14920 1735 14922
rect 0 14864 1674 14920
rect 1730 14864 1735 14920
rect 0 14862 1735 14864
rect 0 14832 480 14862
rect 1669 14859 1735 14862
rect 3969 14922 4035 14925
rect 7097 14922 7163 14925
rect 9029 14922 9095 14925
rect 3969 14920 9095 14922
rect 3969 14864 3974 14920
rect 4030 14864 7102 14920
rect 7158 14864 9034 14920
rect 9090 14864 9095 14920
rect 3969 14862 9095 14864
rect 3969 14859 4035 14862
rect 7097 14859 7163 14862
rect 9029 14859 9095 14862
rect 7808 14720 8128 14721
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 2497 14650 2563 14653
rect 5993 14650 6059 14653
rect 2497 14648 6059 14650
rect 2497 14592 2502 14648
rect 2558 14592 5998 14648
rect 6054 14592 6059 14648
rect 2497 14590 6059 14592
rect 2497 14587 2563 14590
rect 5993 14587 6059 14590
rect 0 14514 480 14544
rect 3325 14514 3391 14517
rect 0 14512 3391 14514
rect 0 14456 3330 14512
rect 3386 14456 3391 14512
rect 0 14454 3391 14456
rect 0 14424 480 14454
rect 3325 14451 3391 14454
rect 6177 14514 6243 14517
rect 11053 14514 11119 14517
rect 6177 14512 11119 14514
rect 6177 14456 6182 14512
rect 6238 14456 11058 14512
rect 11114 14456 11119 14512
rect 6177 14454 11119 14456
rect 6177 14451 6243 14454
rect 11053 14451 11119 14454
rect 8937 14378 9003 14381
rect 12985 14378 13051 14381
rect 8937 14376 13051 14378
rect 8937 14320 8942 14376
rect 8998 14320 12990 14376
rect 13046 14320 13051 14376
rect 8937 14318 13051 14320
rect 8937 14315 9003 14318
rect 12985 14315 13051 14318
rect 4376 14176 4696 14177
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 5441 14106 5507 14109
rect 9213 14106 9279 14109
rect 5441 14104 9279 14106
rect 5441 14048 5446 14104
rect 5502 14048 9218 14104
rect 9274 14048 9279 14104
rect 5441 14046 9279 14048
rect 5441 14043 5507 14046
rect 9213 14043 9279 14046
rect 9857 14106 9923 14109
rect 9857 14104 10058 14106
rect 9857 14048 9862 14104
rect 9918 14048 10058 14104
rect 9857 14046 10058 14048
rect 9857 14043 9923 14046
rect 0 13970 480 14000
rect 2957 13970 3023 13973
rect 0 13968 3023 13970
rect 0 13912 2962 13968
rect 3018 13912 3023 13968
rect 0 13910 3023 13912
rect 0 13880 480 13910
rect 2957 13907 3023 13910
rect 5993 13834 6059 13837
rect 8753 13834 8819 13837
rect 5993 13832 8819 13834
rect 5993 13776 5998 13832
rect 6054 13776 8758 13832
rect 8814 13776 8819 13832
rect 5993 13774 8819 13776
rect 9998 13834 10058 14046
rect 10133 13834 10199 13837
rect 9998 13832 10199 13834
rect 9998 13776 10138 13832
rect 10194 13776 10199 13832
rect 9998 13774 10199 13776
rect 5993 13771 6059 13774
rect 8753 13771 8819 13774
rect 10133 13771 10199 13774
rect 10409 13834 10475 13837
rect 15377 13834 15443 13837
rect 10409 13832 15443 13834
rect 10409 13776 10414 13832
rect 10470 13776 15382 13832
rect 15438 13776 15443 13832
rect 10409 13774 15443 13776
rect 10409 13771 10475 13774
rect 15377 13771 15443 13774
rect 7808 13632 8128 13633
rect 0 13562 480 13592
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 13567 14992 13568
rect 4061 13562 4127 13565
rect 11329 13562 11395 13565
rect 0 13560 4127 13562
rect 0 13504 4066 13560
rect 4122 13504 4127 13560
rect 0 13502 4127 13504
rect 0 13472 480 13502
rect 4061 13499 4127 13502
rect 9814 13560 11395 13562
rect 9814 13504 11334 13560
rect 11390 13504 11395 13560
rect 9814 13502 11395 13504
rect 9814 13429 9874 13502
rect 11329 13499 11395 13502
rect 9765 13424 9874 13429
rect 9765 13368 9770 13424
rect 9826 13368 9874 13424
rect 9765 13366 9874 13368
rect 10133 13426 10199 13429
rect 15745 13426 15811 13429
rect 10133 13424 15811 13426
rect 10133 13368 10138 13424
rect 10194 13368 15750 13424
rect 15806 13368 15811 13424
rect 10133 13366 15811 13368
rect 9765 13363 9831 13366
rect 10133 13363 10199 13366
rect 15745 13363 15811 13366
rect 11053 13290 11119 13293
rect 12433 13290 12499 13293
rect 11053 13288 12499 13290
rect 11053 13232 11058 13288
rect 11114 13232 12438 13288
rect 12494 13232 12499 13288
rect 11053 13230 12499 13232
rect 11053 13227 11119 13230
rect 12433 13227 12499 13230
rect 4376 13088 4696 13089
rect 0 13018 480 13048
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 0 12958 4216 13018
rect 0 12928 480 12958
rect 4156 12882 4216 12958
rect 12065 12882 12131 12885
rect 4156 12880 12131 12882
rect 4156 12824 12070 12880
rect 12126 12824 12131 12880
rect 4156 12822 12131 12824
rect 12065 12819 12131 12822
rect 12709 12882 12775 12885
rect 15837 12882 15903 12885
rect 12709 12880 15903 12882
rect 12709 12824 12714 12880
rect 12770 12824 15842 12880
rect 15898 12824 15903 12880
rect 12709 12822 15903 12824
rect 12709 12819 12775 12822
rect 15837 12819 15903 12822
rect 9673 12746 9739 12749
rect 13905 12746 13971 12749
rect 9673 12744 13971 12746
rect 9673 12688 9678 12744
rect 9734 12688 13910 12744
rect 13966 12688 13971 12744
rect 9673 12686 13971 12688
rect 9673 12683 9739 12686
rect 13905 12683 13971 12686
rect 0 12610 480 12640
rect 3969 12610 4035 12613
rect 4889 12610 4955 12613
rect 0 12608 4035 12610
rect 0 12552 3974 12608
rect 4030 12552 4035 12608
rect 0 12550 4035 12552
rect 0 12520 480 12550
rect 3969 12547 4035 12550
rect 4846 12608 4955 12610
rect 4846 12552 4894 12608
rect 4950 12552 4955 12608
rect 4846 12547 4955 12552
rect 6177 12610 6243 12613
rect 6913 12610 6979 12613
rect 6177 12608 6979 12610
rect 6177 12552 6182 12608
rect 6238 12552 6918 12608
rect 6974 12552 6979 12608
rect 6177 12550 6979 12552
rect 6177 12547 6243 12550
rect 6913 12547 6979 12550
rect 4429 12338 4495 12341
rect 4846 12338 4906 12547
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 9029 12338 9095 12341
rect 4429 12336 9095 12338
rect 4429 12280 4434 12336
rect 4490 12280 9034 12336
rect 9090 12280 9095 12336
rect 4429 12278 9095 12280
rect 4429 12275 4495 12278
rect 9029 12275 9095 12278
rect 3509 12202 3575 12205
rect 8753 12202 8819 12205
rect 3509 12200 8819 12202
rect 3509 12144 3514 12200
rect 3570 12144 8758 12200
rect 8814 12144 8819 12200
rect 3509 12142 8819 12144
rect 3509 12139 3575 12142
rect 8753 12139 8819 12142
rect 0 12066 480 12096
rect 3601 12066 3667 12069
rect 0 12064 3667 12066
rect 0 12008 3606 12064
rect 3662 12008 3667 12064
rect 0 12006 3667 12008
rect 0 11976 480 12006
rect 3601 12003 3667 12006
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 9121 11794 9187 11797
rect 9305 11794 9371 11797
rect 9857 11794 9923 11797
rect 12433 11794 12499 11797
rect 9121 11792 9644 11794
rect 9121 11736 9126 11792
rect 9182 11736 9310 11792
rect 9366 11763 9644 11792
rect 9857 11792 12499 11794
rect 9366 11758 9647 11763
rect 9366 11736 9586 11758
rect 9121 11734 9586 11736
rect 9121 11731 9187 11734
rect 9305 11731 9371 11734
rect 9581 11702 9586 11734
rect 9642 11702 9647 11758
rect 9857 11736 9862 11792
rect 9918 11736 12438 11792
rect 12494 11736 12499 11792
rect 9857 11734 12499 11736
rect 9857 11731 9923 11734
rect 12433 11731 12499 11734
rect 9581 11697 9647 11702
rect 0 11658 480 11688
rect 4153 11658 4219 11661
rect 0 11656 4219 11658
rect 0 11600 4158 11656
rect 4214 11600 4219 11656
rect 0 11598 4219 11600
rect 0 11568 480 11598
rect 4153 11595 4219 11598
rect 7808 11456 8128 11457
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 8753 11386 8819 11389
rect 12709 11386 12775 11389
rect 13629 11386 13695 11389
rect 8753 11384 10012 11386
rect 8753 11328 8758 11384
rect 8814 11328 10012 11384
rect 8753 11326 10012 11328
rect 8753 11323 8819 11326
rect 9765 11250 9831 11253
rect 9952 11250 10012 11326
rect 12709 11384 13695 11386
rect 12709 11328 12714 11384
rect 12770 11328 13634 11384
rect 13690 11328 13695 11384
rect 12709 11326 13695 11328
rect 12709 11323 12775 11326
rect 13629 11323 13695 11326
rect 14641 11250 14707 11253
rect 9765 11248 9874 11250
rect 9765 11192 9770 11248
rect 9826 11192 9874 11248
rect 9765 11187 9874 11192
rect 9952 11248 14707 11250
rect 9952 11192 14646 11248
rect 14702 11192 14707 11248
rect 9952 11190 14707 11192
rect 14641 11187 14707 11190
rect 0 11114 480 11144
rect 8477 11114 8543 11117
rect 0 11112 8543 11114
rect 0 11056 8482 11112
rect 8538 11056 8543 11112
rect 0 11054 8543 11056
rect 9814 11114 9874 11187
rect 9949 11114 10015 11117
rect 9814 11112 10015 11114
rect 9814 11056 9954 11112
rect 10010 11056 10015 11112
rect 9814 11054 10015 11056
rect 0 11024 480 11054
rect 8477 11051 8543 11054
rect 9949 11051 10015 11054
rect 4376 10912 4696 10913
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 9857 10842 9923 10845
rect 9990 10842 9996 10844
rect 9857 10840 9996 10842
rect 9857 10784 9862 10840
rect 9918 10784 9996 10840
rect 9857 10782 9996 10784
rect 9857 10779 9923 10782
rect 9990 10780 9996 10782
rect 10060 10780 10066 10844
rect 0 10706 480 10736
rect 1393 10706 1459 10709
rect 0 10704 1459 10706
rect 0 10648 1398 10704
rect 1454 10648 1459 10704
rect 0 10646 1459 10648
rect 0 10616 480 10646
rect 1393 10643 1459 10646
rect 8569 10570 8635 10573
rect 10501 10570 10567 10573
rect 13169 10570 13235 10573
rect 8569 10568 13235 10570
rect 8569 10512 8574 10568
rect 8630 10512 10506 10568
rect 10562 10512 13174 10568
rect 13230 10512 13235 10568
rect 8569 10510 13235 10512
rect 8569 10507 8635 10510
rect 10501 10507 10567 10510
rect 13169 10507 13235 10510
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 10303 14992 10304
rect 0 10162 480 10192
rect 3969 10162 4035 10165
rect 0 10160 4035 10162
rect 0 10104 3974 10160
rect 4030 10104 4035 10160
rect 0 10102 4035 10104
rect 0 10072 480 10102
rect 3969 10099 4035 10102
rect 10501 10162 10567 10165
rect 12249 10162 12315 10165
rect 13261 10162 13327 10165
rect 10501 10160 13327 10162
rect 10501 10104 10506 10160
rect 10562 10104 12254 10160
rect 12310 10104 13266 10160
rect 13322 10104 13327 10160
rect 10501 10102 13327 10104
rect 10501 10099 10567 10102
rect 12249 10099 12315 10102
rect 13261 10099 13327 10102
rect 7598 9828 7604 9892
rect 7668 9890 7674 9892
rect 9489 9890 9555 9893
rect 7668 9888 9555 9890
rect 7668 9832 9494 9888
rect 9550 9832 9555 9888
rect 7668 9830 9555 9832
rect 7668 9828 7674 9830
rect 9489 9827 9555 9830
rect 4376 9824 4696 9825
rect 0 9754 480 9784
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 4061 9754 4127 9757
rect 0 9752 4127 9754
rect 0 9696 4066 9752
rect 4122 9696 4127 9752
rect 0 9694 4127 9696
rect 0 9664 480 9694
rect 4061 9691 4127 9694
rect 7414 9556 7420 9620
rect 7484 9618 7490 9620
rect 12893 9618 12959 9621
rect 7484 9616 12959 9618
rect 7484 9560 12898 9616
rect 12954 9560 12959 9616
rect 7484 9558 12959 9560
rect 7484 9556 7490 9558
rect 12893 9555 12959 9558
rect 2814 9420 2820 9484
rect 2884 9482 2890 9484
rect 2957 9482 3023 9485
rect 2884 9480 3023 9482
rect 2884 9424 2962 9480
rect 3018 9424 3023 9480
rect 2884 9422 3023 9424
rect 2884 9420 2890 9422
rect 2957 9419 3023 9422
rect 4981 9482 5047 9485
rect 5993 9482 6059 9485
rect 4981 9480 6059 9482
rect 4981 9424 4986 9480
rect 5042 9424 5998 9480
rect 6054 9424 6059 9480
rect 4981 9422 6059 9424
rect 4981 9419 5047 9422
rect 5993 9419 6059 9422
rect 6729 9482 6795 9485
rect 10041 9482 10107 9485
rect 6729 9480 10107 9482
rect 6729 9424 6734 9480
rect 6790 9424 10046 9480
rect 10102 9424 10107 9480
rect 6729 9422 10107 9424
rect 6729 9419 6795 9422
rect 10041 9419 10107 9422
rect 11421 9482 11487 9485
rect 15193 9482 15259 9485
rect 11421 9480 15259 9482
rect 11421 9424 11426 9480
rect 11482 9424 15198 9480
rect 15254 9424 15259 9480
rect 11421 9422 15259 9424
rect 11421 9419 11487 9422
rect 15193 9419 15259 9422
rect 9397 9346 9463 9349
rect 13813 9346 13879 9349
rect 9397 9344 13879 9346
rect 9397 9288 9402 9344
rect 9458 9288 13818 9344
rect 13874 9288 13879 9344
rect 9397 9286 13879 9288
rect 9397 9283 9463 9286
rect 13813 9283 13879 9286
rect 7808 9280 8128 9281
rect 0 9210 480 9240
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 0 9150 4906 9210
rect 0 9120 480 9150
rect 4846 9074 4906 9150
rect 7230 9148 7236 9212
rect 7300 9210 7306 9212
rect 7465 9210 7531 9213
rect 7300 9208 7531 9210
rect 7300 9152 7470 9208
rect 7526 9152 7531 9208
rect 7300 9150 7531 9152
rect 7300 9148 7306 9150
rect 7465 9147 7531 9150
rect 8293 9210 8359 9213
rect 12709 9210 12775 9213
rect 8293 9208 12775 9210
rect 8293 9152 8298 9208
rect 8354 9152 12714 9208
rect 12770 9152 12775 9208
rect 8293 9150 12775 9152
rect 8293 9147 8359 9150
rect 12709 9147 12775 9150
rect 8385 9074 8451 9077
rect 4846 9072 8451 9074
rect 4846 9016 8390 9072
rect 8446 9016 8451 9072
rect 4846 9014 8451 9016
rect 8385 9011 8451 9014
rect 11513 9074 11579 9077
rect 12525 9074 12591 9077
rect 11513 9072 12634 9074
rect 11513 9016 11518 9072
rect 11574 9016 12530 9072
rect 12586 9016 12634 9072
rect 11513 9014 12634 9016
rect 11513 9011 11579 9014
rect 12525 9011 12634 9014
rect 12574 8941 12634 9011
rect 3417 8938 3483 8941
rect 7465 8940 7531 8941
rect 3417 8936 7298 8938
rect 3417 8880 3422 8936
rect 3478 8880 7298 8936
rect 3417 8878 7298 8880
rect 3417 8875 3483 8878
rect 0 8802 480 8832
rect 3969 8802 4035 8805
rect 0 8800 4035 8802
rect 0 8744 3974 8800
rect 4030 8744 4035 8800
rect 0 8742 4035 8744
rect 7238 8802 7298 8878
rect 7414 8876 7420 8940
rect 7484 8938 7531 8940
rect 7484 8936 7576 8938
rect 7526 8880 7576 8936
rect 7484 8878 7576 8880
rect 12574 8936 12683 8941
rect 12574 8880 12622 8936
rect 12678 8880 12683 8936
rect 12574 8878 12683 8880
rect 7484 8876 7531 8878
rect 7465 8875 7531 8876
rect 12617 8875 12683 8878
rect 7598 8802 7604 8804
rect 7238 8742 7604 8802
rect 0 8712 480 8742
rect 3969 8739 4035 8742
rect 7598 8740 7604 8742
rect 7668 8802 7674 8804
rect 7925 8802 7991 8805
rect 7668 8800 7991 8802
rect 7668 8744 7930 8800
rect 7986 8744 7991 8800
rect 7668 8742 7991 8744
rect 7668 8740 7674 8742
rect 7925 8739 7991 8742
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 8671 18424 8672
rect 7230 8604 7236 8668
rect 7300 8666 7306 8668
rect 8109 8666 8175 8669
rect 7300 8664 8175 8666
rect 7300 8608 8114 8664
rect 8170 8608 8175 8664
rect 7300 8606 8175 8608
rect 7300 8604 7306 8606
rect 8109 8603 8175 8606
rect 9673 8530 9739 8533
rect 14273 8530 14339 8533
rect 9673 8528 14339 8530
rect 9673 8472 9678 8528
rect 9734 8472 14278 8528
rect 14334 8472 14339 8528
rect 9673 8470 14339 8472
rect 9673 8467 9739 8470
rect 14273 8467 14339 8470
rect 0 8258 480 8288
rect 4061 8258 4127 8261
rect 0 8256 4127 8258
rect 0 8200 4066 8256
rect 4122 8200 4127 8256
rect 0 8198 4127 8200
rect 0 8168 480 8198
rect 4061 8195 4127 8198
rect 8661 8258 8727 8261
rect 9765 8258 9831 8261
rect 8661 8256 9831 8258
rect 8661 8200 8666 8256
rect 8722 8200 9770 8256
rect 9826 8200 9831 8256
rect 8661 8198 9831 8200
rect 8661 8195 8727 8198
rect 9765 8195 9831 8198
rect 7808 8192 8128 8193
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 8385 7986 8451 7989
rect 13169 7986 13235 7989
rect 8385 7984 13235 7986
rect 8385 7928 8390 7984
rect 8446 7928 13174 7984
rect 13230 7928 13235 7984
rect 8385 7926 13235 7928
rect 8385 7923 8451 7926
rect 13169 7923 13235 7926
rect 0 7850 480 7880
rect 4061 7850 4127 7853
rect 0 7848 4127 7850
rect 0 7792 4066 7848
rect 4122 7792 4127 7848
rect 0 7790 4127 7792
rect 0 7760 480 7790
rect 4061 7787 4127 7790
rect 11605 7850 11671 7853
rect 13353 7850 13419 7853
rect 11605 7848 13419 7850
rect 11605 7792 11610 7848
rect 11666 7792 13358 7848
rect 13414 7792 13419 7848
rect 11605 7790 13419 7792
rect 11605 7787 11671 7790
rect 13353 7787 13419 7790
rect 9857 7714 9923 7717
rect 10174 7714 10180 7716
rect 9857 7712 10180 7714
rect 9857 7656 9862 7712
rect 9918 7656 10180 7712
rect 9857 7654 10180 7656
rect 9857 7651 9923 7654
rect 10174 7652 10180 7654
rect 10244 7652 10250 7716
rect 4376 7648 4696 7649
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 13118 7516 13124 7580
rect 13188 7578 13194 7580
rect 14365 7578 14431 7581
rect 13188 7576 14431 7578
rect 13188 7520 14370 7576
rect 14426 7520 14431 7576
rect 13188 7518 14431 7520
rect 13188 7516 13194 7518
rect 14365 7515 14431 7518
rect 8201 7442 8267 7445
rect 10041 7442 10107 7445
rect 8201 7440 10107 7442
rect 8201 7384 8206 7440
rect 8262 7384 10046 7440
rect 10102 7384 10107 7440
rect 8201 7382 10107 7384
rect 8201 7379 8267 7382
rect 10041 7379 10107 7382
rect 0 7306 480 7336
rect 2497 7306 2563 7309
rect 0 7304 2563 7306
rect 0 7248 2502 7304
rect 2558 7248 2563 7304
rect 0 7246 2563 7248
rect 0 7216 480 7246
rect 2497 7243 2563 7246
rect 9857 7306 9923 7309
rect 15009 7306 15075 7309
rect 9857 7304 15075 7306
rect 9857 7248 9862 7304
rect 9918 7248 15014 7304
rect 15070 7248 15075 7304
rect 9857 7246 15075 7248
rect 9857 7243 9923 7246
rect 15009 7243 15075 7246
rect 10685 7170 10751 7173
rect 11605 7170 11671 7173
rect 10685 7168 11671 7170
rect 10685 7112 10690 7168
rect 10746 7112 11610 7168
rect 11666 7112 11671 7168
rect 10685 7110 11671 7112
rect 10685 7107 10751 7110
rect 11605 7107 11671 7110
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 7039 14992 7040
rect 10685 7034 10751 7037
rect 12249 7034 12315 7037
rect 10685 7032 12315 7034
rect 10685 6976 10690 7032
rect 10746 6976 12254 7032
rect 12310 6976 12315 7032
rect 10685 6974 12315 6976
rect 10685 6971 10751 6974
rect 12249 6971 12315 6974
rect 0 6898 480 6928
rect 3601 6898 3667 6901
rect 0 6896 3667 6898
rect 0 6840 3606 6896
rect 3662 6840 3667 6896
rect 0 6838 3667 6840
rect 0 6808 480 6838
rect 3601 6835 3667 6838
rect 11697 6898 11763 6901
rect 13813 6898 13879 6901
rect 11697 6896 13879 6898
rect 11697 6840 11702 6896
rect 11758 6840 13818 6896
rect 13874 6840 13879 6896
rect 11697 6838 13879 6840
rect 11697 6835 11763 6838
rect 13813 6835 13879 6838
rect 13169 6762 13235 6765
rect 16573 6762 16639 6765
rect 13169 6760 16639 6762
rect 13169 6704 13174 6760
rect 13230 6704 16578 6760
rect 16634 6704 16639 6760
rect 13169 6702 16639 6704
rect 13169 6699 13235 6702
rect 16573 6699 16639 6702
rect 9121 6626 9187 6629
rect 9078 6624 9187 6626
rect 9078 6568 9126 6624
rect 9182 6568 9187 6624
rect 9078 6563 9187 6568
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 0 6354 480 6384
rect 8661 6354 8727 6357
rect 0 6352 8727 6354
rect 0 6296 8666 6352
rect 8722 6296 8727 6352
rect 0 6294 8727 6296
rect 0 6264 480 6294
rect 8661 6291 8727 6294
rect 6913 6218 6979 6221
rect 9078 6218 9138 6563
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 10225 6354 10291 6357
rect 14089 6354 14155 6357
rect 10225 6352 14155 6354
rect 10225 6296 10230 6352
rect 10286 6296 14094 6352
rect 14150 6296 14155 6352
rect 10225 6294 14155 6296
rect 10225 6291 10291 6294
rect 14089 6291 14155 6294
rect 17033 6218 17099 6221
rect 6913 6216 17099 6218
rect 6913 6160 6918 6216
rect 6974 6160 17038 6216
rect 17094 6160 17099 6216
rect 6913 6158 17099 6160
rect 6913 6155 6979 6158
rect 17033 6155 17099 6158
rect 7808 6016 8128 6017
rect 0 5946 480 5976
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 9581 5946 9647 5949
rect 13905 5946 13971 5949
rect 0 5886 2882 5946
rect 0 5856 480 5886
rect 2822 5674 2882 5886
rect 9581 5944 13971 5946
rect 9581 5888 9586 5944
rect 9642 5888 13910 5944
rect 13966 5888 13971 5944
rect 9581 5886 13971 5888
rect 9581 5883 9647 5886
rect 13905 5883 13971 5886
rect 2957 5810 3023 5813
rect 17953 5810 18019 5813
rect 2957 5808 18019 5810
rect 2957 5752 2962 5808
rect 3018 5752 17958 5808
rect 18014 5752 18019 5808
rect 2957 5750 18019 5752
rect 2957 5747 3023 5750
rect 17953 5747 18019 5750
rect 18689 5810 18755 5813
rect 22320 5810 22800 5840
rect 18689 5808 22800 5810
rect 18689 5752 18694 5808
rect 18750 5752 22800 5808
rect 18689 5750 22800 5752
rect 18689 5747 18755 5750
rect 22320 5720 22800 5750
rect 8201 5674 8267 5677
rect 2822 5672 8267 5674
rect 2822 5616 8206 5672
rect 8262 5616 8267 5672
rect 2822 5614 8267 5616
rect 8201 5611 8267 5614
rect 4376 5472 4696 5473
rect 0 5402 480 5432
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 0 5342 4170 5402
rect 0 5312 480 5342
rect 4110 5266 4170 5342
rect 8477 5266 8543 5269
rect 8753 5266 8819 5269
rect 4110 5264 8819 5266
rect 4110 5208 8482 5264
rect 8538 5208 8758 5264
rect 8814 5208 8819 5264
rect 4110 5206 8819 5208
rect 8477 5203 8543 5206
rect 8753 5203 8819 5206
rect 10501 5266 10567 5269
rect 13997 5266 14063 5269
rect 10501 5264 14063 5266
rect 10501 5208 10506 5264
rect 10562 5208 14002 5264
rect 14058 5208 14063 5264
rect 10501 5206 14063 5208
rect 10501 5203 10567 5206
rect 13997 5203 14063 5206
rect 0 4994 480 5024
rect 4797 4994 4863 4997
rect 0 4992 4863 4994
rect 0 4936 4802 4992
rect 4858 4936 4863 4992
rect 0 4934 4863 4936
rect 0 4904 480 4934
rect 4797 4931 4863 4934
rect 7808 4928 8128 4929
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 11513 4858 11579 4861
rect 13169 4858 13235 4861
rect 11513 4856 13235 4858
rect 11513 4800 11518 4856
rect 11574 4800 13174 4856
rect 13230 4800 13235 4856
rect 11513 4798 13235 4800
rect 11513 4795 11579 4798
rect 13169 4795 13235 4798
rect 0 4450 480 4480
rect 4061 4450 4127 4453
rect 0 4448 4127 4450
rect 0 4392 4066 4448
rect 4122 4392 4127 4448
rect 0 4390 4127 4392
rect 0 4360 480 4390
rect 4061 4387 4127 4390
rect 4376 4384 4696 4385
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 5717 4314 5783 4317
rect 8753 4314 8819 4317
rect 5717 4312 8819 4314
rect 5717 4256 5722 4312
rect 5778 4256 8758 4312
rect 8814 4256 8819 4312
rect 5717 4254 8819 4256
rect 5717 4251 5783 4254
rect 8753 4251 8819 4254
rect 5993 4176 6059 4181
rect 5993 4120 5998 4176
rect 6054 4120 6059 4176
rect 5993 4115 6059 4120
rect 0 4042 480 4072
rect 2773 4042 2839 4045
rect 0 4040 2839 4042
rect 0 3984 2778 4040
rect 2834 3984 2839 4040
rect 0 3982 2839 3984
rect 0 3952 480 3982
rect 2773 3979 2839 3982
rect 5349 4042 5415 4045
rect 5996 4042 6056 4115
rect 9857 4042 9923 4045
rect 5349 4040 9923 4042
rect 5349 3984 5354 4040
rect 5410 3984 9862 4040
rect 9918 3984 9923 4040
rect 5349 3982 9923 3984
rect 5349 3979 5415 3982
rect 9857 3979 9923 3982
rect 10133 4042 10199 4045
rect 13169 4042 13235 4045
rect 10133 4040 13235 4042
rect 10133 3984 10138 4040
rect 10194 3984 13174 4040
rect 13230 3984 13235 4040
rect 10133 3982 13235 3984
rect 10133 3979 10199 3982
rect 13169 3979 13235 3982
rect 4613 3906 4679 3909
rect 4981 3906 5047 3909
rect 4613 3904 5047 3906
rect 4613 3848 4618 3904
rect 4674 3848 4986 3904
rect 5042 3848 5047 3904
rect 4613 3846 5047 3848
rect 4613 3843 4679 3846
rect 4981 3843 5047 3846
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 3775 14992 3776
rect 3785 3634 3851 3637
rect 4889 3634 4955 3637
rect 3785 3632 4955 3634
rect 3785 3576 3790 3632
rect 3846 3576 4894 3632
rect 4950 3576 4955 3632
rect 3785 3574 4955 3576
rect 3785 3571 3851 3574
rect 4889 3571 4955 3574
rect 6177 3634 6243 3637
rect 15653 3634 15719 3637
rect 6177 3632 15719 3634
rect 6177 3576 6182 3632
rect 6238 3576 15658 3632
rect 15714 3576 15719 3632
rect 6177 3574 15719 3576
rect 6177 3571 6243 3574
rect 15653 3571 15719 3574
rect 0 3498 480 3528
rect 3693 3498 3759 3501
rect 0 3496 3759 3498
rect 0 3440 3698 3496
rect 3754 3440 3759 3496
rect 0 3438 3759 3440
rect 0 3408 480 3438
rect 3693 3435 3759 3438
rect 9765 3498 9831 3501
rect 10777 3498 10843 3501
rect 11513 3498 11579 3501
rect 9765 3496 11579 3498
rect 9765 3440 9770 3496
rect 9826 3440 10782 3496
rect 10838 3440 11518 3496
rect 11574 3440 11579 3496
rect 9765 3438 11579 3440
rect 9765 3435 9831 3438
rect 10777 3435 10843 3438
rect 11513 3435 11579 3438
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 9489 3226 9555 3229
rect 10685 3226 10751 3229
rect 9489 3224 10751 3226
rect 9489 3168 9494 3224
rect 9550 3168 10690 3224
rect 10746 3168 10751 3224
rect 9489 3166 10751 3168
rect 9489 3163 9555 3166
rect 10685 3163 10751 3166
rect 11697 3226 11763 3229
rect 16021 3226 16087 3229
rect 11697 3224 16087 3226
rect 11697 3168 11702 3224
rect 11758 3168 16026 3224
rect 16082 3168 16087 3224
rect 11697 3166 16087 3168
rect 11697 3163 11763 3166
rect 16021 3163 16087 3166
rect 0 3090 480 3120
rect 2589 3090 2655 3093
rect 0 3088 2655 3090
rect 0 3032 2594 3088
rect 2650 3032 2655 3088
rect 0 3030 2655 3032
rect 0 3000 480 3030
rect 2589 3027 2655 3030
rect 3417 3090 3483 3093
rect 4337 3090 4403 3093
rect 10225 3092 10291 3093
rect 3417 3088 4403 3090
rect 3417 3032 3422 3088
rect 3478 3032 4342 3088
rect 4398 3032 4403 3088
rect 3417 3030 4403 3032
rect 3417 3027 3483 3030
rect 4337 3027 4403 3030
rect 10174 3028 10180 3092
rect 10244 3090 10291 3092
rect 13813 3090 13879 3093
rect 10244 3088 13879 3090
rect 10286 3032 13818 3088
rect 13874 3032 13879 3088
rect 10244 3030 13879 3032
rect 10244 3028 10291 3030
rect 10225 3027 10291 3028
rect 13813 3027 13879 3030
rect 7414 2892 7420 2956
rect 7484 2954 7490 2956
rect 7557 2954 7623 2957
rect 7484 2952 7623 2954
rect 7484 2896 7562 2952
rect 7618 2896 7623 2952
rect 7484 2894 7623 2896
rect 7484 2892 7490 2894
rect 7557 2891 7623 2894
rect 9857 2954 9923 2957
rect 10501 2954 10567 2957
rect 10685 2954 10751 2957
rect 9857 2952 10751 2954
rect 9857 2896 9862 2952
rect 9918 2896 10506 2952
rect 10562 2896 10690 2952
rect 10746 2896 10751 2952
rect 9857 2894 10751 2896
rect 9857 2891 9923 2894
rect 10501 2891 10567 2894
rect 10685 2891 10751 2894
rect 12709 2954 12775 2957
rect 13118 2954 13124 2956
rect 12709 2952 13124 2954
rect 12709 2896 12714 2952
rect 12770 2896 13124 2952
rect 12709 2894 13124 2896
rect 12709 2891 12775 2894
rect 13118 2892 13124 2894
rect 13188 2892 13194 2956
rect 1945 2818 2011 2821
rect 3141 2818 3207 2821
rect 1945 2816 3207 2818
rect 1945 2760 1950 2816
rect 2006 2760 3146 2816
rect 3202 2760 3207 2816
rect 1945 2758 3207 2760
rect 1945 2755 2011 2758
rect 3141 2755 3207 2758
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 2681 2682 2747 2685
rect 2814 2682 2820 2684
rect 2681 2680 2820 2682
rect 2681 2624 2686 2680
rect 2742 2624 2820 2680
rect 2681 2622 2820 2624
rect 2681 2619 2747 2622
rect 2814 2620 2820 2622
rect 2884 2620 2890 2684
rect 0 2546 480 2576
rect 4061 2546 4127 2549
rect 0 2544 4127 2546
rect 0 2488 4066 2544
rect 4122 2488 4127 2544
rect 0 2486 4127 2488
rect 0 2456 480 2486
rect 4061 2483 4127 2486
rect 4376 2208 4696 2209
rect 0 2138 480 2168
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 2681 2138 2747 2141
rect 0 2136 2747 2138
rect 0 2080 2686 2136
rect 2742 2080 2747 2136
rect 0 2078 2747 2080
rect 0 2048 480 2078
rect 2681 2075 2747 2078
rect 0 1594 480 1624
rect 4061 1594 4127 1597
rect 0 1592 4127 1594
rect 0 1536 4066 1592
rect 4122 1536 4127 1592
rect 0 1534 4127 1536
rect 0 1504 480 1534
rect 4061 1531 4127 1534
rect 0 1186 480 1216
rect 2773 1186 2839 1189
rect 0 1184 2839 1186
rect 0 1128 2778 1184
rect 2834 1128 2839 1184
rect 0 1126 2839 1128
rect 0 1096 480 1126
rect 2773 1123 2839 1126
rect 0 642 480 672
rect 3509 642 3575 645
rect 0 640 3575 642
rect 0 584 3514 640
rect 3570 584 3575 640
rect 0 582 3575 584
rect 0 552 480 582
rect 3509 579 3575 582
rect 0 234 480 264
rect 2865 234 2931 237
rect 0 232 2931 234
rect 0 176 2870 232
rect 2926 176 2931 232
rect 0 174 2931 176
rect 0 144 480 174
rect 2865 171 2931 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 9996 16552 10060 16556
rect 9996 16496 10010 16552
rect 10010 16496 10060 16552
rect 9996 16492 10060 16496
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 9996 10780 10060 10844
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 7604 9828 7668 9892
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 7420 9556 7484 9620
rect 2820 9420 2884 9484
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 7236 9148 7300 9212
rect 7420 8936 7484 8940
rect 7420 8880 7470 8936
rect 7470 8880 7484 8936
rect 7420 8876 7484 8880
rect 7604 8740 7668 8804
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 7236 8604 7300 8668
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 10180 7652 10244 7716
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 13124 7516 13188 7580
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 10180 3088 10244 3092
rect 10180 3032 10230 3088
rect 10230 3032 10244 3088
rect 10180 3028 10244 3032
rect 7420 2892 7484 2956
rect 13124 2892 13188 2956
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 2820 2620 2884 2684
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 9995 16556 10061 16557
rect 9995 16492 9996 16556
rect 10060 16492 10061 16556
rect 9995 16491 10061 16492
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 9998 10845 10058 16491
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 9995 10844 10061 10845
rect 9995 10780 9996 10844
rect 10060 10780 10061 10844
rect 9995 10779 10061 10780
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7603 9892 7669 9893
rect 7603 9828 7604 9892
rect 7668 9828 7669 9892
rect 7603 9827 7669 9828
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 2819 9484 2885 9485
rect 2819 9420 2820 9484
rect 2884 9420 2885 9484
rect 2819 9419 2885 9420
rect 2822 2685 2882 9419
rect 4376 8736 4696 9760
rect 7419 9620 7485 9621
rect 7419 9556 7420 9620
rect 7484 9556 7485 9620
rect 7419 9555 7485 9556
rect 7235 9212 7301 9213
rect 7235 9148 7236 9212
rect 7300 9148 7301 9212
rect 7235 9147 7301 9148
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 7238 8669 7298 9147
rect 7422 8941 7482 9555
rect 7419 8940 7485 8941
rect 7419 8876 7420 8940
rect 7484 8876 7485 8940
rect 7419 8875 7485 8876
rect 7235 8668 7301 8669
rect 7235 8604 7236 8668
rect 7300 8604 7301 8668
rect 7235 8603 7301 8604
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 2819 2684 2885 2685
rect 2819 2620 2820 2684
rect 2884 2620 2885 2684
rect 2819 2619 2885 2620
rect 4376 2208 4696 3232
rect 7422 2957 7482 8875
rect 7606 8805 7666 9827
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7603 8804 7669 8805
rect 7603 8740 7604 8804
rect 7668 8740 7669 8804
rect 7603 8739 7669 8740
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 11240 9824 11560 10848
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 10179 7716 10245 7717
rect 10179 7652 10180 7716
rect 10244 7652 10245 7716
rect 10179 7651 10245 7652
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7419 2956 7485 2957
rect 7419 2892 7420 2956
rect 7484 2892 7485 2956
rect 7419 2891 7485 2892
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 2752 8128 3776
rect 10182 3093 10242 7651
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 13123 7580 13189 7581
rect 13123 7516 13124 7580
rect 13188 7516 13189 7580
rect 13123 7515 13189 7516
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 10179 3092 10245 3093
rect 10179 3028 10180 3092
rect 10244 3028 10245 3092
rect 10179 3027 10245 3028
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 2208 11560 3232
rect 13126 2957 13186 7515
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 13123 2956 13189 2957
rect 13123 2892 13124 2956
rect 13188 2892 13189 2956
rect 13123 2891 13189 2892
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 2668 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1606821651
transform 1 0 2300 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1606821651
transform 1 0 1656 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606821651
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 2116 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp 1606821651
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_15
timestamp 1606821651
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1606821651
transform 1 0 3680 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1606821651
transform 1 0 4692 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_2_
timestamp 1606821651
transform 1 0 4324 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22
timestamp 1606821651
transform 1 0 3128 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3864 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32
timestamp 1606821651
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_26
timestamp 1606821651
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_37
timestamp 1606821651
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_48
timestamp 1606821651
transform 1 0 5520 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44
timestamp 1606821651
transform 1 0 5152 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5336 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1606821651
transform 1 0 5704 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1606821651
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1606821651
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 6164 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606821651
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_62
timestamp 1606821651
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606821651
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 8188 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 6900 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1606821651
transform 1 0 7084 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1606821651
transform 1 0 7636 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1606821651
transform 1 0 8648 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69
timestamp 1606821651
transform 1 0 7452 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_80
timestamp 1606821651
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_74
timestamp 1606821651
transform 1 0 7912 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9844 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1606821651
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606821651
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1606821651
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1606821651
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_93
timestamp 1606821651
transform 1 0 9660 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_104
timestamp 1606821651
transform 1 0 10672 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114
timestamp 1606821651
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1606821651
transform 1 0 10764 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10856 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1606821651
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_115
timestamp 1606821651
transform 1 0 11684 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1606821651
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606821651
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 11776 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1606821651
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606821651
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _087_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 13340 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1606821651
transform 1 0 13892 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1606821651
transform 1 0 14168 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 13432 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_131
timestamp 1606821651
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_137
timestamp 1606821651
transform 1 0 13708 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_143 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_132
timestamp 1606821651
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_140
timestamp 1606821651
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_152
timestamp 1606821651
transform 1 0 15088 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_146
timestamp 1606821651
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_152
timestamp 1606821651
transform 1 0 15088 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_147
timestamp 1606821651
transform 1 0 14628 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1606821651
transform 1 0 14720 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1606821651
transform 1 0 14720 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_158
timestamp 1606821651
transform 1 0 15640 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156
timestamp 1606821651
transform 1 0 15456 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606821651
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1606821651
transform 1 0 15640 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1606821651
transform 1 0 15272 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_162
timestamp 1606821651
transform 1 0 16008 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_162
timestamp 1606821651
transform 1 0 16008 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1606821651
transform 1 0 16100 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_177
timestamp 1606821651
transform 1 0 17388 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_167
timestamp 1606821651
transform 1 0 16468 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_172
timestamp 1606821651
transform 1 0 16928 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1606821651
transform 1 0 16560 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1606821651
transform 1 0 17020 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_184
timestamp 1606821651
transform 1 0 18032 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_182
timestamp 1606821651
transform 1 0 17848 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606821651
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606821651
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1606821651
transform 1 0 17480 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1606821651
transform 1 0 18308 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1606821651
transform 1 0 19136 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1606821651
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_191
timestamp 1606821651
transform 1 0 18676 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_195
timestamp 1606821651
transform 1 0 19044 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_200
timestamp 1606821651
transform 1 0 19504 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606821651
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606821651
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606821651
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1606821651
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1606821651
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_212
timestamp 1606821651
transform 1 0 20608 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 1748 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606821651
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1606821651
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _044_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3404 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4140 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606821651
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_23
timestamp 1606821651
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_28
timestamp 1606821651
transform 1 0 3680 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_32
timestamp 1606821651
transform 1 0 4048 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_3_
timestamp 1606821651
transform 1 0 5796 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_49
timestamp 1606821651
transform 1 0 5612 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_60
timestamp 1606821651
transform 1 0 6624 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7084 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_2_64
timestamp 1606821651
transform 1 0 6992 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_81
timestamp 1606821651
transform 1 0 8556 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1606821651
transform 1 0 9108 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 9844 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606821651
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1606821651
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1606821651
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 11500 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_111
timestamp 1606821651
transform 1 0 11316 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1606821651
transform 1 0 14168 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13156 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_129
timestamp 1606821651
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_140
timestamp 1606821651
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1606821651
transform 1 0 16008 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 15272 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606821651
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_146
timestamp 1606821651
transform 1 0 14536 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_152
timestamp 1606821651
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_160
timestamp 1606821651
transform 1 0 15824 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1606821651
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1606821651
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1606821651
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1606821651
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606821651
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606821651
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1606821651
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1606821651
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 1748 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606821651
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1606821651
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 3404 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_23
timestamp 1606821651
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_41
timestamp 1606821651
transform 1 0 4876 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1606821651
transform 1 0 5152 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1606821651
transform 1 0 5612 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606821651
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_47
timestamp 1606821651
transform 1 0 5428 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_58
timestamp 1606821651
transform 1 0 6440 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_62
timestamp 1606821651
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_4_
timestamp 1606821651
transform 1 0 7084 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_5_
timestamp 1606821651
transform 1 0 8096 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_74
timestamp 1606821651
transform 1 0 7912 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1606821651
transform 1 0 10304 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1606821651
transform 1 0 9292 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_85
timestamp 1606821651
transform 1 0 8924 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_98
timestamp 1606821651
transform 1 0 10120 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_104
timestamp 1606821651
transform 1 0 10672 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 12420 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1606821651
transform 1 0 10856 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606821651
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_115
timestamp 1606821651
transform 1 0 11684 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1606821651
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1606821651
transform 1 0 14076 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_139
timestamp 1606821651
transform 1 0 13892 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1606821651
transform 1 0 15088 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_150
timestamp 1606821651
transform 1 0 14904 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_156
timestamp 1606821651
transform 1 0 15456 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606821651
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_168
timestamp 1606821651
transform 1 0 16560 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_180
timestamp 1606821651
transform 1 0 17664 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1606821651
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1606821651
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1606821651
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606821651
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1606821651
transform 1 0 2852 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1606821651
transform 1 0 1840 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606821651
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1606821651
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1606821651
transform 1 0 1748 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_17
timestamp 1606821651
transform 1 0 2668 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 4140 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606821651
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_28
timestamp 1606821651
transform 1 0 3680 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_32
timestamp 1606821651
transform 1 0 4048 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1606821651
transform 1 0 6164 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_4_49
timestamp 1606821651
transform 1 0 5612 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1606821651
transform 1 0 7360 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8372 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_64
timestamp 1606821651
transform 1 0 6992 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_77
timestamp 1606821651
transform 1 0 8188 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1606821651
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606821651
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_88
timestamp 1606821651
transform 1 0 9200 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_102
timestamp 1606821651
transform 1 0 10488 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 11224 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1606821651
transform 1 0 14168 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12880 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_126
timestamp 1606821651
transform 1 0 12696 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_137
timestamp 1606821651
transform 1 0 13708 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_141
timestamp 1606821651
transform 1 0 14076 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1606821651
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606821651
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 1606821651
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_163
timestamp 1606821651
transform 1 0 16100 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1606821651
transform 1 0 17848 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_175
timestamp 1606821651
transform 1 0 17204 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_181
timestamp 1606821651
transform 1 0 17756 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_186
timestamp 1606821651
transform 1 0 18216 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_198
timestamp 1606821651
transform 1 0 19320 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606821651
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606821651
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_210
timestamp 1606821651
transform 1 0 20424 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1606821651
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1606821651
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 2024 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606821651
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1606821651
transform 1 0 1380 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_9
timestamp 1606821651
transform 1 0 1932 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4600 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 3680 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_26
timestamp 1606821651
transform 1 0 3496 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_34
timestamp 1606821651
transform 1 0 4232 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6808 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606821651
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_54
timestamp 1606821651
transform 1 0 6072 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_60
timestamp 1606821651
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1606821651
transform 1 0 8464 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_78
timestamp 1606821651
transform 1 0 8280 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1606821651
transform 1 0 9844 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_5_89
timestamp 1606821651
transform 1 0 9292 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_104
timestamp 1606821651
transform 1 0 10672 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1606821651
transform 1 0 12512 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1606821651
transform 1 0 11316 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606821651
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_110
timestamp 1606821651
transform 1 0 11224 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1606821651
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_123
timestamp 1606821651
transform 1 0 12420 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1606821651
transform 1 0 13524 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1606821651
transform 1 0 14168 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_139
timestamp 1606821651
transform 1 0 13892 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1606821651
transform 1 0 15180 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_151
timestamp 1606821651
transform 1 0 14996 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_162
timestamp 1606821651
transform 1 0 16008 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 16928 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606821651
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_170
timestamp 1606821651
transform 1 0 16744 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_178
timestamp 1606821651
transform 1 0 17480 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_182
timestamp 1606821651
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1606821651
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1606821651
transform 1 0 19780 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_196
timestamp 1606821651
transform 1 0 19136 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_202
timestamp 1606821651
transform 1 0 19688 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_207
timestamp 1606821651
transform 1 0 20148 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606821651
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_219
timestamp 1606821651
transform 1 0 21252 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 1564 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1606821651
transform 1 0 2576 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1606821651
transform 1 0 1564 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606821651
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606821651
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1606821651
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_14
timestamp 1606821651
transform 1 0 2392 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1606821651
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4692 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1606821651
transform 1 0 4232 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1606821651
transform 1 0 3220 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606821651
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_25
timestamp 1606821651
transform 1 0 3404 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_32
timestamp 1606821651
transform 1 0 4048 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_38
timestamp 1606821651
transform 1 0 4600 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_21
timestamp 1606821651
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_32
timestamp 1606821651
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1606821651
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1606821651
transform 1 0 5704 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606821651
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 5244 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_55
timestamp 1606821651
transform 1 0 6164 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_43
timestamp 1606821651
transform 1 0 5060 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_48
timestamp 1606821651
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1606821651
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 7820 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 7268 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_6_83
timestamp 1606821651
transform 1 0 8740 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_71
timestamp 1606821651
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1606821651
transform 1 0 10028 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1606821651
transform 1 0 10580 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606821651
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1606821651
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_93
timestamp 1606821651
transform 1 0 9660 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_101
timestamp 1606821651
transform 1 0 10396 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_89
timestamp 1606821651
transform 1 0 9292 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 11592 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1606821651
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1606821651
transform 1 0 11316 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606821651
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_112
timestamp 1606821651
transform 1 0 11408 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_106
timestamp 1606821651
transform 1 0 10856 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_110
timestamp 1606821651
transform 1 0 11224 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1606821651
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1606821651
transform 1 0 13248 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 13524 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1606821651
transform 1 0 14168 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_130
timestamp 1606821651
transform 1 0 13064 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_135
timestamp 1606821651
transform 1 0 13524 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_141
timestamp 1606821651
transform 1 0 14076 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_132
timestamp 1606821651
transform 1 0 13248 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 15180 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 15272 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606821651
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1606821651
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_151
timestamp 1606821651
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1606821651
transform 1 0 16928 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606821651
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_170
timestamp 1606821651
transform 1 0 16744 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_181
timestamp 1606821651
transform 1 0 17756 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1606821651
transform 1 0 16652 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1606821651
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1606821651
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 18860 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_199
timestamp 1606821651
transform 1 0 19412 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1606821651
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1606821651
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606821651
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606821651
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606821651
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_211
timestamp 1606821651
transform 1 0 20516 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1606821651
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1606821651
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 1656 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606821651
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1606821651
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1606821651
transform 1 0 3312 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 4048 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606821651
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_22
timestamp 1606821651
transform 1 0 3128 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1606821651
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 5888 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_48
timestamp 1606821651
transform 1 0 5520 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8556 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1606821651
transform 1 0 7544 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_68
timestamp 1606821651
transform 1 0 7360 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_79
timestamp 1606821651
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9660 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606821651
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1606821651
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 11592 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_109
timestamp 1606821651
transform 1 0 11132 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_113
timestamp 1606821651
transform 1 0 11500 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1606821651
transform 1 0 13248 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_130
timestamp 1606821651
transform 1 0 13064 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_141
timestamp 1606821651
transform 1 0 14076 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1606821651
transform 1 0 14720 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1606821651
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606821651
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_147
timestamp 1606821651
transform 1 0 14628 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1606821651
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_163
timestamp 1606821651
transform 1 0 16100 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_175
timestamp 1606821651
transform 1 0 17204 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_187
timestamp 1606821651
transform 1 0 18308 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_199
timestamp 1606821651
transform 1 0 19412 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606821651
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606821651
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_211
timestamp 1606821651
transform 1 0 20516 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1606821651
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1606821651
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1606821651
transform 1 0 1932 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1606821651
transform 1 0 2944 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606821651
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1606821651
transform 1 0 1380 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_18
timestamp 1606821651
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1606821651
transform 1 0 4140 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 4600 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_29
timestamp 1606821651
transform 1 0 3772 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_36
timestamp 1606821651
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1606821651
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606821651
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 6256 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1606821651
transform 1 0 6072 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1606821651
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1606821651
transform 1 0 8096 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1606821651
transform 1 0 8556 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_71
timestamp 1606821651
transform 1 0 7636 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_75
timestamp 1606821651
transform 1 0 8004 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_79
timestamp 1606821651
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1606821651
transform 1 0 9568 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 10580 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_90
timestamp 1606821651
transform 1 0 9384 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_101
timestamp 1606821651
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1606821651
transform 1 0 11316 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606821651
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_106
timestamp 1606821651
transform 1 0 10856 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_110
timestamp 1606821651
transform 1 0 11224 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1606821651
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1606821651
transform 1 0 14444 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1606821651
transform 1 0 13432 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_132
timestamp 1606821651
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_143
timestamp 1606821651
transform 1 0 14260 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_154
timestamp 1606821651
transform 1 0 15272 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_166
timestamp 1606821651
transform 1 0 16376 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606821651
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_178
timestamp 1606821651
transform 1 0 17480 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1606821651
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1606821651
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1606821651
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1606821651
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606821651
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1606821651
transform 1 0 2116 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606821651
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1606821651
transform 1 0 1380 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_20
timestamp 1606821651
transform 1 0 2944 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1606821651
transform 1 0 3128 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1606821651
transform 1 0 4232 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606821651
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_25
timestamp 1606821651
transform 1 0 3404 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_32
timestamp 1606821651
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1606821651
transform 1 0 5336 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1606821651
transform 1 0 6348 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_10_43
timestamp 1606821651
transform 1 0 5060 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_55
timestamp 1606821651
transform 1 0 6164 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8556 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1606821651
transform 1 0 7360 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_66
timestamp 1606821651
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_77
timestamp 1606821651
transform 1 0 8188 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 9660 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606821651
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1606821651
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 11684 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_10_109
timestamp 1606821651
transform 1 0 11132 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13340 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_131
timestamp 1606821651
transform 1 0 13156 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606821651
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_149
timestamp 1606821651
transform 1 0 14812 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1606821651
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1606821651
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_178
timestamp 1606821651
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_190
timestamp 1606821651
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_202
timestamp 1606821651
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606821651
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606821651
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1606821651
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1606821651
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 1380 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606821651
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_19
timestamp 1606821651
transform 1 0 2852 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1606821651
transform 1 0 4048 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1606821651
transform 1 0 3036 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_30
timestamp 1606821651
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_41
timestamp 1606821651
transform 1 0 4876 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 5060 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606821651
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1606821651
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_62
timestamp 1606821651
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6992 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 8648 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_80
timestamp 1606821651
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10672 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 10304 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_98
timestamp 1606821651
transform 1 0 10120 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_103
timestamp 1606821651
transform 1 0 10580 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1606821651
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606821651
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1606821651
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1606821651
transform 1 0 13432 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1606821651
transform 1 0 14444 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_132
timestamp 1606821651
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_143
timestamp 1606821651
transform 1 0 14260 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_154
timestamp 1606821651
transform 1 0 15272 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_166
timestamp 1606821651
transform 1 0 16376 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606821651
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_178
timestamp 1606821651
transform 1 0 17480 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1606821651
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1606821651
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1606821651
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1606821651
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606821651
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 2024 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606821651
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1606821651
transform 1 0 1380 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_9
timestamp 1606821651
transform 1 0 1932 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1606821651
transform 1 0 4416 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606821651
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 3680 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1606821651
transform 1 0 3496 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_32
timestamp 1606821651
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1606821651
transform 1 0 5428 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1606821651
transform 1 0 6440 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_45
timestamp 1606821651
transform 1 0 5244 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_56
timestamp 1606821651
transform 1 0 6256 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1606821651
transform 1 0 7452 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1606821651
transform 1 0 8464 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_67
timestamp 1606821651
transform 1 0 7268 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_78
timestamp 1606821651
transform 1 0 8280 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1606821651
transform 1 0 10672 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_6_
timestamp 1606821651
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606821651
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_89
timestamp 1606821651
transform 1 0 9292 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_102
timestamp 1606821651
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_3_
timestamp 1606821651
transform 1 0 11684 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_113
timestamp 1606821651
transform 1 0 11500 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_124
timestamp 1606821651
transform 1 0 12512 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1606821651
transform 1 0 12696 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1606821651
transform 1 0 13708 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_135
timestamp 1606821651
transform 1 0 13524 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606821651
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_146
timestamp 1606821651
transform 1 0 14536 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1606821651
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1606821651
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1606821651
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1606821651
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1606821651
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1606821651
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606821651
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606821651
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1606821651
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1606821651
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1606821651
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1606821651
transform 1 0 1380 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606821651
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606821651
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1564 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1606821651
transform 1 0 1932 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_11
timestamp 1606821651
transform 1 0 2116 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_18
timestamp 1606821651
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1606821651
transform 1 0 2944 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 2300 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1606821651
transform 1 0 3956 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1606821651
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606821651
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_29
timestamp 1606821651
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_40
timestamp 1606821651
transform 1 0 4784 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1606821651
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_41
timestamp 1606821651
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6348 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 5060 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1606821651
transform 1 0 5060 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_3_
timestamp 1606821651
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606821651
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1606821651
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_52
timestamp 1606821651
transform 1 0 5888 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_56
timestamp 1606821651
transform 1 0 6256 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8096 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8188 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 7820 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_71
timestamp 1606821651
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_73
timestamp 1606821651
transform 1 0 7820 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_93
timestamp 1606821651
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_86
timestamp 1606821651
transform 1 0 9016 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_90
timestamp 1606821651
transform 1 0 9384 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_85
timestamp 1606821651
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606821651
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1606821651
transform 1 0 9568 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1606821651
transform 1 0 9108 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_101
timestamp 1606821651
transform 1 0 10396 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_101
timestamp 1606821651
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 9844 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_3_
timestamp 1606821651
transform 1 0 10580 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1606821651
transform 1 0 10120 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 10580 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1606821651
transform 1 0 12420 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1606821651
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1606821651
transform 1 0 11408 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606821651
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1606821651
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_119
timestamp 1606821651
transform 1 0 12052 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1606821651
transform 1 0 13248 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1606821651
transform 1 0 14076 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1606821651
transform 1 0 13248 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1606821651
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606821651
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_150
timestamp 1606821651
transform 1 0 14904 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_162
timestamp 1606821651
transform 1 0 16008 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1606821651
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_166
timestamp 1606821651
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606821651
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_174
timestamp 1606821651
transform 1 0 17112 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1606821651
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1606821651
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_178
timestamp 1606821651
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1606821651
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1606821651
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_190
timestamp 1606821651
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_202
timestamp 1606821651
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606821651
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606821651
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606821651
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1606821651
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1606821651
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 2024 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606821651
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1606821651
transform 1 0 1380 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_9
timestamp 1606821651
transform 1 0 1932 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1606821651
transform 1 0 3680 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4416 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_26
timestamp 1606821651
transform 1 0 3496 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_31
timestamp 1606821651
transform 1 0 3956 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_35
timestamp 1606821651
transform 1 0 4324 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1606821651
transform 1 0 6072 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1606821651
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606821651
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_52
timestamp 1606821651
transform 1 0 5888 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1606821651
transform 1 0 6348 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7544 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_65
timestamp 1606821651
transform 1 0 7084 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_69
timestamp 1606821651
transform 1 0 7452 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1606821651
transform 1 0 9200 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9660 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_86
timestamp 1606821651
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_91
timestamp 1606821651
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1606821651
transform 1 0 11960 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1606821651
transform 1 0 11132 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606821651
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1606821651
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_123
timestamp 1606821651
transform 1 0 12420 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1606821651
transform 1 0 14444 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1606821651
transform 1 0 13432 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1606821651
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_131
timestamp 1606821651
transform 1 0 13156 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_143
timestamp 1606821651
transform 1 0 14260 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_148
timestamp 1606821651
transform 1 0 14720 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_160
timestamp 1606821651
transform 1 0 15824 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606821651
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_172
timestamp 1606821651
transform 1 0 16928 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_180
timestamp 1606821651
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1606821651
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1606821651
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1606821651
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606821651
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 1380 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606821651
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_19
timestamp 1606821651
transform 1 0 2852 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1606821651
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 4784 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 3036 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606821651
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1606821651
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_35
timestamp 1606821651
transform 1 0 4324 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_39
timestamp 1606821651
transform 1 0 4692 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_56
timestamp 1606821651
transform 1 0 6256 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_62
timestamp 1606821651
transform 1 0 6808 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 7912 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l3_in_0_
timestamp 1606821651
transform 1 0 6900 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_72
timestamp 1606821651
transform 1 0 7728 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 9660 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606821651
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1606821651
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 11408 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_16_109
timestamp 1606821651
transform 1 0 11132 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1606821651
transform 1 0 13064 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1606821651
transform 1 0 14076 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_128
timestamp 1606821651
transform 1 0 12880 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_139
timestamp 1606821651
transform 1 0 13892 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606821651
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_150
timestamp 1606821651
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1606821651
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_166
timestamp 1606821651
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_178
timestamp 1606821651
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_190
timestamp 1606821651
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_202
timestamp 1606821651
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606821651
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606821651
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1606821651
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1606821651
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 2300 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1564 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606821651
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1606821651
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_11
timestamp 1606821651
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1606821651
transform 1 0 3956 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_29
timestamp 1606821651
transform 1 0 3772 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_40
timestamp 1606821651
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1606821651
transform 1 0 4968 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1606821651
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606821651
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1606821651
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1606821651
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 8372 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_17_71
timestamp 1606821651
transform 1 0 7636 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_99
timestamp 1606821651
transform 1 0 10212 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 12420 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10856 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606821651
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_105
timestamp 1606821651
transform 1 0 10764 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_115
timestamp 1606821651
transform 1 0 11684 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1606821651
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1606821651
transform 1 0 14076 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_139
timestamp 1606821651
transform 1 0 13892 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_150
timestamp 1606821651
transform 1 0 14904 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_162
timestamp 1606821651
transform 1 0 16008 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 16652 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1606821651
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_168
timestamp 1606821651
transform 1 0 16560 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_175
timestamp 1606821651
transform 1 0 17204 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1606821651
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1606821651
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1606821651
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606821651
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1606821651
transform 1 0 2760 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1606821651
transform 1 0 1748 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606821651
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1606821651
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_16
timestamp 1606821651
transform 1 0 2576 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1606821651
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1606821651
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1606821651
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_41
timestamp 1606821651
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1606821651
transform 1 0 5060 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 5888 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_47
timestamp 1606821651
transform 1 0 5428 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_51
timestamp 1606821651
transform 1 0 5796 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_1_
timestamp 1606821651
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_18_68
timestamp 1606821651
transform 1 0 7360 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_74
timestamp 1606821651
transform 1 0 7912 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1606821651
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10212 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1606821651
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_84
timestamp 1606821651
transform 1 0 8832 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_96
timestamp 1606821651
transform 1 0 9936 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1606821651
transform 1 0 11868 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_115
timestamp 1606821651
transform 1 0 11684 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13432 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_18_126
timestamp 1606821651
transform 1 0 12696 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1606821651
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_150
timestamp 1606821651
transform 1 0 14904 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1606821651
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_166
timestamp 1606821651
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1606821651
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_190
timestamp 1606821651
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_202
timestamp 1606821651
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606821651
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1606821651
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1606821651
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1606821651
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_9
timestamp 1606821651
transform 1 0 1932 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1606821651
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606821651
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606821651
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1380 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1606821651
transform 1 0 1748 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_16
timestamp 1606821651
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1606821651
transform 1 0 2116 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1606821651
transform 1 0 2760 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_20
timestamp 1606821651
transform 1 0 2944 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1606821651
transform 1 0 3128 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1606821651
transform 1 0 3772 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4048 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4692 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1606821651
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_27
timestamp 1606821651
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_33
timestamp 1606821651
transform 1 0 4140 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_26
timestamp 1606821651
transform 1 0 3496 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_30
timestamp 1606821651
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 5704 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1606821651
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1606821651
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_55
timestamp 1606821651
transform 1 0 6164 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_48
timestamp 1606821651
transform 1 0 5520 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 7360 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7912 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_19_71
timestamp 1606821651
transform 1 0 7636 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_66
timestamp 1606821651
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_84
timestamp 1606821651
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_90
timestamp 1606821651
transform 1 0 9384 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1606821651
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1606821651
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 9016 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l3_in_0_
timestamp 1606821651
transform 1 0 9660 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_102
timestamp 1606821651
transform 1 0 10488 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_102
timestamp 1606821651
transform 1 0 10488 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_1_
timestamp 1606821651
transform 1 0 10580 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 10672 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1606821651
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1606821651
transform 1 0 11592 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1606821651
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1606821651
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_112
timestamp 1606821651
transform 1 0 11408 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_123
timestamp 1606821651
transform 1 0 12420 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 12880 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12880 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1606821651
transform 1 0 13892 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_126
timestamp 1606821651
transform 1 0 12696 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_144
timestamp 1606821651
transform 1 0 14352 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_127
timestamp 1606821651
transform 1 0 12788 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_137
timestamp 1606821651
transform 1 0 13708 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1606821651
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_148
timestamp 1606821651
transform 1 0 14720 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_155
timestamp 1606821651
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1606821651
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1606821651
transform 1 0 14536 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_5_
timestamp 1606821651
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_163
timestamp 1606821651
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1606821651
transform 1 0 15548 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_6_
timestamp 1606821651
transform 1 0 16284 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_19_166
timestamp 1606821651
transform 1 0 16376 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1606821651
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_178
timestamp 1606821651
transform 1 0 17480 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_182
timestamp 1606821651
transform 1 0 17848 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1606821651
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_174
timestamp 1606821651
transform 1 0 17112 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_186
timestamp 1606821651
transform 1 0 18216 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1606821651
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1606821651
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_198
timestamp 1606821651
transform 1 0 19320 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606821651
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606821651
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1606821651
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_210
timestamp 1606821651
transform 1 0 20424 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1606821651
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1606821651
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 2484 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1606821651
transform 1 0 1472 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606821651
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 1606821651
transform 1 0 1380 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_13
timestamp 1606821651
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1606821651
transform 1 0 4048 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1606821651
transform 1 0 4876 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_31
timestamp 1606821651
transform 1 0 3956 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1606821651
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1606821651
transform 1 0 5704 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1606821651
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1606821651
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8556 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1606821651
transform 1 0 7544 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_65
timestamp 1606821651
transform 1 0 7084 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_69
timestamp 1606821651
transform 1 0 7452 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_79
timestamp 1606821651
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1606821651
transform 1 0 9384 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1606821651
transform 1 0 10212 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 12420 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1606821651
transform 1 0 11040 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1606821651
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 12052 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_117
timestamp 1606821651
transform 1 0 11868 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_139
timestamp 1606821651
transform 1 0 13892 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 14720 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_21_147
timestamp 1606821651
transform 1 0 14628 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_164
timestamp 1606821651
transform 1 0 16192 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1606821651
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_176
timestamp 1606821651
transform 1 0 17296 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp 1606821651
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1606821651
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1606821651
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1606821651
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606821651
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1606821651
transform 1 0 1472 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 2024 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606821651
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1606821651
transform 1 0 1380 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_8
timestamp 1606821651
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1606821651
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1606821651
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_26
timestamp 1606821651
transform 1 0 3496 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_30
timestamp 1606821651
transform 1 0 3864 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_32
timestamp 1606821651
transform 1 0 4048 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_40
timestamp 1606821651
transform 1 0 4784 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1606821651
transform 1 0 5060 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1606821651
transform 1 0 6348 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 5888 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_55
timestamp 1606821651
transform 1 0 6164 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1606821651
transform 1 0 7452 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1606821651
transform 1 0 8280 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_22_66
timestamp 1606821651
transform 1 0 7176 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1606821651
transform 1 0 10672 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1606821651
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 9292 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_87
timestamp 1606821651
transform 1 0 9108 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_102
timestamp 1606821651
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 11132 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_107
timestamp 1606821651
transform 1 0 10948 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_125
timestamp 1606821651
transform 1 0 12604 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 12788 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_22_143
timestamp 1606821651
transform 1 0 14260 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_4_
timestamp 1606821651
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1606821651
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1606821651
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_163
timestamp 1606821651
transform 1 0 16100 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_175
timestamp 1606821651
transform 1 0 17204 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_187
timestamp 1606821651
transform 1 0 18308 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_199
timestamp 1606821651
transform 1 0 19412 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606821651
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1606821651
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_211
timestamp 1606821651
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1606821651
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1606821651
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1472 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1606821651
transform 1 0 2208 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606821651
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_3
timestamp 1606821651
transform 1 0 1380 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_10
timestamp 1606821651
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1606821651
transform 1 0 3220 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 3956 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_21
timestamp 1606821651
transform 1 0 3036 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_27
timestamp 1606821651
transform 1 0 3588 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6808 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5704 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1606821651
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_47
timestamp 1606821651
transform 1 0 5428 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1606821651
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1606821651
transform 1 0 8464 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_78
timestamp 1606821651
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1606821651
transform 1 0 9476 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10304 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 10028 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_89
timestamp 1606821651
transform 1 0 9292 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_94
timestamp 1606821651
transform 1 0 9752 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1606821651
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1606821651
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_116
timestamp 1606821651
transform 1 0 11776 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12788 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1606821651
transform 1 0 13984 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1606821651
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_126
timestamp 1606821651
transform 1 0 12696 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_136
timestamp 1606821651
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1606821651
transform 1 0 14996 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_149
timestamp 1606821651
transform 1 0 14812 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_160
timestamp 1606821651
transform 1 0 15824 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1606821651
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_172
timestamp 1606821651
transform 1 0 16928 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_180
timestamp 1606821651
transform 1 0 17664 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1606821651
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1606821651
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1606821651
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606821651
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1606821651
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1606821651
transform 1 0 2944 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1606821651
transform 1 0 1932 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606821651
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_7
timestamp 1606821651
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_18
timestamp 1606821651
transform 1 0 2760 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1606821651
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1606821651
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_41
timestamp 1606821651
transform 1 0 4876 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1606821651
transform 1 0 5060 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1606821651
transform 1 0 6072 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_52
timestamp 1606821651
transform 1 0 5888 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1606821651
transform 1 0 7084 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 7912 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 7544 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_63
timestamp 1606821651
transform 1 0 6900 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_68
timestamp 1606821651
transform 1 0 7360 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_73
timestamp 1606821651
transform 1 0 7820 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 9660 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1606821651
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1606821651
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 12604 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l3_in_0_
timestamp 1606821651
transform 1 0 11592 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_109
timestamp 1606821651
transform 1 0 11132 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_113
timestamp 1606821651
transform 1 0 11500 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_123
timestamp 1606821651
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1606821651
transform 1 0 14260 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1606821651
transform 1 0 14076 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1606821651
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_146
timestamp 1606821651
transform 1 0 14536 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1606821651
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1606821651
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1606821651
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1606821651
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1606821651
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1606821651
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606821651
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1606821651
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1606821651
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1606821651
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1606821651
transform 1 0 2300 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1606821651
transform 1 0 1748 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1606821651
transform 1 0 2944 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606821651
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1606821651
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_11
timestamp 1606821651
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_17
timestamp 1606821651
transform 1 0 2668 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 3956 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_29
timestamp 1606821651
transform 1 0 3772 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_40
timestamp 1606821651
transform 1 0 4784 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1606821651
transform 1 0 6164 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1606821651
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1606821651
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1606821651
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_53
timestamp 1606821651
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1606821651
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1606821651
transform 1 0 7912 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_25_71
timestamp 1606821651
transform 1 0 7636 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_83
timestamp 1606821651
transform 1 0 8740 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1606821651
transform 1 0 9108 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1606821651
transform 1 0 10120 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_96
timestamp 1606821651
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_1_
timestamp 1606821651
transform 1 0 12604 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1606821651
transform 1 0 11132 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1606821651
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_107
timestamp 1606821651
transform 1 0 10948 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_118
timestamp 1606821651
transform 1 0 11960 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_123
timestamp 1606821651
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 13616 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_134
timestamp 1606821651
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_142
timestamp 1606821651
transform 1 0 14168 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_154
timestamp 1606821651
transform 1 0 15272 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_166
timestamp 1606821651
transform 1 0 16376 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1606821651
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_178
timestamp 1606821651
transform 1 0 17480 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1606821651
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1606821651
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1606821651
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1606821651
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606821651
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_9
timestamp 1606821651
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1606821651
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1606821651
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606821651
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606821651
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1606821651
transform 1 0 1656 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1606821651
transform 1 0 1564 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_17
timestamp 1606821651
transform 1 0 2668 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_18
timestamp 1606821651
transform 1 0 2760 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_10
timestamp 1606821651
transform 1 0 2024 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2116 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2208 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1606821651
transform 1 0 2944 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1606821651
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4600 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 3220 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1606821651
transform 1 0 4876 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1606821651
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1606821651
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_36
timestamp 1606821651
transform 1 0 4416 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_39
timestamp 1606821651
transform 1 0 4692 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1606821651
transform 1 0 5888 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6256 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6808 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1606821651
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 6440 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_54
timestamp 1606821651
transform 1 0 6072 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_50
timestamp 1606821651
transform 1 0 5704 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_56
timestamp 1606821651
transform 1 0 6256 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 8648 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8096 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_26_72
timestamp 1606821651
transform 1 0 7728 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_78
timestamp 1606821651
transform 1 0 8280 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1606821651
transform 1 0 9108 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10304 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9936 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1606821651
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1606821651
transform 1 0 8924 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_90
timestamp 1606821651
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_93
timestamp 1606821651
transform 1 0 9660 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_98
timestamp 1606821651
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_105
timestamp 1606821651
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_1_
timestamp 1606821651
transform 1 0 10948 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_121
timestamp 1606821651
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_116
timestamp 1606821651
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_122
timestamp 1606821651
transform 1 0 12328 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_116
timestamp 1606821651
transform 1 0 11776 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 11960 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1606821651
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1606821651
transform 1 0 11960 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 12604 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1606821651
transform 1 0 13984 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1606821651
transform 1 0 13432 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 14260 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1606821651
transform 1 0 14076 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_132
timestamp 1606821651
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_138
timestamp 1606821651
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_144
timestamp 1606821651
transform 1 0 14352 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1606821651
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_149
timestamp 1606821651
transform 1 0 14812 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1606821651
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1606821651
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_156
timestamp 1606821651
transform 1 0 15456 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1606821651
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1606821651
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_168
timestamp 1606821651
transform 1 0 16560 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_180
timestamp 1606821651
transform 1 0 17664 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1606821651
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1606821651
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_202
timestamp 1606821651
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1606821651
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1606821651
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606821651
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606821651
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1606821651
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1606821651
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1606821651
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1472 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1606821651
transform 1 0 2944 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2208 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606821651
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_3
timestamp 1606821651
transform 1 0 1380 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_10
timestamp 1606821651
transform 1 0 2024 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_18
timestamp 1606821651
transform 1 0 2760 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4048 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1606821651
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1606821651
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_1_
timestamp 1606821651
transform 1 0 6440 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 5704 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_48
timestamp 1606821651
transform 1 0 5520 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_56
timestamp 1606821651
transform 1 0 6256 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7452 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_67
timestamp 1606821651
transform 1 0 7268 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1606821651
transform 1 0 9108 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_1_
timestamp 1606821651
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1606821651
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1606821651
transform 1 0 8924 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_90
timestamp 1606821651
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_102
timestamp 1606821651
transform 1 0 10488 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10856 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 12512 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_122
timestamp 1606821651
transform 1 0 12328 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1606821651
transform 1 0 14260 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_140
timestamp 1606821651
transform 1 0 13984 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1606821651
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_147
timestamp 1606821651
transform 1 0 14628 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1606821651
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1606821651
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1606821651
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1606821651
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1606821651
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606821651
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1606821651
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1606821651
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1606821651
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1606821651
transform 1 0 1472 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2024 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2760 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606821651
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_3
timestamp 1606821651
transform 1 0 1380 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_8
timestamp 1606821651
transform 1 0 1840 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_16
timestamp 1606821651
transform 1 0 2576 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 3496 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_24
timestamp 1606821651
transform 1 0 3312 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1606821651
transform 1 0 6164 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1606821651
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1606821651
transform 1 0 5152 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1606821651
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_42
timestamp 1606821651
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_53
timestamp 1606821651
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1606821651
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1606821651
transform 1 0 7912 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_29_71
timestamp 1606821651
transform 1 0 7636 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_83
timestamp 1606821651
transform 1 0 8740 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1606821651
transform 1 0 9016 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 10028 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_95
timestamp 1606821651
transform 1 0 9844 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_103
timestamp 1606821651
transform 1 0 10580 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1606821651
transform 1 0 11868 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10856 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1606821651
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_115
timestamp 1606821651
transform 1 0 11684 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1606821651
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1606821651
transform 1 0 14444 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1606821651
transform 1 0 13432 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_132
timestamp 1606821651
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_143
timestamp 1606821651
transform 1 0 14260 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_149
timestamp 1606821651
transform 1 0 14812 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_161
timestamp 1606821651
transform 1 0 15916 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1606821651
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_173
timestamp 1606821651
transform 1 0 17020 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1606821651
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1606821651
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1606821651
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1606821651
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606821651
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1606821651
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1606821651
transform 1 0 1932 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1606821651
transform 1 0 2944 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606821651
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_7
timestamp 1606821651
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_18
timestamp 1606821651
transform 1 0 2760 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1606821651
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1606821651
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1606821651
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_41
timestamp 1606821651
transform 1 0 4876 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1606821651
transform 1 0 6808 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 5152 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_60
timestamp 1606821651
transform 1 0 6624 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7452 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_30_66
timestamp 1606821651
transform 1 0 7176 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1606821651
transform 1 0 9108 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1606821651
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1606821651
transform 1 0 8924 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1606821651
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_102
timestamp 1606821651
transform 1 0 10488 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 11960 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10948 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_30_106
timestamp 1606821651
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_116
timestamp 1606821651
transform 1 0 11776 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 13616 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 14352 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_134
timestamp 1606821651
transform 1 0 13432 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_142
timestamp 1606821651
transform 1 0 14168 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 15272 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1606821651
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_150
timestamp 1606821651
transform 1 0 14904 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_160
timestamp 1606821651
transform 1 0 15824 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_172
timestamp 1606821651
transform 1 0 16928 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_184
timestamp 1606821651
transform 1 0 18032 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 18492 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_188
timestamp 1606821651
transform 1 0 18400 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_195
timestamp 1606821651
transform 1 0 19044 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_207
timestamp 1606821651
transform 1 0 20148 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606821651
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1606821651
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_213
timestamp 1606821651
transform 1 0 20700 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1606821651
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1606821651
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1606821651
transform 1 0 1564 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 2944 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2116 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606821651
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1606821651
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_9
timestamp 1606821651
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_17
timestamp 1606821651
transform 1 0 2668 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1606821651
transform 1 0 4600 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_36
timestamp 1606821651
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_41
timestamp 1606821651
transform 1 0 4876 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 5060 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1606821651
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1606821651
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1606821651
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 8004 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_31_71
timestamp 1606821651
transform 1 0 7636 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9660 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_91
timestamp 1606821651
transform 1 0 9476 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 12420 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1606821651
transform 1 0 11316 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1606821651
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_109
timestamp 1606821651
transform 1 0 11132 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_120
timestamp 1606821651
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1606821651
transform 1 0 14076 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_139
timestamp 1606821651
transform 1 0 13892 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_145
timestamp 1606821651
transform 1 0 14444 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1606821651
transform 1 0 16008 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 14720 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_160
timestamp 1606821651
transform 1 0 15824 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1606821651
transform 1 0 16376 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1606821651
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1606821651
transform 1 0 17112 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1606821651
transform 1 0 16560 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1606821651
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_172
timestamp 1606821651
transform 1 0 16928 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_178
timestamp 1606821651
transform 1 0 17480 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_182
timestamp 1606821651
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1606821651
transform 1 0 19412 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1606821651
transform 1 0 18584 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_188
timestamp 1606821651
transform 1 0 18400 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_194
timestamp 1606821651
transform 1 0 18952 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_198
timestamp 1606821651
transform 1 0 19320 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_203
timestamp 1606821651
transform 1 0 19780 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606821651
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1606821651
transform 1 0 20884 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_219
timestamp 1606821651
transform 1 0 21252 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1606821651
transform 1 0 1656 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2208 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606821651
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_3
timestamp 1606821651
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_10
timestamp 1606821651
transform 1 0 2024 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_18
timestamp 1606821651
transform 1 0 2760 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 3036 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1606821651
transform 1 0 4048 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1606821651
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1606821651
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_41
timestamp 1606821651
transform 1 0 4876 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 5152 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1606821651
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_60
timestamp 1606821651
transform 1 0 6624 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1606821651
transform 1 0 6900 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7360 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_32_66
timestamp 1606821651
transform 1 0 7176 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1606821651
transform 1 0 9016 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1606821651
transform 1 0 9752 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10304 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1606821651
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_84
timestamp 1606821651
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_90
timestamp 1606821651
transform 1 0 9384 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_98
timestamp 1606821651
transform 1 0 10120 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1606821651
transform 1 0 12052 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1606821651
transform 1 0 12604 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 11316 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1606821651
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_109
timestamp 1606821651
transform 1 0 11132 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_117
timestamp 1606821651
transform 1 0 11868 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_122
timestamp 1606821651
transform 1 0 12328 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1606821651
transform 1 0 14168 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1606821651
transform 1 0 13156 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_129
timestamp 1606821651
transform 1 0 12972 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_135
timestamp 1606821651
transform 1 0 13524 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_141
timestamp 1606821651
transform 1 0 14076 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1606821651
transform 1 0 16008 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1606821651
transform 1 0 15456 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1606821651
transform 1 0 14720 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1606821651
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_146
timestamp 1606821651
transform 1 0 14536 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_152
timestamp 1606821651
transform 1 0 15088 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_160
timestamp 1606821651
transform 1 0 15824 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_166
timestamp 1606821651
transform 1 0 16376 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1606821651
transform 1 0 17020 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1606821651
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_172
timestamp 1606821651
transform 1 0 16928 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_177
timestamp 1606821651
transform 1 0 17388 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_185
timestamp 1606821651
transform 1 0 18124 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_187
timestamp 1606821651
transform 1 0 18308 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_199
timestamp 1606821651
transform 1 0 19412 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606821651
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1606821651
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_211
timestamp 1606821651
transform 1 0 20516 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1606821651
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
<< labels >>
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_42_
port 0 nsew default input
rlabel metal2 s 662 0 718 480 6 bottom_left_grid_pin_43_
port 1 nsew default input
rlabel metal2 s 1122 0 1178 480 6 bottom_left_grid_pin_44_
port 2 nsew default input
rlabel metal2 s 1582 0 1638 480 6 bottom_left_grid_pin_45_
port 3 nsew default input
rlabel metal2 s 2042 0 2098 480 6 bottom_left_grid_pin_46_
port 4 nsew default input
rlabel metal2 s 2502 0 2558 480 6 bottom_left_grid_pin_47_
port 5 nsew default input
rlabel metal2 s 2962 0 3018 480 6 bottom_left_grid_pin_48_
port 6 nsew default input
rlabel metal2 s 3422 0 3478 480 6 bottom_left_grid_pin_49_
port 7 nsew default input
rlabel metal2 s 22466 0 22522 480 6 bottom_right_grid_pin_1_
port 8 nsew default input
rlabel metal3 s 22320 5720 22800 5840 6 ccff_head
port 9 nsew default input
rlabel metal3 s 22320 17144 22800 17264 6 ccff_tail
port 10 nsew default tristate
rlabel metal3 s 0 3952 480 4072 6 chanx_left_in[0]
port 11 nsew default input
rlabel metal3 s 0 8712 480 8832 6 chanx_left_in[10]
port 12 nsew default input
rlabel metal3 s 0 9120 480 9240 6 chanx_left_in[11]
port 13 nsew default input
rlabel metal3 s 0 9664 480 9784 6 chanx_left_in[12]
port 14 nsew default input
rlabel metal3 s 0 10072 480 10192 6 chanx_left_in[13]
port 15 nsew default input
rlabel metal3 s 0 10616 480 10736 6 chanx_left_in[14]
port 16 nsew default input
rlabel metal3 s 0 11024 480 11144 6 chanx_left_in[15]
port 17 nsew default input
rlabel metal3 s 0 11568 480 11688 6 chanx_left_in[16]
port 18 nsew default input
rlabel metal3 s 0 11976 480 12096 6 chanx_left_in[17]
port 19 nsew default input
rlabel metal3 s 0 12520 480 12640 6 chanx_left_in[18]
port 20 nsew default input
rlabel metal3 s 0 12928 480 13048 6 chanx_left_in[19]
port 21 nsew default input
rlabel metal3 s 0 4360 480 4480 6 chanx_left_in[1]
port 22 nsew default input
rlabel metal3 s 0 4904 480 5024 6 chanx_left_in[2]
port 23 nsew default input
rlabel metal3 s 0 5312 480 5432 6 chanx_left_in[3]
port 24 nsew default input
rlabel metal3 s 0 5856 480 5976 6 chanx_left_in[4]
port 25 nsew default input
rlabel metal3 s 0 6264 480 6384 6 chanx_left_in[5]
port 26 nsew default input
rlabel metal3 s 0 6808 480 6928 6 chanx_left_in[6]
port 27 nsew default input
rlabel metal3 s 0 7216 480 7336 6 chanx_left_in[7]
port 28 nsew default input
rlabel metal3 s 0 7760 480 7880 6 chanx_left_in[8]
port 29 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_in[9]
port 30 nsew default input
rlabel metal3 s 0 13472 480 13592 6 chanx_left_out[0]
port 31 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 chanx_left_out[10]
port 32 nsew default tristate
rlabel metal3 s 0 18640 480 18760 6 chanx_left_out[11]
port 33 nsew default tristate
rlabel metal3 s 0 19184 480 19304 6 chanx_left_out[12]
port 34 nsew default tristate
rlabel metal3 s 0 19592 480 19712 6 chanx_left_out[13]
port 35 nsew default tristate
rlabel metal3 s 0 20136 480 20256 6 chanx_left_out[14]
port 36 nsew default tristate
rlabel metal3 s 0 20544 480 20664 6 chanx_left_out[15]
port 37 nsew default tristate
rlabel metal3 s 0 21088 480 21208 6 chanx_left_out[16]
port 38 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[17]
port 39 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 chanx_left_out[18]
port 40 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chanx_left_out[19]
port 41 nsew default tristate
rlabel metal3 s 0 13880 480 14000 6 chanx_left_out[1]
port 42 nsew default tristate
rlabel metal3 s 0 14424 480 14544 6 chanx_left_out[2]
port 43 nsew default tristate
rlabel metal3 s 0 14832 480 14952 6 chanx_left_out[3]
port 44 nsew default tristate
rlabel metal3 s 0 15376 480 15496 6 chanx_left_out[4]
port 45 nsew default tristate
rlabel metal3 s 0 15784 480 15904 6 chanx_left_out[5]
port 46 nsew default tristate
rlabel metal3 s 0 16328 480 16448 6 chanx_left_out[6]
port 47 nsew default tristate
rlabel metal3 s 0 16736 480 16856 6 chanx_left_out[7]
port 48 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[8]
port 49 nsew default tristate
rlabel metal3 s 0 17688 480 17808 6 chanx_left_out[9]
port 50 nsew default tristate
rlabel metal2 s 3882 0 3938 480 6 chany_bottom_in[0]
port 51 nsew default input
rlabel metal2 s 8574 0 8630 480 6 chany_bottom_in[10]
port 52 nsew default input
rlabel metal2 s 9034 0 9090 480 6 chany_bottom_in[11]
port 53 nsew default input
rlabel metal2 s 9494 0 9550 480 6 chany_bottom_in[12]
port 54 nsew default input
rlabel metal2 s 9954 0 10010 480 6 chany_bottom_in[13]
port 55 nsew default input
rlabel metal2 s 10414 0 10470 480 6 chany_bottom_in[14]
port 56 nsew default input
rlabel metal2 s 10874 0 10930 480 6 chany_bottom_in[15]
port 57 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[16]
port 58 nsew default input
rlabel metal2 s 11794 0 11850 480 6 chany_bottom_in[17]
port 59 nsew default input
rlabel metal2 s 12254 0 12310 480 6 chany_bottom_in[18]
port 60 nsew default input
rlabel metal2 s 12714 0 12770 480 6 chany_bottom_in[19]
port 61 nsew default input
rlabel metal2 s 4342 0 4398 480 6 chany_bottom_in[1]
port 62 nsew default input
rlabel metal2 s 4802 0 4858 480 6 chany_bottom_in[2]
port 63 nsew default input
rlabel metal2 s 5262 0 5318 480 6 chany_bottom_in[3]
port 64 nsew default input
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_in[4]
port 65 nsew default input
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_in[5]
port 66 nsew default input
rlabel metal2 s 6642 0 6698 480 6 chany_bottom_in[6]
port 67 nsew default input
rlabel metal2 s 7102 0 7158 480 6 chany_bottom_in[7]
port 68 nsew default input
rlabel metal2 s 7562 0 7618 480 6 chany_bottom_in[8]
port 69 nsew default input
rlabel metal2 s 8114 0 8170 480 6 chany_bottom_in[9]
port 70 nsew default input
rlabel metal2 s 13174 0 13230 480 6 chany_bottom_out[0]
port 71 nsew default tristate
rlabel metal2 s 17866 0 17922 480 6 chany_bottom_out[10]
port 72 nsew default tristate
rlabel metal2 s 18326 0 18382 480 6 chany_bottom_out[11]
port 73 nsew default tristate
rlabel metal2 s 18786 0 18842 480 6 chany_bottom_out[12]
port 74 nsew default tristate
rlabel metal2 s 19246 0 19302 480 6 chany_bottom_out[13]
port 75 nsew default tristate
rlabel metal2 s 19706 0 19762 480 6 chany_bottom_out[14]
port 76 nsew default tristate
rlabel metal2 s 20166 0 20222 480 6 chany_bottom_out[15]
port 77 nsew default tristate
rlabel metal2 s 20626 0 20682 480 6 chany_bottom_out[16]
port 78 nsew default tristate
rlabel metal2 s 21086 0 21142 480 6 chany_bottom_out[17]
port 79 nsew default tristate
rlabel metal2 s 21546 0 21602 480 6 chany_bottom_out[18]
port 80 nsew default tristate
rlabel metal2 s 22006 0 22062 480 6 chany_bottom_out[19]
port 81 nsew default tristate
rlabel metal2 s 13634 0 13690 480 6 chany_bottom_out[1]
port 82 nsew default tristate
rlabel metal2 s 14094 0 14150 480 6 chany_bottom_out[2]
port 83 nsew default tristate
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_out[3]
port 84 nsew default tristate
rlabel metal2 s 15014 0 15070 480 6 chany_bottom_out[4]
port 85 nsew default tristate
rlabel metal2 s 15566 0 15622 480 6 chany_bottom_out[5]
port 86 nsew default tristate
rlabel metal2 s 16026 0 16082 480 6 chany_bottom_out[6]
port 87 nsew default tristate
rlabel metal2 s 16486 0 16542 480 6 chany_bottom_out[7]
port 88 nsew default tristate
rlabel metal2 s 16946 0 17002 480 6 chany_bottom_out[8]
port 89 nsew default tristate
rlabel metal2 s 17406 0 17462 480 6 chany_bottom_out[9]
port 90 nsew default tristate
rlabel metal2 s 3790 22320 3846 22800 6 chany_top_in[0]
port 91 nsew default input
rlabel metal2 s 8390 22320 8446 22800 6 chany_top_in[10]
port 92 nsew default input
rlabel metal2 s 8850 22320 8906 22800 6 chany_top_in[11]
port 93 nsew default input
rlabel metal2 s 9310 22320 9366 22800 6 chany_top_in[12]
port 94 nsew default input
rlabel metal2 s 9770 22320 9826 22800 6 chany_top_in[13]
port 95 nsew default input
rlabel metal2 s 10230 22320 10286 22800 6 chany_top_in[14]
port 96 nsew default input
rlabel metal2 s 10690 22320 10746 22800 6 chany_top_in[15]
port 97 nsew default input
rlabel metal2 s 11150 22320 11206 22800 6 chany_top_in[16]
port 98 nsew default input
rlabel metal2 s 11610 22320 11666 22800 6 chany_top_in[17]
port 99 nsew default input
rlabel metal2 s 11978 22320 12034 22800 6 chany_top_in[18]
port 100 nsew default input
rlabel metal2 s 12438 22320 12494 22800 6 chany_top_in[19]
port 101 nsew default input
rlabel metal2 s 4250 22320 4306 22800 6 chany_top_in[1]
port 102 nsew default input
rlabel metal2 s 4710 22320 4766 22800 6 chany_top_in[2]
port 103 nsew default input
rlabel metal2 s 5170 22320 5226 22800 6 chany_top_in[3]
port 104 nsew default input
rlabel metal2 s 5630 22320 5686 22800 6 chany_top_in[4]
port 105 nsew default input
rlabel metal2 s 6090 22320 6146 22800 6 chany_top_in[5]
port 106 nsew default input
rlabel metal2 s 6550 22320 6606 22800 6 chany_top_in[6]
port 107 nsew default input
rlabel metal2 s 7010 22320 7066 22800 6 chany_top_in[7]
port 108 nsew default input
rlabel metal2 s 7470 22320 7526 22800 6 chany_top_in[8]
port 109 nsew default input
rlabel metal2 s 7930 22320 7986 22800 6 chany_top_in[9]
port 110 nsew default input
rlabel metal2 s 12898 22320 12954 22800 6 chany_top_out[0]
port 111 nsew default tristate
rlabel metal2 s 17498 22320 17554 22800 6 chany_top_out[10]
port 112 nsew default tristate
rlabel metal2 s 17958 22320 18014 22800 6 chany_top_out[11]
port 113 nsew default tristate
rlabel metal2 s 18418 22320 18474 22800 6 chany_top_out[12]
port 114 nsew default tristate
rlabel metal2 s 18878 22320 18934 22800 6 chany_top_out[13]
port 115 nsew default tristate
rlabel metal2 s 19338 22320 19394 22800 6 chany_top_out[14]
port 116 nsew default tristate
rlabel metal2 s 19798 22320 19854 22800 6 chany_top_out[15]
port 117 nsew default tristate
rlabel metal2 s 20258 22320 20314 22800 6 chany_top_out[16]
port 118 nsew default tristate
rlabel metal2 s 20718 22320 20774 22800 6 chany_top_out[17]
port 119 nsew default tristate
rlabel metal2 s 21178 22320 21234 22800 6 chany_top_out[18]
port 120 nsew default tristate
rlabel metal2 s 21638 22320 21694 22800 6 chany_top_out[19]
port 121 nsew default tristate
rlabel metal2 s 13358 22320 13414 22800 6 chany_top_out[1]
port 122 nsew default tristate
rlabel metal2 s 13818 22320 13874 22800 6 chany_top_out[2]
port 123 nsew default tristate
rlabel metal2 s 14278 22320 14334 22800 6 chany_top_out[3]
port 124 nsew default tristate
rlabel metal2 s 14738 22320 14794 22800 6 chany_top_out[4]
port 125 nsew default tristate
rlabel metal2 s 15198 22320 15254 22800 6 chany_top_out[5]
port 126 nsew default tristate
rlabel metal2 s 15658 22320 15714 22800 6 chany_top_out[6]
port 127 nsew default tristate
rlabel metal2 s 16118 22320 16174 22800 6 chany_top_out[7]
port 128 nsew default tristate
rlabel metal2 s 16578 22320 16634 22800 6 chany_top_out[8]
port 129 nsew default tristate
rlabel metal2 s 17038 22320 17094 22800 6 chany_top_out[9]
port 130 nsew default tristate
rlabel metal3 s 0 144 480 264 6 left_bottom_grid_pin_34_
port 131 nsew default input
rlabel metal3 s 0 552 480 672 6 left_bottom_grid_pin_35_
port 132 nsew default input
rlabel metal3 s 0 1096 480 1216 6 left_bottom_grid_pin_36_
port 133 nsew default input
rlabel metal3 s 0 1504 480 1624 6 left_bottom_grid_pin_37_
port 134 nsew default input
rlabel metal3 s 0 2048 480 2168 6 left_bottom_grid_pin_38_
port 135 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_39_
port 136 nsew default input
rlabel metal3 s 0 3000 480 3120 6 left_bottom_grid_pin_40_
port 137 nsew default input
rlabel metal3 s 0 3408 480 3528 6 left_bottom_grid_pin_41_
port 138 nsew default input
rlabel metal2 s 22098 22320 22154 22800 6 prog_clk_0_N_in
port 139 nsew default input
rlabel metal2 s 202 22320 258 22800 6 top_left_grid_pin_42_
port 140 nsew default input
rlabel metal2 s 570 22320 626 22800 6 top_left_grid_pin_43_
port 141 nsew default input
rlabel metal2 s 1030 22320 1086 22800 6 top_left_grid_pin_44_
port 142 nsew default input
rlabel metal2 s 1490 22320 1546 22800 6 top_left_grid_pin_45_
port 143 nsew default input
rlabel metal2 s 1950 22320 2006 22800 6 top_left_grid_pin_46_
port 144 nsew default input
rlabel metal2 s 2410 22320 2466 22800 6 top_left_grid_pin_47_
port 145 nsew default input
rlabel metal2 s 2870 22320 2926 22800 6 top_left_grid_pin_48_
port 146 nsew default input
rlabel metal2 s 3330 22320 3386 22800 6 top_left_grid_pin_49_
port 147 nsew default input
rlabel metal2 s 22558 22320 22614 22800 6 top_right_grid_pin_1_
port 148 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 149 nsew default input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 150 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22800
<< end >>
