magic
tech sky130A
magscale 1 2
timestamp 1606930023
<< locali >>
rect 12817 18071 12851 18309
rect 16589 15963 16623 16133
rect 11161 14331 11195 14501
rect 14289 13787 14323 13957
rect 17877 13719 17911 13889
rect 15117 13311 15151 13481
rect 18705 13175 18739 13481
rect 16681 9911 16715 10081
rect 19533 8415 19567 8517
rect 14289 6171 14323 6341
rect 15025 5695 15059 5865
<< viali >>
rect 10333 20009 10367 20043
rect 11897 20009 11931 20043
rect 11989 20009 12023 20043
rect 12817 20009 12851 20043
rect 13737 20009 13771 20043
rect 14289 20009 14323 20043
rect 14841 20009 14875 20043
rect 16313 20009 16347 20043
rect 16865 20009 16899 20043
rect 17417 20009 17451 20043
rect 18521 20009 18555 20043
rect 19073 20009 19107 20043
rect 19625 20009 19659 20043
rect 20177 20009 20211 20043
rect 20729 20009 20763 20043
rect 10425 19941 10459 19975
rect 10977 19873 11011 19907
rect 12633 19873 12667 19907
rect 13553 19873 13587 19907
rect 14105 19873 14139 19907
rect 14657 19873 14691 19907
rect 15577 19873 15611 19907
rect 16129 19873 16163 19907
rect 16681 19873 16715 19907
rect 17233 19873 17267 19907
rect 18337 19873 18371 19907
rect 18889 19873 18923 19907
rect 19441 19873 19475 19907
rect 19993 19873 20027 19907
rect 20545 19873 20579 19907
rect 10609 19805 10643 19839
rect 12081 19805 12115 19839
rect 11161 19737 11195 19771
rect 9965 19669 9999 19703
rect 11529 19669 11563 19703
rect 15761 19669 15795 19703
rect 10149 19329 10183 19363
rect 12449 19329 12483 19363
rect 16405 19329 16439 19363
rect 8493 19261 8527 19295
rect 11805 19261 11839 19295
rect 14105 19261 14139 19295
rect 14749 19261 14783 19295
rect 15025 19261 15059 19295
rect 17049 19261 17083 19295
rect 18245 19261 18279 19295
rect 18521 19261 18555 19295
rect 19073 19261 19107 19295
rect 19717 19261 19751 19295
rect 8760 19193 8794 19227
rect 10416 19193 10450 19227
rect 12694 19193 12728 19227
rect 17325 19193 17359 19227
rect 20545 19193 20579 19227
rect 9873 19125 9907 19159
rect 11529 19125 11563 19159
rect 11989 19125 12023 19159
rect 13829 19125 13863 19159
rect 14289 19125 14323 19159
rect 15761 19125 15795 19159
rect 16129 19125 16163 19159
rect 16221 19125 16255 19159
rect 19257 19125 19291 19159
rect 9137 18921 9171 18955
rect 11897 18921 11931 18955
rect 16681 18921 16715 18955
rect 17141 18921 17175 18955
rect 17969 18921 18003 18955
rect 18797 18921 18831 18955
rect 10784 18853 10818 18887
rect 12992 18853 13026 18887
rect 15546 18853 15580 18887
rect 19993 18853 20027 18887
rect 7757 18785 7791 18819
rect 8024 18785 8058 18819
rect 9965 18785 9999 18819
rect 10517 18785 10551 18819
rect 12173 18785 12207 18819
rect 12725 18785 12759 18819
rect 14381 18785 14415 18819
rect 14657 18785 14691 18819
rect 16957 18785 16991 18819
rect 17785 18785 17819 18819
rect 18613 18785 18647 18819
rect 19165 18785 19199 18819
rect 19717 18785 19751 18819
rect 15301 18717 15335 18751
rect 10149 18649 10183 18683
rect 12357 18581 12391 18615
rect 14105 18581 14139 18615
rect 19349 18581 19383 18615
rect 12909 18377 12943 18411
rect 15761 18377 15795 18411
rect 19441 18377 19475 18411
rect 8861 18309 8895 18343
rect 9965 18309 9999 18343
rect 12817 18309 12851 18343
rect 17693 18309 17727 18343
rect 9413 18241 9447 18275
rect 10425 18241 10459 18275
rect 10609 18241 10643 18275
rect 12449 18241 12483 18275
rect 9229 18173 9263 18207
rect 9321 18173 9355 18207
rect 10977 18173 11011 18207
rect 11805 18173 11839 18207
rect 10333 18105 10367 18139
rect 11253 18105 11287 18139
rect 13553 18241 13587 18275
rect 16313 18241 16347 18275
rect 18797 18241 18831 18275
rect 19993 18241 20027 18275
rect 13921 18173 13955 18207
rect 14188 18173 14222 18207
rect 15577 18173 15611 18207
rect 19257 18173 19291 18207
rect 19809 18173 19843 18207
rect 20545 18173 20579 18207
rect 16580 18105 16614 18139
rect 18521 18105 18555 18139
rect 20821 18105 20855 18139
rect 11989 18037 12023 18071
rect 12817 18037 12851 18071
rect 13277 18037 13311 18071
rect 13369 18037 13403 18071
rect 15301 18037 15335 18071
rect 18153 18037 18187 18071
rect 18613 18037 18647 18071
rect 8953 17833 8987 17867
rect 9689 17833 9723 17867
rect 10057 17833 10091 17867
rect 13001 17833 13035 17867
rect 15761 17833 15795 17867
rect 16773 17833 16807 17867
rect 19165 17833 19199 17867
rect 19257 17833 19291 17867
rect 19809 17833 19843 17867
rect 20913 17833 20947 17867
rect 17408 17765 17442 17799
rect 7573 17697 7607 17731
rect 7840 17697 7874 17731
rect 10149 17697 10183 17731
rect 10793 17697 10827 17731
rect 11897 17697 11931 17731
rect 11989 17697 12023 17731
rect 12541 17697 12575 17731
rect 13369 17697 13403 17731
rect 14565 17697 14599 17731
rect 15301 17697 15335 17731
rect 16129 17697 16163 17731
rect 16957 17697 16991 17731
rect 17141 17697 17175 17731
rect 20177 17697 20211 17731
rect 10333 17629 10367 17663
rect 11069 17629 11103 17663
rect 12081 17629 12115 17663
rect 13461 17629 13495 17663
rect 13553 17629 13587 17663
rect 14657 17629 14691 17663
rect 14841 17629 14875 17663
rect 16221 17629 16255 17663
rect 16313 17629 16347 17663
rect 19441 17629 19475 17663
rect 20269 17629 20303 17663
rect 20361 17629 20395 17663
rect 18521 17561 18555 17595
rect 11529 17493 11563 17527
rect 14197 17493 14231 17527
rect 18797 17493 18831 17527
rect 8401 17289 8435 17323
rect 12541 17289 12575 17323
rect 14749 17289 14783 17323
rect 15761 17289 15795 17323
rect 11989 17221 12023 17255
rect 13737 17221 13771 17255
rect 17049 17221 17083 17255
rect 9229 17153 9263 17187
rect 10241 17153 10275 17187
rect 11345 17153 11379 17187
rect 13001 17153 13035 17187
rect 13185 17153 13219 17187
rect 14381 17153 14415 17187
rect 15393 17153 15427 17187
rect 16313 17153 16347 17187
rect 19993 17153 20027 17187
rect 7021 17085 7055 17119
rect 11805 17085 11839 17119
rect 14197 17085 14231 17119
rect 16865 17085 16899 17119
rect 17417 17085 17451 17119
rect 18061 17085 18095 17119
rect 19717 17085 19751 17119
rect 20453 17085 20487 17119
rect 7288 17017 7322 17051
rect 10057 17017 10091 17051
rect 11161 17017 11195 17051
rect 15117 17017 15151 17051
rect 18328 17017 18362 17051
rect 20729 17017 20763 17051
rect 8677 16949 8711 16983
rect 9045 16949 9079 16983
rect 9137 16949 9171 16983
rect 9689 16949 9723 16983
rect 10149 16949 10183 16983
rect 10793 16949 10827 16983
rect 11253 16949 11287 16983
rect 12909 16949 12943 16983
rect 14105 16949 14139 16983
rect 15209 16949 15243 16983
rect 16129 16949 16163 16983
rect 16221 16949 16255 16983
rect 17601 16949 17635 16983
rect 19441 16949 19475 16983
rect 7389 16745 7423 16779
rect 7481 16745 7515 16779
rect 8217 16745 8251 16779
rect 11805 16745 11839 16779
rect 12081 16745 12115 16779
rect 17141 16745 17175 16779
rect 17969 16745 18003 16779
rect 18521 16745 18555 16779
rect 18981 16745 19015 16779
rect 19533 16745 19567 16779
rect 8677 16677 8711 16711
rect 9965 16677 9999 16711
rect 12449 16677 12483 16711
rect 13093 16677 13127 16711
rect 13820 16677 13854 16711
rect 15301 16677 15335 16711
rect 17877 16677 17911 16711
rect 19993 16677 20027 16711
rect 8585 16609 8619 16643
rect 9505 16609 9539 16643
rect 9689 16609 9723 16643
rect 10692 16609 10726 16643
rect 13553 16609 13587 16643
rect 16129 16609 16163 16643
rect 16221 16609 16255 16643
rect 16957 16609 16991 16643
rect 18889 16609 18923 16643
rect 19901 16609 19935 16643
rect 7665 16541 7699 16575
rect 8769 16541 8803 16575
rect 10425 16541 10459 16575
rect 12541 16541 12575 16575
rect 12633 16541 12667 16575
rect 16405 16541 16439 16575
rect 18153 16541 18187 16575
rect 19165 16541 19199 16575
rect 20085 16541 20119 16575
rect 7021 16473 7055 16507
rect 9321 16473 9355 16507
rect 17509 16473 17543 16507
rect 14933 16405 14967 16439
rect 15761 16405 15795 16439
rect 8217 16201 8251 16235
rect 13829 16201 13863 16235
rect 15485 16133 15519 16167
rect 16589 16133 16623 16167
rect 16773 16133 16807 16167
rect 9505 16065 9539 16099
rect 11713 16065 11747 16099
rect 12449 16065 12483 16099
rect 16221 16065 16255 16099
rect 16313 16065 16347 16099
rect 6837 15997 6871 16031
rect 8769 15997 8803 16031
rect 14105 15997 14139 16031
rect 17417 16065 17451 16099
rect 18061 16065 18095 16099
rect 20361 16065 20395 16099
rect 17141 15997 17175 16031
rect 20821 15997 20855 16031
rect 7104 15929 7138 15963
rect 9045 15929 9079 15963
rect 9772 15929 9806 15963
rect 11621 15929 11655 15963
rect 12716 15929 12750 15963
rect 14372 15929 14406 15963
rect 16129 15929 16163 15963
rect 16589 15929 16623 15963
rect 18328 15929 18362 15963
rect 20177 15929 20211 15963
rect 10885 15861 10919 15895
rect 11161 15861 11195 15895
rect 11529 15861 11563 15895
rect 15761 15861 15795 15895
rect 17233 15861 17267 15895
rect 19441 15861 19475 15895
rect 19809 15861 19843 15895
rect 20269 15861 20303 15895
rect 21005 15861 21039 15895
rect 7941 15657 7975 15691
rect 10517 15657 10551 15691
rect 10885 15657 10919 15691
rect 13001 15657 13035 15691
rect 13461 15657 13495 15691
rect 15669 15657 15703 15691
rect 17785 15657 17819 15691
rect 20453 15657 20487 15691
rect 6368 15589 6402 15623
rect 12265 15589 12299 15623
rect 13369 15589 13403 15623
rect 15761 15589 15795 15623
rect 18766 15589 18800 15623
rect 6101 15521 6135 15555
rect 8769 15521 8803 15555
rect 9689 15521 9723 15555
rect 14565 15521 14599 15555
rect 14657 15521 14691 15555
rect 16405 15521 16439 15555
rect 16672 15521 16706 15555
rect 18061 15521 18095 15555
rect 20269 15521 20303 15555
rect 8861 15453 8895 15487
rect 9045 15453 9079 15487
rect 9965 15453 9999 15487
rect 10977 15453 11011 15487
rect 11069 15453 11103 15487
rect 12357 15453 12391 15487
rect 12541 15453 12575 15487
rect 13553 15453 13587 15487
rect 14841 15453 14875 15487
rect 15853 15453 15887 15487
rect 18521 15453 18555 15487
rect 7481 15317 7515 15351
rect 8401 15317 8435 15351
rect 11897 15317 11931 15351
rect 14197 15317 14231 15351
rect 15301 15317 15335 15351
rect 19901 15317 19935 15351
rect 5733 15113 5767 15147
rect 8861 15113 8895 15147
rect 10333 15113 10367 15147
rect 11345 15113 11379 15147
rect 13829 15113 13863 15147
rect 18153 15113 18187 15147
rect 21005 15113 21039 15147
rect 15761 15045 15795 15079
rect 16405 15045 16439 15079
rect 6193 14977 6227 15011
rect 6377 14977 6411 15011
rect 9689 14977 9723 15011
rect 10885 14977 10919 15011
rect 11805 14977 11839 15011
rect 11989 14977 12023 15011
rect 14381 14977 14415 15011
rect 17325 14977 17359 15011
rect 18705 14977 18739 15011
rect 19165 14977 19199 15011
rect 6101 14909 6135 14943
rect 7481 14909 7515 14943
rect 7748 14909 7782 14943
rect 10701 14909 10735 14943
rect 11713 14909 11747 14943
rect 12449 14909 12483 14943
rect 14289 14909 14323 14943
rect 14648 14909 14682 14943
rect 16221 14909 16255 14943
rect 18521 14909 18555 14943
rect 20821 14909 20855 14943
rect 9505 14841 9539 14875
rect 12716 14841 12750 14875
rect 17141 14841 17175 14875
rect 19432 14841 19466 14875
rect 9137 14773 9171 14807
rect 9597 14773 9631 14807
rect 10793 14773 10827 14807
rect 14105 14773 14139 14807
rect 16773 14773 16807 14807
rect 17233 14773 17267 14807
rect 18613 14773 18647 14807
rect 20545 14773 20579 14807
rect 8769 14569 8803 14603
rect 11345 14569 11379 14603
rect 13829 14569 13863 14603
rect 19257 14569 19291 14603
rect 20085 14569 20119 14603
rect 7012 14501 7046 14535
rect 8861 14501 8895 14535
rect 11161 14501 11195 14535
rect 14657 14501 14691 14535
rect 16396 14501 16430 14535
rect 6745 14433 6779 14467
rect 9689 14433 9723 14467
rect 9956 14433 9990 14467
rect 8953 14365 8987 14399
rect 11529 14433 11563 14467
rect 11980 14433 12014 14467
rect 13737 14433 13771 14467
rect 14381 14433 14415 14467
rect 15301 14433 15335 14467
rect 16129 14433 16163 14467
rect 18153 14433 18187 14467
rect 18245 14433 18279 14467
rect 19073 14433 19107 14467
rect 19993 14433 20027 14467
rect 11713 14365 11747 14399
rect 13921 14365 13955 14399
rect 15577 14365 15611 14399
rect 18337 14365 18371 14399
rect 20177 14365 20211 14399
rect 20913 14365 20947 14399
rect 8125 14297 8159 14331
rect 11161 14297 11195 14331
rect 19625 14297 19659 14331
rect 8401 14229 8435 14263
rect 11069 14229 11103 14263
rect 13093 14229 13127 14263
rect 13369 14229 13403 14263
rect 17509 14229 17543 14263
rect 17785 14229 17819 14263
rect 12449 14025 12483 14059
rect 15945 14025 15979 14059
rect 17693 14025 17727 14059
rect 18061 14025 18095 14059
rect 19809 14025 19843 14059
rect 21005 14025 21039 14059
rect 14289 13957 14323 13991
rect 14473 13957 14507 13991
rect 15485 13957 15519 13991
rect 8769 13889 8803 13923
rect 9505 13889 9539 13923
rect 11621 13889 11655 13923
rect 11713 13889 11747 13923
rect 13001 13889 13035 13923
rect 13921 13889 13955 13923
rect 14013 13889 14047 13923
rect 9772 13821 9806 13855
rect 12817 13821 12851 13855
rect 14933 13889 14967 13923
rect 15025 13889 15059 13923
rect 17877 13889 17911 13923
rect 18613 13889 18647 13923
rect 19257 13889 19291 13923
rect 20361 13889 20395 13923
rect 15669 13821 15703 13855
rect 15761 13821 15795 13855
rect 16313 13821 16347 13855
rect 13829 13753 13863 13787
rect 14289 13753 14323 13787
rect 16580 13753 16614 13787
rect 19073 13821 19107 13855
rect 20821 13821 20855 13855
rect 18429 13753 18463 13787
rect 20177 13753 20211 13787
rect 10885 13685 10919 13719
rect 11161 13685 11195 13719
rect 11529 13685 11563 13719
rect 12909 13685 12943 13719
rect 13461 13685 13495 13719
rect 14841 13685 14875 13719
rect 17877 13685 17911 13719
rect 18521 13685 18555 13719
rect 20269 13685 20303 13719
rect 9321 13481 9355 13515
rect 9873 13481 9907 13515
rect 10333 13481 10367 13515
rect 10885 13481 10919 13515
rect 11345 13481 11379 13515
rect 12817 13481 12851 13515
rect 14197 13481 14231 13515
rect 15117 13481 15151 13515
rect 16497 13481 16531 13515
rect 17049 13481 17083 13515
rect 17141 13481 17175 13515
rect 17877 13481 17911 13515
rect 18705 13481 18739 13515
rect 18889 13481 18923 13515
rect 19809 13481 19843 13515
rect 12357 13413 12391 13447
rect 14657 13413 14691 13447
rect 9505 13345 9539 13379
rect 10241 13345 10275 13379
rect 11253 13345 11287 13379
rect 12081 13345 12115 13379
rect 13001 13345 13035 13379
rect 13185 13345 13219 13379
rect 14565 13345 14599 13379
rect 15761 13413 15795 13447
rect 15669 13345 15703 13379
rect 16313 13345 16347 13379
rect 18245 13345 18279 13379
rect 10425 13277 10459 13311
rect 11437 13277 11471 13311
rect 13461 13277 13495 13311
rect 14841 13277 14875 13311
rect 15117 13277 15151 13311
rect 15853 13277 15887 13311
rect 17325 13277 17359 13311
rect 17693 13277 17727 13311
rect 18337 13277 18371 13311
rect 18521 13277 18555 13311
rect 16681 13209 16715 13243
rect 19717 13345 19751 13379
rect 19993 13277 20027 13311
rect 15301 13141 15335 13175
rect 18705 13141 18739 13175
rect 19349 13141 19383 13175
rect 10425 12937 10459 12971
rect 12449 12937 12483 12971
rect 16497 12937 16531 12971
rect 16773 12937 16807 12971
rect 8769 12801 8803 12835
rect 10977 12801 11011 12835
rect 13001 12801 13035 12835
rect 17417 12801 17451 12835
rect 18337 12801 18371 12835
rect 20637 12801 20671 12835
rect 9036 12733 9070 12767
rect 13461 12733 13495 12767
rect 15117 12733 15151 12767
rect 17233 12733 17267 12767
rect 18061 12733 18095 12767
rect 18797 12733 18831 12767
rect 19064 12733 19098 12767
rect 20453 12733 20487 12767
rect 10793 12665 10827 12699
rect 11437 12665 11471 12699
rect 12817 12665 12851 12699
rect 13728 12665 13762 12699
rect 15362 12665 15396 12699
rect 17141 12665 17175 12699
rect 10149 12597 10183 12631
rect 10885 12597 10919 12631
rect 12909 12597 12943 12631
rect 14841 12597 14875 12631
rect 20177 12597 20211 12631
rect 12725 12393 12759 12427
rect 14381 12393 14415 12427
rect 14657 12393 14691 12427
rect 17601 12393 17635 12427
rect 19993 12393 20027 12427
rect 20453 12393 20487 12427
rect 8024 12325 8058 12359
rect 13246 12325 13280 12359
rect 16120 12325 16154 12359
rect 20913 12325 20947 12359
rect 7757 12257 7791 12291
rect 9689 12257 9723 12291
rect 11612 12257 11646 12291
rect 13001 12257 13035 12291
rect 17969 12257 18003 12291
rect 18613 12257 18647 12291
rect 18880 12257 18914 12291
rect 20269 12257 20303 12291
rect 9965 12189 9999 12223
rect 11345 12189 11379 12223
rect 15301 12189 15335 12223
rect 15853 12189 15887 12223
rect 18061 12189 18095 12223
rect 18245 12189 18279 12223
rect 9137 12053 9171 12087
rect 17233 12053 17267 12087
rect 11529 11849 11563 11883
rect 12633 11849 12667 11883
rect 14381 11849 14415 11883
rect 15577 11849 15611 11883
rect 19349 11849 19383 11883
rect 21097 11849 21131 11883
rect 13553 11781 13587 11815
rect 12081 11713 12115 11747
rect 13185 11713 13219 11747
rect 14197 11713 14231 11747
rect 14933 11713 14967 11747
rect 16037 11713 16071 11747
rect 16221 11713 16255 11747
rect 17601 11713 17635 11747
rect 18613 11713 18647 11747
rect 8217 11645 8251 11679
rect 14013 11645 14047 11679
rect 19165 11645 19199 11679
rect 19717 11645 19751 11679
rect 8484 11577 8518 11611
rect 11253 11577 11287 11611
rect 11897 11577 11931 11611
rect 13093 11577 13127 11611
rect 15945 11577 15979 11611
rect 18429 11577 18463 11611
rect 19984 11577 20018 11611
rect 9597 11509 9631 11543
rect 9873 11509 9907 11543
rect 11989 11509 12023 11543
rect 13001 11509 13035 11543
rect 13921 11509 13955 11543
rect 14749 11509 14783 11543
rect 14841 11509 14875 11543
rect 16957 11509 16991 11543
rect 17325 11509 17359 11543
rect 17417 11509 17451 11543
rect 18061 11509 18095 11543
rect 18521 11509 18555 11543
rect 9689 11305 9723 11339
rect 10057 11305 10091 11339
rect 12357 11305 12391 11339
rect 14197 11305 14231 11339
rect 15577 11305 15611 11339
rect 8953 11237 8987 11271
rect 16856 11237 16890 11271
rect 18705 11237 18739 11271
rect 19993 11237 20027 11271
rect 10977 11169 11011 11203
rect 11244 11169 11278 11203
rect 12909 11169 12943 11203
rect 15945 11169 15979 11203
rect 18613 11169 18647 11203
rect 19901 11169 19935 11203
rect 9045 11101 9079 11135
rect 9137 11101 9171 11135
rect 10149 11101 10183 11135
rect 10241 11101 10275 11135
rect 16037 11101 16071 11135
rect 16129 11101 16163 11135
rect 16589 11101 16623 11135
rect 18797 11101 18831 11135
rect 20085 11101 20119 11135
rect 8585 11033 8619 11067
rect 17969 11033 18003 11067
rect 18245 11033 18279 11067
rect 19533 10965 19567 10999
rect 12449 10761 12483 10795
rect 13461 10761 13495 10795
rect 15393 10761 15427 10795
rect 18613 10761 18647 10795
rect 11345 10693 11379 10727
rect 11897 10625 11931 10659
rect 13093 10625 13127 10659
rect 14105 10625 14139 10659
rect 15117 10625 15151 10659
rect 15853 10625 15887 10659
rect 16037 10625 16071 10659
rect 18061 10625 18095 10659
rect 19257 10625 19291 10659
rect 8033 10557 8067 10591
rect 8300 10557 8334 10591
rect 9689 10557 9723 10591
rect 10609 10557 10643 10591
rect 11713 10557 11747 10591
rect 12909 10557 12943 10591
rect 13829 10557 13863 10591
rect 13921 10557 13955 10591
rect 15025 10557 15059 10591
rect 15761 10557 15795 10591
rect 16313 10557 16347 10591
rect 16580 10557 16614 10591
rect 18981 10557 19015 10591
rect 19625 10557 19659 10591
rect 9965 10489 9999 10523
rect 14933 10489 14967 10523
rect 19892 10489 19926 10523
rect 9413 10421 9447 10455
rect 10425 10421 10459 10455
rect 11805 10421 11839 10455
rect 12817 10421 12851 10455
rect 14565 10421 14599 10455
rect 17693 10421 17727 10455
rect 19073 10421 19107 10455
rect 21005 10421 21039 10455
rect 9689 10217 9723 10251
rect 12081 10217 12115 10251
rect 13645 10217 13679 10251
rect 14197 10217 14231 10251
rect 14657 10217 14691 10251
rect 15301 10217 15335 10251
rect 16773 10217 16807 10251
rect 17233 10217 17267 10251
rect 18061 10217 18095 10251
rect 20453 10217 20487 10251
rect 20913 10217 20947 10251
rect 10968 10149 11002 10183
rect 12633 10149 12667 10183
rect 13553 10149 13587 10183
rect 15761 10149 15795 10183
rect 16405 10149 16439 10183
rect 17141 10149 17175 10183
rect 19340 10149 19374 10183
rect 9137 10081 9171 10115
rect 10057 10081 10091 10115
rect 12357 10081 12391 10115
rect 14565 10081 14599 10115
rect 15669 10081 15703 10115
rect 16129 10081 16163 10115
rect 16681 10081 16715 10115
rect 18429 10081 18463 10115
rect 10149 10013 10183 10047
rect 10241 10013 10275 10047
rect 10701 10013 10735 10047
rect 13737 10013 13771 10047
rect 14749 10013 14783 10047
rect 15945 10013 15979 10047
rect 17417 10013 17451 10047
rect 18521 10013 18555 10047
rect 18705 10013 18739 10047
rect 19073 10013 19107 10047
rect 13185 9877 13219 9911
rect 16681 9877 16715 9911
rect 17417 9673 17451 9707
rect 11437 9605 11471 9639
rect 16129 9605 16163 9639
rect 14473 9537 14507 9571
rect 16681 9537 16715 9571
rect 18061 9537 18095 9571
rect 20545 9537 20579 9571
rect 20637 9537 20671 9571
rect 8217 9469 8251 9503
rect 8484 9469 8518 9503
rect 10057 9469 10091 9503
rect 12449 9469 12483 9503
rect 12716 9469 12750 9503
rect 14289 9469 14323 9503
rect 14740 9469 14774 9503
rect 16589 9469 16623 9503
rect 17601 9469 17635 9503
rect 10324 9401 10358 9435
rect 16957 9401 16991 9435
rect 18306 9401 18340 9435
rect 20453 9401 20487 9435
rect 9597 9333 9631 9367
rect 11713 9333 11747 9367
rect 13829 9333 13863 9367
rect 14105 9333 14139 9367
rect 15853 9333 15887 9367
rect 16497 9333 16531 9367
rect 19441 9333 19475 9367
rect 20085 9333 20119 9367
rect 8585 9129 8619 9163
rect 11069 9129 11103 9163
rect 11345 9129 11379 9163
rect 17141 9129 17175 9163
rect 17601 9129 17635 9163
rect 19993 9129 20027 9163
rect 9045 9061 9079 9095
rect 13268 9061 13302 9095
rect 17969 9061 18003 9095
rect 18880 9061 18914 9095
rect 8953 8993 8987 9027
rect 9689 8993 9723 9027
rect 9956 8993 9990 9027
rect 11713 8993 11747 9027
rect 13001 8993 13035 9027
rect 15761 8993 15795 9027
rect 16028 8993 16062 9027
rect 18613 8993 18647 9027
rect 9229 8925 9263 8959
rect 11805 8925 11839 8959
rect 11897 8925 11931 8959
rect 18061 8925 18095 8959
rect 18245 8925 18279 8959
rect 14381 8789 14415 8823
rect 10609 8585 10643 8619
rect 10885 8585 10919 8619
rect 11897 8585 11931 8619
rect 15209 8585 15243 8619
rect 18705 8585 18739 8619
rect 12449 8517 12483 8551
rect 16773 8517 16807 8551
rect 19533 8517 19567 8551
rect 19717 8517 19751 8551
rect 11437 8449 11471 8483
rect 13001 8449 13035 8483
rect 14381 8449 14415 8483
rect 16405 8449 16439 8483
rect 17417 8449 17451 8483
rect 19349 8449 19383 8483
rect 20177 8449 20211 8483
rect 20361 8449 20395 8483
rect 9229 8381 9263 8415
rect 11253 8381 11287 8415
rect 12081 8381 12115 8415
rect 15393 8381 15427 8415
rect 17233 8381 17267 8415
rect 19165 8381 19199 8415
rect 19533 8381 19567 8415
rect 9496 8313 9530 8347
rect 11345 8313 11379 8347
rect 12817 8313 12851 8347
rect 14289 8313 14323 8347
rect 16129 8313 16163 8347
rect 16221 8313 16255 8347
rect 17141 8313 17175 8347
rect 19073 8313 19107 8347
rect 12909 8245 12943 8279
rect 13829 8245 13863 8279
rect 14197 8245 14231 8279
rect 15761 8245 15795 8279
rect 20085 8245 20119 8279
rect 10057 8041 10091 8075
rect 12449 8041 12483 8075
rect 12909 8041 12943 8075
rect 13369 8041 13403 8075
rect 13921 8041 13955 8075
rect 14289 8041 14323 8075
rect 15761 8041 15795 8075
rect 16221 8041 16255 8075
rect 20361 8041 20395 8075
rect 20913 8041 20947 8075
rect 9137 7973 9171 8007
rect 13277 7973 13311 8007
rect 19248 7973 19282 8007
rect 8861 7905 8895 7939
rect 10425 7905 10459 7939
rect 11325 7905 11359 7939
rect 14381 7905 14415 7939
rect 16129 7905 16163 7939
rect 16773 7905 16807 7939
rect 17040 7905 17074 7939
rect 18981 7905 19015 7939
rect 10517 7837 10551 7871
rect 10701 7837 10735 7871
rect 11069 7837 11103 7871
rect 13461 7837 13495 7871
rect 14473 7837 14507 7871
rect 16405 7837 16439 7871
rect 18153 7701 18187 7735
rect 9781 7497 9815 7531
rect 10333 7497 10367 7531
rect 11345 7497 11379 7531
rect 12817 7497 12851 7531
rect 15209 7497 15243 7531
rect 16957 7497 16991 7531
rect 10885 7361 10919 7395
rect 11897 7361 11931 7395
rect 13369 7361 13403 7395
rect 17233 7361 17267 7395
rect 18613 7361 18647 7395
rect 20453 7361 20487 7395
rect 8401 7293 8435 7327
rect 10793 7293 10827 7327
rect 13829 7293 13863 7327
rect 14096 7293 14130 7327
rect 15577 7293 15611 7327
rect 15844 7293 15878 7327
rect 18429 7293 18463 7327
rect 20361 7293 20395 7327
rect 8668 7225 8702 7259
rect 11713 7225 11747 7259
rect 20269 7225 20303 7259
rect 10701 7157 10735 7191
rect 11805 7157 11839 7191
rect 13185 7157 13219 7191
rect 13277 7157 13311 7191
rect 18061 7157 18095 7191
rect 18521 7157 18555 7191
rect 19901 7157 19935 7191
rect 9689 6953 9723 6987
rect 13461 6953 13495 6987
rect 13921 6953 13955 6987
rect 15669 6953 15703 6987
rect 16313 6953 16347 6987
rect 17325 6953 17359 6987
rect 17877 6953 17911 6987
rect 18245 6953 18279 6987
rect 20545 6953 20579 6987
rect 11069 6885 11103 6919
rect 14289 6885 14323 6919
rect 17233 6885 17267 6919
rect 10057 6817 10091 6851
rect 12072 6817 12106 6851
rect 15761 6817 15795 6851
rect 16497 6817 16531 6851
rect 19432 6817 19466 6851
rect 9137 6749 9171 6783
rect 10149 6749 10183 6783
rect 10241 6749 10275 6783
rect 11161 6749 11195 6783
rect 11253 6749 11287 6783
rect 11805 6749 11839 6783
rect 14381 6749 14415 6783
rect 14473 6749 14507 6783
rect 15853 6749 15887 6783
rect 17509 6749 17543 6783
rect 18337 6749 18371 6783
rect 18521 6749 18555 6783
rect 19165 6749 19199 6783
rect 16865 6681 16899 6715
rect 10701 6613 10735 6647
rect 13185 6613 13219 6647
rect 15301 6613 15335 6647
rect 9873 6409 9907 6443
rect 10149 6409 10183 6443
rect 18245 6409 18279 6443
rect 20637 6409 20671 6443
rect 14289 6341 14323 6375
rect 10701 6273 10735 6307
rect 11713 6273 11747 6307
rect 13093 6273 13127 6307
rect 14105 6273 14139 6307
rect 6837 6205 6871 6239
rect 8493 6205 8527 6239
rect 10517 6205 10551 6239
rect 11621 6205 11655 6239
rect 13829 6205 13863 6239
rect 15025 6273 15059 6307
rect 16313 6273 16347 6307
rect 17233 6273 17267 6307
rect 18889 6273 18923 6307
rect 16129 6205 16163 6239
rect 17141 6205 17175 6239
rect 19257 6205 19291 6239
rect 19524 6205 19558 6239
rect 7082 6137 7116 6171
rect 8738 6137 8772 6171
rect 11529 6137 11563 6171
rect 12817 6137 12851 6171
rect 13921 6137 13955 6171
rect 14289 6137 14323 6171
rect 14933 6137 14967 6171
rect 16037 6137 16071 6171
rect 18613 6137 18647 6171
rect 8217 6069 8251 6103
rect 10609 6069 10643 6103
rect 11161 6069 11195 6103
rect 12449 6069 12483 6103
rect 12909 6069 12943 6103
rect 13461 6069 13495 6103
rect 14473 6069 14507 6103
rect 14841 6069 14875 6103
rect 15669 6069 15703 6103
rect 16681 6069 16715 6103
rect 17049 6069 17083 6103
rect 18705 6069 18739 6103
rect 9781 5865 9815 5899
rect 10149 5865 10183 5899
rect 13001 5865 13035 5899
rect 14197 5865 14231 5899
rect 14565 5865 14599 5899
rect 15025 5865 15059 5899
rect 16681 5865 16715 5899
rect 18613 5865 18647 5899
rect 20913 5865 20947 5899
rect 11152 5797 11186 5831
rect 10885 5729 10919 5763
rect 12909 5729 12943 5763
rect 14657 5729 14691 5763
rect 15568 5797 15602 5831
rect 19134 5797 19168 5831
rect 15301 5729 15335 5763
rect 17233 5729 17267 5763
rect 17500 5729 17534 5763
rect 10241 5661 10275 5695
rect 10333 5661 10367 5695
rect 13185 5661 13219 5695
rect 14841 5661 14875 5695
rect 15025 5661 15059 5695
rect 18889 5661 18923 5695
rect 12265 5593 12299 5627
rect 12541 5525 12575 5559
rect 20269 5525 20303 5559
rect 10333 5321 10367 5355
rect 11345 5321 11379 5355
rect 12449 5321 12483 5355
rect 15025 5321 15059 5355
rect 17233 5321 17267 5355
rect 19901 5321 19935 5355
rect 10793 5185 10827 5219
rect 10977 5185 11011 5219
rect 13093 5185 13127 5219
rect 15853 5185 15887 5219
rect 18521 5185 18555 5219
rect 20729 5185 20763 5219
rect 11529 5117 11563 5151
rect 13645 5117 13679 5151
rect 16120 5117 16154 5151
rect 18788 5117 18822 5151
rect 11897 5049 11931 5083
rect 12817 5049 12851 5083
rect 13890 5049 13924 5083
rect 20545 5049 20579 5083
rect 10701 4981 10735 5015
rect 12909 4981 12943 5015
rect 15301 4981 15335 5015
rect 18061 4981 18095 5015
rect 20177 4981 20211 5015
rect 20637 4981 20671 5015
rect 13461 4777 13495 4811
rect 15301 4777 15335 4811
rect 16313 4777 16347 4811
rect 17785 4777 17819 4811
rect 18153 4777 18187 4811
rect 19165 4777 19199 4811
rect 20177 4777 20211 4811
rect 12081 4641 12115 4675
rect 12348 4641 12382 4675
rect 13737 4641 13771 4675
rect 14565 4641 14599 4675
rect 15669 4641 15703 4675
rect 19257 4641 19291 4675
rect 15761 4573 15795 4607
rect 15853 4573 15887 4607
rect 16957 4573 16991 4607
rect 18245 4573 18279 4607
rect 18337 4573 18371 4607
rect 19441 4573 19475 4607
rect 20269 4573 20303 4607
rect 20361 4573 20395 4607
rect 13921 4437 13955 4471
rect 14749 4437 14783 4471
rect 18797 4437 18831 4471
rect 19809 4437 19843 4471
rect 19717 4233 19751 4267
rect 9137 4097 9171 4131
rect 11437 4097 11471 4131
rect 13369 4097 13403 4131
rect 14565 4097 14599 4131
rect 20177 4097 20211 4131
rect 20269 4097 20303 4131
rect 15025 4029 15059 4063
rect 15761 4029 15795 4063
rect 16497 4029 16531 4063
rect 17417 4029 17451 4063
rect 18061 4029 18095 4063
rect 20085 4029 20119 4063
rect 20729 4029 20763 4063
rect 9404 3961 9438 3995
rect 11161 3961 11195 3995
rect 11805 3961 11839 3995
rect 13277 3961 13311 3995
rect 14381 3961 14415 3995
rect 16037 3961 16071 3995
rect 18328 3961 18362 3995
rect 10517 3893 10551 3927
rect 10793 3893 10827 3927
rect 11253 3893 11287 3927
rect 12817 3893 12851 3927
rect 13185 3893 13219 3927
rect 14013 3893 14047 3927
rect 14473 3893 14507 3927
rect 15209 3893 15243 3927
rect 16681 3893 16715 3927
rect 17601 3893 17635 3927
rect 19441 3893 19475 3927
rect 20913 3893 20947 3927
rect 11437 3689 11471 3723
rect 14749 3689 14783 3723
rect 17049 3689 17083 3723
rect 18705 3689 18739 3723
rect 11958 3621 11992 3655
rect 15936 3621 15970 3655
rect 17570 3621 17604 3655
rect 10057 3553 10091 3587
rect 10324 3553 10358 3587
rect 13369 3553 13403 3587
rect 13625 3553 13659 3587
rect 15669 3553 15703 3587
rect 17325 3553 17359 3587
rect 19073 3553 19107 3587
rect 19809 3553 19843 3587
rect 11713 3485 11747 3519
rect 19349 3485 19383 3519
rect 20085 3485 20119 3519
rect 13093 3417 13127 3451
rect 10425 3145 10459 3179
rect 13369 3145 13403 3179
rect 16589 3145 16623 3179
rect 18061 3145 18095 3179
rect 16221 3077 16255 3111
rect 19625 3077 19659 3111
rect 10977 3009 11011 3043
rect 13921 3009 13955 3043
rect 14381 3009 14415 3043
rect 17233 3009 17267 3043
rect 18521 3009 18555 3043
rect 18705 3009 18739 3043
rect 11621 2941 11655 2975
rect 12449 2941 12483 2975
rect 13829 2941 13863 2975
rect 16037 2941 16071 2975
rect 16957 2941 16991 2975
rect 18429 2941 18463 2975
rect 18889 2941 18923 2975
rect 19441 2941 19475 2975
rect 19993 2941 20027 2975
rect 20545 2941 20579 2975
rect 11897 2873 11931 2907
rect 12725 2873 12759 2907
rect 14626 2873 14660 2907
rect 10793 2805 10827 2839
rect 10885 2805 10919 2839
rect 13737 2805 13771 2839
rect 15761 2805 15795 2839
rect 17049 2805 17083 2839
rect 20177 2805 20211 2839
rect 20729 2805 20763 2839
rect 16037 2601 16071 2635
rect 13737 2533 13771 2567
rect 11345 2465 11379 2499
rect 11897 2465 11931 2499
rect 12725 2465 12759 2499
rect 13461 2465 13495 2499
rect 14197 2465 14231 2499
rect 14749 2465 14783 2499
rect 15945 2465 15979 2499
rect 16589 2465 16623 2499
rect 17325 2465 17359 2499
rect 18429 2465 18463 2499
rect 18981 2465 19015 2499
rect 19533 2465 19567 2499
rect 20361 2465 20395 2499
rect 12909 2397 12943 2431
rect 16129 2397 16163 2431
rect 11529 2329 11563 2363
rect 14933 2329 14967 2363
rect 15577 2329 15611 2363
rect 19717 2329 19751 2363
rect 12081 2261 12115 2295
rect 14381 2261 14415 2295
rect 16773 2261 16807 2295
rect 17509 2261 17543 2295
rect 18613 2261 18647 2295
rect 19165 2261 19199 2295
rect 20545 2261 20579 2295
<< metal1 >>
rect 7466 20204 7472 20256
rect 7524 20244 7530 20256
rect 12066 20244 12072 20256
rect 7524 20216 12072 20244
rect 7524 20204 7530 20216
rect 12066 20204 12072 20216
rect 12124 20204 12130 20256
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 10321 20043 10379 20049
rect 10321 20009 10333 20043
rect 10367 20040 10379 20043
rect 11146 20040 11152 20052
rect 10367 20012 11152 20040
rect 10367 20009 10379 20012
rect 10321 20003 10379 20009
rect 11146 20000 11152 20012
rect 11204 20000 11210 20052
rect 11330 20000 11336 20052
rect 11388 20040 11394 20052
rect 11885 20043 11943 20049
rect 11885 20040 11897 20043
rect 11388 20012 11897 20040
rect 11388 20000 11394 20012
rect 11885 20009 11897 20012
rect 11931 20009 11943 20043
rect 11885 20003 11943 20009
rect 11977 20043 12035 20049
rect 11977 20009 11989 20043
rect 12023 20040 12035 20043
rect 12066 20040 12072 20052
rect 12023 20012 12072 20040
rect 12023 20009 12035 20012
rect 11977 20003 12035 20009
rect 12066 20000 12072 20012
rect 12124 20040 12130 20052
rect 12342 20040 12348 20052
rect 12124 20012 12348 20040
rect 12124 20000 12130 20012
rect 12342 20000 12348 20012
rect 12400 20000 12406 20052
rect 12805 20043 12863 20049
rect 12805 20009 12817 20043
rect 12851 20040 12863 20043
rect 13078 20040 13084 20052
rect 12851 20012 13084 20040
rect 12851 20009 12863 20012
rect 12805 20003 12863 20009
rect 13078 20000 13084 20012
rect 13136 20000 13142 20052
rect 13725 20043 13783 20049
rect 13725 20009 13737 20043
rect 13771 20009 13783 20043
rect 13725 20003 13783 20009
rect 10413 19975 10471 19981
rect 10413 19941 10425 19975
rect 10459 19972 10471 19975
rect 10778 19972 10784 19984
rect 10459 19944 10784 19972
rect 10459 19941 10471 19944
rect 10413 19935 10471 19941
rect 10778 19932 10784 19944
rect 10836 19972 10842 19984
rect 13740 19972 13768 20003
rect 14182 20000 14188 20052
rect 14240 20040 14246 20052
rect 14277 20043 14335 20049
rect 14277 20040 14289 20043
rect 14240 20012 14289 20040
rect 14240 20000 14246 20012
rect 14277 20009 14289 20012
rect 14323 20009 14335 20043
rect 14277 20003 14335 20009
rect 14550 20000 14556 20052
rect 14608 20040 14614 20052
rect 14829 20043 14887 20049
rect 14829 20040 14841 20043
rect 14608 20012 14841 20040
rect 14608 20000 14614 20012
rect 14829 20009 14841 20012
rect 14875 20009 14887 20043
rect 14829 20003 14887 20009
rect 15286 20000 15292 20052
rect 15344 20040 15350 20052
rect 16301 20043 16359 20049
rect 16301 20040 16313 20043
rect 15344 20012 16313 20040
rect 15344 20000 15350 20012
rect 16301 20009 16313 20012
rect 16347 20009 16359 20043
rect 16301 20003 16359 20009
rect 16574 20000 16580 20052
rect 16632 20040 16638 20052
rect 16853 20043 16911 20049
rect 16853 20040 16865 20043
rect 16632 20012 16865 20040
rect 16632 20000 16638 20012
rect 16853 20009 16865 20012
rect 16899 20009 16911 20043
rect 16853 20003 16911 20009
rect 17405 20043 17463 20049
rect 17405 20009 17417 20043
rect 17451 20040 17463 20043
rect 17494 20040 17500 20052
rect 17451 20012 17500 20040
rect 17451 20009 17463 20012
rect 17405 20003 17463 20009
rect 17494 20000 17500 20012
rect 17552 20000 17558 20052
rect 18046 20000 18052 20052
rect 18104 20040 18110 20052
rect 18509 20043 18567 20049
rect 18509 20040 18521 20043
rect 18104 20012 18521 20040
rect 18104 20000 18110 20012
rect 18509 20009 18521 20012
rect 18555 20009 18567 20043
rect 18509 20003 18567 20009
rect 19061 20043 19119 20049
rect 19061 20009 19073 20043
rect 19107 20040 19119 20043
rect 19150 20040 19156 20052
rect 19107 20012 19156 20040
rect 19107 20009 19119 20012
rect 19061 20003 19119 20009
rect 19150 20000 19156 20012
rect 19208 20000 19214 20052
rect 19613 20043 19671 20049
rect 19613 20009 19625 20043
rect 19659 20040 19671 20043
rect 19702 20040 19708 20052
rect 19659 20012 19708 20040
rect 19659 20009 19671 20012
rect 19613 20003 19671 20009
rect 19702 20000 19708 20012
rect 19760 20000 19766 20052
rect 20162 20040 20168 20052
rect 20123 20012 20168 20040
rect 20162 20000 20168 20012
rect 20220 20000 20226 20052
rect 20622 20000 20628 20052
rect 20680 20040 20686 20052
rect 20717 20043 20775 20049
rect 20717 20040 20729 20043
rect 20680 20012 20729 20040
rect 20680 20000 20686 20012
rect 20717 20009 20729 20012
rect 20763 20009 20775 20043
rect 20717 20003 20775 20009
rect 20254 19972 20260 19984
rect 10836 19944 12940 19972
rect 13740 19944 20260 19972
rect 10836 19932 10842 19944
rect 10870 19864 10876 19916
rect 10928 19904 10934 19916
rect 10965 19907 11023 19913
rect 10965 19904 10977 19907
rect 10928 19876 10977 19904
rect 10928 19864 10934 19876
rect 10965 19873 10977 19876
rect 11011 19873 11023 19907
rect 12618 19904 12624 19916
rect 12579 19876 12624 19904
rect 10965 19867 11023 19873
rect 12618 19864 12624 19876
rect 12676 19864 12682 19916
rect 10597 19839 10655 19845
rect 10597 19805 10609 19839
rect 10643 19836 10655 19839
rect 10686 19836 10692 19848
rect 10643 19808 10692 19836
rect 10643 19805 10655 19808
rect 10597 19799 10655 19805
rect 10686 19796 10692 19808
rect 10744 19796 10750 19848
rect 12066 19836 12072 19848
rect 12027 19808 12072 19836
rect 12066 19796 12072 19808
rect 12124 19796 12130 19848
rect 11149 19771 11207 19777
rect 11149 19737 11161 19771
rect 11195 19768 11207 19771
rect 11882 19768 11888 19780
rect 11195 19740 11888 19768
rect 11195 19737 11207 19740
rect 11149 19731 11207 19737
rect 11882 19728 11888 19740
rect 11940 19728 11946 19780
rect 12912 19768 12940 19944
rect 20254 19932 20260 19944
rect 20312 19932 20318 19984
rect 13078 19864 13084 19916
rect 13136 19904 13142 19916
rect 13541 19907 13599 19913
rect 13541 19904 13553 19907
rect 13136 19876 13553 19904
rect 13136 19864 13142 19876
rect 13541 19873 13553 19876
rect 13587 19873 13599 19907
rect 14090 19904 14096 19916
rect 14051 19876 14096 19904
rect 13541 19867 13599 19873
rect 14090 19864 14096 19876
rect 14148 19864 14154 19916
rect 14645 19907 14703 19913
rect 14645 19873 14657 19907
rect 14691 19873 14703 19907
rect 14645 19867 14703 19873
rect 13906 19796 13912 19848
rect 13964 19836 13970 19848
rect 14660 19836 14688 19867
rect 15010 19864 15016 19916
rect 15068 19904 15074 19916
rect 15565 19907 15623 19913
rect 15565 19904 15577 19907
rect 15068 19876 15577 19904
rect 15068 19864 15074 19876
rect 15565 19873 15577 19876
rect 15611 19873 15623 19907
rect 15565 19867 15623 19873
rect 16117 19907 16175 19913
rect 16117 19873 16129 19907
rect 16163 19873 16175 19907
rect 16117 19867 16175 19873
rect 16669 19907 16727 19913
rect 16669 19873 16681 19907
rect 16715 19873 16727 19907
rect 16669 19867 16727 19873
rect 13964 19808 14688 19836
rect 13964 19796 13970 19808
rect 15378 19796 15384 19848
rect 15436 19836 15442 19848
rect 16132 19836 16160 19867
rect 15436 19808 16160 19836
rect 16684 19836 16712 19867
rect 17126 19864 17132 19916
rect 17184 19904 17190 19916
rect 17221 19907 17279 19913
rect 17221 19904 17233 19907
rect 17184 19876 17233 19904
rect 17184 19864 17190 19876
rect 17221 19873 17233 19876
rect 17267 19873 17279 19907
rect 17221 19867 17279 19873
rect 18325 19907 18383 19913
rect 18325 19873 18337 19907
rect 18371 19873 18383 19907
rect 18325 19867 18383 19873
rect 17402 19836 17408 19848
rect 16684 19808 17408 19836
rect 15436 19796 15442 19808
rect 17402 19796 17408 19808
rect 17460 19796 17466 19848
rect 18340 19768 18368 19867
rect 18690 19864 18696 19916
rect 18748 19904 18754 19916
rect 18877 19907 18935 19913
rect 18877 19904 18889 19907
rect 18748 19876 18889 19904
rect 18748 19864 18754 19876
rect 18877 19873 18889 19876
rect 18923 19873 18935 19907
rect 19426 19904 19432 19916
rect 19387 19876 19432 19904
rect 18877 19867 18935 19873
rect 19426 19864 19432 19876
rect 19484 19864 19490 19916
rect 19978 19904 19984 19916
rect 19939 19876 19984 19904
rect 19978 19864 19984 19876
rect 20036 19864 20042 19916
rect 20162 19864 20168 19916
rect 20220 19904 20226 19916
rect 20533 19907 20591 19913
rect 20533 19904 20545 19907
rect 20220 19876 20545 19904
rect 20220 19864 20226 19876
rect 20533 19873 20545 19876
rect 20579 19873 20591 19907
rect 20533 19867 20591 19873
rect 12912 19740 18368 19768
rect 9953 19703 10011 19709
rect 9953 19669 9965 19703
rect 9999 19700 10011 19703
rect 10318 19700 10324 19712
rect 9999 19672 10324 19700
rect 9999 19669 10011 19672
rect 9953 19663 10011 19669
rect 10318 19660 10324 19672
rect 10376 19660 10382 19712
rect 11517 19703 11575 19709
rect 11517 19669 11529 19703
rect 11563 19700 11575 19703
rect 12158 19700 12164 19712
rect 11563 19672 12164 19700
rect 11563 19669 11575 19672
rect 11517 19663 11575 19669
rect 12158 19660 12164 19672
rect 12216 19660 12222 19712
rect 15749 19703 15807 19709
rect 15749 19669 15761 19703
rect 15795 19700 15807 19703
rect 17954 19700 17960 19712
rect 15795 19672 17960 19700
rect 15795 19669 15807 19672
rect 15749 19663 15807 19669
rect 17954 19660 17960 19672
rect 18012 19660 18018 19712
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 8478 19456 8484 19508
rect 8536 19496 8542 19508
rect 10502 19496 10508 19508
rect 8536 19468 10508 19496
rect 8536 19456 8542 19468
rect 10152 19369 10180 19468
rect 10502 19456 10508 19468
rect 10560 19496 10566 19508
rect 10560 19468 11100 19496
rect 10560 19456 10566 19468
rect 11072 19428 11100 19468
rect 11072 19400 12480 19428
rect 12452 19369 12480 19400
rect 13464 19400 14964 19428
rect 10137 19363 10195 19369
rect 10137 19329 10149 19363
rect 10183 19329 10195 19363
rect 10137 19323 10195 19329
rect 12437 19363 12495 19369
rect 12437 19329 12449 19363
rect 12483 19329 12495 19363
rect 12437 19323 12495 19329
rect 7742 19252 7748 19304
rect 7800 19292 7806 19304
rect 8478 19292 8484 19304
rect 7800 19264 8484 19292
rect 7800 19252 7806 19264
rect 8478 19252 8484 19264
rect 8536 19252 8542 19304
rect 11790 19292 11796 19304
rect 8680 19264 10548 19292
rect 11751 19264 11796 19292
rect 8202 19184 8208 19236
rect 8260 19224 8266 19236
rect 8680 19224 8708 19264
rect 8260 19196 8708 19224
rect 8748 19227 8806 19233
rect 8260 19184 8266 19196
rect 8748 19193 8760 19227
rect 8794 19224 8806 19227
rect 8938 19224 8944 19236
rect 8794 19196 8944 19224
rect 8794 19193 8806 19196
rect 8748 19187 8806 19193
rect 8938 19184 8944 19196
rect 8996 19184 9002 19236
rect 10404 19227 10462 19233
rect 10404 19193 10416 19227
rect 10450 19193 10462 19227
rect 10520 19224 10548 19264
rect 11790 19252 11796 19264
rect 11848 19252 11854 19304
rect 11882 19224 11888 19236
rect 10520 19196 11888 19224
rect 10404 19187 10462 19193
rect 6362 19116 6368 19168
rect 6420 19156 6426 19168
rect 9306 19156 9312 19168
rect 6420 19128 9312 19156
rect 6420 19116 6426 19128
rect 9306 19116 9312 19128
rect 9364 19116 9370 19168
rect 9861 19159 9919 19165
rect 9861 19125 9873 19159
rect 9907 19156 9919 19159
rect 10428 19156 10456 19187
rect 11882 19184 11888 19196
rect 11940 19184 11946 19236
rect 12066 19184 12072 19236
rect 12124 19224 12130 19236
rect 12682 19227 12740 19233
rect 12682 19224 12694 19227
rect 12124 19196 12694 19224
rect 12124 19184 12130 19196
rect 12682 19193 12694 19196
rect 12728 19193 12740 19227
rect 12682 19187 12740 19193
rect 10686 19156 10692 19168
rect 9907 19128 10692 19156
rect 9907 19125 9919 19128
rect 9861 19119 9919 19125
rect 10686 19116 10692 19128
rect 10744 19116 10750 19168
rect 11514 19156 11520 19168
rect 11475 19128 11520 19156
rect 11514 19116 11520 19128
rect 11572 19116 11578 19168
rect 11977 19159 12035 19165
rect 11977 19125 11989 19159
rect 12023 19156 12035 19159
rect 12526 19156 12532 19168
rect 12023 19128 12532 19156
rect 12023 19125 12035 19128
rect 11977 19119 12035 19125
rect 12526 19116 12532 19128
rect 12584 19116 12590 19168
rect 12802 19116 12808 19168
rect 12860 19156 12866 19168
rect 13464 19156 13492 19400
rect 14936 19360 14964 19400
rect 16393 19363 16451 19369
rect 14936 19332 15148 19360
rect 14093 19295 14151 19301
rect 14093 19261 14105 19295
rect 14139 19292 14151 19295
rect 14182 19292 14188 19304
rect 14139 19264 14188 19292
rect 14139 19261 14151 19264
rect 14093 19255 14151 19261
rect 14182 19252 14188 19264
rect 14240 19252 14246 19304
rect 14274 19252 14280 19304
rect 14332 19292 14338 19304
rect 14737 19295 14795 19301
rect 14737 19292 14749 19295
rect 14332 19264 14749 19292
rect 14332 19252 14338 19264
rect 14737 19261 14749 19264
rect 14783 19261 14795 19295
rect 15010 19292 15016 19304
rect 14971 19264 15016 19292
rect 14737 19255 14795 19261
rect 15010 19252 15016 19264
rect 15068 19252 15074 19304
rect 15120 19292 15148 19332
rect 16393 19329 16405 19363
rect 16439 19360 16451 19363
rect 16666 19360 16672 19372
rect 16439 19332 16672 19360
rect 16439 19329 16451 19332
rect 16393 19323 16451 19329
rect 16666 19320 16672 19332
rect 16724 19320 16730 19372
rect 16776 19332 17172 19360
rect 16776 19292 16804 19332
rect 15120 19264 16804 19292
rect 16850 19252 16856 19304
rect 16908 19292 16914 19304
rect 17037 19295 17095 19301
rect 17037 19292 17049 19295
rect 16908 19264 17049 19292
rect 16908 19252 16914 19264
rect 17037 19261 17049 19264
rect 17083 19261 17095 19295
rect 17144 19292 17172 19332
rect 17144 19264 17540 19292
rect 17037 19255 17095 19261
rect 13630 19184 13636 19236
rect 13688 19224 13694 19236
rect 13688 19196 14320 19224
rect 13688 19184 13694 19196
rect 13814 19156 13820 19168
rect 12860 19128 13492 19156
rect 13775 19128 13820 19156
rect 12860 19116 12866 19128
rect 13814 19116 13820 19128
rect 13872 19116 13878 19168
rect 14292 19165 14320 19196
rect 15764 19196 17264 19224
rect 15764 19165 15792 19196
rect 14277 19159 14335 19165
rect 14277 19125 14289 19159
rect 14323 19125 14335 19159
rect 14277 19119 14335 19125
rect 15749 19159 15807 19165
rect 15749 19125 15761 19159
rect 15795 19125 15807 19159
rect 16114 19156 16120 19168
rect 16075 19128 16120 19156
rect 15749 19119 15807 19125
rect 16114 19116 16120 19128
rect 16172 19116 16178 19168
rect 16206 19116 16212 19168
rect 16264 19156 16270 19168
rect 17236 19156 17264 19196
rect 17310 19184 17316 19236
rect 17368 19224 17374 19236
rect 17512 19224 17540 19264
rect 17862 19252 17868 19304
rect 17920 19292 17926 19304
rect 18233 19295 18291 19301
rect 18233 19292 18245 19295
rect 17920 19264 18245 19292
rect 17920 19252 17926 19264
rect 18233 19261 18245 19264
rect 18279 19261 18291 19295
rect 18233 19255 18291 19261
rect 18509 19295 18567 19301
rect 18509 19261 18521 19295
rect 18555 19292 18567 19295
rect 19061 19295 19119 19301
rect 19061 19292 19073 19295
rect 18555 19264 19073 19292
rect 18555 19261 18567 19264
rect 18509 19255 18567 19261
rect 19061 19261 19073 19264
rect 19107 19261 19119 19295
rect 19061 19255 19119 19261
rect 19150 19252 19156 19304
rect 19208 19292 19214 19304
rect 19705 19295 19763 19301
rect 19705 19292 19717 19295
rect 19208 19264 19717 19292
rect 19208 19252 19214 19264
rect 19705 19261 19717 19264
rect 19751 19261 19763 19295
rect 19705 19255 19763 19261
rect 20070 19224 20076 19236
rect 17368 19196 17413 19224
rect 17512 19196 20076 19224
rect 17368 19184 17374 19196
rect 20070 19184 20076 19196
rect 20128 19184 20134 19236
rect 20530 19224 20536 19236
rect 20491 19196 20536 19224
rect 20530 19184 20536 19196
rect 20588 19184 20594 19236
rect 19058 19156 19064 19168
rect 16264 19128 16309 19156
rect 17236 19128 19064 19156
rect 16264 19116 16270 19128
rect 19058 19116 19064 19128
rect 19116 19116 19122 19168
rect 19242 19156 19248 19168
rect 19203 19128 19248 19156
rect 19242 19116 19248 19128
rect 19300 19116 19306 19168
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 290 18912 296 18964
rect 348 18952 354 18964
rect 348 18924 8892 18952
rect 348 18912 354 18924
rect 8864 18884 8892 18924
rect 8938 18912 8944 18964
rect 8996 18952 9002 18964
rect 9125 18955 9183 18961
rect 9125 18952 9137 18955
rect 8996 18924 9137 18952
rect 8996 18912 9002 18924
rect 9125 18921 9137 18924
rect 9171 18921 9183 18955
rect 9125 18915 9183 18921
rect 11885 18955 11943 18961
rect 11885 18921 11897 18955
rect 11931 18952 11943 18955
rect 12066 18952 12072 18964
rect 11931 18924 12072 18952
rect 11931 18921 11943 18924
rect 11885 18915 11943 18921
rect 12066 18912 12072 18924
rect 12124 18912 12130 18964
rect 13538 18952 13544 18964
rect 12995 18924 13544 18952
rect 9858 18884 9864 18896
rect 8864 18856 9864 18884
rect 9858 18844 9864 18856
rect 9916 18844 9922 18896
rect 10594 18844 10600 18896
rect 10652 18884 10658 18896
rect 10772 18887 10830 18893
rect 10772 18884 10784 18887
rect 10652 18856 10784 18884
rect 10652 18844 10658 18856
rect 10772 18853 10784 18856
rect 10818 18884 10830 18887
rect 11514 18884 11520 18896
rect 10818 18856 11520 18884
rect 10818 18853 10830 18856
rect 10772 18847 10830 18853
rect 11514 18844 11520 18856
rect 11572 18844 11578 18896
rect 12995 18893 13023 18924
rect 13538 18912 13544 18924
rect 13596 18952 13602 18964
rect 13814 18952 13820 18964
rect 13596 18924 13820 18952
rect 13596 18912 13602 18924
rect 13814 18912 13820 18924
rect 13872 18912 13878 18964
rect 16666 18952 16672 18964
rect 16627 18924 16672 18952
rect 16666 18912 16672 18924
rect 16724 18912 16730 18964
rect 16942 18912 16948 18964
rect 17000 18952 17006 18964
rect 17129 18955 17187 18961
rect 17129 18952 17141 18955
rect 17000 18924 17141 18952
rect 17000 18912 17006 18924
rect 17129 18921 17141 18924
rect 17175 18921 17187 18955
rect 17129 18915 17187 18921
rect 17957 18955 18015 18961
rect 17957 18921 17969 18955
rect 18003 18952 18015 18955
rect 18506 18952 18512 18964
rect 18003 18924 18512 18952
rect 18003 18921 18015 18924
rect 17957 18915 18015 18921
rect 18506 18912 18512 18924
rect 18564 18912 18570 18964
rect 18598 18912 18604 18964
rect 18656 18952 18662 18964
rect 18785 18955 18843 18961
rect 18785 18952 18797 18955
rect 18656 18924 18797 18952
rect 18656 18912 18662 18924
rect 18785 18921 18797 18924
rect 18831 18921 18843 18955
rect 18785 18915 18843 18921
rect 18874 18912 18880 18964
rect 18932 18952 18938 18964
rect 21910 18952 21916 18964
rect 18932 18924 21916 18952
rect 18932 18912 18938 18924
rect 21910 18912 21916 18924
rect 21968 18912 21974 18964
rect 12980 18887 13038 18893
rect 12980 18853 12992 18887
rect 13026 18853 13038 18887
rect 13630 18884 13636 18896
rect 12980 18847 13038 18853
rect 13096 18856 13636 18884
rect 7742 18816 7748 18828
rect 7703 18788 7748 18816
rect 7742 18776 7748 18788
rect 7800 18776 7806 18828
rect 8012 18819 8070 18825
rect 8012 18785 8024 18819
rect 8058 18816 8070 18819
rect 8846 18816 8852 18828
rect 8058 18788 8852 18816
rect 8058 18785 8070 18788
rect 8012 18779 8070 18785
rect 8846 18776 8852 18788
rect 8904 18776 8910 18828
rect 9953 18819 10011 18825
rect 9953 18785 9965 18819
rect 9999 18816 10011 18819
rect 10226 18816 10232 18828
rect 9999 18788 10232 18816
rect 9999 18785 10011 18788
rect 9953 18779 10011 18785
rect 10226 18776 10232 18788
rect 10284 18776 10290 18828
rect 10502 18816 10508 18828
rect 10463 18788 10508 18816
rect 10502 18776 10508 18788
rect 10560 18776 10566 18828
rect 12066 18776 12072 18828
rect 12124 18816 12130 18828
rect 12161 18819 12219 18825
rect 12161 18816 12173 18819
rect 12124 18788 12173 18816
rect 12124 18776 12130 18788
rect 12161 18785 12173 18788
rect 12207 18785 12219 18819
rect 12161 18779 12219 18785
rect 12713 18819 12771 18825
rect 12713 18785 12725 18819
rect 12759 18816 12771 18819
rect 13096 18816 13124 18856
rect 13630 18844 13636 18856
rect 13688 18884 13694 18896
rect 15286 18884 15292 18896
rect 13688 18856 15292 18884
rect 13688 18844 13694 18856
rect 15286 18844 15292 18856
rect 15344 18844 15350 18896
rect 15470 18844 15476 18896
rect 15528 18893 15534 18896
rect 15528 18887 15592 18893
rect 15528 18853 15546 18887
rect 15580 18853 15592 18887
rect 19978 18884 19984 18896
rect 19939 18856 19984 18884
rect 15528 18847 15592 18853
rect 15528 18844 15534 18847
rect 19978 18844 19984 18856
rect 20036 18844 20042 18896
rect 12759 18788 13124 18816
rect 12759 18785 12771 18788
rect 12713 18779 12771 18785
rect 13262 18776 13268 18828
rect 13320 18816 13326 18828
rect 14369 18819 14427 18825
rect 14369 18816 14381 18819
rect 13320 18788 14381 18816
rect 13320 18776 13326 18788
rect 14369 18785 14381 18788
rect 14415 18785 14427 18819
rect 14369 18779 14427 18785
rect 14645 18819 14703 18825
rect 14645 18785 14657 18819
rect 14691 18816 14703 18819
rect 14691 18788 16528 18816
rect 14691 18785 14703 18788
rect 14645 18779 14703 18785
rect 9674 18708 9680 18760
rect 9732 18748 9738 18760
rect 10410 18748 10416 18760
rect 9732 18720 10416 18748
rect 9732 18708 9738 18720
rect 10410 18708 10416 18720
rect 10468 18708 10474 18760
rect 14182 18708 14188 18760
rect 14240 18748 14246 18760
rect 15102 18748 15108 18760
rect 14240 18720 15108 18748
rect 14240 18708 14246 18720
rect 15102 18708 15108 18720
rect 15160 18708 15166 18760
rect 15286 18748 15292 18760
rect 15247 18720 15292 18748
rect 15286 18708 15292 18720
rect 15344 18708 15350 18760
rect 16500 18748 16528 18788
rect 16574 18776 16580 18828
rect 16632 18816 16638 18828
rect 16945 18819 17003 18825
rect 16945 18816 16957 18819
rect 16632 18788 16957 18816
rect 16632 18776 16638 18788
rect 16945 18785 16957 18788
rect 16991 18785 17003 18819
rect 16945 18779 17003 18785
rect 17310 18776 17316 18828
rect 17368 18816 17374 18828
rect 17773 18819 17831 18825
rect 17773 18816 17785 18819
rect 17368 18788 17785 18816
rect 17368 18776 17374 18788
rect 17773 18785 17785 18788
rect 17819 18785 17831 18819
rect 17773 18779 17831 18785
rect 18601 18819 18659 18825
rect 18601 18785 18613 18819
rect 18647 18816 18659 18819
rect 18782 18816 18788 18828
rect 18647 18788 18788 18816
rect 18647 18785 18659 18788
rect 18601 18779 18659 18785
rect 18782 18776 18788 18788
rect 18840 18776 18846 18828
rect 19153 18819 19211 18825
rect 19153 18785 19165 18819
rect 19199 18816 19211 18819
rect 19518 18816 19524 18828
rect 19199 18788 19524 18816
rect 19199 18785 19211 18788
rect 19153 18779 19211 18785
rect 19518 18776 19524 18788
rect 19576 18776 19582 18828
rect 19702 18816 19708 18828
rect 19663 18788 19708 18816
rect 19702 18776 19708 18788
rect 19760 18776 19766 18828
rect 16758 18748 16764 18760
rect 16500 18720 16764 18748
rect 16758 18708 16764 18720
rect 16816 18708 16822 18760
rect 17034 18708 17040 18760
rect 17092 18748 17098 18760
rect 21358 18748 21364 18760
rect 17092 18720 21364 18748
rect 17092 18708 17098 18720
rect 21358 18708 21364 18720
rect 21416 18708 21422 18760
rect 3050 18640 3056 18692
rect 3108 18680 3114 18692
rect 3108 18652 7788 18680
rect 3108 18640 3114 18652
rect 4706 18572 4712 18624
rect 4764 18612 4770 18624
rect 6178 18612 6184 18624
rect 4764 18584 6184 18612
rect 4764 18572 4770 18584
rect 6178 18572 6184 18584
rect 6236 18572 6242 18624
rect 7760 18612 7788 18652
rect 9766 18640 9772 18692
rect 9824 18680 9830 18692
rect 10137 18683 10195 18689
rect 10137 18680 10149 18683
rect 9824 18652 10149 18680
rect 9824 18640 9830 18652
rect 10137 18649 10149 18652
rect 10183 18649 10195 18683
rect 20806 18680 20812 18692
rect 10137 18643 10195 18649
rect 14016 18652 14320 18680
rect 12250 18612 12256 18624
rect 7760 18584 12256 18612
rect 12250 18572 12256 18584
rect 12308 18572 12314 18624
rect 12345 18615 12403 18621
rect 12345 18581 12357 18615
rect 12391 18612 12403 18615
rect 14016 18612 14044 18652
rect 12391 18584 14044 18612
rect 14093 18615 14151 18621
rect 12391 18581 12403 18584
rect 12345 18575 12403 18581
rect 14093 18581 14105 18615
rect 14139 18612 14151 18615
rect 14182 18612 14188 18624
rect 14139 18584 14188 18612
rect 14139 18581 14151 18584
rect 14093 18575 14151 18581
rect 14182 18572 14188 18584
rect 14240 18572 14246 18624
rect 14292 18612 14320 18652
rect 16592 18652 20812 18680
rect 16592 18612 16620 18652
rect 20806 18640 20812 18652
rect 20864 18640 20870 18692
rect 14292 18584 16620 18612
rect 19242 18572 19248 18624
rect 19300 18612 19306 18624
rect 19337 18615 19395 18621
rect 19337 18612 19349 18615
rect 19300 18584 19349 18612
rect 19300 18572 19306 18584
rect 19337 18581 19349 18584
rect 19383 18581 19395 18615
rect 19337 18575 19395 18581
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 9582 18368 9588 18420
rect 9640 18408 9646 18420
rect 11974 18408 11980 18420
rect 9640 18380 11980 18408
rect 9640 18368 9646 18380
rect 11974 18368 11980 18380
rect 12032 18368 12038 18420
rect 12897 18411 12955 18417
rect 12897 18377 12909 18411
rect 12943 18408 12955 18411
rect 13262 18408 13268 18420
rect 12943 18380 13268 18408
rect 12943 18377 12955 18380
rect 12897 18371 12955 18377
rect 13262 18368 13268 18380
rect 13320 18368 13326 18420
rect 15749 18411 15807 18417
rect 13372 18380 14872 18408
rect 8849 18343 8907 18349
rect 8849 18309 8861 18343
rect 8895 18340 8907 18343
rect 9950 18340 9956 18352
rect 8895 18312 9812 18340
rect 9911 18312 9956 18340
rect 8895 18309 8907 18312
rect 8849 18303 8907 18309
rect 3602 18232 3608 18284
rect 3660 18272 3666 18284
rect 8202 18272 8208 18284
rect 3660 18244 8208 18272
rect 3660 18232 3666 18244
rect 8202 18232 8208 18244
rect 8260 18232 8266 18284
rect 8938 18232 8944 18284
rect 8996 18272 9002 18284
rect 9401 18275 9459 18281
rect 9401 18272 9413 18275
rect 8996 18244 9413 18272
rect 8996 18232 9002 18244
rect 9401 18241 9413 18244
rect 9447 18241 9459 18275
rect 9784 18272 9812 18312
rect 9950 18300 9956 18312
rect 10008 18300 10014 18352
rect 10502 18300 10508 18352
rect 10560 18340 10566 18352
rect 10686 18340 10692 18352
rect 10560 18312 10692 18340
rect 10560 18300 10566 18312
rect 10686 18300 10692 18312
rect 10744 18300 10750 18352
rect 12805 18343 12863 18349
rect 12805 18309 12817 18343
rect 12851 18340 12863 18343
rect 13372 18340 13400 18380
rect 12851 18312 13400 18340
rect 14844 18340 14872 18380
rect 15749 18377 15761 18411
rect 15795 18408 15807 18411
rect 15838 18408 15844 18420
rect 15795 18380 15844 18408
rect 15795 18377 15807 18380
rect 15749 18371 15807 18377
rect 15838 18368 15844 18380
rect 15896 18368 15902 18420
rect 17034 18408 17040 18420
rect 15948 18380 17040 18408
rect 15948 18340 15976 18380
rect 17034 18368 17040 18380
rect 17092 18368 17098 18420
rect 19150 18368 19156 18420
rect 19208 18408 19214 18420
rect 19429 18411 19487 18417
rect 19429 18408 19441 18411
rect 19208 18380 19441 18408
rect 19208 18368 19214 18380
rect 19429 18377 19441 18380
rect 19475 18377 19487 18411
rect 19429 18371 19487 18377
rect 14844 18312 15976 18340
rect 17681 18343 17739 18349
rect 12851 18309 12863 18312
rect 12805 18303 12863 18309
rect 17681 18309 17693 18343
rect 17727 18309 17739 18343
rect 17681 18303 17739 18309
rect 10134 18272 10140 18284
rect 9784 18244 10140 18272
rect 9401 18235 9459 18241
rect 10134 18232 10140 18244
rect 10192 18232 10198 18284
rect 10410 18272 10416 18284
rect 10371 18244 10416 18272
rect 10410 18232 10416 18244
rect 10468 18232 10474 18284
rect 10594 18272 10600 18284
rect 10555 18244 10600 18272
rect 10594 18232 10600 18244
rect 10652 18232 10658 18284
rect 11146 18232 11152 18284
rect 11204 18272 11210 18284
rect 12437 18275 12495 18281
rect 12437 18272 12449 18275
rect 11204 18244 12449 18272
rect 11204 18232 11210 18244
rect 12437 18241 12449 18244
rect 12483 18241 12495 18275
rect 12437 18235 12495 18241
rect 13541 18275 13599 18281
rect 13541 18241 13553 18275
rect 13587 18272 13599 18275
rect 13587 18244 14044 18272
rect 13587 18241 13599 18244
rect 13541 18235 13599 18241
rect 9122 18164 9128 18216
rect 9180 18204 9186 18216
rect 9217 18207 9275 18213
rect 9217 18204 9229 18207
rect 9180 18176 9229 18204
rect 9180 18164 9186 18176
rect 9217 18173 9229 18176
rect 9263 18173 9275 18207
rect 9217 18167 9275 18173
rect 9306 18164 9312 18216
rect 9364 18204 9370 18216
rect 10965 18207 11023 18213
rect 9364 18176 9409 18204
rect 9364 18164 9370 18176
rect 10965 18173 10977 18207
rect 11011 18173 11023 18207
rect 10965 18167 11023 18173
rect 11793 18207 11851 18213
rect 11793 18173 11805 18207
rect 11839 18204 11851 18207
rect 13170 18204 13176 18216
rect 11839 18176 13176 18204
rect 11839 18173 11851 18176
rect 11793 18167 11851 18173
rect 4154 18096 4160 18148
rect 4212 18136 4218 18148
rect 9490 18136 9496 18148
rect 4212 18108 9496 18136
rect 4212 18096 4218 18108
rect 9490 18096 9496 18108
rect 9548 18096 9554 18148
rect 10318 18136 10324 18148
rect 10279 18108 10324 18136
rect 10318 18096 10324 18108
rect 10376 18096 10382 18148
rect 5810 18028 5816 18080
rect 5868 18068 5874 18080
rect 7466 18068 7472 18080
rect 5868 18040 7472 18068
rect 5868 18028 5874 18040
rect 7466 18028 7472 18040
rect 7524 18028 7530 18080
rect 10594 18028 10600 18080
rect 10652 18068 10658 18080
rect 10980 18068 11008 18167
rect 13170 18164 13176 18176
rect 13228 18164 13234 18216
rect 13630 18164 13636 18216
rect 13688 18204 13694 18216
rect 13909 18207 13967 18213
rect 13909 18204 13921 18207
rect 13688 18176 13921 18204
rect 13688 18164 13694 18176
rect 13909 18173 13921 18176
rect 13955 18173 13967 18207
rect 14016 18204 14044 18244
rect 15286 18232 15292 18284
rect 15344 18272 15350 18284
rect 16298 18272 16304 18284
rect 15344 18244 16304 18272
rect 15344 18232 15350 18244
rect 16298 18232 16304 18244
rect 16356 18232 16362 18284
rect 17696 18272 17724 18303
rect 17954 18300 17960 18352
rect 18012 18340 18018 18352
rect 18012 18312 20024 18340
rect 18012 18300 18018 18312
rect 18785 18275 18843 18281
rect 18785 18272 18797 18275
rect 17696 18244 18797 18272
rect 18785 18241 18797 18244
rect 18831 18272 18843 18275
rect 18874 18272 18880 18284
rect 18831 18244 18880 18272
rect 18831 18241 18843 18244
rect 18785 18235 18843 18241
rect 18874 18232 18880 18244
rect 18932 18232 18938 18284
rect 19058 18232 19064 18284
rect 19116 18272 19122 18284
rect 19996 18281 20024 18312
rect 19981 18275 20039 18281
rect 19116 18244 19840 18272
rect 19116 18232 19122 18244
rect 14182 18213 14188 18216
rect 14176 18204 14188 18213
rect 14016 18176 14188 18204
rect 13909 18167 13967 18173
rect 14176 18167 14188 18176
rect 14182 18164 14188 18167
rect 14240 18164 14246 18216
rect 15565 18207 15623 18213
rect 15565 18173 15577 18207
rect 15611 18204 15623 18207
rect 15746 18204 15752 18216
rect 15611 18176 15752 18204
rect 15611 18173 15623 18176
rect 15565 18167 15623 18173
rect 15746 18164 15752 18176
rect 15804 18164 15810 18216
rect 19812 18213 19840 18244
rect 19981 18241 19993 18275
rect 20027 18241 20039 18275
rect 19981 18235 20039 18241
rect 19245 18207 19303 18213
rect 19245 18204 19257 18207
rect 15856 18176 19257 18204
rect 11241 18139 11299 18145
rect 11241 18105 11253 18139
rect 11287 18136 11299 18139
rect 15856 18136 15884 18176
rect 19245 18173 19257 18176
rect 19291 18173 19303 18207
rect 19245 18167 19303 18173
rect 19797 18207 19855 18213
rect 19797 18173 19809 18207
rect 19843 18173 19855 18207
rect 19797 18167 19855 18173
rect 20533 18207 20591 18213
rect 20533 18173 20545 18207
rect 20579 18173 20591 18207
rect 20533 18167 20591 18173
rect 11287 18108 15884 18136
rect 16568 18139 16626 18145
rect 11287 18105 11299 18108
rect 11241 18099 11299 18105
rect 16568 18105 16580 18139
rect 16614 18136 16626 18139
rect 16666 18136 16672 18148
rect 16614 18108 16672 18136
rect 16614 18105 16626 18108
rect 16568 18099 16626 18105
rect 16666 18096 16672 18108
rect 16724 18096 16730 18148
rect 18509 18139 18567 18145
rect 18509 18105 18521 18139
rect 18555 18136 18567 18139
rect 19978 18136 19984 18148
rect 18555 18108 19984 18136
rect 18555 18105 18567 18108
rect 18509 18099 18567 18105
rect 19978 18096 19984 18108
rect 20036 18096 20042 18148
rect 10652 18040 11008 18068
rect 11977 18071 12035 18077
rect 10652 18028 10658 18040
rect 11977 18037 11989 18071
rect 12023 18068 12035 18071
rect 12805 18071 12863 18077
rect 12805 18068 12817 18071
rect 12023 18040 12817 18068
rect 12023 18037 12035 18040
rect 11977 18031 12035 18037
rect 12805 18037 12817 18040
rect 12851 18037 12863 18071
rect 13262 18068 13268 18080
rect 13223 18040 13268 18068
rect 12805 18031 12863 18037
rect 13262 18028 13268 18040
rect 13320 18028 13326 18080
rect 13354 18028 13360 18080
rect 13412 18068 13418 18080
rect 15289 18071 15347 18077
rect 13412 18040 13457 18068
rect 13412 18028 13418 18040
rect 15289 18037 15301 18071
rect 15335 18068 15347 18071
rect 15470 18068 15476 18080
rect 15335 18040 15476 18068
rect 15335 18037 15347 18040
rect 15289 18031 15347 18037
rect 15470 18028 15476 18040
rect 15528 18068 15534 18080
rect 16298 18068 16304 18080
rect 15528 18040 16304 18068
rect 15528 18028 15534 18040
rect 16298 18028 16304 18040
rect 16356 18028 16362 18080
rect 18138 18068 18144 18080
rect 18099 18040 18144 18068
rect 18138 18028 18144 18040
rect 18196 18028 18202 18080
rect 18598 18068 18604 18080
rect 18559 18040 18604 18068
rect 18598 18028 18604 18040
rect 18656 18028 18662 18080
rect 18690 18028 18696 18080
rect 18748 18068 18754 18080
rect 20548 18068 20576 18167
rect 20806 18136 20812 18148
rect 20767 18108 20812 18136
rect 20806 18096 20812 18108
rect 20864 18096 20870 18148
rect 18748 18040 20576 18068
rect 18748 18028 18754 18040
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 7742 17824 7748 17876
rect 7800 17864 7806 17876
rect 8662 17864 8668 17876
rect 7800 17836 8668 17864
rect 7800 17824 7806 17836
rect 8662 17824 8668 17836
rect 8720 17824 8726 17876
rect 8846 17824 8852 17876
rect 8904 17864 8910 17876
rect 8941 17867 8999 17873
rect 8941 17864 8953 17867
rect 8904 17836 8953 17864
rect 8904 17824 8910 17836
rect 8941 17833 8953 17836
rect 8987 17833 8999 17867
rect 9674 17864 9680 17876
rect 9635 17836 9680 17864
rect 8941 17827 8999 17833
rect 9674 17824 9680 17836
rect 9732 17824 9738 17876
rect 10045 17867 10103 17873
rect 10045 17833 10057 17867
rect 10091 17864 10103 17867
rect 12894 17864 12900 17876
rect 10091 17836 12900 17864
rect 10091 17833 10103 17836
rect 10045 17827 10103 17833
rect 12894 17824 12900 17836
rect 12952 17824 12958 17876
rect 12989 17867 13047 17873
rect 12989 17833 13001 17867
rect 13035 17864 13047 17867
rect 13262 17864 13268 17876
rect 13035 17836 13268 17864
rect 13035 17833 13047 17836
rect 12989 17827 13047 17833
rect 13262 17824 13268 17836
rect 13320 17824 13326 17876
rect 15749 17867 15807 17873
rect 15749 17833 15761 17867
rect 15795 17864 15807 17867
rect 16114 17864 16120 17876
rect 15795 17836 16120 17864
rect 15795 17833 15807 17836
rect 15749 17827 15807 17833
rect 16114 17824 16120 17836
rect 16172 17824 16178 17876
rect 16390 17824 16396 17876
rect 16448 17864 16454 17876
rect 16761 17867 16819 17873
rect 16761 17864 16773 17867
rect 16448 17836 16773 17864
rect 16448 17824 16454 17836
rect 16761 17833 16773 17836
rect 16807 17833 16819 17867
rect 16761 17827 16819 17833
rect 842 17756 848 17808
rect 900 17796 906 17808
rect 8478 17796 8484 17808
rect 900 17768 8484 17796
rect 900 17756 906 17768
rect 8478 17756 8484 17768
rect 8536 17756 8542 17808
rect 9950 17756 9956 17808
rect 10008 17796 10014 17808
rect 16776 17796 16804 17827
rect 18138 17824 18144 17876
rect 18196 17864 18202 17876
rect 19153 17867 19211 17873
rect 19153 17864 19165 17867
rect 18196 17836 19165 17864
rect 18196 17824 18202 17836
rect 19153 17833 19165 17836
rect 19199 17833 19211 17867
rect 19153 17827 19211 17833
rect 19245 17867 19303 17873
rect 19245 17833 19257 17867
rect 19291 17864 19303 17867
rect 19797 17867 19855 17873
rect 19797 17864 19809 17867
rect 19291 17836 19809 17864
rect 19291 17833 19303 17836
rect 19245 17827 19303 17833
rect 19797 17833 19809 17836
rect 19843 17833 19855 17867
rect 19797 17827 19855 17833
rect 19978 17824 19984 17876
rect 20036 17864 20042 17876
rect 20901 17867 20959 17873
rect 20901 17864 20913 17867
rect 20036 17836 20913 17864
rect 20036 17824 20042 17836
rect 20901 17833 20913 17836
rect 20947 17833 20959 17867
rect 20901 17827 20959 17833
rect 17396 17799 17454 17805
rect 10008 17768 10824 17796
rect 16776 17768 17172 17796
rect 10008 17756 10014 17768
rect 7561 17731 7619 17737
rect 7561 17697 7573 17731
rect 7607 17728 7619 17731
rect 7650 17728 7656 17740
rect 7607 17700 7656 17728
rect 7607 17697 7619 17700
rect 7561 17691 7619 17697
rect 7650 17688 7656 17700
rect 7708 17688 7714 17740
rect 7828 17731 7886 17737
rect 7828 17697 7840 17731
rect 7874 17728 7886 17731
rect 8386 17728 8392 17740
rect 7874 17700 8392 17728
rect 7874 17697 7886 17700
rect 7828 17691 7886 17697
rect 8386 17688 8392 17700
rect 8444 17688 8450 17740
rect 10134 17728 10140 17740
rect 10095 17700 10140 17728
rect 10134 17688 10140 17700
rect 10192 17688 10198 17740
rect 10796 17737 10824 17768
rect 10781 17731 10839 17737
rect 10781 17697 10793 17731
rect 10827 17697 10839 17731
rect 11882 17728 11888 17740
rect 11843 17700 11888 17728
rect 10781 17691 10839 17697
rect 11882 17688 11888 17700
rect 11940 17688 11946 17740
rect 11977 17731 12035 17737
rect 11977 17697 11989 17731
rect 12023 17728 12035 17731
rect 12529 17731 12587 17737
rect 12023 17700 12480 17728
rect 12023 17697 12035 17700
rect 11977 17691 12035 17697
rect 10318 17660 10324 17672
rect 10279 17632 10324 17660
rect 10318 17620 10324 17632
rect 10376 17620 10382 17672
rect 11057 17663 11115 17669
rect 11057 17629 11069 17663
rect 11103 17629 11115 17663
rect 11057 17623 11115 17629
rect 11072 17592 11100 17623
rect 11606 17620 11612 17672
rect 11664 17660 11670 17672
rect 12069 17663 12127 17669
rect 12069 17660 12081 17663
rect 11664 17632 12081 17660
rect 11664 17620 11670 17632
rect 12069 17629 12081 17632
rect 12115 17629 12127 17663
rect 12452 17660 12480 17700
rect 12529 17697 12541 17731
rect 12575 17728 12587 17731
rect 13357 17731 13415 17737
rect 13357 17728 13369 17731
rect 12575 17700 13369 17728
rect 12575 17697 12587 17700
rect 12529 17691 12587 17697
rect 13357 17697 13369 17700
rect 13403 17697 13415 17731
rect 14550 17728 14556 17740
rect 14511 17700 14556 17728
rect 13357 17691 13415 17697
rect 14550 17688 14556 17700
rect 14608 17688 14614 17740
rect 15289 17731 15347 17737
rect 15289 17697 15301 17731
rect 15335 17728 15347 17731
rect 16117 17731 16175 17737
rect 16117 17728 16129 17731
rect 15335 17700 16129 17728
rect 15335 17697 15347 17700
rect 15289 17691 15347 17697
rect 16117 17697 16129 17700
rect 16163 17697 16175 17731
rect 16117 17691 16175 17697
rect 16224 17700 16620 17728
rect 12986 17660 12992 17672
rect 12452 17632 12992 17660
rect 12069 17623 12127 17629
rect 12986 17620 12992 17632
rect 13044 17620 13050 17672
rect 13446 17660 13452 17672
rect 13407 17632 13452 17660
rect 13446 17620 13452 17632
rect 13504 17620 13510 17672
rect 13538 17620 13544 17672
rect 13596 17660 13602 17672
rect 13596 17632 13641 17660
rect 13596 17620 13602 17632
rect 13998 17620 14004 17672
rect 14056 17660 14062 17672
rect 14645 17663 14703 17669
rect 14645 17660 14657 17663
rect 14056 17632 14657 17660
rect 14056 17620 14062 17632
rect 14645 17629 14657 17632
rect 14691 17629 14703 17663
rect 14645 17623 14703 17629
rect 14829 17663 14887 17669
rect 14829 17629 14841 17663
rect 14875 17660 14887 17663
rect 15010 17660 15016 17672
rect 14875 17632 15016 17660
rect 14875 17629 14887 17632
rect 14829 17623 14887 17629
rect 15010 17620 15016 17632
rect 15068 17620 15074 17672
rect 15930 17620 15936 17672
rect 15988 17660 15994 17672
rect 16224 17669 16252 17700
rect 16209 17663 16267 17669
rect 16209 17660 16221 17663
rect 15988 17632 16221 17660
rect 15988 17620 15994 17632
rect 16209 17629 16221 17632
rect 16255 17629 16267 17663
rect 16209 17623 16267 17629
rect 16298 17620 16304 17672
rect 16356 17660 16362 17672
rect 16592 17660 16620 17700
rect 16666 17688 16672 17740
rect 16724 17728 16730 17740
rect 17144 17737 17172 17768
rect 17396 17765 17408 17799
rect 17442 17796 17454 17799
rect 18874 17796 18880 17808
rect 17442 17768 18880 17796
rect 17442 17765 17454 17768
rect 17396 17759 17454 17765
rect 18874 17756 18880 17768
rect 18932 17796 18938 17808
rect 18932 17768 20392 17796
rect 18932 17756 18938 17768
rect 16945 17731 17003 17737
rect 16945 17728 16957 17731
rect 16724 17700 16957 17728
rect 16724 17688 16730 17700
rect 16945 17697 16957 17700
rect 16991 17697 17003 17731
rect 16945 17691 17003 17697
rect 17129 17731 17187 17737
rect 17129 17697 17141 17731
rect 17175 17697 17187 17731
rect 19150 17728 19156 17740
rect 17129 17691 17187 17697
rect 17236 17700 19156 17728
rect 17236 17660 17264 17700
rect 19150 17688 19156 17700
rect 19208 17688 19214 17740
rect 20165 17731 20223 17737
rect 20165 17728 20177 17731
rect 19352 17700 20177 17728
rect 19352 17660 19380 17700
rect 20165 17697 20177 17700
rect 20211 17697 20223 17731
rect 20165 17691 20223 17697
rect 16356 17632 16401 17660
rect 16592 17632 17264 17660
rect 18156 17632 19380 17660
rect 19429 17663 19487 17669
rect 16356 17620 16362 17632
rect 16942 17592 16948 17604
rect 11072 17564 16948 17592
rect 16942 17552 16948 17564
rect 17000 17552 17006 17604
rect 11054 17484 11060 17536
rect 11112 17524 11118 17536
rect 11517 17527 11575 17533
rect 11517 17524 11529 17527
rect 11112 17496 11529 17524
rect 11112 17484 11118 17496
rect 11517 17493 11529 17496
rect 11563 17493 11575 17527
rect 11517 17487 11575 17493
rect 14185 17527 14243 17533
rect 14185 17493 14197 17527
rect 14231 17524 14243 17527
rect 15562 17524 15568 17536
rect 14231 17496 15568 17524
rect 14231 17493 14243 17496
rect 14185 17487 14243 17493
rect 15562 17484 15568 17496
rect 15620 17484 15626 17536
rect 16482 17484 16488 17536
rect 16540 17524 16546 17536
rect 18156 17524 18184 17632
rect 19429 17629 19441 17663
rect 19475 17629 19487 17663
rect 19429 17623 19487 17629
rect 18506 17592 18512 17604
rect 18419 17564 18512 17592
rect 18506 17552 18512 17564
rect 18564 17592 18570 17604
rect 19444 17592 19472 17623
rect 19610 17620 19616 17672
rect 19668 17660 19674 17672
rect 20364 17669 20392 17768
rect 20257 17663 20315 17669
rect 20257 17660 20269 17663
rect 19668 17632 20269 17660
rect 19668 17620 19674 17632
rect 20257 17629 20269 17632
rect 20303 17629 20315 17663
rect 20257 17623 20315 17629
rect 20349 17663 20407 17669
rect 20349 17629 20361 17663
rect 20395 17629 20407 17663
rect 20349 17623 20407 17629
rect 18564 17564 19472 17592
rect 18564 17552 18570 17564
rect 16540 17496 18184 17524
rect 18785 17527 18843 17533
rect 16540 17484 16546 17496
rect 18785 17493 18797 17527
rect 18831 17524 18843 17527
rect 19426 17524 19432 17536
rect 18831 17496 19432 17524
rect 18831 17493 18843 17496
rect 18785 17487 18843 17493
rect 19426 17484 19432 17496
rect 19484 17484 19490 17536
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 8386 17320 8392 17332
rect 8347 17292 8392 17320
rect 8386 17280 8392 17292
rect 8444 17280 8450 17332
rect 8478 17280 8484 17332
rect 8536 17320 8542 17332
rect 12529 17323 12587 17329
rect 8536 17292 11928 17320
rect 8536 17280 8542 17292
rect 8404 17184 8432 17280
rect 8846 17212 8852 17264
rect 8904 17252 8910 17264
rect 8904 17224 10272 17252
rect 8904 17212 8910 17224
rect 8754 17184 8760 17196
rect 8404 17156 8760 17184
rect 8754 17144 8760 17156
rect 8812 17184 8818 17196
rect 10244 17193 10272 17224
rect 9217 17187 9275 17193
rect 9217 17184 9229 17187
rect 8812 17156 9229 17184
rect 8812 17144 8818 17156
rect 9217 17153 9229 17156
rect 9263 17153 9275 17187
rect 9217 17147 9275 17153
rect 10229 17187 10287 17193
rect 10229 17153 10241 17187
rect 10275 17153 10287 17187
rect 10229 17147 10287 17153
rect 10686 17144 10692 17196
rect 10744 17184 10750 17196
rect 11333 17187 11391 17193
rect 11333 17184 11345 17187
rect 10744 17156 11345 17184
rect 10744 17144 10750 17156
rect 11333 17153 11345 17156
rect 11379 17184 11391 17187
rect 11698 17184 11704 17196
rect 11379 17156 11704 17184
rect 11379 17153 11391 17156
rect 11333 17147 11391 17153
rect 11698 17144 11704 17156
rect 11756 17144 11762 17196
rect 7009 17119 7067 17125
rect 7009 17085 7021 17119
rect 7055 17116 7067 17119
rect 8662 17116 8668 17128
rect 7055 17088 8668 17116
rect 7055 17085 7067 17088
rect 7009 17079 7067 17085
rect 8662 17076 8668 17088
rect 8720 17076 8726 17128
rect 9306 17076 9312 17128
rect 9364 17116 9370 17128
rect 9364 17088 10548 17116
rect 9364 17076 9370 17088
rect 7276 17051 7334 17057
rect 7276 17017 7288 17051
rect 7322 17048 7334 17051
rect 7650 17048 7656 17060
rect 7322 17020 7656 17048
rect 7322 17017 7334 17020
rect 7276 17011 7334 17017
rect 7650 17008 7656 17020
rect 7708 17008 7714 17060
rect 10045 17051 10103 17057
rect 10045 17048 10057 17051
rect 8680 17020 10057 17048
rect 8680 16989 8708 17020
rect 10045 17017 10057 17020
rect 10091 17017 10103 17051
rect 10520 17048 10548 17088
rect 10594 17076 10600 17128
rect 10652 17116 10658 17128
rect 11514 17116 11520 17128
rect 10652 17088 11520 17116
rect 10652 17076 10658 17088
rect 11514 17076 11520 17088
rect 11572 17076 11578 17128
rect 11606 17076 11612 17128
rect 11664 17116 11670 17128
rect 11793 17119 11851 17125
rect 11793 17116 11805 17119
rect 11664 17088 11805 17116
rect 11664 17076 11670 17088
rect 11793 17085 11805 17088
rect 11839 17085 11851 17119
rect 11900 17116 11928 17292
rect 12529 17289 12541 17323
rect 12575 17320 12587 17323
rect 13354 17320 13360 17332
rect 12575 17292 13360 17320
rect 12575 17289 12587 17292
rect 12529 17283 12587 17289
rect 13354 17280 13360 17292
rect 13412 17280 13418 17332
rect 13648 17292 14504 17320
rect 11977 17255 12035 17261
rect 11977 17221 11989 17255
rect 12023 17252 12035 17255
rect 13648 17252 13676 17292
rect 12023 17224 13676 17252
rect 13725 17255 13783 17261
rect 12023 17221 12035 17224
rect 11977 17215 12035 17221
rect 13725 17221 13737 17255
rect 13771 17252 13783 17255
rect 13998 17252 14004 17264
rect 13771 17224 14004 17252
rect 13771 17221 13783 17224
rect 13725 17215 13783 17221
rect 13998 17212 14004 17224
rect 14056 17212 14062 17264
rect 14476 17252 14504 17292
rect 14550 17280 14556 17332
rect 14608 17320 14614 17332
rect 14737 17323 14795 17329
rect 14737 17320 14749 17323
rect 14608 17292 14749 17320
rect 14608 17280 14614 17292
rect 14737 17289 14749 17292
rect 14783 17289 14795 17323
rect 14737 17283 14795 17289
rect 15749 17323 15807 17329
rect 15749 17289 15761 17323
rect 15795 17320 15807 17323
rect 16206 17320 16212 17332
rect 15795 17292 16212 17320
rect 15795 17289 15807 17292
rect 15749 17283 15807 17289
rect 16206 17280 16212 17292
rect 16264 17280 16270 17332
rect 22462 17320 22468 17332
rect 16316 17292 22468 17320
rect 16316 17252 16344 17292
rect 22462 17280 22468 17292
rect 22520 17280 22526 17332
rect 14476 17224 16344 17252
rect 17037 17255 17095 17261
rect 17037 17221 17049 17255
rect 17083 17252 17095 17255
rect 18046 17252 18052 17264
rect 17083 17224 18052 17252
rect 17083 17221 17095 17224
rect 17037 17215 17095 17221
rect 18046 17212 18052 17224
rect 18104 17212 18110 17264
rect 12158 17144 12164 17196
rect 12216 17184 12222 17196
rect 12989 17187 13047 17193
rect 12989 17184 13001 17187
rect 12216 17156 13001 17184
rect 12216 17144 12222 17156
rect 12989 17153 13001 17156
rect 13035 17153 13047 17187
rect 12989 17147 13047 17153
rect 13173 17187 13231 17193
rect 13173 17153 13185 17187
rect 13219 17184 13231 17187
rect 13538 17184 13544 17196
rect 13219 17156 13544 17184
rect 13219 17153 13231 17156
rect 13173 17147 13231 17153
rect 13538 17144 13544 17156
rect 13596 17144 13602 17196
rect 14369 17187 14427 17193
rect 14369 17153 14381 17187
rect 14415 17184 14427 17187
rect 14458 17184 14464 17196
rect 14415 17156 14464 17184
rect 14415 17153 14427 17156
rect 14369 17147 14427 17153
rect 14458 17144 14464 17156
rect 14516 17184 14522 17196
rect 15381 17187 15439 17193
rect 15381 17184 15393 17187
rect 14516 17156 15393 17184
rect 14516 17144 14522 17156
rect 15381 17153 15393 17156
rect 15427 17153 15439 17187
rect 16298 17184 16304 17196
rect 16259 17156 16304 17184
rect 15381 17147 15439 17153
rect 14185 17119 14243 17125
rect 14185 17116 14197 17119
rect 11900 17088 14197 17116
rect 11793 17079 11851 17085
rect 14185 17085 14197 17088
rect 14231 17085 14243 17119
rect 15396 17116 15424 17147
rect 16298 17144 16304 17156
rect 16356 17144 16362 17196
rect 19981 17187 20039 17193
rect 19981 17153 19993 17187
rect 20027 17184 20039 17187
rect 20714 17184 20720 17196
rect 20027 17156 20720 17184
rect 20027 17153 20039 17156
rect 19981 17147 20039 17153
rect 20714 17144 20720 17156
rect 20772 17144 20778 17196
rect 16390 17116 16396 17128
rect 15396 17088 16396 17116
rect 14185 17079 14243 17085
rect 16390 17076 16396 17088
rect 16448 17076 16454 17128
rect 16758 17076 16764 17128
rect 16816 17116 16822 17128
rect 16853 17119 16911 17125
rect 16853 17116 16865 17119
rect 16816 17088 16865 17116
rect 16816 17076 16822 17088
rect 16853 17085 16865 17088
rect 16899 17085 16911 17119
rect 16853 17079 16911 17085
rect 17405 17119 17463 17125
rect 17405 17085 17417 17119
rect 17451 17116 17463 17119
rect 17954 17116 17960 17128
rect 17451 17088 17960 17116
rect 17451 17085 17463 17088
rect 17405 17079 17463 17085
rect 17954 17076 17960 17088
rect 18012 17076 18018 17128
rect 18049 17119 18107 17125
rect 18049 17085 18061 17119
rect 18095 17085 18107 17119
rect 18049 17079 18107 17085
rect 11149 17051 11207 17057
rect 10520 17020 10916 17048
rect 10045 17011 10103 17017
rect 8665 16983 8723 16989
rect 8665 16949 8677 16983
rect 8711 16949 8723 16983
rect 9030 16980 9036 16992
rect 8991 16952 9036 16980
rect 8665 16943 8723 16949
rect 9030 16940 9036 16952
rect 9088 16940 9094 16992
rect 9125 16983 9183 16989
rect 9125 16949 9137 16983
rect 9171 16980 9183 16983
rect 9306 16980 9312 16992
rect 9171 16952 9312 16980
rect 9171 16949 9183 16952
rect 9125 16943 9183 16949
rect 9306 16940 9312 16952
rect 9364 16940 9370 16992
rect 9677 16983 9735 16989
rect 9677 16949 9689 16983
rect 9723 16980 9735 16983
rect 9766 16980 9772 16992
rect 9723 16952 9772 16980
rect 9723 16949 9735 16952
rect 9677 16943 9735 16949
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 9858 16940 9864 16992
rect 9916 16980 9922 16992
rect 10137 16983 10195 16989
rect 10137 16980 10149 16983
rect 9916 16952 10149 16980
rect 9916 16940 9922 16952
rect 10137 16949 10149 16952
rect 10183 16949 10195 16983
rect 10778 16980 10784 16992
rect 10739 16952 10784 16980
rect 10137 16943 10195 16949
rect 10778 16940 10784 16952
rect 10836 16940 10842 16992
rect 10888 16980 10916 17020
rect 11149 17017 11161 17051
rect 11195 17048 11207 17051
rect 15105 17051 15163 17057
rect 15105 17048 15117 17051
rect 11195 17020 12940 17048
rect 11195 17017 11207 17020
rect 11149 17011 11207 17017
rect 11238 16980 11244 16992
rect 10888 16952 11244 16980
rect 11238 16940 11244 16952
rect 11296 16940 11302 16992
rect 12912 16989 12940 17020
rect 13464 17020 15117 17048
rect 13464 16992 13492 17020
rect 15105 17017 15117 17020
rect 15151 17017 15163 17051
rect 15105 17011 15163 17017
rect 15654 17008 15660 17060
rect 15712 17048 15718 17060
rect 15712 17020 16252 17048
rect 15712 17008 15718 17020
rect 12897 16983 12955 16989
rect 12897 16949 12909 16983
rect 12943 16980 12955 16983
rect 13446 16980 13452 16992
rect 12943 16952 13452 16980
rect 12943 16949 12955 16952
rect 12897 16943 12955 16949
rect 13446 16940 13452 16952
rect 13504 16940 13510 16992
rect 13814 16940 13820 16992
rect 13872 16980 13878 16992
rect 14093 16983 14151 16989
rect 14093 16980 14105 16983
rect 13872 16952 14105 16980
rect 13872 16940 13878 16952
rect 14093 16949 14105 16952
rect 14139 16980 14151 16983
rect 14182 16980 14188 16992
rect 14139 16952 14188 16980
rect 14139 16949 14151 16952
rect 14093 16943 14151 16949
rect 14182 16940 14188 16952
rect 14240 16940 14246 16992
rect 14366 16940 14372 16992
rect 14424 16980 14430 16992
rect 15197 16983 15255 16989
rect 15197 16980 15209 16983
rect 14424 16952 15209 16980
rect 14424 16940 14430 16952
rect 15197 16949 15209 16952
rect 15243 16949 15255 16983
rect 15197 16943 15255 16949
rect 15470 16940 15476 16992
rect 15528 16980 15534 16992
rect 16224 16989 16252 17020
rect 17770 17008 17776 17060
rect 17828 17048 17834 17060
rect 18064 17048 18092 17079
rect 19426 17076 19432 17128
rect 19484 17116 19490 17128
rect 19705 17119 19763 17125
rect 19705 17116 19717 17119
rect 19484 17088 19717 17116
rect 19484 17076 19490 17088
rect 19705 17085 19717 17088
rect 19751 17085 19763 17119
rect 20438 17116 20444 17128
rect 20399 17088 20444 17116
rect 19705 17079 19763 17085
rect 20438 17076 20444 17088
rect 20496 17076 20502 17128
rect 17828 17020 18092 17048
rect 18316 17051 18374 17057
rect 17828 17008 17834 17020
rect 18316 17017 18328 17051
rect 18362 17048 18374 17051
rect 18506 17048 18512 17060
rect 18362 17020 18512 17048
rect 18362 17017 18374 17020
rect 18316 17011 18374 17017
rect 18506 17008 18512 17020
rect 18564 17008 18570 17060
rect 19518 17008 19524 17060
rect 19576 17048 19582 17060
rect 20717 17051 20775 17057
rect 20717 17048 20729 17051
rect 19576 17020 20729 17048
rect 19576 17008 19582 17020
rect 20717 17017 20729 17020
rect 20763 17017 20775 17051
rect 20717 17011 20775 17017
rect 16117 16983 16175 16989
rect 16117 16980 16129 16983
rect 15528 16952 16129 16980
rect 15528 16940 15534 16952
rect 16117 16949 16129 16952
rect 16163 16949 16175 16983
rect 16117 16943 16175 16949
rect 16209 16983 16267 16989
rect 16209 16949 16221 16983
rect 16255 16980 16267 16983
rect 16298 16980 16304 16992
rect 16255 16952 16304 16980
rect 16255 16949 16267 16952
rect 16209 16943 16267 16949
rect 16298 16940 16304 16952
rect 16356 16940 16362 16992
rect 17589 16983 17647 16989
rect 17589 16949 17601 16983
rect 17635 16980 17647 16983
rect 17954 16980 17960 16992
rect 17635 16952 17960 16980
rect 17635 16949 17647 16952
rect 17589 16943 17647 16949
rect 17954 16940 17960 16952
rect 18012 16940 18018 16992
rect 19334 16940 19340 16992
rect 19392 16980 19398 16992
rect 19429 16983 19487 16989
rect 19429 16980 19441 16983
rect 19392 16952 19441 16980
rect 19392 16940 19398 16952
rect 19429 16949 19441 16952
rect 19475 16949 19487 16983
rect 19429 16943 19487 16949
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 6914 16736 6920 16788
rect 6972 16776 6978 16788
rect 7377 16779 7435 16785
rect 7377 16776 7389 16779
rect 6972 16748 7389 16776
rect 6972 16736 6978 16748
rect 7377 16745 7389 16748
rect 7423 16745 7435 16779
rect 7377 16739 7435 16745
rect 7466 16736 7472 16788
rect 7524 16776 7530 16788
rect 7742 16776 7748 16788
rect 7524 16748 7748 16776
rect 7524 16736 7530 16748
rect 7742 16736 7748 16748
rect 7800 16736 7806 16788
rect 8205 16779 8263 16785
rect 8205 16745 8217 16779
rect 8251 16776 8263 16779
rect 9858 16776 9864 16788
rect 8251 16748 9864 16776
rect 8251 16745 8263 16748
rect 8205 16739 8263 16745
rect 9858 16736 9864 16748
rect 9916 16736 9922 16788
rect 9968 16748 11100 16776
rect 9968 16717 9996 16748
rect 8665 16711 8723 16717
rect 8665 16708 8677 16711
rect 7024 16680 8677 16708
rect 7024 16513 7052 16680
rect 8665 16677 8677 16680
rect 8711 16677 8723 16711
rect 8665 16671 8723 16677
rect 9953 16711 10011 16717
rect 9953 16677 9965 16711
rect 9999 16677 10011 16711
rect 11072 16708 11100 16748
rect 11514 16736 11520 16788
rect 11572 16776 11578 16788
rect 11793 16779 11851 16785
rect 11793 16776 11805 16779
rect 11572 16748 11805 16776
rect 11572 16736 11578 16748
rect 11793 16745 11805 16748
rect 11839 16745 11851 16779
rect 11793 16739 11851 16745
rect 11882 16736 11888 16788
rect 11940 16776 11946 16788
rect 12069 16779 12127 16785
rect 12069 16776 12081 16779
rect 11940 16748 12081 16776
rect 11940 16736 11946 16748
rect 12069 16745 12081 16748
rect 12115 16745 12127 16779
rect 16206 16776 16212 16788
rect 12069 16739 12127 16745
rect 12176 16748 16212 16776
rect 12176 16708 12204 16748
rect 16206 16736 16212 16748
rect 16264 16736 16270 16788
rect 17129 16779 17187 16785
rect 17129 16745 17141 16779
rect 17175 16776 17187 16779
rect 17957 16779 18015 16785
rect 17175 16748 17816 16776
rect 17175 16745 17187 16748
rect 17129 16739 17187 16745
rect 11072 16680 12204 16708
rect 12437 16711 12495 16717
rect 9953 16671 10011 16677
rect 12437 16677 12449 16711
rect 12483 16708 12495 16711
rect 13081 16711 13139 16717
rect 13081 16708 13093 16711
rect 12483 16680 13093 16708
rect 12483 16677 12495 16680
rect 12437 16671 12495 16677
rect 13081 16677 13093 16680
rect 13127 16677 13139 16711
rect 13081 16671 13139 16677
rect 13808 16711 13866 16717
rect 13808 16677 13820 16711
rect 13854 16708 13866 16711
rect 14458 16708 14464 16720
rect 13854 16680 14464 16708
rect 13854 16677 13866 16680
rect 13808 16671 13866 16677
rect 14458 16668 14464 16680
rect 14516 16668 14522 16720
rect 15289 16711 15347 16717
rect 15289 16677 15301 16711
rect 15335 16708 15347 16711
rect 17034 16708 17040 16720
rect 15335 16680 17040 16708
rect 15335 16677 15347 16680
rect 15289 16671 15347 16677
rect 17034 16668 17040 16680
rect 17092 16668 17098 16720
rect 8573 16643 8631 16649
rect 8573 16609 8585 16643
rect 8619 16640 8631 16643
rect 9214 16640 9220 16652
rect 8619 16612 9220 16640
rect 8619 16609 8631 16612
rect 8573 16603 8631 16609
rect 9214 16600 9220 16612
rect 9272 16600 9278 16652
rect 9490 16640 9496 16652
rect 9451 16612 9496 16640
rect 9490 16600 9496 16612
rect 9548 16600 9554 16652
rect 9674 16640 9680 16652
rect 9635 16612 9680 16640
rect 9674 16600 9680 16612
rect 9732 16600 9738 16652
rect 10686 16649 10692 16652
rect 10680 16603 10692 16649
rect 10744 16640 10750 16652
rect 13541 16643 13599 16649
rect 10744 16612 10780 16640
rect 10686 16600 10692 16603
rect 10744 16600 10750 16612
rect 13541 16609 13553 16643
rect 13587 16640 13599 16643
rect 13630 16640 13636 16652
rect 13587 16612 13636 16640
rect 13587 16609 13599 16612
rect 13541 16603 13599 16609
rect 13630 16600 13636 16612
rect 13688 16600 13694 16652
rect 16114 16640 16120 16652
rect 15120 16612 16120 16640
rect 7650 16572 7656 16584
rect 7563 16544 7656 16572
rect 7650 16532 7656 16544
rect 7708 16572 7714 16584
rect 8202 16572 8208 16584
rect 7708 16544 8208 16572
rect 7708 16532 7714 16544
rect 8202 16532 8208 16544
rect 8260 16532 8266 16584
rect 8754 16572 8760 16584
rect 8715 16544 8760 16572
rect 8754 16532 8760 16544
rect 8812 16532 8818 16584
rect 10318 16532 10324 16584
rect 10376 16572 10382 16584
rect 10413 16575 10471 16581
rect 10413 16572 10425 16575
rect 10376 16544 10425 16572
rect 10376 16532 10382 16544
rect 10413 16541 10425 16544
rect 10459 16541 10471 16575
rect 10413 16535 10471 16541
rect 7009 16507 7067 16513
rect 7009 16473 7021 16507
rect 7055 16473 7067 16507
rect 7009 16467 7067 16473
rect 8662 16464 8668 16516
rect 8720 16504 8726 16516
rect 9309 16507 9367 16513
rect 9309 16504 9321 16507
rect 8720 16476 9321 16504
rect 8720 16464 8726 16476
rect 9309 16473 9321 16476
rect 9355 16504 9367 16507
rect 9398 16504 9404 16516
rect 9355 16476 9404 16504
rect 9355 16473 9367 16476
rect 9309 16467 9367 16473
rect 9398 16464 9404 16476
rect 9456 16464 9462 16516
rect 10428 16436 10456 16535
rect 12250 16532 12256 16584
rect 12308 16572 12314 16584
rect 12529 16575 12587 16581
rect 12529 16572 12541 16575
rect 12308 16544 12541 16572
rect 12308 16532 12314 16544
rect 12529 16541 12541 16544
rect 12575 16541 12587 16575
rect 12529 16535 12587 16541
rect 12621 16575 12679 16581
rect 12621 16541 12633 16575
rect 12667 16541 12679 16575
rect 15120 16572 15148 16612
rect 16114 16600 16120 16612
rect 16172 16600 16178 16652
rect 16209 16643 16267 16649
rect 16209 16609 16221 16643
rect 16255 16640 16267 16643
rect 16482 16640 16488 16652
rect 16255 16612 16488 16640
rect 16255 16609 16267 16612
rect 16209 16603 16267 16609
rect 12621 16535 12679 16541
rect 14568 16544 15148 16572
rect 12342 16464 12348 16516
rect 12400 16504 12406 16516
rect 12636 16504 12664 16535
rect 12400 16476 12664 16504
rect 12400 16464 12406 16476
rect 12434 16436 12440 16448
rect 10428 16408 12440 16436
rect 12434 16396 12440 16408
rect 12492 16396 12498 16448
rect 13722 16396 13728 16448
rect 13780 16436 13786 16448
rect 14568 16436 14596 16544
rect 15194 16532 15200 16584
rect 15252 16572 15258 16584
rect 16022 16572 16028 16584
rect 15252 16544 16028 16572
rect 15252 16532 15258 16544
rect 16022 16532 16028 16544
rect 16080 16572 16086 16584
rect 16224 16572 16252 16603
rect 16482 16600 16488 16612
rect 16540 16600 16546 16652
rect 16942 16640 16948 16652
rect 16903 16612 16948 16640
rect 16942 16600 16948 16612
rect 17000 16600 17006 16652
rect 17788 16640 17816 16748
rect 17957 16745 17969 16779
rect 18003 16776 18015 16779
rect 18509 16779 18567 16785
rect 18509 16776 18521 16779
rect 18003 16748 18521 16776
rect 18003 16745 18015 16748
rect 17957 16739 18015 16745
rect 18509 16745 18521 16748
rect 18555 16745 18567 16779
rect 18966 16776 18972 16788
rect 18927 16748 18972 16776
rect 18509 16739 18567 16745
rect 18966 16736 18972 16748
rect 19024 16736 19030 16788
rect 19521 16779 19579 16785
rect 19521 16745 19533 16779
rect 19567 16745 19579 16779
rect 19521 16739 19579 16745
rect 17865 16711 17923 16717
rect 17865 16677 17877 16711
rect 17911 16708 17923 16711
rect 19536 16708 19564 16739
rect 19981 16711 20039 16717
rect 19981 16708 19993 16711
rect 17911 16680 19564 16708
rect 19628 16680 19993 16708
rect 17911 16677 17923 16680
rect 17865 16671 17923 16677
rect 17954 16640 17960 16652
rect 17788 16612 17960 16640
rect 17954 16600 17960 16612
rect 18012 16600 18018 16652
rect 18598 16640 18604 16652
rect 18064 16612 18604 16640
rect 16390 16572 16396 16584
rect 16080 16544 16252 16572
rect 16351 16544 16396 16572
rect 16080 16532 16086 16544
rect 16390 16532 16396 16544
rect 16448 16532 16454 16584
rect 17497 16507 17555 16513
rect 17497 16473 17509 16507
rect 17543 16504 17555 16507
rect 18064 16504 18092 16612
rect 18598 16600 18604 16612
rect 18656 16600 18662 16652
rect 18877 16643 18935 16649
rect 18877 16609 18889 16643
rect 18923 16609 18935 16643
rect 18877 16603 18935 16609
rect 18141 16575 18199 16581
rect 18141 16541 18153 16575
rect 18187 16572 18199 16575
rect 18690 16572 18696 16584
rect 18187 16544 18696 16572
rect 18187 16541 18199 16544
rect 18141 16535 18199 16541
rect 18690 16532 18696 16544
rect 18748 16532 18754 16584
rect 17543 16476 18092 16504
rect 17543 16473 17555 16476
rect 17497 16467 17555 16473
rect 13780 16408 14596 16436
rect 14921 16439 14979 16445
rect 13780 16396 13786 16408
rect 14921 16405 14933 16439
rect 14967 16436 14979 16439
rect 15010 16436 15016 16448
rect 14967 16408 15016 16436
rect 14967 16405 14979 16408
rect 14921 16399 14979 16405
rect 15010 16396 15016 16408
rect 15068 16396 15074 16448
rect 15746 16436 15752 16448
rect 15707 16408 15752 16436
rect 15746 16396 15752 16408
rect 15804 16396 15810 16448
rect 16942 16396 16948 16448
rect 17000 16436 17006 16448
rect 18892 16436 18920 16603
rect 19058 16600 19064 16652
rect 19116 16640 19122 16652
rect 19628 16640 19656 16680
rect 19981 16677 19993 16680
rect 20027 16677 20039 16711
rect 19981 16671 20039 16677
rect 19886 16640 19892 16652
rect 19116 16612 19656 16640
rect 19847 16612 19892 16640
rect 19116 16600 19122 16612
rect 19886 16600 19892 16612
rect 19944 16600 19950 16652
rect 19153 16575 19211 16581
rect 19153 16541 19165 16575
rect 19199 16572 19211 16575
rect 19334 16572 19340 16584
rect 19199 16544 19340 16572
rect 19199 16541 19211 16544
rect 19153 16535 19211 16541
rect 19334 16532 19340 16544
rect 19392 16532 19398 16584
rect 20073 16575 20131 16581
rect 20073 16541 20085 16575
rect 20119 16541 20131 16575
rect 20073 16535 20131 16541
rect 19352 16504 19380 16532
rect 20088 16504 20116 16535
rect 19352 16476 20116 16504
rect 17000 16408 18920 16436
rect 17000 16396 17006 16408
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 8202 16232 8208 16244
rect 8163 16204 8208 16232
rect 8202 16192 8208 16204
rect 8260 16192 8266 16244
rect 9766 16232 9772 16244
rect 9232 16204 9772 16232
rect 8662 16056 8668 16108
rect 8720 16056 8726 16108
rect 6825 16031 6883 16037
rect 6825 15997 6837 16031
rect 6871 16028 6883 16031
rect 7558 16028 7564 16040
rect 6871 16000 7564 16028
rect 6871 15997 6883 16000
rect 6825 15991 6883 15997
rect 7558 15988 7564 16000
rect 7616 16028 7622 16040
rect 8680 16028 8708 16056
rect 7616 16000 8708 16028
rect 8757 16031 8815 16037
rect 7616 15988 7622 16000
rect 8757 15997 8769 16031
rect 8803 16028 8815 16031
rect 9232 16028 9260 16204
rect 9766 16192 9772 16204
rect 9824 16192 9830 16244
rect 11698 16192 11704 16244
rect 11756 16232 11762 16244
rect 12342 16232 12348 16244
rect 11756 16204 12348 16232
rect 11756 16192 11762 16204
rect 12342 16192 12348 16204
rect 12400 16232 12406 16244
rect 13538 16232 13544 16244
rect 12400 16204 13544 16232
rect 12400 16192 12406 16204
rect 13538 16192 13544 16204
rect 13596 16232 13602 16244
rect 13817 16235 13875 16241
rect 13817 16232 13829 16235
rect 13596 16204 13829 16232
rect 13596 16192 13602 16204
rect 13817 16201 13829 16204
rect 13863 16201 13875 16235
rect 13817 16195 13875 16201
rect 15010 16192 15016 16244
rect 15068 16232 15074 16244
rect 15068 16204 16344 16232
rect 15068 16192 15074 16204
rect 15473 16167 15531 16173
rect 15473 16133 15485 16167
rect 15519 16164 15531 16167
rect 15838 16164 15844 16176
rect 15519 16136 15844 16164
rect 15519 16133 15531 16136
rect 15473 16127 15531 16133
rect 15838 16124 15844 16136
rect 15896 16124 15902 16176
rect 9398 16056 9404 16108
rect 9456 16096 9462 16108
rect 9493 16099 9551 16105
rect 9493 16096 9505 16099
rect 9456 16068 9505 16096
rect 9456 16056 9462 16068
rect 9493 16065 9505 16068
rect 9539 16065 9551 16099
rect 9493 16059 9551 16065
rect 10686 16056 10692 16108
rect 10744 16096 10750 16108
rect 10962 16096 10968 16108
rect 10744 16068 10968 16096
rect 10744 16056 10750 16068
rect 10962 16056 10968 16068
rect 11020 16056 11026 16108
rect 11698 16096 11704 16108
rect 11659 16068 11704 16096
rect 11698 16056 11704 16068
rect 11756 16056 11762 16108
rect 12434 16096 12440 16108
rect 12395 16068 12440 16096
rect 12434 16056 12440 16068
rect 12492 16056 12498 16108
rect 13630 16056 13636 16108
rect 13688 16096 13694 16108
rect 13688 16068 14044 16096
rect 13688 16056 13694 16068
rect 14016 16040 14044 16068
rect 15746 16056 15752 16108
rect 15804 16096 15810 16108
rect 16316 16105 16344 16204
rect 16482 16192 16488 16244
rect 16540 16232 16546 16244
rect 17770 16232 17776 16244
rect 16540 16204 17776 16232
rect 16540 16192 16546 16204
rect 17770 16192 17776 16204
rect 17828 16232 17834 16244
rect 17828 16204 17908 16232
rect 17828 16192 17834 16204
rect 16577 16167 16635 16173
rect 16577 16133 16589 16167
rect 16623 16164 16635 16167
rect 16761 16167 16819 16173
rect 16761 16164 16773 16167
rect 16623 16136 16773 16164
rect 16623 16133 16635 16136
rect 16577 16127 16635 16133
rect 16761 16133 16773 16136
rect 16807 16133 16819 16167
rect 16761 16127 16819 16133
rect 16209 16099 16267 16105
rect 16209 16096 16221 16099
rect 15804 16068 16221 16096
rect 15804 16056 15810 16068
rect 16209 16065 16221 16068
rect 16255 16065 16267 16099
rect 16209 16059 16267 16065
rect 16301 16099 16359 16105
rect 16301 16065 16313 16099
rect 16347 16065 16359 16099
rect 16301 16059 16359 16065
rect 16390 16056 16396 16108
rect 16448 16096 16454 16108
rect 17405 16099 17463 16105
rect 17405 16096 17417 16099
rect 16448 16068 17417 16096
rect 16448 16056 16454 16068
rect 17405 16065 17417 16068
rect 17451 16096 17463 16099
rect 17770 16096 17776 16108
rect 17451 16068 17776 16096
rect 17451 16065 17463 16068
rect 17405 16059 17463 16065
rect 17770 16056 17776 16068
rect 17828 16056 17834 16108
rect 17880 16096 17908 16204
rect 18046 16096 18052 16108
rect 17880 16068 18052 16096
rect 18046 16056 18052 16068
rect 18104 16056 18110 16108
rect 20346 16096 20352 16108
rect 20307 16068 20352 16096
rect 20346 16056 20352 16068
rect 20404 16056 20410 16108
rect 8803 16000 9260 16028
rect 9692 16000 13952 16028
rect 8803 15997 8815 16000
rect 8757 15991 8815 15997
rect 7092 15963 7150 15969
rect 7092 15929 7104 15963
rect 7138 15960 7150 15963
rect 8662 15960 8668 15972
rect 7138 15932 8668 15960
rect 7138 15929 7150 15932
rect 7092 15923 7150 15929
rect 8662 15920 8668 15932
rect 8720 15920 8726 15972
rect 9033 15963 9091 15969
rect 9033 15929 9045 15963
rect 9079 15960 9091 15963
rect 9692 15960 9720 16000
rect 9079 15932 9720 15960
rect 9760 15963 9818 15969
rect 9079 15929 9091 15932
rect 9033 15923 9091 15929
rect 9760 15929 9772 15963
rect 9806 15960 9818 15963
rect 10594 15960 10600 15972
rect 9806 15932 10600 15960
rect 9806 15929 9818 15932
rect 9760 15923 9818 15929
rect 10594 15920 10600 15932
rect 10652 15920 10658 15972
rect 12710 15969 12716 15972
rect 11609 15963 11667 15969
rect 11609 15960 11621 15963
rect 10704 15932 11621 15960
rect 10042 15852 10048 15904
rect 10100 15892 10106 15904
rect 10704 15892 10732 15932
rect 11609 15929 11621 15932
rect 11655 15929 11667 15963
rect 12704 15960 12716 15969
rect 12671 15932 12716 15960
rect 11609 15923 11667 15929
rect 12704 15923 12716 15932
rect 12710 15920 12716 15923
rect 12768 15920 12774 15972
rect 13924 15960 13952 16000
rect 13998 15988 14004 16040
rect 14056 16028 14062 16040
rect 14093 16031 14151 16037
rect 14093 16028 14105 16031
rect 14056 16000 14105 16028
rect 14056 15988 14062 16000
rect 14093 15997 14105 16000
rect 14139 15997 14151 16031
rect 14093 15991 14151 15997
rect 14200 16000 16896 16028
rect 14200 15960 14228 16000
rect 13924 15932 14228 15960
rect 14360 15963 14418 15969
rect 14360 15929 14372 15963
rect 14406 15960 14418 15963
rect 15010 15960 15016 15972
rect 14406 15932 15016 15960
rect 14406 15929 14418 15932
rect 14360 15923 14418 15929
rect 15010 15920 15016 15932
rect 15068 15920 15074 15972
rect 16117 15963 16175 15969
rect 15304 15932 15884 15960
rect 10100 15864 10732 15892
rect 10873 15895 10931 15901
rect 10100 15852 10106 15864
rect 10873 15861 10885 15895
rect 10919 15892 10931 15895
rect 10962 15892 10968 15904
rect 10919 15864 10968 15892
rect 10919 15861 10931 15864
rect 10873 15855 10931 15861
rect 10962 15852 10968 15864
rect 11020 15852 11026 15904
rect 11146 15892 11152 15904
rect 11107 15864 11152 15892
rect 11146 15852 11152 15864
rect 11204 15852 11210 15904
rect 11517 15895 11575 15901
rect 11517 15861 11529 15895
rect 11563 15892 11575 15895
rect 12526 15892 12532 15904
rect 11563 15864 12532 15892
rect 11563 15861 11575 15864
rect 11517 15855 11575 15861
rect 12526 15852 12532 15864
rect 12584 15892 12590 15904
rect 13262 15892 13268 15904
rect 12584 15864 13268 15892
rect 12584 15852 12590 15864
rect 13262 15852 13268 15864
rect 13320 15852 13326 15904
rect 13814 15852 13820 15904
rect 13872 15892 13878 15904
rect 15304 15892 15332 15932
rect 13872 15864 15332 15892
rect 13872 15852 13878 15864
rect 15654 15852 15660 15904
rect 15712 15892 15718 15904
rect 15749 15895 15807 15901
rect 15749 15892 15761 15895
rect 15712 15864 15761 15892
rect 15712 15852 15718 15864
rect 15749 15861 15761 15864
rect 15795 15861 15807 15895
rect 15856 15892 15884 15932
rect 16117 15929 16129 15963
rect 16163 15960 16175 15963
rect 16577 15963 16635 15969
rect 16577 15960 16589 15963
rect 16163 15932 16589 15960
rect 16163 15929 16175 15932
rect 16117 15923 16175 15929
rect 16577 15929 16589 15932
rect 16623 15929 16635 15963
rect 16868 15960 16896 16000
rect 17034 15988 17040 16040
rect 17092 16028 17098 16040
rect 17129 16031 17187 16037
rect 17129 16028 17141 16031
rect 17092 16000 17141 16028
rect 17092 15988 17098 16000
rect 17129 15997 17141 16000
rect 17175 15997 17187 16031
rect 20809 16031 20867 16037
rect 20809 16028 20821 16031
rect 17129 15991 17187 15997
rect 17236 16000 20821 16028
rect 17236 15960 17264 16000
rect 20809 15997 20821 16000
rect 20855 15997 20867 16031
rect 20809 15991 20867 15997
rect 16868 15932 17264 15960
rect 18316 15963 18374 15969
rect 16577 15923 16635 15929
rect 18316 15929 18328 15963
rect 18362 15960 18374 15963
rect 19334 15960 19340 15972
rect 18362 15932 19340 15960
rect 18362 15929 18374 15932
rect 18316 15923 18374 15929
rect 19334 15920 19340 15932
rect 19392 15920 19398 15972
rect 19610 15920 19616 15972
rect 19668 15960 19674 15972
rect 20162 15960 20168 15972
rect 19668 15932 19932 15960
rect 20075 15932 20168 15960
rect 19668 15920 19674 15932
rect 17221 15895 17279 15901
rect 17221 15892 17233 15895
rect 15856 15864 17233 15892
rect 15749 15855 15807 15861
rect 17221 15861 17233 15864
rect 17267 15861 17279 15895
rect 17221 15855 17279 15861
rect 18690 15852 18696 15904
rect 18748 15892 18754 15904
rect 19429 15895 19487 15901
rect 19429 15892 19441 15895
rect 18748 15864 19441 15892
rect 18748 15852 18754 15864
rect 19429 15861 19441 15864
rect 19475 15861 19487 15895
rect 19794 15892 19800 15904
rect 19755 15864 19800 15892
rect 19429 15855 19487 15861
rect 19794 15852 19800 15864
rect 19852 15852 19858 15904
rect 19904 15892 19932 15932
rect 20162 15920 20168 15932
rect 20220 15960 20226 15972
rect 20898 15960 20904 15972
rect 20220 15932 20904 15960
rect 20220 15920 20226 15932
rect 20898 15920 20904 15932
rect 20956 15920 20962 15972
rect 20070 15892 20076 15904
rect 19904 15864 20076 15892
rect 20070 15852 20076 15864
rect 20128 15892 20134 15904
rect 20257 15895 20315 15901
rect 20257 15892 20269 15895
rect 20128 15864 20269 15892
rect 20128 15852 20134 15864
rect 20257 15861 20269 15864
rect 20303 15861 20315 15895
rect 20990 15892 20996 15904
rect 20951 15864 20996 15892
rect 20257 15855 20315 15861
rect 20990 15852 20996 15864
rect 21048 15852 21054 15904
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 7929 15691 7987 15697
rect 7929 15657 7941 15691
rect 7975 15688 7987 15691
rect 9030 15688 9036 15700
rect 7975 15660 9036 15688
rect 7975 15657 7987 15660
rect 7929 15651 7987 15657
rect 9030 15648 9036 15660
rect 9088 15648 9094 15700
rect 9674 15648 9680 15700
rect 9732 15688 9738 15700
rect 10505 15691 10563 15697
rect 10505 15688 10517 15691
rect 9732 15660 10517 15688
rect 9732 15648 9738 15660
rect 10505 15657 10517 15660
rect 10551 15657 10563 15691
rect 10505 15651 10563 15657
rect 10873 15691 10931 15697
rect 10873 15657 10885 15691
rect 10919 15688 10931 15691
rect 11054 15688 11060 15700
rect 10919 15660 11060 15688
rect 10919 15657 10931 15660
rect 10873 15651 10931 15657
rect 11054 15648 11060 15660
rect 11112 15648 11118 15700
rect 12986 15688 12992 15700
rect 12947 15660 12992 15688
rect 12986 15648 12992 15660
rect 13044 15648 13050 15700
rect 13449 15691 13507 15697
rect 13449 15657 13461 15691
rect 13495 15688 13507 15691
rect 15194 15688 15200 15700
rect 13495 15660 15200 15688
rect 13495 15657 13507 15660
rect 13449 15651 13507 15657
rect 15194 15648 15200 15660
rect 15252 15648 15258 15700
rect 15654 15688 15660 15700
rect 15615 15660 15660 15688
rect 15654 15648 15660 15660
rect 15712 15648 15718 15700
rect 17770 15688 17776 15700
rect 17731 15660 17776 15688
rect 17770 15648 17776 15660
rect 17828 15648 17834 15700
rect 17880 15660 18911 15688
rect 6356 15623 6414 15629
rect 6356 15589 6368 15623
rect 6402 15620 6414 15623
rect 10962 15620 10968 15632
rect 6402 15592 10968 15620
rect 6402 15589 6414 15592
rect 6356 15583 6414 15589
rect 10962 15580 10968 15592
rect 11020 15580 11026 15632
rect 12253 15623 12311 15629
rect 12253 15589 12265 15623
rect 12299 15620 12311 15623
rect 12434 15620 12440 15632
rect 12299 15592 12440 15620
rect 12299 15589 12311 15592
rect 12253 15583 12311 15589
rect 12434 15580 12440 15592
rect 12492 15580 12498 15632
rect 13357 15623 13415 15629
rect 13357 15589 13369 15623
rect 13403 15620 13415 15623
rect 13722 15620 13728 15632
rect 13403 15592 13728 15620
rect 13403 15589 13415 15592
rect 13357 15583 13415 15589
rect 13722 15580 13728 15592
rect 13780 15580 13786 15632
rect 13998 15580 14004 15632
rect 14056 15620 14062 15632
rect 14056 15592 15516 15620
rect 14056 15580 14062 15592
rect 6089 15555 6147 15561
rect 6089 15521 6101 15555
rect 6135 15552 6147 15555
rect 7558 15552 7564 15564
rect 6135 15524 7564 15552
rect 6135 15521 6147 15524
rect 6089 15515 6147 15521
rect 7558 15512 7564 15524
rect 7616 15512 7622 15564
rect 8757 15555 8815 15561
rect 8757 15521 8769 15555
rect 8803 15552 8815 15555
rect 9674 15552 9680 15564
rect 8803 15524 9536 15552
rect 9635 15524 9680 15552
rect 8803 15521 8815 15524
rect 8757 15515 8815 15521
rect 8110 15444 8116 15496
rect 8168 15484 8174 15496
rect 8849 15487 8907 15493
rect 8849 15484 8861 15487
rect 8168 15456 8861 15484
rect 8168 15444 8174 15456
rect 8849 15453 8861 15456
rect 8895 15453 8907 15487
rect 9030 15484 9036 15496
rect 8991 15456 9036 15484
rect 8849 15447 8907 15453
rect 9030 15444 9036 15456
rect 9088 15444 9094 15496
rect 7466 15348 7472 15360
rect 7427 15320 7472 15348
rect 7466 15308 7472 15320
rect 7524 15308 7530 15360
rect 8389 15351 8447 15357
rect 8389 15317 8401 15351
rect 8435 15348 8447 15351
rect 8846 15348 8852 15360
rect 8435 15320 8852 15348
rect 8435 15317 8447 15320
rect 8389 15311 8447 15317
rect 8846 15308 8852 15320
rect 8904 15308 8910 15360
rect 9508 15348 9536 15524
rect 9674 15512 9680 15524
rect 9732 15512 9738 15564
rect 10980 15552 11008 15580
rect 14550 15552 14556 15564
rect 10980 15524 11100 15552
rect 14511 15524 14556 15552
rect 9953 15487 10011 15493
rect 9953 15453 9965 15487
rect 9999 15453 10011 15487
rect 10962 15484 10968 15496
rect 10923 15456 10968 15484
rect 9953 15447 10011 15453
rect 9968 15416 9996 15447
rect 10962 15444 10968 15456
rect 11020 15444 11026 15496
rect 11072 15493 11100 15524
rect 14550 15512 14556 15524
rect 14608 15512 14614 15564
rect 14645 15555 14703 15561
rect 14645 15521 14657 15555
rect 14691 15552 14703 15555
rect 15488 15552 15516 15592
rect 15562 15580 15568 15632
rect 15620 15620 15626 15632
rect 15749 15623 15807 15629
rect 15749 15620 15761 15623
rect 15620 15592 15761 15620
rect 15620 15580 15626 15592
rect 15749 15589 15761 15592
rect 15795 15589 15807 15623
rect 15749 15583 15807 15589
rect 16114 15580 16120 15632
rect 16172 15620 16178 15632
rect 17880 15620 17908 15660
rect 16172 15592 17908 15620
rect 16172 15580 16178 15592
rect 18690 15580 18696 15632
rect 18748 15629 18754 15632
rect 18748 15623 18812 15629
rect 18748 15589 18766 15623
rect 18800 15589 18812 15623
rect 18883 15620 18911 15660
rect 19242 15648 19248 15700
rect 19300 15688 19306 15700
rect 20441 15691 20499 15697
rect 20441 15688 20453 15691
rect 19300 15660 20453 15688
rect 19300 15648 19306 15660
rect 20441 15657 20453 15660
rect 20487 15657 20499 15691
rect 20441 15651 20499 15657
rect 20162 15620 20168 15632
rect 18883 15592 20168 15620
rect 18748 15583 18812 15589
rect 18748 15580 18754 15583
rect 20162 15580 20168 15592
rect 20220 15580 20226 15632
rect 16393 15555 16451 15561
rect 16393 15552 16405 15555
rect 14691 15524 15424 15552
rect 15488 15524 16405 15552
rect 14691 15521 14703 15524
rect 14645 15515 14703 15521
rect 11057 15487 11115 15493
rect 11057 15453 11069 15487
rect 11103 15453 11115 15487
rect 12342 15484 12348 15496
rect 12303 15456 12348 15484
rect 11057 15447 11115 15453
rect 12342 15444 12348 15456
rect 12400 15444 12406 15496
rect 12529 15487 12587 15493
rect 12529 15453 12541 15487
rect 12575 15484 12587 15487
rect 13078 15484 13084 15496
rect 12575 15456 13084 15484
rect 12575 15453 12587 15456
rect 12529 15447 12587 15453
rect 13078 15444 13084 15456
rect 13136 15444 13142 15496
rect 13538 15444 13544 15496
rect 13596 15484 13602 15496
rect 14829 15487 14887 15493
rect 13596 15456 13641 15484
rect 13596 15444 13602 15456
rect 14829 15453 14841 15487
rect 14875 15484 14887 15487
rect 15010 15484 15016 15496
rect 14875 15456 15016 15484
rect 14875 15453 14887 15456
rect 14829 15447 14887 15453
rect 15010 15444 15016 15456
rect 15068 15444 15074 15496
rect 15396 15484 15424 15524
rect 16393 15521 16405 15524
rect 16439 15552 16451 15555
rect 16482 15552 16488 15564
rect 16439 15524 16488 15552
rect 16439 15521 16451 15524
rect 16393 15515 16451 15521
rect 16482 15512 16488 15524
rect 16540 15512 16546 15564
rect 16660 15555 16718 15561
rect 16660 15521 16672 15555
rect 16706 15552 16718 15555
rect 17494 15552 17500 15564
rect 16706 15524 17500 15552
rect 16706 15521 16718 15524
rect 16660 15515 16718 15521
rect 17494 15512 17500 15524
rect 17552 15512 17558 15564
rect 18049 15555 18107 15561
rect 18049 15521 18061 15555
rect 18095 15552 18107 15555
rect 19886 15552 19892 15564
rect 18095 15524 19892 15552
rect 18095 15521 18107 15524
rect 18049 15515 18107 15521
rect 19886 15512 19892 15524
rect 19944 15512 19950 15564
rect 20257 15555 20315 15561
rect 20257 15521 20269 15555
rect 20303 15552 20315 15555
rect 20806 15552 20812 15564
rect 20303 15524 20812 15552
rect 20303 15521 20315 15524
rect 20257 15515 20315 15521
rect 20806 15512 20812 15524
rect 20864 15512 20870 15564
rect 15562 15484 15568 15496
rect 15396 15456 15568 15484
rect 15562 15444 15568 15456
rect 15620 15444 15626 15496
rect 15838 15444 15844 15496
rect 15896 15484 15902 15496
rect 15896 15456 15941 15484
rect 15896 15444 15902 15456
rect 18138 15444 18144 15496
rect 18196 15484 18202 15496
rect 18509 15487 18567 15493
rect 18509 15484 18521 15487
rect 18196 15456 18521 15484
rect 18196 15444 18202 15456
rect 18509 15453 18521 15456
rect 18555 15453 18567 15487
rect 18509 15447 18567 15453
rect 9968 15388 15792 15416
rect 11698 15348 11704 15360
rect 9508 15320 11704 15348
rect 11698 15308 11704 15320
rect 11756 15308 11762 15360
rect 11885 15351 11943 15357
rect 11885 15317 11897 15351
rect 11931 15348 11943 15351
rect 12802 15348 12808 15360
rect 11931 15320 12808 15348
rect 11931 15317 11943 15320
rect 11885 15311 11943 15317
rect 12802 15308 12808 15320
rect 12860 15308 12866 15360
rect 13906 15308 13912 15360
rect 13964 15348 13970 15360
rect 14185 15351 14243 15357
rect 14185 15348 14197 15351
rect 13964 15320 14197 15348
rect 13964 15308 13970 15320
rect 14185 15317 14197 15320
rect 14231 15317 14243 15351
rect 15286 15348 15292 15360
rect 15247 15320 15292 15348
rect 14185 15311 14243 15317
rect 15286 15308 15292 15320
rect 15344 15308 15350 15360
rect 15764 15348 15792 15388
rect 17328 15388 17908 15416
rect 17328 15348 17356 15388
rect 15764 15320 17356 15348
rect 17880 15348 17908 15388
rect 19150 15348 19156 15360
rect 17880 15320 19156 15348
rect 19150 15308 19156 15320
rect 19208 15308 19214 15360
rect 19426 15308 19432 15360
rect 19484 15348 19490 15360
rect 19889 15351 19947 15357
rect 19889 15348 19901 15351
rect 19484 15320 19901 15348
rect 19484 15308 19490 15320
rect 19889 15317 19901 15320
rect 19935 15348 19947 15351
rect 20346 15348 20352 15360
rect 19935 15320 20352 15348
rect 19935 15317 19947 15320
rect 19889 15311 19947 15317
rect 20346 15308 20352 15320
rect 20404 15308 20410 15360
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 5721 15147 5779 15153
rect 5721 15113 5733 15147
rect 5767 15144 5779 15147
rect 8110 15144 8116 15156
rect 5767 15116 8116 15144
rect 5767 15113 5779 15116
rect 5721 15107 5779 15113
rect 8110 15104 8116 15116
rect 8168 15104 8174 15156
rect 8202 15104 8208 15156
rect 8260 15144 8266 15156
rect 8260 15116 8616 15144
rect 8260 15104 8266 15116
rect 7466 15076 7472 15088
rect 6380 15048 7472 15076
rect 6178 15008 6184 15020
rect 6139 14980 6184 15008
rect 6178 14968 6184 14980
rect 6236 14968 6242 15020
rect 6380 15017 6408 15048
rect 7466 15036 7472 15048
rect 7524 15036 7530 15088
rect 8588 15076 8616 15116
rect 8662 15104 8668 15156
rect 8720 15144 8726 15156
rect 8849 15147 8907 15153
rect 8849 15144 8861 15147
rect 8720 15116 8861 15144
rect 8720 15104 8726 15116
rect 8849 15113 8861 15116
rect 8895 15113 8907 15147
rect 8849 15107 8907 15113
rect 10321 15147 10379 15153
rect 10321 15113 10333 15147
rect 10367 15144 10379 15147
rect 10962 15144 10968 15156
rect 10367 15116 10968 15144
rect 10367 15113 10379 15116
rect 10321 15107 10379 15113
rect 10962 15104 10968 15116
rect 11020 15104 11026 15156
rect 11333 15147 11391 15153
rect 11333 15113 11345 15147
rect 11379 15144 11391 15147
rect 12342 15144 12348 15156
rect 11379 15116 12348 15144
rect 11379 15113 11391 15116
rect 11333 15107 11391 15113
rect 12342 15104 12348 15116
rect 12400 15104 12406 15156
rect 12710 15104 12716 15156
rect 12768 15144 12774 15156
rect 13630 15144 13636 15156
rect 12768 15116 13636 15144
rect 12768 15104 12774 15116
rect 13630 15104 13636 15116
rect 13688 15144 13694 15156
rect 13817 15147 13875 15153
rect 13817 15144 13829 15147
rect 13688 15116 13829 15144
rect 13688 15104 13694 15116
rect 13817 15113 13829 15116
rect 13863 15113 13875 15147
rect 13817 15107 13875 15113
rect 15010 15104 15016 15156
rect 15068 15144 15074 15156
rect 15068 15116 15332 15144
rect 15068 15104 15074 15116
rect 15304 15076 15332 15116
rect 15470 15104 15476 15156
rect 15528 15144 15534 15156
rect 15930 15144 15936 15156
rect 15528 15116 15936 15144
rect 15528 15104 15534 15116
rect 15930 15104 15936 15116
rect 15988 15104 15994 15156
rect 18141 15147 18199 15153
rect 18141 15113 18153 15147
rect 18187 15144 18199 15147
rect 19518 15144 19524 15156
rect 18187 15116 19524 15144
rect 18187 15113 18199 15116
rect 18141 15107 18199 15113
rect 19518 15104 19524 15116
rect 19576 15104 19582 15156
rect 20993 15147 21051 15153
rect 20993 15113 21005 15147
rect 21039 15144 21051 15147
rect 21174 15144 21180 15156
rect 21039 15116 21180 15144
rect 21039 15113 21051 15116
rect 20993 15107 21051 15113
rect 21174 15104 21180 15116
rect 21232 15104 21238 15156
rect 15749 15079 15807 15085
rect 15749 15076 15761 15079
rect 8588 15048 11008 15076
rect 15304 15048 15761 15076
rect 6365 15011 6423 15017
rect 6365 14977 6377 15011
rect 6411 14977 6423 15011
rect 6365 14971 6423 14977
rect 9030 14968 9036 15020
rect 9088 15008 9094 15020
rect 9677 15011 9735 15017
rect 9677 15008 9689 15011
rect 9088 14980 9689 15008
rect 9088 14968 9094 14980
rect 9677 14977 9689 14980
rect 9723 14977 9735 15011
rect 9677 14971 9735 14977
rect 10594 14968 10600 15020
rect 10652 15008 10658 15020
rect 10873 15011 10931 15017
rect 10873 15008 10885 15011
rect 10652 14980 10885 15008
rect 10652 14968 10658 14980
rect 10873 14977 10885 14980
rect 10919 14977 10931 15011
rect 10873 14971 10931 14977
rect 5534 14900 5540 14952
rect 5592 14940 5598 14952
rect 6086 14940 6092 14952
rect 5592 14912 6092 14940
rect 5592 14900 5598 14912
rect 6086 14900 6092 14912
rect 6144 14900 6150 14952
rect 7469 14943 7527 14949
rect 7469 14909 7481 14943
rect 7515 14940 7527 14943
rect 7558 14940 7564 14952
rect 7515 14912 7564 14940
rect 7515 14909 7527 14912
rect 7469 14903 7527 14909
rect 7558 14900 7564 14912
rect 7616 14900 7622 14952
rect 7736 14943 7794 14949
rect 7736 14909 7748 14943
rect 7782 14940 7794 14943
rect 9048 14940 9076 14968
rect 7782 14912 9076 14940
rect 10689 14943 10747 14949
rect 7782 14909 7794 14912
rect 7736 14903 7794 14909
rect 10689 14909 10701 14943
rect 10735 14940 10747 14943
rect 10778 14940 10784 14952
rect 10735 14912 10784 14940
rect 10735 14909 10747 14912
rect 10689 14903 10747 14909
rect 10778 14900 10784 14912
rect 10836 14900 10842 14952
rect 10980 14940 11008 15048
rect 15749 15045 15761 15048
rect 15795 15045 15807 15079
rect 15749 15039 15807 15045
rect 16393 15079 16451 15085
rect 16393 15045 16405 15079
rect 16439 15076 16451 15079
rect 17954 15076 17960 15088
rect 16439 15048 17960 15076
rect 16439 15045 16451 15048
rect 16393 15039 16451 15045
rect 17954 15036 17960 15048
rect 18012 15036 18018 15088
rect 11793 15011 11851 15017
rect 11793 14977 11805 15011
rect 11839 15008 11851 15011
rect 11882 15008 11888 15020
rect 11839 14980 11888 15008
rect 11839 14977 11851 14980
rect 11793 14971 11851 14977
rect 11882 14968 11888 14980
rect 11940 14968 11946 15020
rect 11974 14968 11980 15020
rect 12032 15008 12038 15020
rect 14369 15011 14427 15017
rect 14369 15008 14381 15011
rect 12032 14980 12077 15008
rect 14200 14980 14381 15008
rect 12032 14968 12038 14980
rect 11701 14943 11759 14949
rect 11701 14940 11713 14943
rect 10980 14912 11713 14940
rect 11701 14909 11713 14912
rect 11747 14940 11759 14943
rect 12437 14943 12495 14949
rect 11747 14912 11928 14940
rect 11747 14909 11759 14912
rect 11701 14903 11759 14909
rect 11900 14884 11928 14912
rect 12437 14909 12449 14943
rect 12483 14940 12495 14943
rect 13998 14940 14004 14952
rect 12483 14912 14004 14940
rect 12483 14909 12495 14912
rect 12437 14903 12495 14909
rect 13998 14900 14004 14912
rect 14056 14940 14062 14952
rect 14200 14940 14228 14980
rect 14369 14977 14381 14980
rect 14415 14977 14427 15011
rect 17310 15008 17316 15020
rect 17271 14980 17316 15008
rect 14369 14971 14427 14977
rect 17310 14968 17316 14980
rect 17368 14968 17374 15020
rect 18598 14968 18604 15020
rect 18656 15008 18662 15020
rect 18693 15011 18751 15017
rect 18693 15008 18705 15011
rect 18656 14980 18705 15008
rect 18656 14968 18662 14980
rect 18693 14977 18705 14980
rect 18739 14977 18751 15011
rect 18693 14971 18751 14977
rect 18966 14968 18972 15020
rect 19024 15008 19030 15020
rect 19153 15011 19211 15017
rect 19153 15008 19165 15011
rect 19024 14980 19165 15008
rect 19024 14968 19030 14980
rect 19153 14977 19165 14980
rect 19199 14977 19211 15011
rect 19153 14971 19211 14977
rect 14056 14912 14228 14940
rect 14277 14943 14335 14949
rect 14056 14900 14062 14912
rect 14277 14909 14289 14943
rect 14323 14909 14335 14943
rect 14277 14903 14335 14909
rect 14636 14943 14694 14949
rect 14636 14909 14648 14943
rect 14682 14940 14694 14943
rect 15838 14940 15844 14952
rect 14682 14912 15844 14940
rect 14682 14909 14694 14912
rect 14636 14903 14694 14909
rect 8754 14832 8760 14884
rect 8812 14872 8818 14884
rect 9493 14875 9551 14881
rect 9493 14872 9505 14875
rect 8812 14844 9505 14872
rect 8812 14832 8818 14844
rect 9493 14841 9505 14844
rect 9539 14841 9551 14875
rect 9493 14835 9551 14841
rect 11882 14832 11888 14884
rect 11940 14832 11946 14884
rect 12704 14875 12762 14881
rect 12704 14841 12716 14875
rect 12750 14872 12762 14875
rect 13078 14872 13084 14884
rect 12750 14844 13084 14872
rect 12750 14841 12762 14844
rect 12704 14835 12762 14841
rect 13078 14832 13084 14844
rect 13136 14832 13142 14884
rect 14292 14872 14320 14903
rect 15838 14900 15844 14912
rect 15896 14900 15902 14952
rect 16206 14940 16212 14952
rect 16167 14912 16212 14940
rect 16206 14900 16212 14912
rect 16264 14900 16270 14952
rect 18509 14943 18567 14949
rect 18509 14909 18521 14943
rect 18555 14940 18567 14943
rect 18555 14912 19104 14940
rect 18555 14909 18567 14912
rect 18509 14903 18567 14909
rect 15654 14872 15660 14884
rect 13188 14844 14320 14872
rect 14936 14844 15660 14872
rect 9122 14804 9128 14816
rect 9083 14776 9128 14804
rect 9122 14764 9128 14776
rect 9180 14764 9186 14816
rect 9582 14804 9588 14816
rect 9543 14776 9588 14804
rect 9582 14764 9588 14776
rect 9640 14764 9646 14816
rect 10781 14807 10839 14813
rect 10781 14773 10793 14807
rect 10827 14804 10839 14807
rect 11146 14804 11152 14816
rect 10827 14776 11152 14804
rect 10827 14773 10839 14776
rect 10781 14767 10839 14773
rect 11146 14764 11152 14776
rect 11204 14764 11210 14816
rect 12618 14764 12624 14816
rect 12676 14804 12682 14816
rect 13188 14804 13216 14844
rect 12676 14776 13216 14804
rect 14093 14807 14151 14813
rect 12676 14764 12682 14776
rect 14093 14773 14105 14807
rect 14139 14804 14151 14807
rect 14936 14804 14964 14844
rect 15654 14832 15660 14844
rect 15712 14832 15718 14884
rect 17129 14875 17187 14881
rect 17129 14841 17141 14875
rect 17175 14872 17187 14875
rect 18874 14872 18880 14884
rect 17175 14844 18880 14872
rect 17175 14841 17187 14844
rect 17129 14835 17187 14841
rect 18874 14832 18880 14844
rect 18932 14832 18938 14884
rect 16758 14804 16764 14816
rect 14139 14776 14964 14804
rect 16719 14776 16764 14804
rect 14139 14773 14151 14776
rect 14093 14767 14151 14773
rect 16758 14764 16764 14776
rect 16816 14764 16822 14816
rect 17218 14804 17224 14816
rect 17179 14776 17224 14804
rect 17218 14764 17224 14776
rect 17276 14764 17282 14816
rect 18601 14807 18659 14813
rect 18601 14773 18613 14807
rect 18647 14804 18659 14807
rect 18690 14804 18696 14816
rect 18647 14776 18696 14804
rect 18647 14773 18659 14776
rect 18601 14767 18659 14773
rect 18690 14764 18696 14776
rect 18748 14764 18754 14816
rect 19076 14804 19104 14912
rect 20714 14900 20720 14952
rect 20772 14940 20778 14952
rect 20809 14943 20867 14949
rect 20809 14940 20821 14943
rect 20772 14912 20821 14940
rect 20772 14900 20778 14912
rect 20809 14909 20821 14912
rect 20855 14909 20867 14943
rect 20809 14903 20867 14909
rect 19426 14881 19432 14884
rect 19420 14872 19432 14881
rect 19387 14844 19432 14872
rect 19420 14835 19432 14844
rect 19426 14832 19432 14835
rect 19484 14832 19490 14884
rect 19886 14804 19892 14816
rect 19076 14776 19892 14804
rect 19886 14764 19892 14776
rect 19944 14764 19950 14816
rect 20162 14764 20168 14816
rect 20220 14804 20226 14816
rect 20533 14807 20591 14813
rect 20533 14804 20545 14807
rect 20220 14776 20545 14804
rect 20220 14764 20226 14776
rect 20533 14773 20545 14776
rect 20579 14773 20591 14807
rect 20533 14767 20591 14773
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 8757 14603 8815 14609
rect 8757 14569 8769 14603
rect 8803 14600 8815 14603
rect 9122 14600 9128 14612
rect 8803 14572 9128 14600
rect 8803 14569 8815 14572
rect 8757 14563 8815 14569
rect 9122 14560 9128 14572
rect 9180 14560 9186 14612
rect 9490 14560 9496 14612
rect 9548 14600 9554 14612
rect 11333 14603 11391 14609
rect 11333 14600 11345 14603
rect 9548 14572 11345 14600
rect 9548 14560 9554 14572
rect 11333 14569 11345 14572
rect 11379 14569 11391 14603
rect 12618 14600 12624 14612
rect 11333 14563 11391 14569
rect 11532 14572 12624 14600
rect 7000 14535 7058 14541
rect 7000 14501 7012 14535
rect 7046 14532 7058 14535
rect 7466 14532 7472 14544
rect 7046 14504 7472 14532
rect 7046 14501 7058 14504
rect 7000 14495 7058 14501
rect 7466 14492 7472 14504
rect 7524 14492 7530 14544
rect 8846 14532 8852 14544
rect 8807 14504 8852 14532
rect 8846 14492 8852 14504
rect 8904 14492 8910 14544
rect 11149 14535 11207 14541
rect 11149 14532 11161 14535
rect 9692 14504 11161 14532
rect 6733 14467 6791 14473
rect 6733 14433 6745 14467
rect 6779 14464 6791 14467
rect 9398 14464 9404 14476
rect 6779 14436 9404 14464
rect 6779 14433 6791 14436
rect 6733 14427 6791 14433
rect 9398 14424 9404 14436
rect 9456 14464 9462 14476
rect 9692 14473 9720 14504
rect 11149 14501 11161 14504
rect 11195 14501 11207 14535
rect 11149 14495 11207 14501
rect 11532 14473 11560 14572
rect 12618 14560 12624 14572
rect 12676 14560 12682 14612
rect 12802 14560 12808 14612
rect 12860 14600 12866 14612
rect 13817 14603 13875 14609
rect 13817 14600 13829 14603
rect 12860 14572 13829 14600
rect 12860 14560 12866 14572
rect 13817 14569 13829 14572
rect 13863 14569 13875 14603
rect 19242 14600 19248 14612
rect 13817 14563 13875 14569
rect 14016 14572 17448 14600
rect 19203 14572 19248 14600
rect 14016 14532 14044 14572
rect 11615 14504 14044 14532
rect 9677 14467 9735 14473
rect 9677 14464 9689 14467
rect 9456 14436 9689 14464
rect 9456 14424 9462 14436
rect 9677 14433 9689 14436
rect 9723 14433 9735 14467
rect 9677 14427 9735 14433
rect 9944 14467 10002 14473
rect 9944 14433 9956 14467
rect 9990 14464 10002 14467
rect 11517 14467 11575 14473
rect 9990 14436 11468 14464
rect 9990 14433 10002 14436
rect 9944 14427 10002 14433
rect 8662 14356 8668 14408
rect 8720 14396 8726 14408
rect 8941 14399 8999 14405
rect 8941 14396 8953 14399
rect 8720 14368 8953 14396
rect 8720 14356 8726 14368
rect 8941 14365 8953 14368
rect 8987 14365 8999 14399
rect 11440 14396 11468 14436
rect 11517 14433 11529 14467
rect 11563 14433 11575 14467
rect 11517 14427 11575 14433
rect 11615 14396 11643 14504
rect 14090 14492 14096 14544
rect 14148 14532 14154 14544
rect 14645 14535 14703 14541
rect 14645 14532 14657 14535
rect 14148 14504 14657 14532
rect 14148 14492 14154 14504
rect 14645 14501 14657 14504
rect 14691 14501 14703 14535
rect 14645 14495 14703 14501
rect 15654 14492 15660 14544
rect 15712 14532 15718 14544
rect 16384 14535 16442 14541
rect 15712 14504 16344 14532
rect 15712 14492 15718 14504
rect 11974 14473 11980 14476
rect 11968 14464 11980 14473
rect 11935 14436 11980 14464
rect 11968 14427 11980 14436
rect 11974 14424 11980 14427
rect 12032 14424 12038 14476
rect 13446 14424 13452 14476
rect 13504 14464 13510 14476
rect 13725 14467 13783 14473
rect 13725 14464 13737 14467
rect 13504 14436 13737 14464
rect 13504 14424 13510 14436
rect 13725 14433 13737 14436
rect 13771 14433 13783 14467
rect 14366 14464 14372 14476
rect 14327 14436 14372 14464
rect 13725 14427 13783 14433
rect 14366 14424 14372 14436
rect 14424 14424 14430 14476
rect 15286 14464 15292 14476
rect 15247 14436 15292 14464
rect 15286 14424 15292 14436
rect 15344 14424 15350 14476
rect 16117 14467 16175 14473
rect 16117 14433 16129 14467
rect 16163 14464 16175 14467
rect 16206 14464 16212 14476
rect 16163 14436 16212 14464
rect 16163 14433 16175 14436
rect 16117 14427 16175 14433
rect 16206 14424 16212 14436
rect 16264 14424 16270 14476
rect 16316 14464 16344 14504
rect 16384 14501 16396 14535
rect 16430 14532 16442 14535
rect 17310 14532 17316 14544
rect 16430 14504 17316 14532
rect 16430 14501 16442 14504
rect 16384 14495 16442 14501
rect 17310 14492 17316 14504
rect 17368 14492 17374 14544
rect 17420 14532 17448 14572
rect 19242 14560 19248 14572
rect 19300 14560 19306 14612
rect 19794 14560 19800 14612
rect 19852 14600 19858 14612
rect 20073 14603 20131 14609
rect 20073 14600 20085 14603
rect 19852 14572 20085 14600
rect 19852 14560 19858 14572
rect 20073 14569 20085 14572
rect 20119 14569 20131 14603
rect 20073 14563 20131 14569
rect 17420 14504 18644 14532
rect 16666 14464 16672 14476
rect 16316 14436 16672 14464
rect 16666 14424 16672 14436
rect 16724 14424 16730 14476
rect 17954 14424 17960 14476
rect 18012 14464 18018 14476
rect 18141 14467 18199 14473
rect 18141 14464 18153 14467
rect 18012 14436 18153 14464
rect 18012 14424 18018 14436
rect 18141 14433 18153 14436
rect 18187 14433 18199 14467
rect 18141 14427 18199 14433
rect 18233 14467 18291 14473
rect 18233 14433 18245 14467
rect 18279 14464 18291 14467
rect 18506 14464 18512 14476
rect 18279 14436 18512 14464
rect 18279 14433 18291 14436
rect 18233 14427 18291 14433
rect 18506 14424 18512 14436
rect 18564 14424 18570 14476
rect 11440 14368 11643 14396
rect 11701 14399 11759 14405
rect 8941 14359 8999 14365
rect 11701 14365 11713 14399
rect 11747 14365 11759 14399
rect 11701 14359 11759 14365
rect 8113 14331 8171 14337
rect 8113 14297 8125 14331
rect 8159 14328 8171 14331
rect 9030 14328 9036 14340
rect 8159 14300 9036 14328
rect 8159 14297 8171 14300
rect 8113 14291 8171 14297
rect 9030 14288 9036 14300
rect 9088 14288 9094 14340
rect 11149 14331 11207 14337
rect 11149 14297 11161 14331
rect 11195 14328 11207 14331
rect 11716 14328 11744 14359
rect 13630 14356 13636 14408
rect 13688 14396 13694 14408
rect 13909 14399 13967 14405
rect 13909 14396 13921 14399
rect 13688 14368 13921 14396
rect 13688 14356 13694 14368
rect 13909 14365 13921 14368
rect 13955 14365 13967 14399
rect 13909 14359 13967 14365
rect 14090 14356 14096 14408
rect 14148 14396 14154 14408
rect 14274 14396 14280 14408
rect 14148 14368 14280 14396
rect 14148 14356 14154 14368
rect 14274 14356 14280 14368
rect 14332 14356 14338 14408
rect 15565 14399 15623 14405
rect 15565 14365 15577 14399
rect 15611 14396 15623 14399
rect 16022 14396 16028 14408
rect 15611 14368 16028 14396
rect 15611 14365 15623 14368
rect 15565 14359 15623 14365
rect 16022 14356 16028 14368
rect 16080 14356 16086 14408
rect 17310 14356 17316 14408
rect 17368 14396 17374 14408
rect 18325 14399 18383 14405
rect 18325 14396 18337 14399
rect 17368 14368 18337 14396
rect 17368 14356 17374 14368
rect 18325 14365 18337 14368
rect 18371 14365 18383 14399
rect 18616 14396 18644 14504
rect 19061 14467 19119 14473
rect 19061 14433 19073 14467
rect 19107 14464 19119 14467
rect 19150 14464 19156 14476
rect 19107 14436 19156 14464
rect 19107 14433 19119 14436
rect 19061 14427 19119 14433
rect 19150 14424 19156 14436
rect 19208 14424 19214 14476
rect 19794 14424 19800 14476
rect 19852 14464 19858 14476
rect 19981 14467 20039 14473
rect 19981 14464 19993 14467
rect 19852 14436 19993 14464
rect 19852 14424 19858 14436
rect 19981 14433 19993 14436
rect 20027 14433 20039 14467
rect 19981 14427 20039 14433
rect 20162 14396 20168 14408
rect 18616 14368 20168 14396
rect 18325 14359 18383 14365
rect 20162 14356 20168 14368
rect 20220 14356 20226 14408
rect 20346 14356 20352 14408
rect 20404 14396 20410 14408
rect 20901 14399 20959 14405
rect 20901 14396 20913 14399
rect 20404 14368 20913 14396
rect 20404 14356 20410 14368
rect 20901 14365 20913 14368
rect 20947 14365 20959 14399
rect 20901 14359 20959 14365
rect 11195 14300 11744 14328
rect 11195 14297 11207 14300
rect 11149 14291 11207 14297
rect 17678 14288 17684 14340
rect 17736 14328 17742 14340
rect 19334 14328 19340 14340
rect 17736 14300 19340 14328
rect 17736 14288 17742 14300
rect 19334 14288 19340 14300
rect 19392 14288 19398 14340
rect 19613 14331 19671 14337
rect 19613 14297 19625 14331
rect 19659 14328 19671 14331
rect 20438 14328 20444 14340
rect 19659 14300 20444 14328
rect 19659 14297 19671 14300
rect 19613 14291 19671 14297
rect 20438 14288 20444 14300
rect 20496 14288 20502 14340
rect 8389 14263 8447 14269
rect 8389 14229 8401 14263
rect 8435 14260 8447 14263
rect 9674 14260 9680 14272
rect 8435 14232 9680 14260
rect 8435 14229 8447 14232
rect 8389 14223 8447 14229
rect 9674 14220 9680 14232
rect 9732 14220 9738 14272
rect 11054 14260 11060 14272
rect 11015 14232 11060 14260
rect 11054 14220 11060 14232
rect 11112 14220 11118 14272
rect 13078 14260 13084 14272
rect 13039 14232 13084 14260
rect 13078 14220 13084 14232
rect 13136 14220 13142 14272
rect 13170 14220 13176 14272
rect 13228 14260 13234 14272
rect 13357 14263 13415 14269
rect 13357 14260 13369 14263
rect 13228 14232 13369 14260
rect 13228 14220 13234 14232
rect 13357 14229 13369 14232
rect 13403 14229 13415 14263
rect 13357 14223 13415 14229
rect 13998 14220 14004 14272
rect 14056 14260 14062 14272
rect 15378 14260 15384 14272
rect 14056 14232 15384 14260
rect 14056 14220 14062 14232
rect 15378 14220 15384 14232
rect 15436 14220 15442 14272
rect 17494 14260 17500 14272
rect 17455 14232 17500 14260
rect 17494 14220 17500 14232
rect 17552 14220 17558 14272
rect 17770 14260 17776 14272
rect 17731 14232 17776 14260
rect 17770 14220 17776 14232
rect 17828 14220 17834 14272
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 6086 14016 6092 14068
rect 6144 14056 6150 14068
rect 6144 14028 12388 14056
rect 6144 14016 6150 14028
rect 12360 13988 12388 14028
rect 12434 14016 12440 14068
rect 12492 14056 12498 14068
rect 15286 14056 15292 14068
rect 12492 14028 12537 14056
rect 12636 14028 15292 14056
rect 12492 14016 12498 14028
rect 12636 13988 12664 14028
rect 15286 14016 15292 14028
rect 15344 14016 15350 14068
rect 15933 14059 15991 14065
rect 15933 14025 15945 14059
rect 15979 14056 15991 14059
rect 15979 14028 17264 14056
rect 15979 14025 15991 14028
rect 15933 14019 15991 14025
rect 12360 13960 12664 13988
rect 13078 13948 13084 14000
rect 13136 13988 13142 14000
rect 14277 13991 14335 13997
rect 13136 13960 14044 13988
rect 13136 13948 13142 13960
rect 8754 13920 8760 13932
rect 8715 13892 8760 13920
rect 8754 13880 8760 13892
rect 8812 13880 8818 13932
rect 9398 13880 9404 13932
rect 9456 13920 9462 13932
rect 9493 13923 9551 13929
rect 9493 13920 9505 13923
rect 9456 13892 9505 13920
rect 9456 13880 9462 13892
rect 9493 13889 9505 13892
rect 9539 13889 9551 13923
rect 9493 13883 9551 13889
rect 10686 13880 10692 13932
rect 10744 13920 10750 13932
rect 11514 13920 11520 13932
rect 10744 13892 11520 13920
rect 10744 13880 10750 13892
rect 11514 13880 11520 13892
rect 11572 13920 11578 13932
rect 11609 13923 11667 13929
rect 11609 13920 11621 13923
rect 11572 13892 11621 13920
rect 11572 13880 11578 13892
rect 11609 13889 11621 13892
rect 11655 13889 11667 13923
rect 11609 13883 11667 13889
rect 11701 13923 11759 13929
rect 11701 13889 11713 13923
rect 11747 13889 11759 13923
rect 11701 13883 11759 13889
rect 9760 13855 9818 13861
rect 9760 13821 9772 13855
rect 9806 13852 9818 13855
rect 11054 13852 11060 13864
rect 9806 13824 11060 13852
rect 9806 13821 9818 13824
rect 9760 13815 9818 13821
rect 11054 13812 11060 13824
rect 11112 13852 11118 13864
rect 11716 13852 11744 13883
rect 11974 13880 11980 13932
rect 12032 13920 12038 13932
rect 12989 13923 13047 13929
rect 12989 13920 13001 13923
rect 12032 13892 13001 13920
rect 12032 13880 12038 13892
rect 12989 13889 13001 13892
rect 13035 13889 13047 13923
rect 13906 13920 13912 13932
rect 13867 13892 13912 13920
rect 12989 13883 13047 13889
rect 11112 13824 11744 13852
rect 11112 13812 11118 13824
rect 12526 13812 12532 13864
rect 12584 13852 12590 13864
rect 12805 13855 12863 13861
rect 12805 13852 12817 13855
rect 12584 13824 12817 13852
rect 12584 13812 12590 13824
rect 12805 13821 12817 13824
rect 12851 13852 12863 13855
rect 12894 13852 12900 13864
rect 12851 13824 12900 13852
rect 12851 13821 12863 13824
rect 12805 13815 12863 13821
rect 12894 13812 12900 13824
rect 12952 13812 12958 13864
rect 13004 13852 13032 13883
rect 13906 13880 13912 13892
rect 13964 13880 13970 13932
rect 14016 13929 14044 13960
rect 14277 13957 14289 13991
rect 14323 13988 14335 13991
rect 14461 13991 14519 13997
rect 14461 13988 14473 13991
rect 14323 13960 14473 13988
rect 14323 13957 14335 13960
rect 14277 13951 14335 13957
rect 14461 13957 14473 13960
rect 14507 13957 14519 13991
rect 15378 13988 15384 14000
rect 14461 13951 14519 13957
rect 14936 13960 15384 13988
rect 14936 13929 14964 13960
rect 15378 13948 15384 13960
rect 15436 13948 15442 14000
rect 15473 13991 15531 13997
rect 15473 13957 15485 13991
rect 15519 13988 15531 13991
rect 16206 13988 16212 14000
rect 15519 13960 16212 13988
rect 15519 13957 15531 13960
rect 15473 13951 15531 13957
rect 16206 13948 16212 13960
rect 16264 13948 16270 14000
rect 17236 13988 17264 14028
rect 17310 14016 17316 14068
rect 17368 14056 17374 14068
rect 17681 14059 17739 14065
rect 17681 14056 17693 14059
rect 17368 14028 17693 14056
rect 17368 14016 17374 14028
rect 17681 14025 17693 14028
rect 17727 14025 17739 14059
rect 17681 14019 17739 14025
rect 17954 14016 17960 14068
rect 18012 14056 18018 14068
rect 18049 14059 18107 14065
rect 18049 14056 18061 14059
rect 18012 14028 18061 14056
rect 18012 14016 18018 14028
rect 18049 14025 18061 14028
rect 18095 14025 18107 14059
rect 18049 14019 18107 14025
rect 18598 14016 18604 14068
rect 18656 14016 18662 14068
rect 19794 14056 19800 14068
rect 19755 14028 19800 14056
rect 19794 14016 19800 14028
rect 19852 14016 19858 14068
rect 20622 14016 20628 14068
rect 20680 14056 20686 14068
rect 20993 14059 21051 14065
rect 20993 14056 21005 14059
rect 20680 14028 21005 14056
rect 20680 14016 20686 14028
rect 20993 14025 21005 14028
rect 21039 14025 21051 14059
rect 20993 14019 21051 14025
rect 17586 13988 17592 14000
rect 17236 13960 17592 13988
rect 17586 13948 17592 13960
rect 17644 13948 17650 14000
rect 18616 13988 18644 14016
rect 18064 13960 18644 13988
rect 18064 13932 18092 13960
rect 14001 13923 14059 13929
rect 14001 13889 14013 13923
rect 14047 13889 14059 13923
rect 14001 13883 14059 13889
rect 14921 13923 14979 13929
rect 14921 13889 14933 13923
rect 14967 13889 14979 13923
rect 14921 13883 14979 13889
rect 15010 13880 15016 13932
rect 15068 13920 15074 13932
rect 15068 13892 15113 13920
rect 15764 13892 16436 13920
rect 15068 13880 15074 13892
rect 15028 13852 15056 13880
rect 15654 13852 15660 13864
rect 13004 13824 15056 13852
rect 15615 13824 15660 13852
rect 15654 13812 15660 13824
rect 15712 13812 15718 13864
rect 15764 13861 15792 13892
rect 15749 13855 15807 13861
rect 15749 13821 15761 13855
rect 15795 13821 15807 13855
rect 15749 13815 15807 13821
rect 16206 13812 16212 13864
rect 16264 13852 16270 13864
rect 16301 13855 16359 13861
rect 16301 13852 16313 13855
rect 16264 13824 16313 13852
rect 16264 13812 16270 13824
rect 16301 13821 16313 13824
rect 16347 13821 16359 13855
rect 16408 13852 16436 13892
rect 17310 13880 17316 13932
rect 17368 13920 17374 13932
rect 17865 13923 17923 13929
rect 17865 13920 17877 13923
rect 17368 13892 17877 13920
rect 17368 13880 17374 13892
rect 17865 13889 17877 13892
rect 17911 13889 17923 13923
rect 17865 13883 17923 13889
rect 18046 13880 18052 13932
rect 18104 13880 18110 13932
rect 18414 13880 18420 13932
rect 18472 13920 18478 13932
rect 18601 13923 18659 13929
rect 18601 13920 18613 13923
rect 18472 13892 18613 13920
rect 18472 13880 18478 13892
rect 18601 13889 18613 13892
rect 18647 13889 18659 13923
rect 19245 13923 19303 13929
rect 19245 13920 19257 13923
rect 18601 13883 18659 13889
rect 18708 13892 19257 13920
rect 18708 13852 18736 13892
rect 19245 13889 19257 13892
rect 19291 13889 19303 13923
rect 19245 13883 19303 13889
rect 19426 13880 19432 13932
rect 19484 13920 19490 13932
rect 20349 13923 20407 13929
rect 20349 13920 20361 13923
rect 19484 13892 20361 13920
rect 19484 13880 19490 13892
rect 20349 13889 20361 13892
rect 20395 13889 20407 13923
rect 20349 13883 20407 13889
rect 19058 13852 19064 13864
rect 16408 13824 18736 13852
rect 19019 13824 19064 13852
rect 16301 13815 16359 13821
rect 19058 13812 19064 13824
rect 19116 13812 19122 13864
rect 19334 13812 19340 13864
rect 19392 13852 19398 13864
rect 19794 13852 19800 13864
rect 19392 13824 19800 13852
rect 19392 13812 19398 13824
rect 19794 13812 19800 13824
rect 19852 13812 19858 13864
rect 20806 13852 20812 13864
rect 20767 13824 20812 13852
rect 20806 13812 20812 13824
rect 20864 13812 20870 13864
rect 1394 13744 1400 13796
rect 1452 13784 1458 13796
rect 13817 13787 13875 13793
rect 1452 13756 8892 13784
rect 1452 13744 1458 13756
rect 8864 13716 8892 13756
rect 9876 13756 13768 13784
rect 9876 13716 9904 13756
rect 10870 13716 10876 13728
rect 8864 13688 9904 13716
rect 10831 13688 10876 13716
rect 10870 13676 10876 13688
rect 10928 13676 10934 13728
rect 11146 13716 11152 13728
rect 11107 13688 11152 13716
rect 11146 13676 11152 13688
rect 11204 13676 11210 13728
rect 11517 13719 11575 13725
rect 11517 13685 11529 13719
rect 11563 13716 11575 13719
rect 11698 13716 11704 13728
rect 11563 13688 11704 13716
rect 11563 13685 11575 13688
rect 11517 13679 11575 13685
rect 11698 13676 11704 13688
rect 11756 13716 11762 13728
rect 12897 13719 12955 13725
rect 12897 13716 12909 13719
rect 11756 13688 12909 13716
rect 11756 13676 11762 13688
rect 12897 13685 12909 13688
rect 12943 13716 12955 13719
rect 13078 13716 13084 13728
rect 12943 13688 13084 13716
rect 12943 13685 12955 13688
rect 12897 13679 12955 13685
rect 13078 13676 13084 13688
rect 13136 13676 13142 13728
rect 13446 13716 13452 13728
rect 13407 13688 13452 13716
rect 13446 13676 13452 13688
rect 13504 13676 13510 13728
rect 13740 13716 13768 13756
rect 13817 13753 13829 13787
rect 13863 13784 13875 13787
rect 14277 13787 14335 13793
rect 14277 13784 14289 13787
rect 13863 13756 14289 13784
rect 13863 13753 13875 13756
rect 13817 13747 13875 13753
rect 14277 13753 14289 13756
rect 14323 13753 14335 13787
rect 16568 13787 16626 13793
rect 14277 13747 14335 13753
rect 14476 13756 14964 13784
rect 14476 13716 14504 13756
rect 13740 13688 14504 13716
rect 14550 13676 14556 13728
rect 14608 13716 14614 13728
rect 14829 13719 14887 13725
rect 14829 13716 14841 13719
rect 14608 13688 14841 13716
rect 14608 13676 14614 13688
rect 14829 13685 14841 13688
rect 14875 13685 14887 13719
rect 14936 13716 14964 13756
rect 16568 13753 16580 13787
rect 16614 13784 16626 13787
rect 18322 13784 18328 13796
rect 16614 13756 18328 13784
rect 16614 13753 16626 13756
rect 16568 13747 16626 13753
rect 18322 13744 18328 13756
rect 18380 13744 18386 13796
rect 18417 13787 18475 13793
rect 18417 13753 18429 13787
rect 18463 13784 18475 13787
rect 18598 13784 18604 13796
rect 18463 13756 18604 13784
rect 18463 13753 18475 13756
rect 18417 13747 18475 13753
rect 18598 13744 18604 13756
rect 18656 13744 18662 13796
rect 20165 13787 20223 13793
rect 20165 13753 20177 13787
rect 20211 13784 20223 13787
rect 20346 13784 20352 13796
rect 20211 13756 20352 13784
rect 20211 13753 20223 13756
rect 20165 13747 20223 13753
rect 20346 13744 20352 13756
rect 20404 13744 20410 13796
rect 17678 13716 17684 13728
rect 14936 13688 17684 13716
rect 14829 13679 14887 13685
rect 17678 13676 17684 13688
rect 17736 13676 17742 13728
rect 17865 13719 17923 13725
rect 17865 13685 17877 13719
rect 17911 13716 17923 13719
rect 18509 13719 18567 13725
rect 18509 13716 18521 13719
rect 17911 13688 18521 13716
rect 17911 13685 17923 13688
rect 17865 13679 17923 13685
rect 18509 13685 18521 13688
rect 18555 13685 18567 13719
rect 18509 13679 18567 13685
rect 19242 13676 19248 13728
rect 19300 13716 19306 13728
rect 20257 13719 20315 13725
rect 20257 13716 20269 13719
rect 19300 13688 20269 13716
rect 19300 13676 19306 13688
rect 20257 13685 20269 13688
rect 20303 13685 20315 13719
rect 20257 13679 20315 13685
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 9309 13515 9367 13521
rect 9309 13481 9321 13515
rect 9355 13512 9367 13515
rect 9398 13512 9404 13524
rect 9355 13484 9404 13512
rect 9355 13481 9367 13484
rect 9309 13475 9367 13481
rect 9398 13472 9404 13484
rect 9456 13472 9462 13524
rect 9861 13515 9919 13521
rect 9861 13481 9873 13515
rect 9907 13481 9919 13515
rect 9861 13475 9919 13481
rect 10321 13515 10379 13521
rect 10321 13481 10333 13515
rect 10367 13512 10379 13515
rect 10873 13515 10931 13521
rect 10873 13512 10885 13515
rect 10367 13484 10885 13512
rect 10367 13481 10379 13484
rect 10321 13475 10379 13481
rect 10873 13481 10885 13484
rect 10919 13481 10931 13515
rect 10873 13475 10931 13481
rect 9876 13444 9904 13475
rect 11146 13472 11152 13524
rect 11204 13512 11210 13524
rect 11333 13515 11391 13521
rect 11333 13512 11345 13515
rect 11204 13484 11345 13512
rect 11204 13472 11210 13484
rect 11333 13481 11345 13484
rect 11379 13481 11391 13515
rect 11333 13475 11391 13481
rect 12618 13472 12624 13524
rect 12676 13512 12682 13524
rect 12805 13515 12863 13521
rect 12805 13512 12817 13515
rect 12676 13484 12817 13512
rect 12676 13472 12682 13484
rect 12805 13481 12817 13484
rect 12851 13481 12863 13515
rect 12805 13475 12863 13481
rect 14185 13515 14243 13521
rect 14185 13481 14197 13515
rect 14231 13512 14243 13515
rect 14366 13512 14372 13524
rect 14231 13484 14372 13512
rect 14231 13481 14243 13484
rect 14185 13475 14243 13481
rect 14366 13472 14372 13484
rect 14424 13472 14430 13524
rect 15105 13515 15163 13521
rect 15105 13481 15117 13515
rect 15151 13512 15163 13515
rect 16390 13512 16396 13524
rect 15151 13484 16396 13512
rect 15151 13481 15163 13484
rect 15105 13475 15163 13481
rect 16390 13472 16396 13484
rect 16448 13472 16454 13524
rect 16485 13515 16543 13521
rect 16485 13481 16497 13515
rect 16531 13481 16543 13515
rect 16485 13475 16543 13481
rect 10502 13444 10508 13456
rect 9876 13416 10508 13444
rect 10502 13404 10508 13416
rect 10560 13404 10566 13456
rect 12345 13447 12403 13453
rect 12345 13413 12357 13447
rect 12391 13444 12403 13447
rect 12710 13444 12716 13456
rect 12391 13416 12716 13444
rect 12391 13413 12403 13416
rect 12345 13407 12403 13413
rect 12710 13404 12716 13416
rect 12768 13404 12774 13456
rect 14645 13447 14703 13453
rect 13004 13416 14228 13444
rect 9490 13376 9496 13388
rect 9451 13348 9496 13376
rect 9490 13336 9496 13348
rect 9548 13336 9554 13388
rect 10226 13376 10232 13388
rect 10187 13348 10232 13376
rect 10226 13336 10232 13348
rect 10284 13336 10290 13388
rect 11241 13379 11299 13385
rect 11241 13345 11253 13379
rect 11287 13376 11299 13379
rect 11606 13376 11612 13388
rect 11287 13348 11612 13376
rect 11287 13345 11299 13348
rect 11241 13339 11299 13345
rect 11606 13336 11612 13348
rect 11664 13376 11670 13388
rect 12069 13379 12127 13385
rect 11664 13348 12020 13376
rect 11664 13336 11670 13348
rect 10413 13311 10471 13317
rect 10413 13277 10425 13311
rect 10459 13277 10471 13311
rect 10413 13271 10471 13277
rect 9490 13200 9496 13252
rect 9548 13240 9554 13252
rect 10428 13240 10456 13271
rect 10870 13268 10876 13320
rect 10928 13308 10934 13320
rect 11425 13311 11483 13317
rect 11425 13308 11437 13311
rect 10928 13280 11437 13308
rect 10928 13268 10934 13280
rect 11425 13277 11437 13280
rect 11471 13277 11483 13311
rect 11992 13308 12020 13348
rect 12069 13345 12081 13379
rect 12115 13376 12127 13379
rect 12434 13376 12440 13388
rect 12115 13348 12440 13376
rect 12115 13345 12127 13348
rect 12069 13339 12127 13345
rect 12434 13336 12440 13348
rect 12492 13336 12498 13388
rect 13004 13385 13032 13416
rect 14200 13388 14228 13416
rect 14645 13413 14657 13447
rect 14691 13444 14703 13447
rect 15562 13444 15568 13456
rect 14691 13416 15568 13444
rect 14691 13413 14703 13416
rect 14645 13407 14703 13413
rect 15562 13404 15568 13416
rect 15620 13404 15626 13456
rect 15746 13444 15752 13456
rect 15707 13416 15752 13444
rect 15746 13404 15752 13416
rect 15804 13404 15810 13456
rect 16500 13444 16528 13475
rect 16758 13472 16764 13524
rect 16816 13512 16822 13524
rect 17037 13515 17095 13521
rect 17037 13512 17049 13515
rect 16816 13484 17049 13512
rect 16816 13472 16822 13484
rect 17037 13481 17049 13484
rect 17083 13481 17095 13515
rect 17037 13475 17095 13481
rect 17129 13515 17187 13521
rect 17129 13481 17141 13515
rect 17175 13512 17187 13515
rect 17770 13512 17776 13524
rect 17175 13484 17776 13512
rect 17175 13481 17187 13484
rect 17129 13475 17187 13481
rect 17770 13472 17776 13484
rect 17828 13472 17834 13524
rect 17865 13515 17923 13521
rect 17865 13481 17877 13515
rect 17911 13512 17923 13515
rect 18506 13512 18512 13524
rect 17911 13484 18512 13512
rect 17911 13481 17923 13484
rect 17865 13475 17923 13481
rect 18506 13472 18512 13484
rect 18564 13472 18570 13524
rect 18598 13472 18604 13524
rect 18656 13512 18662 13524
rect 18693 13515 18751 13521
rect 18693 13512 18705 13515
rect 18656 13484 18705 13512
rect 18656 13472 18662 13484
rect 18693 13481 18705 13484
rect 18739 13481 18751 13515
rect 18874 13512 18880 13524
rect 18835 13484 18880 13512
rect 18693 13475 18751 13481
rect 18874 13472 18880 13484
rect 18932 13472 18938 13524
rect 19518 13472 19524 13524
rect 19576 13512 19582 13524
rect 19797 13515 19855 13521
rect 19797 13512 19809 13515
rect 19576 13484 19809 13512
rect 19576 13472 19582 13484
rect 19797 13481 19809 13484
rect 19843 13481 19855 13515
rect 19797 13475 19855 13481
rect 17954 13444 17960 13456
rect 16500 13416 17960 13444
rect 17954 13404 17960 13416
rect 18012 13404 18018 13456
rect 12989 13379 13047 13385
rect 12989 13345 13001 13379
rect 13035 13345 13047 13379
rect 13170 13376 13176 13388
rect 13131 13348 13176 13376
rect 12989 13339 13047 13345
rect 13170 13336 13176 13348
rect 13228 13336 13234 13388
rect 14182 13336 14188 13388
rect 14240 13336 14246 13388
rect 14553 13379 14611 13385
rect 14553 13345 14565 13379
rect 14599 13376 14611 13379
rect 14918 13376 14924 13388
rect 14599 13348 14924 13376
rect 14599 13345 14611 13348
rect 14553 13339 14611 13345
rect 14918 13336 14924 13348
rect 14976 13336 14982 13388
rect 15194 13336 15200 13388
rect 15252 13376 15258 13388
rect 15657 13379 15715 13385
rect 15657 13376 15669 13379
rect 15252 13348 15669 13376
rect 15252 13336 15258 13348
rect 15657 13345 15669 13348
rect 15703 13345 15715 13379
rect 15657 13339 15715 13345
rect 16022 13336 16028 13388
rect 16080 13376 16086 13388
rect 16301 13379 16359 13385
rect 16301 13376 16313 13379
rect 16080 13348 16313 13376
rect 16080 13336 16086 13348
rect 16301 13345 16313 13348
rect 16347 13345 16359 13379
rect 16301 13339 16359 13345
rect 17770 13336 17776 13388
rect 17828 13376 17834 13388
rect 18233 13379 18291 13385
rect 18233 13376 18245 13379
rect 17828 13348 18245 13376
rect 17828 13336 17834 13348
rect 18233 13345 18245 13348
rect 18279 13345 18291 13379
rect 18233 13339 18291 13345
rect 18598 13336 18604 13388
rect 18656 13376 18662 13388
rect 19705 13379 19763 13385
rect 19705 13376 19717 13379
rect 18656 13348 19717 13376
rect 18656 13336 18662 13348
rect 19705 13345 19717 13348
rect 19751 13345 19763 13379
rect 19705 13339 19763 13345
rect 12250 13308 12256 13320
rect 11992 13280 12256 13308
rect 11425 13271 11483 13277
rect 12250 13268 12256 13280
rect 12308 13268 12314 13320
rect 13449 13311 13507 13317
rect 13449 13277 13461 13311
rect 13495 13308 13507 13311
rect 14458 13308 14464 13320
rect 13495 13280 14464 13308
rect 13495 13277 13507 13280
rect 13449 13271 13507 13277
rect 14458 13268 14464 13280
rect 14516 13268 14522 13320
rect 14829 13311 14887 13317
rect 14829 13277 14841 13311
rect 14875 13308 14887 13311
rect 15105 13311 15163 13317
rect 15105 13308 15117 13311
rect 14875 13280 15117 13308
rect 14875 13277 14887 13280
rect 14829 13271 14887 13277
rect 15105 13277 15117 13280
rect 15151 13277 15163 13311
rect 15841 13311 15899 13317
rect 15841 13308 15853 13311
rect 15105 13271 15163 13277
rect 15212 13280 15853 13308
rect 9548 13212 10456 13240
rect 9548 13200 9554 13212
rect 12526 13132 12532 13184
rect 12584 13172 12590 13184
rect 13722 13172 13728 13184
rect 12584 13144 13728 13172
rect 12584 13132 12590 13144
rect 13722 13132 13728 13144
rect 13780 13132 13786 13184
rect 14366 13132 14372 13184
rect 14424 13172 14430 13184
rect 15212 13172 15240 13280
rect 15841 13277 15853 13280
rect 15887 13277 15899 13311
rect 15841 13271 15899 13277
rect 16758 13268 16764 13320
rect 16816 13308 16822 13320
rect 17218 13308 17224 13320
rect 16816 13280 17224 13308
rect 16816 13268 16822 13280
rect 17218 13268 17224 13280
rect 17276 13268 17282 13320
rect 17313 13311 17371 13317
rect 17313 13277 17325 13311
rect 17359 13308 17371 13311
rect 17494 13308 17500 13320
rect 17359 13280 17500 13308
rect 17359 13277 17371 13280
rect 17313 13271 17371 13277
rect 17494 13268 17500 13280
rect 17552 13268 17558 13320
rect 17678 13308 17684 13320
rect 17639 13280 17684 13308
rect 17678 13268 17684 13280
rect 17736 13308 17742 13320
rect 18325 13311 18383 13317
rect 18325 13308 18337 13311
rect 17736 13280 18337 13308
rect 17736 13268 17742 13280
rect 18325 13277 18337 13280
rect 18371 13277 18383 13311
rect 18506 13308 18512 13320
rect 18467 13280 18512 13308
rect 18325 13271 18383 13277
rect 18506 13268 18512 13280
rect 18564 13268 18570 13320
rect 19978 13308 19984 13320
rect 19939 13280 19984 13308
rect 19978 13268 19984 13280
rect 20036 13268 20042 13320
rect 16669 13243 16727 13249
rect 16669 13209 16681 13243
rect 16715 13240 16727 13243
rect 19058 13240 19064 13252
rect 16715 13212 19064 13240
rect 16715 13209 16727 13212
rect 16669 13203 16727 13209
rect 19058 13200 19064 13212
rect 19116 13200 19122 13252
rect 14424 13144 15240 13172
rect 15289 13175 15347 13181
rect 14424 13132 14430 13144
rect 15289 13141 15301 13175
rect 15335 13172 15347 13175
rect 15838 13172 15844 13184
rect 15335 13144 15844 13172
rect 15335 13141 15347 13144
rect 15289 13135 15347 13141
rect 15838 13132 15844 13144
rect 15896 13132 15902 13184
rect 15930 13132 15936 13184
rect 15988 13172 15994 13184
rect 18693 13175 18751 13181
rect 18693 13172 18705 13175
rect 15988 13144 18705 13172
rect 15988 13132 15994 13144
rect 18693 13141 18705 13144
rect 18739 13141 18751 13175
rect 18693 13135 18751 13141
rect 19337 13175 19395 13181
rect 19337 13141 19349 13175
rect 19383 13172 19395 13175
rect 20438 13172 20444 13184
rect 19383 13144 20444 13172
rect 19383 13141 19395 13144
rect 19337 13135 19395 13141
rect 20438 13132 20444 13144
rect 20496 13132 20502 13184
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 9398 12968 9404 12980
rect 8772 12940 9404 12968
rect 8772 12844 8800 12940
rect 9398 12928 9404 12940
rect 9456 12928 9462 12980
rect 10226 12928 10232 12980
rect 10284 12968 10290 12980
rect 10413 12971 10471 12977
rect 10413 12968 10425 12971
rect 10284 12940 10425 12968
rect 10284 12928 10290 12940
rect 10413 12937 10425 12940
rect 10459 12937 10471 12971
rect 10413 12931 10471 12937
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 12492 12940 12537 12968
rect 13464 12940 16068 12968
rect 12492 12928 12498 12940
rect 12066 12860 12072 12912
rect 12124 12900 12130 12912
rect 13464 12900 13492 12940
rect 12124 12872 13492 12900
rect 16040 12900 16068 12940
rect 16114 12928 16120 12980
rect 16172 12968 16178 12980
rect 16390 12968 16396 12980
rect 16172 12940 16396 12968
rect 16172 12928 16178 12940
rect 16390 12928 16396 12940
rect 16448 12968 16454 12980
rect 16485 12971 16543 12977
rect 16485 12968 16497 12971
rect 16448 12940 16497 12968
rect 16448 12928 16454 12940
rect 16485 12937 16497 12940
rect 16531 12937 16543 12971
rect 16758 12968 16764 12980
rect 16719 12940 16764 12968
rect 16485 12931 16543 12937
rect 16758 12928 16764 12940
rect 16816 12928 16822 12980
rect 16868 12940 20668 12968
rect 16868 12900 16896 12940
rect 18782 12900 18788 12912
rect 16040 12872 16896 12900
rect 18340 12872 18788 12900
rect 12124 12860 12130 12872
rect 8754 12832 8760 12844
rect 8667 12804 8760 12832
rect 8754 12792 8760 12804
rect 8812 12792 8818 12844
rect 10965 12835 11023 12841
rect 10965 12801 10977 12835
rect 11011 12801 11023 12835
rect 12986 12832 12992 12844
rect 12947 12804 12992 12832
rect 10965 12795 11023 12801
rect 9024 12767 9082 12773
rect 9024 12733 9036 12767
rect 9070 12764 9082 12767
rect 10870 12764 10876 12776
rect 9070 12736 10876 12764
rect 9070 12733 9082 12736
rect 9024 12727 9082 12733
rect 10870 12724 10876 12736
rect 10928 12764 10934 12776
rect 10980 12764 11008 12795
rect 12986 12792 12992 12804
rect 13044 12792 13050 12844
rect 16758 12792 16764 12844
rect 16816 12832 16822 12844
rect 17126 12832 17132 12844
rect 16816 12804 17132 12832
rect 16816 12792 16822 12804
rect 17126 12792 17132 12804
rect 17184 12792 17190 12844
rect 18340 12841 18368 12872
rect 18782 12860 18788 12872
rect 18840 12860 18846 12912
rect 20640 12841 20668 12940
rect 17405 12835 17463 12841
rect 17405 12801 17417 12835
rect 17451 12832 17463 12835
rect 18325 12835 18383 12841
rect 17451 12804 17724 12832
rect 17451 12801 17463 12804
rect 17405 12795 17463 12801
rect 10928 12736 11008 12764
rect 10928 12724 10934 12736
rect 13078 12724 13084 12776
rect 13136 12764 13142 12776
rect 13449 12767 13507 12773
rect 13449 12764 13461 12767
rect 13136 12736 13461 12764
rect 13136 12724 13142 12736
rect 13449 12733 13461 12736
rect 13495 12764 13507 12767
rect 15105 12767 15163 12773
rect 15105 12764 15117 12767
rect 13495 12736 15117 12764
rect 13495 12733 13507 12736
rect 13449 12727 13507 12733
rect 15105 12733 15117 12736
rect 15151 12764 15163 12767
rect 15194 12764 15200 12776
rect 15151 12736 15200 12764
rect 15151 12733 15163 12736
rect 15105 12727 15163 12733
rect 15194 12724 15200 12736
rect 15252 12724 15258 12776
rect 16206 12764 16212 12776
rect 15764 12736 16212 12764
rect 10781 12699 10839 12705
rect 10781 12665 10793 12699
rect 10827 12696 10839 12699
rect 11425 12699 11483 12705
rect 11425 12696 11437 12699
rect 10827 12668 11437 12696
rect 10827 12665 10839 12668
rect 10781 12659 10839 12665
rect 11425 12665 11437 12668
rect 11471 12665 11483 12699
rect 11425 12659 11483 12665
rect 12434 12656 12440 12708
rect 12492 12696 12498 12708
rect 12805 12699 12863 12705
rect 12805 12696 12817 12699
rect 12492 12668 12817 12696
rect 12492 12656 12498 12668
rect 12805 12665 12817 12668
rect 12851 12665 12863 12699
rect 12805 12659 12863 12665
rect 13716 12699 13774 12705
rect 13716 12665 13728 12699
rect 13762 12696 13774 12699
rect 14366 12696 14372 12708
rect 13762 12668 14372 12696
rect 13762 12665 13774 12668
rect 13716 12659 13774 12665
rect 14366 12656 14372 12668
rect 14424 12656 14430 12708
rect 15350 12699 15408 12705
rect 15350 12696 15362 12699
rect 14844 12668 15362 12696
rect 9490 12588 9496 12640
rect 9548 12628 9554 12640
rect 10137 12631 10195 12637
rect 10137 12628 10149 12631
rect 9548 12600 10149 12628
rect 9548 12588 9554 12600
rect 10137 12597 10149 12600
rect 10183 12597 10195 12631
rect 10137 12591 10195 12597
rect 10873 12631 10931 12637
rect 10873 12597 10885 12631
rect 10919 12628 10931 12631
rect 11054 12628 11060 12640
rect 10919 12600 11060 12628
rect 10919 12597 10931 12600
rect 10873 12591 10931 12597
rect 11054 12588 11060 12600
rect 11112 12588 11118 12640
rect 12894 12628 12900 12640
rect 12855 12600 12900 12628
rect 12894 12588 12900 12600
rect 12952 12588 12958 12640
rect 14844 12637 14872 12668
rect 15350 12665 15362 12668
rect 15396 12696 15408 12699
rect 15764 12696 15792 12736
rect 16206 12724 16212 12736
rect 16264 12724 16270 12776
rect 16942 12724 16948 12776
rect 17000 12764 17006 12776
rect 17221 12767 17279 12773
rect 17221 12764 17233 12767
rect 17000 12736 17233 12764
rect 17000 12724 17006 12736
rect 17221 12733 17233 12736
rect 17267 12764 17279 12767
rect 17586 12764 17592 12776
rect 17267 12736 17592 12764
rect 17267 12733 17279 12736
rect 17221 12727 17279 12733
rect 17586 12724 17592 12736
rect 17644 12724 17650 12776
rect 17129 12699 17187 12705
rect 17129 12696 17141 12699
rect 15396 12668 15792 12696
rect 15856 12668 17141 12696
rect 15396 12665 15408 12668
rect 15350 12659 15408 12665
rect 14829 12631 14887 12637
rect 14829 12597 14841 12631
rect 14875 12597 14887 12631
rect 14829 12591 14887 12597
rect 15010 12588 15016 12640
rect 15068 12628 15074 12640
rect 15856 12628 15884 12668
rect 17129 12665 17141 12668
rect 17175 12665 17187 12699
rect 17129 12659 17187 12665
rect 15068 12600 15884 12628
rect 15068 12588 15074 12600
rect 16666 12588 16672 12640
rect 16724 12628 16730 12640
rect 17218 12628 17224 12640
rect 16724 12600 17224 12628
rect 16724 12588 16730 12600
rect 17218 12588 17224 12600
rect 17276 12588 17282 12640
rect 17696 12628 17724 12804
rect 18325 12801 18337 12835
rect 18371 12801 18383 12835
rect 18325 12795 18383 12801
rect 20625 12835 20683 12841
rect 20625 12801 20637 12835
rect 20671 12801 20683 12835
rect 20625 12795 20683 12801
rect 18049 12767 18107 12773
rect 18049 12733 18061 12767
rect 18095 12764 18107 12767
rect 18414 12764 18420 12776
rect 18095 12736 18420 12764
rect 18095 12733 18107 12736
rect 18049 12727 18107 12733
rect 18414 12724 18420 12736
rect 18472 12724 18478 12776
rect 18785 12767 18843 12773
rect 18785 12733 18797 12767
rect 18831 12764 18843 12767
rect 18874 12764 18880 12776
rect 18831 12736 18880 12764
rect 18831 12733 18843 12736
rect 18785 12727 18843 12733
rect 18874 12724 18880 12736
rect 18932 12724 18938 12776
rect 19052 12767 19110 12773
rect 19052 12733 19064 12767
rect 19098 12764 19110 12767
rect 19978 12764 19984 12776
rect 19098 12736 19984 12764
rect 19098 12733 19110 12736
rect 19052 12727 19110 12733
rect 19978 12724 19984 12736
rect 20036 12724 20042 12776
rect 20438 12764 20444 12776
rect 20399 12736 20444 12764
rect 20438 12724 20444 12736
rect 20496 12724 20502 12776
rect 18506 12628 18512 12640
rect 17696 12600 18512 12628
rect 18506 12588 18512 12600
rect 18564 12628 18570 12640
rect 20165 12631 20223 12637
rect 20165 12628 20177 12631
rect 18564 12600 20177 12628
rect 18564 12588 18570 12600
rect 20165 12597 20177 12600
rect 20211 12597 20223 12631
rect 20165 12591 20223 12597
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 12713 12427 12771 12433
rect 12713 12393 12725 12427
rect 12759 12393 12771 12427
rect 12713 12387 12771 12393
rect 8012 12359 8070 12365
rect 8012 12325 8024 12359
rect 8058 12356 8070 12359
rect 9490 12356 9496 12368
rect 8058 12328 9496 12356
rect 8058 12325 8070 12328
rect 8012 12319 8070 12325
rect 9490 12316 9496 12328
rect 9548 12316 9554 12368
rect 9582 12316 9588 12368
rect 9640 12356 9646 12368
rect 12728 12356 12756 12387
rect 12986 12384 12992 12436
rect 13044 12384 13050 12436
rect 14366 12424 14372 12436
rect 14327 12396 14372 12424
rect 14366 12384 14372 12396
rect 14424 12384 14430 12436
rect 14550 12384 14556 12436
rect 14608 12424 14614 12436
rect 14645 12427 14703 12433
rect 14645 12424 14657 12427
rect 14608 12396 14657 12424
rect 14608 12384 14614 12396
rect 14645 12393 14657 12396
rect 14691 12393 14703 12427
rect 17402 12424 17408 12436
rect 14645 12387 14703 12393
rect 15948 12396 17408 12424
rect 13004 12356 13032 12384
rect 13234 12359 13292 12365
rect 13234 12356 13246 12359
rect 9640 12328 12664 12356
rect 12728 12328 13246 12356
rect 9640 12316 9646 12328
rect 7745 12291 7803 12297
rect 7745 12257 7757 12291
rect 7791 12288 7803 12291
rect 9674 12288 9680 12300
rect 7791 12260 8800 12288
rect 9635 12260 9680 12288
rect 7791 12257 7803 12260
rect 7745 12251 7803 12257
rect 8772 12232 8800 12260
rect 9674 12248 9680 12260
rect 9732 12248 9738 12300
rect 11600 12291 11658 12297
rect 9784 12260 11008 12288
rect 8754 12180 8760 12232
rect 8812 12220 8818 12232
rect 9784 12220 9812 12260
rect 10980 12232 11008 12260
rect 11600 12257 11612 12291
rect 11646 12288 11658 12291
rect 12066 12288 12072 12300
rect 11646 12260 12072 12288
rect 11646 12257 11658 12260
rect 11600 12251 11658 12257
rect 12066 12248 12072 12260
rect 12124 12248 12130 12300
rect 8812 12192 9812 12220
rect 9953 12223 10011 12229
rect 8812 12180 8818 12192
rect 9953 12189 9965 12223
rect 9999 12189 10011 12223
rect 9953 12183 10011 12189
rect 9122 12084 9128 12096
rect 9083 12056 9128 12084
rect 9122 12044 9128 12056
rect 9180 12044 9186 12096
rect 9968 12084 9996 12183
rect 10962 12180 10968 12232
rect 11020 12220 11026 12232
rect 11333 12223 11391 12229
rect 11333 12220 11345 12223
rect 11020 12192 11345 12220
rect 11020 12180 11026 12192
rect 11333 12189 11345 12192
rect 11379 12189 11391 12223
rect 12636 12220 12664 12328
rect 13234 12325 13246 12328
rect 13280 12325 13292 12359
rect 13234 12319 13292 12325
rect 14734 12316 14740 12368
rect 14792 12356 14798 12368
rect 15948 12356 15976 12396
rect 17402 12384 17408 12396
rect 17460 12384 17466 12436
rect 17589 12427 17647 12433
rect 17589 12393 17601 12427
rect 17635 12424 17647 12427
rect 18506 12424 18512 12436
rect 17635 12396 18512 12424
rect 17635 12393 17647 12396
rect 17589 12387 17647 12393
rect 18506 12384 18512 12396
rect 18564 12384 18570 12436
rect 18874 12424 18880 12436
rect 18616 12396 18880 12424
rect 16114 12365 16120 12368
rect 16108 12356 16120 12365
rect 14792 12328 15976 12356
rect 16075 12328 16120 12356
rect 14792 12316 14798 12328
rect 16108 12319 16120 12328
rect 16114 12316 16120 12319
rect 16172 12316 16178 12368
rect 16574 12356 16580 12368
rect 16224 12328 16580 12356
rect 12986 12288 12992 12300
rect 12947 12260 12992 12288
rect 12986 12248 12992 12260
rect 13044 12248 13050 12300
rect 16224 12288 16252 12328
rect 16574 12316 16580 12328
rect 16632 12316 16638 12368
rect 18616 12297 18644 12396
rect 18874 12384 18880 12396
rect 18932 12384 18938 12436
rect 19978 12424 19984 12436
rect 19939 12396 19984 12424
rect 19978 12384 19984 12396
rect 20036 12384 20042 12436
rect 20346 12384 20352 12436
rect 20404 12424 20410 12436
rect 20441 12427 20499 12433
rect 20441 12424 20453 12427
rect 20404 12396 20453 12424
rect 20404 12384 20410 12396
rect 20441 12393 20453 12396
rect 20487 12393 20499 12427
rect 20441 12387 20499 12393
rect 20901 12359 20959 12365
rect 20901 12356 20913 12359
rect 18708 12328 20913 12356
rect 13096 12260 16252 12288
rect 17957 12291 18015 12297
rect 13096 12220 13124 12260
rect 17957 12257 17969 12291
rect 18003 12288 18015 12291
rect 18601 12291 18659 12297
rect 18003 12260 18552 12288
rect 18003 12257 18015 12260
rect 17957 12251 18015 12257
rect 15286 12220 15292 12232
rect 12636 12192 13124 12220
rect 15247 12192 15292 12220
rect 11333 12183 11391 12189
rect 15286 12180 15292 12192
rect 15344 12180 15350 12232
rect 15746 12180 15752 12232
rect 15804 12220 15810 12232
rect 15841 12223 15899 12229
rect 15841 12220 15853 12223
rect 15804 12192 15853 12220
rect 15804 12180 15810 12192
rect 15841 12189 15853 12192
rect 15887 12189 15899 12223
rect 18046 12220 18052 12232
rect 18007 12192 18052 12220
rect 15841 12183 15899 12189
rect 18046 12180 18052 12192
rect 18104 12180 18110 12232
rect 18233 12223 18291 12229
rect 18233 12189 18245 12223
rect 18279 12189 18291 12223
rect 18524 12220 18552 12260
rect 18601 12257 18613 12291
rect 18647 12257 18659 12291
rect 18601 12251 18659 12257
rect 18708 12220 18736 12328
rect 20901 12325 20913 12328
rect 20947 12325 20959 12359
rect 20901 12319 20959 12325
rect 18874 12297 18880 12300
rect 18868 12288 18880 12297
rect 18835 12260 18880 12288
rect 18868 12251 18880 12260
rect 18874 12248 18880 12251
rect 18932 12248 18938 12300
rect 19426 12248 19432 12300
rect 19484 12288 19490 12300
rect 20257 12291 20315 12297
rect 20257 12288 20269 12291
rect 19484 12260 20269 12288
rect 19484 12248 19490 12260
rect 20257 12257 20269 12260
rect 20303 12257 20315 12291
rect 20257 12251 20315 12257
rect 18524 12192 18736 12220
rect 18233 12183 18291 12189
rect 17954 12112 17960 12164
rect 18012 12152 18018 12164
rect 18248 12152 18276 12183
rect 18012 12124 18644 12152
rect 18012 12112 18018 12124
rect 15746 12084 15752 12096
rect 9968 12056 15752 12084
rect 15746 12044 15752 12056
rect 15804 12044 15810 12096
rect 17218 12084 17224 12096
rect 17179 12056 17224 12084
rect 17218 12044 17224 12056
rect 17276 12044 17282 12096
rect 18616 12084 18644 12124
rect 18874 12084 18880 12096
rect 18616 12056 18880 12084
rect 18874 12044 18880 12056
rect 18932 12044 18938 12096
rect 19702 12044 19708 12096
rect 19760 12084 19766 12096
rect 20346 12084 20352 12096
rect 19760 12056 20352 12084
rect 19760 12044 19766 12056
rect 20346 12044 20352 12056
rect 20404 12044 20410 12096
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 11517 11883 11575 11889
rect 11517 11849 11529 11883
rect 11563 11880 11575 11883
rect 12434 11880 12440 11892
rect 11563 11852 12440 11880
rect 11563 11849 11575 11852
rect 11517 11843 11575 11849
rect 12434 11840 12440 11852
rect 12492 11840 12498 11892
rect 12621 11883 12679 11889
rect 12621 11849 12633 11883
rect 12667 11880 12679 11883
rect 12894 11880 12900 11892
rect 12667 11852 12900 11880
rect 12667 11849 12679 11852
rect 12621 11843 12679 11849
rect 12894 11840 12900 11852
rect 12952 11840 12958 11892
rect 14369 11883 14427 11889
rect 14369 11849 14381 11883
rect 14415 11880 14427 11883
rect 14918 11880 14924 11892
rect 14415 11852 14924 11880
rect 14415 11849 14427 11852
rect 14369 11843 14427 11849
rect 14918 11840 14924 11852
rect 14976 11840 14982 11892
rect 15562 11880 15568 11892
rect 15523 11852 15568 11880
rect 15562 11840 15568 11852
rect 15620 11840 15626 11892
rect 15746 11840 15752 11892
rect 15804 11880 15810 11892
rect 15804 11852 18736 11880
rect 15804 11840 15810 11852
rect 13541 11815 13599 11821
rect 13541 11781 13553 11815
rect 13587 11812 13599 11815
rect 13587 11784 16068 11812
rect 13587 11781 13599 11784
rect 13541 11775 13599 11781
rect 12066 11744 12072 11756
rect 12027 11716 12072 11744
rect 12066 11704 12072 11716
rect 12124 11744 12130 11756
rect 13173 11747 13231 11753
rect 13173 11744 13185 11747
rect 12124 11716 13185 11744
rect 12124 11704 12130 11716
rect 13173 11713 13185 11716
rect 13219 11713 13231 11747
rect 13173 11707 13231 11713
rect 14185 11747 14243 11753
rect 14185 11713 14197 11747
rect 14231 11744 14243 11747
rect 14366 11744 14372 11756
rect 14231 11716 14372 11744
rect 14231 11713 14243 11716
rect 14185 11707 14243 11713
rect 14366 11704 14372 11716
rect 14424 11744 14430 11756
rect 14921 11747 14979 11753
rect 14921 11744 14933 11747
rect 14424 11716 14933 11744
rect 14424 11704 14430 11716
rect 14921 11713 14933 11716
rect 14967 11713 14979 11747
rect 14921 11707 14979 11713
rect 15654 11704 15660 11756
rect 15712 11744 15718 11756
rect 15930 11744 15936 11756
rect 15712 11716 15936 11744
rect 15712 11704 15718 11716
rect 15930 11704 15936 11716
rect 15988 11704 15994 11756
rect 16040 11753 16068 11784
rect 17218 11772 17224 11824
rect 17276 11812 17282 11824
rect 17276 11784 17816 11812
rect 17276 11772 17282 11784
rect 16025 11747 16083 11753
rect 16025 11713 16037 11747
rect 16071 11713 16083 11747
rect 16206 11744 16212 11756
rect 16167 11716 16212 11744
rect 16025 11707 16083 11713
rect 16206 11704 16212 11716
rect 16264 11704 16270 11756
rect 17589 11747 17647 11753
rect 17589 11713 17601 11747
rect 17635 11744 17647 11747
rect 17678 11744 17684 11756
rect 17635 11716 17684 11744
rect 17635 11713 17647 11716
rect 17589 11707 17647 11713
rect 17678 11704 17684 11716
rect 17736 11704 17742 11756
rect 17788 11744 17816 11784
rect 18601 11747 18659 11753
rect 18601 11744 18613 11747
rect 17788 11716 18613 11744
rect 18601 11713 18613 11716
rect 18647 11713 18659 11747
rect 18708 11744 18736 11852
rect 19150 11840 19156 11892
rect 19208 11880 19214 11892
rect 19337 11883 19395 11889
rect 19337 11880 19349 11883
rect 19208 11852 19349 11880
rect 19208 11840 19214 11852
rect 19337 11849 19349 11852
rect 19383 11849 19395 11883
rect 21085 11883 21143 11889
rect 21085 11880 21097 11883
rect 19337 11843 19395 11849
rect 19444 11852 21097 11880
rect 18874 11772 18880 11824
rect 18932 11812 18938 11824
rect 19444 11812 19472 11852
rect 21085 11849 21097 11852
rect 21131 11849 21143 11883
rect 21085 11843 21143 11849
rect 18932 11784 19472 11812
rect 18932 11772 18938 11784
rect 18708 11716 19840 11744
rect 18601 11707 18659 11713
rect 8205 11679 8263 11685
rect 8205 11645 8217 11679
rect 8251 11676 8263 11679
rect 8754 11676 8760 11688
rect 8251 11648 8760 11676
rect 8251 11645 8263 11648
rect 8205 11639 8263 11645
rect 8754 11636 8760 11648
rect 8812 11636 8818 11688
rect 8938 11636 8944 11688
rect 8996 11676 9002 11688
rect 9582 11676 9588 11688
rect 8996 11648 9588 11676
rect 8996 11636 9002 11648
rect 9582 11636 9588 11648
rect 9640 11636 9646 11688
rect 9950 11636 9956 11688
rect 10008 11676 10014 11688
rect 10870 11676 10876 11688
rect 10008 11648 10876 11676
rect 10008 11636 10014 11648
rect 10870 11636 10876 11648
rect 10928 11676 10934 11688
rect 14001 11679 14059 11685
rect 14001 11676 14013 11679
rect 10928 11648 14013 11676
rect 10928 11636 10934 11648
rect 14001 11645 14013 11648
rect 14047 11645 14059 11679
rect 14001 11639 14059 11645
rect 14458 11636 14464 11688
rect 14516 11676 14522 11688
rect 19153 11679 19211 11685
rect 19153 11676 19165 11679
rect 14516 11648 19165 11676
rect 14516 11636 14522 11648
rect 19153 11645 19165 11648
rect 19199 11645 19211 11679
rect 19153 11639 19211 11645
rect 19610 11636 19616 11688
rect 19668 11676 19674 11688
rect 19705 11679 19763 11685
rect 19705 11676 19717 11679
rect 19668 11648 19717 11676
rect 19668 11636 19674 11648
rect 19705 11645 19717 11648
rect 19751 11645 19763 11679
rect 19812 11676 19840 11716
rect 20806 11676 20812 11688
rect 19812 11648 20812 11676
rect 19705 11639 19763 11645
rect 20806 11636 20812 11648
rect 20864 11636 20870 11688
rect 8472 11611 8530 11617
rect 8472 11577 8484 11611
rect 8518 11608 8530 11611
rect 9122 11608 9128 11620
rect 8518 11580 9128 11608
rect 8518 11577 8530 11580
rect 8472 11571 8530 11577
rect 9122 11568 9128 11580
rect 9180 11568 9186 11620
rect 11241 11611 11299 11617
rect 11241 11577 11253 11611
rect 11287 11608 11299 11611
rect 11885 11611 11943 11617
rect 11885 11608 11897 11611
rect 11287 11580 11897 11608
rect 11287 11577 11299 11580
rect 11241 11571 11299 11577
rect 11885 11577 11897 11580
rect 11931 11577 11943 11611
rect 11885 11571 11943 11577
rect 12710 11568 12716 11620
rect 12768 11608 12774 11620
rect 13081 11611 13139 11617
rect 13081 11608 13093 11611
rect 12768 11580 13093 11608
rect 12768 11568 12774 11580
rect 13081 11577 13093 11580
rect 13127 11577 13139 11611
rect 13081 11571 13139 11577
rect 14918 11568 14924 11620
rect 14976 11608 14982 11620
rect 15933 11611 15991 11617
rect 15933 11608 15945 11611
rect 14976 11580 15945 11608
rect 14976 11568 14982 11580
rect 15933 11577 15945 11580
rect 15979 11577 15991 11611
rect 15933 11571 15991 11577
rect 16574 11568 16580 11620
rect 16632 11608 16638 11620
rect 17494 11608 17500 11620
rect 16632 11580 17500 11608
rect 16632 11568 16638 11580
rect 17494 11568 17500 11580
rect 17552 11568 17558 11620
rect 18417 11611 18475 11617
rect 18417 11577 18429 11611
rect 18463 11608 18475 11611
rect 18966 11608 18972 11620
rect 18463 11580 18972 11608
rect 18463 11577 18475 11580
rect 18417 11571 18475 11577
rect 18966 11568 18972 11580
rect 19024 11568 19030 11620
rect 19978 11617 19984 11620
rect 19972 11608 19984 11617
rect 19939 11580 19984 11608
rect 19972 11571 19984 11580
rect 19978 11568 19984 11571
rect 20036 11568 20042 11620
rect 9490 11500 9496 11552
rect 9548 11540 9554 11552
rect 9585 11543 9643 11549
rect 9585 11540 9597 11543
rect 9548 11512 9597 11540
rect 9548 11500 9554 11512
rect 9585 11509 9597 11512
rect 9631 11509 9643 11543
rect 9585 11503 9643 11509
rect 9861 11543 9919 11549
rect 9861 11509 9873 11543
rect 9907 11540 9919 11543
rect 10042 11540 10048 11552
rect 9907 11512 10048 11540
rect 9907 11509 9919 11512
rect 9861 11503 9919 11509
rect 10042 11500 10048 11512
rect 10100 11500 10106 11552
rect 11977 11543 12035 11549
rect 11977 11509 11989 11543
rect 12023 11540 12035 11543
rect 12434 11540 12440 11552
rect 12023 11512 12440 11540
rect 12023 11509 12035 11512
rect 11977 11503 12035 11509
rect 12434 11500 12440 11512
rect 12492 11500 12498 11552
rect 12986 11540 12992 11552
rect 12947 11512 12992 11540
rect 12986 11500 12992 11512
rect 13044 11500 13050 11552
rect 13909 11543 13967 11549
rect 13909 11509 13921 11543
rect 13955 11540 13967 11543
rect 14458 11540 14464 11552
rect 13955 11512 14464 11540
rect 13955 11509 13967 11512
rect 13909 11503 13967 11509
rect 14458 11500 14464 11512
rect 14516 11500 14522 11552
rect 14550 11500 14556 11552
rect 14608 11540 14614 11552
rect 14737 11543 14795 11549
rect 14737 11540 14749 11543
rect 14608 11512 14749 11540
rect 14608 11500 14614 11512
rect 14737 11509 14749 11512
rect 14783 11509 14795 11543
rect 14737 11503 14795 11509
rect 14829 11543 14887 11549
rect 14829 11509 14841 11543
rect 14875 11540 14887 11543
rect 15470 11540 15476 11552
rect 14875 11512 15476 11540
rect 14875 11509 14887 11512
rect 14829 11503 14887 11509
rect 15470 11500 15476 11512
rect 15528 11500 15534 11552
rect 15746 11500 15752 11552
rect 15804 11540 15810 11552
rect 16482 11540 16488 11552
rect 15804 11512 16488 11540
rect 15804 11500 15810 11512
rect 16482 11500 16488 11512
rect 16540 11500 16546 11552
rect 16942 11540 16948 11552
rect 16903 11512 16948 11540
rect 16942 11500 16948 11512
rect 17000 11500 17006 11552
rect 17310 11540 17316 11552
rect 17271 11512 17316 11540
rect 17310 11500 17316 11512
rect 17368 11500 17374 11552
rect 17405 11543 17463 11549
rect 17405 11509 17417 11543
rect 17451 11540 17463 11543
rect 18049 11543 18107 11549
rect 18049 11540 18061 11543
rect 17451 11512 18061 11540
rect 17451 11509 17463 11512
rect 17405 11503 17463 11509
rect 18049 11509 18061 11512
rect 18095 11509 18107 11543
rect 18049 11503 18107 11509
rect 18509 11543 18567 11549
rect 18509 11509 18521 11543
rect 18555 11540 18567 11543
rect 18782 11540 18788 11552
rect 18555 11512 18788 11540
rect 18555 11509 18567 11512
rect 18509 11503 18567 11509
rect 18782 11500 18788 11512
rect 18840 11500 18846 11552
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 9674 11336 9680 11348
rect 9635 11308 9680 11336
rect 9674 11296 9680 11308
rect 9732 11296 9738 11348
rect 10042 11336 10048 11348
rect 10003 11308 10048 11336
rect 10042 11296 10048 11308
rect 10100 11296 10106 11348
rect 12066 11296 12072 11348
rect 12124 11336 12130 11348
rect 12345 11339 12403 11345
rect 12345 11336 12357 11339
rect 12124 11308 12357 11336
rect 12124 11296 12130 11308
rect 12345 11305 12357 11308
rect 12391 11305 12403 11339
rect 14182 11336 14188 11348
rect 14143 11308 14188 11336
rect 12345 11299 12403 11305
rect 14182 11296 14188 11308
rect 14240 11296 14246 11348
rect 15565 11339 15623 11345
rect 15565 11305 15577 11339
rect 15611 11336 15623 11339
rect 17310 11336 17316 11348
rect 15611 11308 17316 11336
rect 15611 11305 15623 11308
rect 15565 11299 15623 11305
rect 17310 11296 17316 11308
rect 17368 11296 17374 11348
rect 19242 11336 19248 11348
rect 18708 11308 19248 11336
rect 8941 11271 8999 11277
rect 8941 11237 8953 11271
rect 8987 11268 8999 11271
rect 9030 11268 9036 11280
rect 8987 11240 9036 11268
rect 8987 11237 8999 11240
rect 8941 11231 8999 11237
rect 9030 11228 9036 11240
rect 9088 11228 9094 11280
rect 12158 11268 12164 11280
rect 9416 11240 12164 11268
rect 9214 11200 9220 11212
rect 9048 11172 9220 11200
rect 9048 11141 9076 11172
rect 9214 11160 9220 11172
rect 9272 11200 9278 11212
rect 9416 11200 9444 11240
rect 12158 11228 12164 11240
rect 12216 11228 12222 11280
rect 16844 11271 16902 11277
rect 16844 11268 16856 11271
rect 16132 11240 16856 11268
rect 9272 11172 9444 11200
rect 9272 11160 9278 11172
rect 9490 11160 9496 11212
rect 9548 11200 9554 11212
rect 10962 11200 10968 11212
rect 9548 11172 10272 11200
rect 10923 11172 10968 11200
rect 9548 11160 9554 11172
rect 9033 11135 9091 11141
rect 9033 11101 9045 11135
rect 9079 11101 9091 11135
rect 9033 11095 9091 11101
rect 9122 11092 9128 11144
rect 9180 11132 9186 11144
rect 10244 11141 10272 11172
rect 10962 11160 10968 11172
rect 11020 11160 11026 11212
rect 11232 11203 11290 11209
rect 11232 11169 11244 11203
rect 11278 11200 11290 11203
rect 11790 11200 11796 11212
rect 11278 11172 11796 11200
rect 11278 11169 11290 11172
rect 11232 11163 11290 11169
rect 11790 11160 11796 11172
rect 11848 11160 11854 11212
rect 12897 11203 12955 11209
rect 12897 11169 12909 11203
rect 12943 11169 12955 11203
rect 12897 11163 12955 11169
rect 10137 11135 10195 11141
rect 9180 11104 9225 11132
rect 9180 11092 9186 11104
rect 10137 11101 10149 11135
rect 10183 11101 10195 11135
rect 10137 11095 10195 11101
rect 10229 11135 10287 11141
rect 10229 11101 10241 11135
rect 10275 11101 10287 11135
rect 12912 11132 12940 11163
rect 15746 11160 15752 11212
rect 15804 11200 15810 11212
rect 15933 11203 15991 11209
rect 15933 11200 15945 11203
rect 15804 11172 15945 11200
rect 15804 11160 15810 11172
rect 15933 11169 15945 11172
rect 15979 11169 15991 11203
rect 15933 11163 15991 11169
rect 16132 11141 16160 11240
rect 16844 11237 16856 11240
rect 16890 11268 16902 11271
rect 17218 11268 17224 11280
rect 16890 11240 17224 11268
rect 16890 11237 16902 11240
rect 16844 11231 16902 11237
rect 17218 11228 17224 11240
rect 17276 11228 17282 11280
rect 18414 11228 18420 11280
rect 18472 11268 18478 11280
rect 18708 11277 18736 11308
rect 19242 11296 19248 11308
rect 19300 11296 19306 11348
rect 18693 11271 18751 11277
rect 18693 11268 18705 11271
rect 18472 11240 18705 11268
rect 18472 11228 18478 11240
rect 18693 11237 18705 11240
rect 18739 11237 18751 11271
rect 18693 11231 18751 11237
rect 19058 11228 19064 11280
rect 19116 11268 19122 11280
rect 19981 11271 20039 11277
rect 19981 11268 19993 11271
rect 19116 11240 19993 11268
rect 19116 11228 19122 11240
rect 19981 11237 19993 11240
rect 20027 11237 20039 11271
rect 19981 11231 20039 11237
rect 17402 11160 17408 11212
rect 17460 11200 17466 11212
rect 17954 11200 17960 11212
rect 17460 11172 17960 11200
rect 17460 11160 17466 11172
rect 17954 11160 17960 11172
rect 18012 11160 18018 11212
rect 18598 11200 18604 11212
rect 18559 11172 18604 11200
rect 18598 11160 18604 11172
rect 18656 11160 18662 11212
rect 19889 11203 19947 11209
rect 19889 11169 19901 11203
rect 19935 11200 19947 11203
rect 20898 11200 20904 11212
rect 19935 11172 20904 11200
rect 19935 11169 19947 11172
rect 19889 11163 19947 11169
rect 20898 11160 20904 11172
rect 20956 11160 20962 11212
rect 16025 11135 16083 11141
rect 12912 11104 15976 11132
rect 10229 11095 10287 11101
rect 8573 11067 8631 11073
rect 8573 11033 8585 11067
rect 8619 11064 8631 11067
rect 10152 11064 10180 11095
rect 8619 11036 10180 11064
rect 8619 11033 8631 11036
rect 8573 11027 8631 11033
rect 14458 11024 14464 11076
rect 14516 11064 14522 11076
rect 15746 11064 15752 11076
rect 14516 11036 15752 11064
rect 14516 11024 14522 11036
rect 15746 11024 15752 11036
rect 15804 11024 15810 11076
rect 13722 10956 13728 11008
rect 13780 10996 13786 11008
rect 14366 10996 14372 11008
rect 13780 10968 14372 10996
rect 13780 10956 13786 10968
rect 14366 10956 14372 10968
rect 14424 10956 14430 11008
rect 15948 10996 15976 11104
rect 16025 11101 16037 11135
rect 16071 11101 16083 11135
rect 16025 11095 16083 11101
rect 16117 11135 16175 11141
rect 16117 11101 16129 11135
rect 16163 11101 16175 11135
rect 16117 11095 16175 11101
rect 16040 11064 16068 11095
rect 16390 11092 16396 11144
rect 16448 11132 16454 11144
rect 16577 11135 16635 11141
rect 16577 11132 16589 11135
rect 16448 11104 16589 11132
rect 16448 11092 16454 11104
rect 16577 11101 16589 11104
rect 16623 11101 16635 11135
rect 18785 11135 18843 11141
rect 18785 11132 18797 11135
rect 16577 11095 16635 11101
rect 17972 11104 18797 11132
rect 16482 11064 16488 11076
rect 16040 11036 16488 11064
rect 16482 11024 16488 11036
rect 16540 11024 16546 11076
rect 17678 11024 17684 11076
rect 17736 11064 17742 11076
rect 17972 11073 18000 11104
rect 18785 11101 18797 11104
rect 18831 11101 18843 11135
rect 18785 11095 18843 11101
rect 20070 11092 20076 11144
rect 20128 11132 20134 11144
rect 20128 11104 20173 11132
rect 20128 11092 20134 11104
rect 17957 11067 18015 11073
rect 17957 11064 17969 11067
rect 17736 11036 17969 11064
rect 17736 11024 17742 11036
rect 17957 11033 17969 11036
rect 18003 11033 18015 11067
rect 17957 11027 18015 11033
rect 18046 11024 18052 11076
rect 18104 11064 18110 11076
rect 18233 11067 18291 11073
rect 18233 11064 18245 11067
rect 18104 11036 18245 11064
rect 18104 11024 18110 11036
rect 18233 11033 18245 11036
rect 18279 11033 18291 11067
rect 20530 11064 20536 11076
rect 18233 11027 18291 11033
rect 18331 11036 20536 11064
rect 18331 10996 18359 11036
rect 20530 11024 20536 11036
rect 20588 11024 20594 11076
rect 15948 10968 18359 10996
rect 19334 10956 19340 11008
rect 19392 10996 19398 11008
rect 19521 10999 19579 11005
rect 19521 10996 19533 10999
rect 19392 10968 19533 10996
rect 19392 10956 19398 10968
rect 19521 10965 19533 10968
rect 19567 10965 19579 10999
rect 19521 10959 19579 10965
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 12434 10752 12440 10804
rect 12492 10792 12498 10804
rect 12492 10764 12537 10792
rect 12492 10752 12498 10764
rect 12986 10752 12992 10804
rect 13044 10792 13050 10804
rect 13449 10795 13507 10801
rect 13449 10792 13461 10795
rect 13044 10764 13461 10792
rect 13044 10752 13050 10764
rect 13449 10761 13461 10764
rect 13495 10761 13507 10795
rect 13449 10755 13507 10761
rect 13556 10764 14136 10792
rect 11333 10727 11391 10733
rect 11333 10693 11345 10727
rect 11379 10724 11391 10727
rect 12710 10724 12716 10736
rect 11379 10696 12716 10724
rect 11379 10693 11391 10696
rect 11333 10687 11391 10693
rect 12710 10684 12716 10696
rect 12768 10684 12774 10736
rect 11790 10616 11796 10668
rect 11848 10656 11854 10668
rect 11885 10659 11943 10665
rect 11885 10656 11897 10659
rect 11848 10628 11897 10656
rect 11848 10616 11854 10628
rect 11885 10625 11897 10628
rect 11931 10656 11943 10659
rect 13081 10659 13139 10665
rect 13081 10656 13093 10659
rect 11931 10628 13093 10656
rect 11931 10625 11943 10628
rect 11885 10619 11943 10625
rect 13081 10625 13093 10628
rect 13127 10656 13139 10659
rect 13556 10656 13584 10764
rect 13998 10724 14004 10736
rect 13127 10628 13584 10656
rect 13648 10696 14004 10724
rect 13127 10625 13139 10628
rect 13081 10619 13139 10625
rect 8021 10591 8079 10597
rect 8021 10557 8033 10591
rect 8067 10557 8079 10591
rect 8021 10551 8079 10557
rect 8288 10591 8346 10597
rect 8288 10557 8300 10591
rect 8334 10588 8346 10591
rect 9490 10588 9496 10600
rect 8334 10560 9496 10588
rect 8334 10557 8346 10560
rect 8288 10551 8346 10557
rect 8036 10520 8064 10551
rect 9490 10548 9496 10560
rect 9548 10548 9554 10600
rect 9674 10588 9680 10600
rect 9635 10560 9680 10588
rect 9674 10548 9680 10560
rect 9732 10548 9738 10600
rect 10597 10591 10655 10597
rect 10597 10557 10609 10591
rect 10643 10588 10655 10591
rect 11606 10588 11612 10600
rect 10643 10560 11612 10588
rect 10643 10557 10655 10560
rect 10597 10551 10655 10557
rect 11606 10548 11612 10560
rect 11664 10548 11670 10600
rect 11701 10591 11759 10597
rect 11701 10557 11713 10591
rect 11747 10588 11759 10591
rect 12434 10588 12440 10600
rect 11747 10560 12440 10588
rect 11747 10557 11759 10560
rect 11701 10551 11759 10557
rect 12434 10548 12440 10560
rect 12492 10548 12498 10600
rect 12710 10548 12716 10600
rect 12768 10588 12774 10600
rect 12897 10591 12955 10597
rect 12897 10588 12909 10591
rect 12768 10560 12909 10588
rect 12768 10548 12774 10560
rect 12897 10557 12909 10560
rect 12943 10588 12955 10591
rect 13648 10588 13676 10696
rect 13998 10684 14004 10696
rect 14056 10684 14062 10736
rect 14108 10665 14136 10764
rect 14366 10752 14372 10804
rect 14424 10792 14430 10804
rect 15102 10792 15108 10804
rect 14424 10764 15108 10792
rect 14424 10752 14430 10764
rect 15102 10752 15108 10764
rect 15160 10752 15166 10804
rect 15378 10792 15384 10804
rect 15339 10764 15384 10792
rect 15378 10752 15384 10764
rect 15436 10752 15442 10804
rect 16482 10792 16488 10804
rect 16316 10764 16488 10792
rect 14093 10659 14151 10665
rect 14093 10625 14105 10659
rect 14139 10625 14151 10659
rect 15102 10656 15108 10668
rect 15063 10628 15108 10656
rect 14093 10619 14151 10625
rect 15102 10616 15108 10628
rect 15160 10616 15166 10668
rect 15838 10656 15844 10668
rect 15799 10628 15844 10656
rect 15838 10616 15844 10628
rect 15896 10616 15902 10668
rect 16025 10659 16083 10665
rect 16025 10625 16037 10659
rect 16071 10656 16083 10659
rect 16206 10656 16212 10668
rect 16071 10628 16212 10656
rect 16071 10625 16083 10628
rect 16025 10619 16083 10625
rect 16206 10616 16212 10628
rect 16264 10616 16270 10668
rect 12943 10560 13676 10588
rect 12943 10557 12955 10560
rect 12897 10551 12955 10557
rect 13722 10548 13728 10600
rect 13780 10588 13786 10600
rect 13817 10591 13875 10597
rect 13817 10588 13829 10591
rect 13780 10560 13829 10588
rect 13780 10548 13786 10560
rect 13817 10557 13829 10560
rect 13863 10557 13875 10591
rect 13817 10551 13875 10557
rect 13909 10591 13967 10597
rect 13909 10557 13921 10591
rect 13955 10588 13967 10591
rect 14458 10588 14464 10600
rect 13955 10560 14464 10588
rect 13955 10557 13967 10560
rect 13909 10551 13967 10557
rect 14458 10548 14464 10560
rect 14516 10548 14522 10600
rect 14550 10548 14556 10600
rect 14608 10588 14614 10600
rect 15013 10591 15071 10597
rect 15013 10588 15025 10591
rect 14608 10560 15025 10588
rect 14608 10548 14614 10560
rect 15013 10557 15025 10560
rect 15059 10557 15071 10591
rect 15013 10551 15071 10557
rect 15286 10548 15292 10600
rect 15344 10588 15350 10600
rect 15749 10591 15807 10597
rect 15749 10588 15761 10591
rect 15344 10560 15761 10588
rect 15344 10548 15350 10560
rect 15749 10557 15761 10560
rect 15795 10557 15807 10591
rect 15749 10551 15807 10557
rect 16114 10548 16120 10600
rect 16172 10588 16178 10600
rect 16316 10597 16344 10764
rect 16482 10752 16488 10764
rect 16540 10752 16546 10804
rect 18506 10752 18512 10804
rect 18564 10792 18570 10804
rect 18601 10795 18659 10801
rect 18601 10792 18613 10795
rect 18564 10764 18613 10792
rect 18564 10752 18570 10764
rect 18601 10761 18613 10764
rect 18647 10761 18659 10795
rect 18601 10755 18659 10761
rect 17586 10684 17592 10736
rect 17644 10724 17650 10736
rect 18322 10724 18328 10736
rect 17644 10696 18328 10724
rect 17644 10684 17650 10696
rect 18322 10684 18328 10696
rect 18380 10684 18386 10736
rect 17678 10616 17684 10668
rect 17736 10616 17742 10668
rect 18049 10659 18107 10665
rect 18049 10625 18061 10659
rect 18095 10656 18107 10659
rect 18598 10656 18604 10668
rect 18095 10628 18604 10656
rect 18095 10625 18107 10628
rect 18049 10619 18107 10625
rect 18598 10616 18604 10628
rect 18656 10616 18662 10668
rect 19245 10659 19303 10665
rect 19245 10625 19257 10659
rect 19291 10656 19303 10659
rect 19291 10628 19564 10656
rect 19291 10625 19303 10628
rect 19245 10619 19303 10625
rect 16301 10591 16359 10597
rect 16301 10588 16313 10591
rect 16172 10560 16313 10588
rect 16172 10548 16178 10560
rect 16301 10557 16313 10560
rect 16347 10557 16359 10591
rect 16301 10551 16359 10557
rect 16568 10591 16626 10597
rect 16568 10557 16580 10591
rect 16614 10588 16626 10591
rect 17696 10588 17724 10616
rect 16614 10560 17724 10588
rect 18969 10591 19027 10597
rect 16614 10557 16626 10560
rect 16568 10551 16626 10557
rect 18969 10557 18981 10591
rect 19015 10588 19027 10591
rect 19334 10588 19340 10600
rect 19015 10560 19340 10588
rect 19015 10557 19027 10560
rect 18969 10551 19027 10557
rect 19334 10548 19340 10560
rect 19392 10548 19398 10600
rect 8202 10520 8208 10532
rect 8036 10492 8208 10520
rect 8202 10480 8208 10492
rect 8260 10480 8266 10532
rect 9953 10523 10011 10529
rect 9953 10489 9965 10523
rect 9999 10520 10011 10523
rect 14921 10523 14979 10529
rect 9999 10492 14872 10520
rect 9999 10489 10011 10492
rect 9953 10483 10011 10489
rect 9214 10412 9220 10464
rect 9272 10452 9278 10464
rect 9401 10455 9459 10461
rect 9401 10452 9413 10455
rect 9272 10424 9413 10452
rect 9272 10412 9278 10424
rect 9401 10421 9413 10424
rect 9447 10421 9459 10455
rect 9401 10415 9459 10421
rect 10413 10455 10471 10461
rect 10413 10421 10425 10455
rect 10459 10452 10471 10455
rect 10686 10452 10692 10464
rect 10459 10424 10692 10452
rect 10459 10421 10471 10424
rect 10413 10415 10471 10421
rect 10686 10412 10692 10424
rect 10744 10412 10750 10464
rect 10870 10412 10876 10464
rect 10928 10452 10934 10464
rect 11793 10455 11851 10461
rect 11793 10452 11805 10455
rect 10928 10424 11805 10452
rect 10928 10412 10934 10424
rect 11793 10421 11805 10424
rect 11839 10421 11851 10455
rect 11793 10415 11851 10421
rect 12618 10412 12624 10464
rect 12676 10452 12682 10464
rect 12802 10452 12808 10464
rect 12676 10424 12808 10452
rect 12676 10412 12682 10424
rect 12802 10412 12808 10424
rect 12860 10412 12866 10464
rect 13998 10412 14004 10464
rect 14056 10452 14062 10464
rect 14553 10455 14611 10461
rect 14553 10452 14565 10455
rect 14056 10424 14565 10452
rect 14056 10412 14062 10424
rect 14553 10421 14565 10424
rect 14599 10421 14611 10455
rect 14844 10452 14872 10492
rect 14921 10489 14933 10523
rect 14967 10520 14979 10523
rect 16390 10520 16396 10532
rect 14967 10492 16396 10520
rect 14967 10489 14979 10492
rect 14921 10483 14979 10489
rect 16390 10480 16396 10492
rect 16448 10480 16454 10532
rect 19426 10520 19432 10532
rect 16500 10492 19432 10520
rect 16500 10452 16528 10492
rect 19426 10480 19432 10492
rect 19484 10480 19490 10532
rect 19536 10520 19564 10628
rect 19610 10548 19616 10600
rect 19668 10588 19674 10600
rect 19668 10560 19713 10588
rect 19668 10548 19674 10560
rect 19880 10523 19938 10529
rect 19880 10520 19892 10523
rect 19536 10492 19892 10520
rect 19880 10489 19892 10492
rect 19926 10520 19938 10523
rect 20438 10520 20444 10532
rect 19926 10492 20444 10520
rect 19926 10489 19938 10492
rect 19880 10483 19938 10489
rect 20438 10480 20444 10492
rect 20496 10480 20502 10532
rect 14844 10424 16528 10452
rect 17681 10455 17739 10461
rect 14553 10415 14611 10421
rect 17681 10421 17693 10455
rect 17727 10452 17739 10455
rect 18046 10452 18052 10464
rect 17727 10424 18052 10452
rect 17727 10421 17739 10424
rect 17681 10415 17739 10421
rect 18046 10412 18052 10424
rect 18104 10412 18110 10464
rect 19058 10452 19064 10464
rect 19019 10424 19064 10452
rect 19058 10412 19064 10424
rect 19116 10412 19122 10464
rect 19334 10412 19340 10464
rect 19392 10452 19398 10464
rect 19978 10452 19984 10464
rect 19392 10424 19984 10452
rect 19392 10412 19398 10424
rect 19978 10412 19984 10424
rect 20036 10452 20042 10464
rect 20993 10455 21051 10461
rect 20993 10452 21005 10455
rect 20036 10424 21005 10452
rect 20036 10412 20042 10424
rect 20993 10421 21005 10424
rect 21039 10421 21051 10455
rect 20993 10415 21051 10421
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 9674 10248 9680 10260
rect 9635 10220 9680 10248
rect 9674 10208 9680 10220
rect 9732 10208 9738 10260
rect 11790 10208 11796 10260
rect 11848 10248 11854 10260
rect 12069 10251 12127 10257
rect 12069 10248 12081 10251
rect 11848 10220 12081 10248
rect 11848 10208 11854 10220
rect 12069 10217 12081 10220
rect 12115 10217 12127 10251
rect 12069 10211 12127 10217
rect 13633 10251 13691 10257
rect 13633 10217 13645 10251
rect 13679 10248 13691 10251
rect 14185 10251 14243 10257
rect 14185 10248 14197 10251
rect 13679 10220 14197 10248
rect 13679 10217 13691 10220
rect 13633 10211 13691 10217
rect 14185 10217 14197 10220
rect 14231 10217 14243 10251
rect 14185 10211 14243 10217
rect 14645 10251 14703 10257
rect 14645 10217 14657 10251
rect 14691 10248 14703 10251
rect 15289 10251 15347 10257
rect 15289 10248 15301 10251
rect 14691 10220 15301 10248
rect 14691 10217 14703 10220
rect 14645 10211 14703 10217
rect 15289 10217 15301 10220
rect 15335 10217 15347 10251
rect 16761 10251 16819 10257
rect 16761 10248 16773 10251
rect 15289 10211 15347 10217
rect 16132 10220 16773 10248
rect 9950 10140 9956 10192
rect 10008 10180 10014 10192
rect 10778 10180 10784 10192
rect 10008 10152 10784 10180
rect 10008 10140 10014 10152
rect 10778 10140 10784 10152
rect 10836 10140 10842 10192
rect 10956 10183 11014 10189
rect 10956 10149 10968 10183
rect 11002 10180 11014 10183
rect 11146 10180 11152 10192
rect 11002 10152 11152 10180
rect 11002 10149 11014 10152
rect 10956 10143 11014 10149
rect 11146 10140 11152 10152
rect 11204 10140 11210 10192
rect 11882 10140 11888 10192
rect 11940 10180 11946 10192
rect 12621 10183 12679 10189
rect 12621 10180 12633 10183
rect 11940 10152 12633 10180
rect 11940 10140 11946 10152
rect 12621 10149 12633 10152
rect 12667 10149 12679 10183
rect 12621 10143 12679 10149
rect 13541 10183 13599 10189
rect 13541 10149 13553 10183
rect 13587 10180 13599 10183
rect 13998 10180 14004 10192
rect 13587 10152 14004 10180
rect 13587 10149 13599 10152
rect 13541 10143 13599 10149
rect 13998 10140 14004 10152
rect 14056 10140 14062 10192
rect 14274 10140 14280 10192
rect 14332 10180 14338 10192
rect 15010 10180 15016 10192
rect 14332 10152 15016 10180
rect 14332 10140 14338 10152
rect 15010 10140 15016 10152
rect 15068 10180 15074 10192
rect 15749 10183 15807 10189
rect 15749 10180 15761 10183
rect 15068 10152 15761 10180
rect 15068 10140 15074 10152
rect 15749 10149 15761 10152
rect 15795 10149 15807 10183
rect 15749 10143 15807 10149
rect 9125 10115 9183 10121
rect 9125 10081 9137 10115
rect 9171 10112 9183 10115
rect 10045 10115 10103 10121
rect 10045 10112 10057 10115
rect 9171 10084 10057 10112
rect 9171 10081 9183 10084
rect 9125 10075 9183 10081
rect 10045 10081 10057 10084
rect 10091 10081 10103 10115
rect 12342 10112 12348 10124
rect 12303 10084 12348 10112
rect 10045 10075 10103 10081
rect 12342 10072 12348 10084
rect 12400 10072 12406 10124
rect 14553 10115 14611 10121
rect 14553 10081 14565 10115
rect 14599 10112 14611 10115
rect 15562 10112 15568 10124
rect 14599 10084 15568 10112
rect 14599 10081 14611 10084
rect 14553 10075 14611 10081
rect 15562 10072 15568 10084
rect 15620 10072 15626 10124
rect 16132 10121 16160 10220
rect 16761 10217 16773 10220
rect 16807 10217 16819 10251
rect 16761 10211 16819 10217
rect 16942 10208 16948 10260
rect 17000 10248 17006 10260
rect 17221 10251 17279 10257
rect 17221 10248 17233 10251
rect 17000 10220 17233 10248
rect 17000 10208 17006 10220
rect 17221 10217 17233 10220
rect 17267 10217 17279 10251
rect 17221 10211 17279 10217
rect 18049 10251 18107 10257
rect 18049 10217 18061 10251
rect 18095 10248 18107 10251
rect 19058 10248 19064 10260
rect 18095 10220 19064 10248
rect 18095 10217 18107 10220
rect 18049 10211 18107 10217
rect 19058 10208 19064 10220
rect 19116 10208 19122 10260
rect 20438 10248 20444 10260
rect 20399 10220 20444 10248
rect 20438 10208 20444 10220
rect 20496 10208 20502 10260
rect 20898 10248 20904 10260
rect 20859 10220 20904 10248
rect 20898 10208 20904 10220
rect 20956 10208 20962 10260
rect 16393 10183 16451 10189
rect 16393 10149 16405 10183
rect 16439 10180 16451 10183
rect 17034 10180 17040 10192
rect 16439 10152 17040 10180
rect 16439 10149 16451 10152
rect 16393 10143 16451 10149
rect 17034 10140 17040 10152
rect 17092 10140 17098 10192
rect 17129 10183 17187 10189
rect 17129 10149 17141 10183
rect 17175 10180 17187 10183
rect 17954 10180 17960 10192
rect 17175 10152 17960 10180
rect 17175 10149 17187 10152
rect 17129 10143 17187 10149
rect 17954 10140 17960 10152
rect 18012 10140 18018 10192
rect 19328 10183 19386 10189
rect 19328 10180 19340 10183
rect 18708 10152 19340 10180
rect 15657 10115 15715 10121
rect 15657 10081 15669 10115
rect 15703 10112 15715 10115
rect 16117 10115 16175 10121
rect 15703 10084 15884 10112
rect 15703 10081 15715 10084
rect 15657 10075 15715 10081
rect 10134 10044 10140 10056
rect 10095 10016 10140 10044
rect 10134 10004 10140 10016
rect 10192 10004 10198 10056
rect 10229 10047 10287 10053
rect 10229 10013 10241 10047
rect 10275 10013 10287 10047
rect 10686 10044 10692 10056
rect 10647 10016 10692 10044
rect 10229 10007 10287 10013
rect 9582 9936 9588 9988
rect 9640 9976 9646 9988
rect 10244 9976 10272 10007
rect 10686 10004 10692 10016
rect 10744 10004 10750 10056
rect 13722 10044 13728 10056
rect 13683 10016 13728 10044
rect 13722 10004 13728 10016
rect 13780 10004 13786 10056
rect 13998 10004 14004 10056
rect 14056 10044 14062 10056
rect 14737 10047 14795 10053
rect 14737 10044 14749 10047
rect 14056 10016 14749 10044
rect 14056 10004 14062 10016
rect 14737 10013 14749 10016
rect 14783 10044 14795 10047
rect 15102 10044 15108 10056
rect 14783 10016 15108 10044
rect 14783 10013 14795 10016
rect 14737 10007 14795 10013
rect 15102 10004 15108 10016
rect 15160 10004 15166 10056
rect 9640 9948 10272 9976
rect 9640 9936 9646 9948
rect 12434 9936 12440 9988
rect 12492 9976 12498 9988
rect 14918 9976 14924 9988
rect 12492 9948 14924 9976
rect 12492 9936 12498 9948
rect 14918 9936 14924 9948
rect 14976 9936 14982 9988
rect 15856 9976 15884 10084
rect 16117 10081 16129 10115
rect 16163 10081 16175 10115
rect 16117 10075 16175 10081
rect 16669 10115 16727 10121
rect 16669 10081 16681 10115
rect 16715 10112 16727 10115
rect 16758 10112 16764 10124
rect 16715 10084 16764 10112
rect 16715 10081 16727 10084
rect 16669 10075 16727 10081
rect 16758 10072 16764 10084
rect 16816 10112 16822 10124
rect 18417 10115 18475 10121
rect 18417 10112 18429 10115
rect 16816 10084 18429 10112
rect 16816 10072 16822 10084
rect 18417 10081 18429 10084
rect 18463 10081 18475 10115
rect 18417 10075 18475 10081
rect 15933 10047 15991 10053
rect 15933 10013 15945 10047
rect 15979 10044 15991 10047
rect 16206 10044 16212 10056
rect 15979 10016 16212 10044
rect 15979 10013 15991 10016
rect 15933 10007 15991 10013
rect 16206 10004 16212 10016
rect 16264 10044 16270 10056
rect 16482 10044 16488 10056
rect 16264 10016 16488 10044
rect 16264 10004 16270 10016
rect 16482 10004 16488 10016
rect 16540 10004 16546 10056
rect 17405 10047 17463 10053
rect 17405 10013 17417 10047
rect 17451 10044 17463 10047
rect 17954 10044 17960 10056
rect 17451 10016 17960 10044
rect 17451 10013 17463 10016
rect 17405 10007 17463 10013
rect 17954 10004 17960 10016
rect 18012 10004 18018 10056
rect 18506 10044 18512 10056
rect 18467 10016 18512 10044
rect 18506 10004 18512 10016
rect 18564 10004 18570 10056
rect 18708 10053 18736 10152
rect 19328 10149 19340 10152
rect 19374 10180 19386 10183
rect 20070 10180 20076 10192
rect 19374 10152 20076 10180
rect 19374 10149 19386 10152
rect 19328 10143 19386 10149
rect 20070 10140 20076 10152
rect 20128 10140 20134 10192
rect 19610 10112 19616 10124
rect 19076 10084 19616 10112
rect 19076 10056 19104 10084
rect 19610 10072 19616 10084
rect 19668 10072 19674 10124
rect 18693 10047 18751 10053
rect 18693 10013 18705 10047
rect 18739 10013 18751 10047
rect 19058 10044 19064 10056
rect 19019 10016 19064 10044
rect 18693 10007 18751 10013
rect 19058 10004 19064 10016
rect 19116 10004 19122 10056
rect 16298 9976 16304 9988
rect 15856 9948 16304 9976
rect 16298 9936 16304 9948
rect 16356 9976 16362 9988
rect 18598 9976 18604 9988
rect 16356 9948 18604 9976
rect 16356 9936 16362 9948
rect 18598 9936 18604 9948
rect 18656 9936 18662 9988
rect 12986 9868 12992 9920
rect 13044 9908 13050 9920
rect 13173 9911 13231 9917
rect 13173 9908 13185 9911
rect 13044 9880 13185 9908
rect 13044 9868 13050 9880
rect 13173 9877 13185 9880
rect 13219 9877 13231 9911
rect 13173 9871 13231 9877
rect 14366 9868 14372 9920
rect 14424 9908 14430 9920
rect 16669 9911 16727 9917
rect 16669 9908 16681 9911
rect 14424 9880 16681 9908
rect 14424 9868 14430 9880
rect 16669 9877 16681 9880
rect 16715 9877 16727 9911
rect 16669 9871 16727 9877
rect 17586 9868 17592 9920
rect 17644 9908 17650 9920
rect 19242 9908 19248 9920
rect 17644 9880 19248 9908
rect 17644 9868 17650 9880
rect 19242 9868 19248 9880
rect 19300 9868 19306 9920
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 9306 9664 9312 9716
rect 9364 9704 9370 9716
rect 14366 9704 14372 9716
rect 9364 9676 14372 9704
rect 9364 9664 9370 9676
rect 14366 9664 14372 9676
rect 14424 9664 14430 9716
rect 15746 9704 15752 9716
rect 14476 9676 15752 9704
rect 11146 9596 11152 9648
rect 11204 9636 11210 9648
rect 11425 9639 11483 9645
rect 11425 9636 11437 9639
rect 11204 9608 11437 9636
rect 11204 9596 11210 9608
rect 11425 9605 11437 9608
rect 11471 9636 11483 9639
rect 11882 9636 11888 9648
rect 11471 9608 11888 9636
rect 11471 9605 11483 9608
rect 11425 9599 11483 9605
rect 11882 9596 11888 9608
rect 11940 9596 11946 9648
rect 14476 9577 14504 9676
rect 15746 9664 15752 9676
rect 15804 9704 15810 9716
rect 16758 9704 16764 9716
rect 15804 9676 16764 9704
rect 15804 9664 15810 9676
rect 16758 9664 16764 9676
rect 16816 9704 16822 9716
rect 17405 9707 17463 9713
rect 17405 9704 17417 9707
rect 16816 9676 17417 9704
rect 16816 9664 16822 9676
rect 17405 9673 17417 9676
rect 17451 9704 17463 9707
rect 19058 9704 19064 9716
rect 17451 9676 19064 9704
rect 17451 9673 17463 9676
rect 17405 9667 17463 9673
rect 15562 9596 15568 9648
rect 15620 9636 15626 9648
rect 16117 9639 16175 9645
rect 16117 9636 16129 9639
rect 15620 9608 16129 9636
rect 15620 9596 15626 9608
rect 16117 9605 16129 9608
rect 16163 9605 16175 9639
rect 16117 9599 16175 9605
rect 16206 9596 16212 9648
rect 16264 9636 16270 9648
rect 16264 9608 17632 9636
rect 16264 9596 16270 9608
rect 14461 9571 14519 9577
rect 14461 9537 14473 9571
rect 14507 9537 14519 9571
rect 14461 9531 14519 9537
rect 15838 9528 15844 9580
rect 15896 9568 15902 9580
rect 15896 9540 16436 9568
rect 15896 9528 15902 9540
rect 8202 9500 8208 9512
rect 8115 9472 8208 9500
rect 8202 9460 8208 9472
rect 8260 9460 8266 9512
rect 8472 9503 8530 9509
rect 8472 9469 8484 9503
rect 8518 9500 8530 9503
rect 9214 9500 9220 9512
rect 8518 9472 9220 9500
rect 8518 9469 8530 9472
rect 8472 9463 8530 9469
rect 9214 9460 9220 9472
rect 9272 9460 9278 9512
rect 9674 9460 9680 9512
rect 9732 9500 9738 9512
rect 10045 9503 10103 9509
rect 10045 9500 10057 9503
rect 9732 9472 10057 9500
rect 9732 9460 9738 9472
rect 10045 9469 10057 9472
rect 10091 9500 10103 9503
rect 10686 9500 10692 9512
rect 10091 9472 10692 9500
rect 10091 9469 10103 9472
rect 10045 9463 10103 9469
rect 10686 9460 10692 9472
rect 10744 9500 10750 9512
rect 12434 9500 12440 9512
rect 10744 9472 12440 9500
rect 10744 9460 10750 9472
rect 12434 9460 12440 9472
rect 12492 9500 12498 9512
rect 12704 9503 12762 9509
rect 12492 9472 12537 9500
rect 12492 9460 12498 9472
rect 12704 9469 12716 9503
rect 12750 9500 12762 9503
rect 13998 9500 14004 9512
rect 12750 9472 14004 9500
rect 12750 9469 12762 9472
rect 12704 9463 12762 9469
rect 13998 9460 14004 9472
rect 14056 9460 14062 9512
rect 14182 9460 14188 9512
rect 14240 9500 14246 9512
rect 14277 9503 14335 9509
rect 14277 9500 14289 9503
rect 14240 9472 14289 9500
rect 14240 9460 14246 9472
rect 14277 9469 14289 9472
rect 14323 9469 14335 9503
rect 14277 9463 14335 9469
rect 14728 9503 14786 9509
rect 14728 9469 14740 9503
rect 14774 9500 14786 9503
rect 16114 9500 16120 9512
rect 14774 9472 16120 9500
rect 14774 9469 14786 9472
rect 14728 9463 14786 9469
rect 16114 9460 16120 9472
rect 16172 9460 16178 9512
rect 16408 9500 16436 9540
rect 16482 9528 16488 9580
rect 16540 9568 16546 9580
rect 16669 9571 16727 9577
rect 16669 9568 16681 9571
rect 16540 9540 16681 9568
rect 16540 9528 16546 9540
rect 16669 9537 16681 9540
rect 16715 9537 16727 9571
rect 16669 9531 16727 9537
rect 17604 9509 17632 9608
rect 18064 9577 18092 9676
rect 19058 9664 19064 9676
rect 19116 9664 19122 9716
rect 20162 9664 20168 9716
rect 20220 9704 20226 9716
rect 20806 9704 20812 9716
rect 20220 9676 20812 9704
rect 20220 9664 20226 9676
rect 20806 9664 20812 9676
rect 20864 9664 20870 9716
rect 18049 9571 18107 9577
rect 18049 9537 18061 9571
rect 18095 9537 18107 9571
rect 20530 9568 20536 9580
rect 20491 9540 20536 9568
rect 18049 9531 18107 9537
rect 20530 9528 20536 9540
rect 20588 9528 20594 9580
rect 20622 9528 20628 9580
rect 20680 9568 20686 9580
rect 20680 9540 20725 9568
rect 20680 9528 20686 9540
rect 16577 9503 16635 9509
rect 16577 9500 16589 9503
rect 16408 9472 16589 9500
rect 16577 9469 16589 9472
rect 16623 9469 16635 9503
rect 16577 9463 16635 9469
rect 17589 9503 17647 9509
rect 17589 9469 17601 9503
rect 17635 9469 17647 9503
rect 17589 9463 17647 9469
rect 18138 9460 18144 9512
rect 18196 9500 18202 9512
rect 20548 9500 20576 9528
rect 18196 9472 20576 9500
rect 18196 9460 18202 9472
rect 8220 9432 8248 9460
rect 9692 9432 9720 9460
rect 10318 9441 10324 9444
rect 10312 9432 10324 9441
rect 8220 9404 9720 9432
rect 10279 9404 10324 9432
rect 10312 9395 10324 9404
rect 10318 9392 10324 9395
rect 10376 9392 10382 9444
rect 14918 9392 14924 9444
rect 14976 9432 14982 9444
rect 15286 9432 15292 9444
rect 14976 9404 15292 9432
rect 14976 9392 14982 9404
rect 15286 9392 15292 9404
rect 15344 9392 15350 9444
rect 15470 9392 15476 9444
rect 15528 9432 15534 9444
rect 15528 9404 16344 9432
rect 15528 9392 15534 9404
rect 16316 9376 16344 9404
rect 16390 9392 16396 9444
rect 16448 9432 16454 9444
rect 16945 9435 17003 9441
rect 16945 9432 16957 9435
rect 16448 9404 16957 9432
rect 16448 9392 16454 9404
rect 16945 9401 16957 9404
rect 16991 9401 17003 9435
rect 16945 9395 17003 9401
rect 17954 9392 17960 9444
rect 18012 9432 18018 9444
rect 18294 9435 18352 9441
rect 18294 9432 18306 9435
rect 18012 9404 18306 9432
rect 18012 9392 18018 9404
rect 18294 9401 18306 9404
rect 18340 9401 18352 9435
rect 18294 9395 18352 9401
rect 20441 9435 20499 9441
rect 20441 9401 20453 9435
rect 20487 9432 20499 9435
rect 20898 9432 20904 9444
rect 20487 9404 20904 9432
rect 20487 9401 20499 9404
rect 20441 9395 20499 9401
rect 20898 9392 20904 9404
rect 20956 9392 20962 9444
rect 9582 9364 9588 9376
rect 9543 9336 9588 9364
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 11698 9364 11704 9376
rect 11659 9336 11704 9364
rect 11698 9324 11704 9336
rect 11756 9324 11762 9376
rect 13722 9324 13728 9376
rect 13780 9364 13786 9376
rect 13817 9367 13875 9373
rect 13817 9364 13829 9367
rect 13780 9336 13829 9364
rect 13780 9324 13786 9336
rect 13817 9333 13829 9336
rect 13863 9333 13875 9367
rect 13817 9327 13875 9333
rect 13998 9324 14004 9376
rect 14056 9364 14062 9376
rect 14093 9367 14151 9373
rect 14093 9364 14105 9367
rect 14056 9336 14105 9364
rect 14056 9324 14062 9336
rect 14093 9333 14105 9336
rect 14139 9333 14151 9367
rect 14093 9327 14151 9333
rect 15102 9324 15108 9376
rect 15160 9364 15166 9376
rect 15841 9367 15899 9373
rect 15841 9364 15853 9367
rect 15160 9336 15853 9364
rect 15160 9324 15166 9336
rect 15841 9333 15853 9336
rect 15887 9333 15899 9367
rect 15841 9327 15899 9333
rect 16298 9324 16304 9376
rect 16356 9364 16362 9376
rect 16485 9367 16543 9373
rect 16485 9364 16497 9367
rect 16356 9336 16497 9364
rect 16356 9324 16362 9336
rect 16485 9333 16497 9336
rect 16531 9333 16543 9367
rect 19426 9364 19432 9376
rect 19387 9336 19432 9364
rect 16485 9327 16543 9333
rect 19426 9324 19432 9336
rect 19484 9324 19490 9376
rect 19518 9324 19524 9376
rect 19576 9364 19582 9376
rect 20073 9367 20131 9373
rect 20073 9364 20085 9367
rect 19576 9336 20085 9364
rect 19576 9324 19582 9336
rect 20073 9333 20085 9336
rect 20119 9333 20131 9367
rect 20073 9327 20131 9333
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 8573 9163 8631 9169
rect 8573 9129 8585 9163
rect 8619 9160 8631 9163
rect 10134 9160 10140 9172
rect 8619 9132 10140 9160
rect 8619 9129 8631 9132
rect 8573 9123 8631 9129
rect 10134 9120 10140 9132
rect 10192 9120 10198 9172
rect 10318 9120 10324 9172
rect 10376 9160 10382 9172
rect 10962 9160 10968 9172
rect 10376 9132 10968 9160
rect 10376 9120 10382 9132
rect 10962 9120 10968 9132
rect 11020 9160 11026 9172
rect 11057 9163 11115 9169
rect 11057 9160 11069 9163
rect 11020 9132 11069 9160
rect 11020 9120 11026 9132
rect 11057 9129 11069 9132
rect 11103 9129 11115 9163
rect 11057 9123 11115 9129
rect 11333 9163 11391 9169
rect 11333 9129 11345 9163
rect 11379 9160 11391 9163
rect 12342 9160 12348 9172
rect 11379 9132 12348 9160
rect 11379 9129 11391 9132
rect 11333 9123 11391 9129
rect 12342 9120 12348 9132
rect 12400 9120 12406 9172
rect 16482 9120 16488 9172
rect 16540 9160 16546 9172
rect 17129 9163 17187 9169
rect 17129 9160 17141 9163
rect 16540 9132 17141 9160
rect 16540 9120 16546 9132
rect 17129 9129 17141 9132
rect 17175 9129 17187 9163
rect 17129 9123 17187 9129
rect 17589 9163 17647 9169
rect 17589 9129 17601 9163
rect 17635 9160 17647 9163
rect 18506 9160 18512 9172
rect 17635 9132 18512 9160
rect 17635 9129 17647 9132
rect 17589 9123 17647 9129
rect 18506 9120 18512 9132
rect 18564 9120 18570 9172
rect 19978 9160 19984 9172
rect 19939 9132 19984 9160
rect 19978 9120 19984 9132
rect 20036 9120 20042 9172
rect 9033 9095 9091 9101
rect 9033 9061 9045 9095
rect 9079 9092 9091 9095
rect 12526 9092 12532 9104
rect 9079 9064 12532 9092
rect 9079 9061 9091 9064
rect 9033 9055 9091 9061
rect 12526 9052 12532 9064
rect 12584 9052 12590 9104
rect 13256 9095 13314 9101
rect 13256 9061 13268 9095
rect 13302 9092 13314 9095
rect 13722 9092 13728 9104
rect 13302 9064 13728 9092
rect 13302 9061 13314 9064
rect 13256 9055 13314 9061
rect 13722 9052 13728 9064
rect 13780 9052 13786 9104
rect 16298 9052 16304 9104
rect 16356 9092 16362 9104
rect 17957 9095 18015 9101
rect 16356 9064 17080 9092
rect 16356 9052 16362 9064
rect 6914 8984 6920 9036
rect 6972 9024 6978 9036
rect 8941 9027 8999 9033
rect 8941 9024 8953 9027
rect 6972 8996 8953 9024
rect 6972 8984 6978 8996
rect 8941 8993 8953 8996
rect 8987 8993 8999 9027
rect 9674 9024 9680 9036
rect 9635 8996 9680 9024
rect 8941 8987 8999 8993
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 9944 9027 10002 9033
rect 9944 8993 9956 9027
rect 9990 9024 10002 9027
rect 10502 9024 10508 9036
rect 9990 8996 10508 9024
rect 9990 8993 10002 8996
rect 9944 8987 10002 8993
rect 10502 8984 10508 8996
rect 10560 8984 10566 9036
rect 10870 8984 10876 9036
rect 10928 9024 10934 9036
rect 11701 9027 11759 9033
rect 11701 9024 11713 9027
rect 10928 8996 11713 9024
rect 10928 8984 10934 8996
rect 11701 8993 11713 8996
rect 11747 8993 11759 9027
rect 11701 8987 11759 8993
rect 11974 8984 11980 9036
rect 12032 9024 12038 9036
rect 12342 9024 12348 9036
rect 12032 8996 12348 9024
rect 12032 8984 12038 8996
rect 12342 8984 12348 8996
rect 12400 8984 12406 9036
rect 12434 8984 12440 9036
rect 12492 9024 12498 9036
rect 12989 9027 13047 9033
rect 12989 9024 13001 9027
rect 12492 8996 13001 9024
rect 12492 8984 12498 8996
rect 12989 8993 13001 8996
rect 13035 8993 13047 9027
rect 15746 9024 15752 9036
rect 15707 8996 15752 9024
rect 12989 8987 13047 8993
rect 15746 8984 15752 8996
rect 15804 8984 15810 9036
rect 16016 9027 16074 9033
rect 16016 8993 16028 9027
rect 16062 9024 16074 9027
rect 16942 9024 16948 9036
rect 16062 8996 16948 9024
rect 16062 8993 16074 8996
rect 16016 8987 16074 8993
rect 16942 8984 16948 8996
rect 17000 8984 17006 9036
rect 17052 9024 17080 9064
rect 17957 9061 17969 9095
rect 18003 9092 18015 9095
rect 18138 9092 18144 9104
rect 18003 9064 18144 9092
rect 18003 9061 18015 9064
rect 17957 9055 18015 9061
rect 18138 9052 18144 9064
rect 18196 9052 18202 9104
rect 18868 9095 18926 9101
rect 18868 9092 18880 9095
rect 18524 9064 18880 9092
rect 18322 9024 18328 9036
rect 17052 8996 18328 9024
rect 18322 8984 18328 8996
rect 18380 8984 18386 9036
rect 9214 8956 9220 8968
rect 9175 8928 9220 8956
rect 9214 8916 9220 8928
rect 9272 8916 9278 8968
rect 11790 8956 11796 8968
rect 11751 8928 11796 8956
rect 11790 8916 11796 8928
rect 11848 8916 11854 8968
rect 11882 8916 11888 8968
rect 11940 8956 11946 8968
rect 18049 8959 18107 8965
rect 11940 8928 11985 8956
rect 11940 8916 11946 8928
rect 18049 8925 18061 8959
rect 18095 8925 18107 8959
rect 18049 8919 18107 8925
rect 18233 8959 18291 8965
rect 18233 8925 18245 8959
rect 18279 8956 18291 8959
rect 18524 8956 18552 9064
rect 18868 9061 18880 9064
rect 18914 9092 18926 9095
rect 19426 9092 19432 9104
rect 18914 9064 19432 9092
rect 18914 9061 18926 9064
rect 18868 9055 18926 9061
rect 19426 9052 19432 9064
rect 19484 9052 19490 9104
rect 18601 9027 18659 9033
rect 18601 8993 18613 9027
rect 18647 9024 18659 9027
rect 19150 9024 19156 9036
rect 18647 8996 19156 9024
rect 18647 8993 18659 8996
rect 18601 8987 18659 8993
rect 19150 8984 19156 8996
rect 19208 8984 19214 9036
rect 18279 8928 18552 8956
rect 18279 8925 18291 8928
rect 18233 8919 18291 8925
rect 12894 8888 12900 8900
rect 11532 8860 12900 8888
rect 8846 8780 8852 8832
rect 8904 8820 8910 8832
rect 11532 8820 11560 8860
rect 12894 8848 12900 8860
rect 12952 8848 12958 8900
rect 15654 8888 15660 8900
rect 13924 8860 15660 8888
rect 8904 8792 11560 8820
rect 8904 8780 8910 8792
rect 11606 8780 11612 8832
rect 11664 8820 11670 8832
rect 11882 8820 11888 8832
rect 11664 8792 11888 8820
rect 11664 8780 11670 8792
rect 11882 8780 11888 8792
rect 11940 8780 11946 8832
rect 11974 8780 11980 8832
rect 12032 8820 12038 8832
rect 13924 8820 13952 8860
rect 15654 8848 15660 8860
rect 15712 8848 15718 8900
rect 18064 8888 18092 8919
rect 18506 8888 18512 8900
rect 18064 8860 18512 8888
rect 18506 8848 18512 8860
rect 18564 8848 18570 8900
rect 14366 8820 14372 8832
rect 12032 8792 13952 8820
rect 14327 8792 14372 8820
rect 12032 8780 12038 8792
rect 14366 8780 14372 8792
rect 14424 8780 14430 8832
rect 14458 8780 14464 8832
rect 14516 8820 14522 8832
rect 17954 8820 17960 8832
rect 14516 8792 17960 8820
rect 14516 8780 14522 8792
rect 17954 8780 17960 8792
rect 18012 8780 18018 8832
rect 18598 8780 18604 8832
rect 18656 8820 18662 8832
rect 19978 8820 19984 8832
rect 18656 8792 19984 8820
rect 18656 8780 18662 8792
rect 19978 8780 19984 8792
rect 20036 8780 20042 8832
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 3418 8576 3424 8628
rect 3476 8616 3482 8628
rect 10318 8616 10324 8628
rect 3476 8588 10324 8616
rect 3476 8576 3482 8588
rect 10318 8576 10324 8588
rect 10376 8576 10382 8628
rect 10502 8576 10508 8628
rect 10560 8616 10566 8628
rect 10597 8619 10655 8625
rect 10597 8616 10609 8619
rect 10560 8588 10609 8616
rect 10560 8576 10566 8588
rect 10597 8585 10609 8588
rect 10643 8585 10655 8619
rect 10870 8616 10876 8628
rect 10831 8588 10876 8616
rect 10597 8579 10655 8585
rect 10870 8576 10876 8588
rect 10928 8576 10934 8628
rect 11882 8616 11888 8628
rect 11843 8588 11888 8616
rect 11882 8576 11888 8588
rect 11940 8576 11946 8628
rect 15197 8619 15255 8625
rect 15197 8585 15209 8619
rect 15243 8616 15255 8619
rect 16206 8616 16212 8628
rect 15243 8588 16212 8616
rect 15243 8585 15255 8588
rect 15197 8579 15255 8585
rect 16206 8576 16212 8588
rect 16264 8576 16270 8628
rect 17218 8616 17224 8628
rect 16684 8588 17224 8616
rect 11606 8508 11612 8560
rect 11664 8548 11670 8560
rect 12437 8551 12495 8557
rect 12437 8548 12449 8551
rect 11664 8520 12449 8548
rect 11664 8508 11670 8520
rect 12437 8517 12449 8520
rect 12483 8517 12495 8551
rect 12437 8511 12495 8517
rect 12894 8508 12900 8560
rect 12952 8548 12958 8560
rect 16684 8548 16712 8588
rect 17218 8576 17224 8588
rect 17276 8616 17282 8628
rect 18598 8616 18604 8628
rect 17276 8588 18604 8616
rect 17276 8576 17282 8588
rect 18598 8576 18604 8588
rect 18656 8576 18662 8628
rect 18693 8619 18751 8625
rect 18693 8585 18705 8619
rect 18739 8616 18751 8619
rect 19610 8616 19616 8628
rect 18739 8588 19616 8616
rect 18739 8585 18751 8588
rect 18693 8579 18751 8585
rect 19610 8576 19616 8588
rect 19668 8576 19674 8628
rect 19978 8576 19984 8628
rect 20036 8616 20042 8628
rect 20036 8588 20208 8616
rect 20036 8576 20042 8588
rect 12952 8520 16712 8548
rect 16761 8551 16819 8557
rect 12952 8508 12958 8520
rect 16761 8517 16773 8551
rect 16807 8548 16819 8551
rect 17034 8548 17040 8560
rect 16807 8520 17040 8548
rect 16807 8517 16819 8520
rect 16761 8511 16819 8517
rect 17034 8508 17040 8520
rect 17092 8508 17098 8560
rect 18322 8508 18328 8560
rect 18380 8548 18386 8560
rect 19521 8551 19579 8557
rect 18380 8520 19380 8548
rect 18380 8508 18386 8520
rect 10962 8440 10968 8492
rect 11020 8480 11026 8492
rect 11425 8483 11483 8489
rect 11425 8480 11437 8483
rect 11020 8452 11437 8480
rect 11020 8440 11026 8452
rect 11425 8449 11437 8452
rect 11471 8449 11483 8483
rect 11425 8443 11483 8449
rect 12526 8440 12532 8492
rect 12584 8480 12590 8492
rect 12989 8483 13047 8489
rect 12989 8480 13001 8483
rect 12584 8452 13001 8480
rect 12584 8440 12590 8452
rect 12989 8449 13001 8452
rect 13035 8449 13047 8483
rect 14366 8480 14372 8492
rect 14327 8452 14372 8480
rect 12989 8443 13047 8449
rect 14366 8440 14372 8452
rect 14424 8440 14430 8492
rect 15838 8440 15844 8492
rect 15896 8480 15902 8492
rect 16298 8480 16304 8492
rect 15896 8452 16304 8480
rect 15896 8440 15902 8452
rect 16298 8440 16304 8452
rect 16356 8440 16362 8492
rect 16393 8483 16451 8489
rect 16393 8449 16405 8483
rect 16439 8480 16451 8483
rect 16574 8480 16580 8492
rect 16439 8452 16580 8480
rect 16439 8449 16451 8452
rect 16393 8443 16451 8449
rect 16574 8440 16580 8452
rect 16632 8440 16638 8492
rect 17402 8480 17408 8492
rect 17363 8452 17408 8480
rect 17402 8440 17408 8452
rect 17460 8440 17466 8492
rect 19352 8489 19380 8520
rect 19521 8517 19533 8551
rect 19567 8548 19579 8551
rect 19705 8551 19763 8557
rect 19705 8548 19717 8551
rect 19567 8520 19717 8548
rect 19567 8517 19579 8520
rect 19521 8511 19579 8517
rect 19705 8517 19717 8520
rect 19751 8517 19763 8551
rect 19705 8511 19763 8517
rect 19337 8483 19395 8489
rect 19337 8449 19349 8483
rect 19383 8480 19395 8483
rect 19978 8480 19984 8492
rect 19383 8452 19984 8480
rect 19383 8449 19395 8452
rect 19337 8443 19395 8449
rect 19978 8440 19984 8452
rect 20036 8440 20042 8492
rect 20180 8489 20208 8588
rect 20165 8483 20223 8489
rect 20165 8449 20177 8483
rect 20211 8449 20223 8483
rect 20165 8443 20223 8449
rect 20349 8483 20407 8489
rect 20349 8449 20361 8483
rect 20395 8480 20407 8483
rect 20622 8480 20628 8492
rect 20395 8452 20628 8480
rect 20395 8449 20407 8452
rect 20349 8443 20407 8449
rect 20622 8440 20628 8452
rect 20680 8440 20686 8492
rect 9217 8415 9275 8421
rect 9217 8381 9229 8415
rect 9263 8412 9275 8415
rect 9858 8412 9864 8424
rect 9263 8384 9864 8412
rect 9263 8381 9275 8384
rect 9217 8375 9275 8381
rect 9858 8372 9864 8384
rect 9916 8372 9922 8424
rect 11241 8415 11299 8421
rect 11241 8381 11253 8415
rect 11287 8412 11299 8415
rect 11698 8412 11704 8424
rect 11287 8384 11704 8412
rect 11287 8381 11299 8384
rect 11241 8375 11299 8381
rect 11698 8372 11704 8384
rect 11756 8372 11762 8424
rect 12069 8415 12127 8421
rect 12069 8381 12081 8415
rect 12115 8412 12127 8415
rect 13998 8412 14004 8424
rect 12115 8384 14004 8412
rect 12115 8381 12127 8384
rect 12069 8375 12127 8381
rect 13998 8372 14004 8384
rect 14056 8412 14062 8424
rect 15381 8415 15439 8421
rect 15381 8412 15393 8415
rect 14056 8384 15393 8412
rect 14056 8372 14062 8384
rect 15381 8381 15393 8384
rect 15427 8381 15439 8415
rect 15381 8375 15439 8381
rect 16482 8372 16488 8424
rect 16540 8412 16546 8424
rect 16540 8384 16712 8412
rect 16540 8372 16546 8384
rect 9484 8347 9542 8353
rect 9484 8313 9496 8347
rect 9530 8344 9542 8347
rect 9766 8344 9772 8356
rect 9530 8316 9772 8344
rect 9530 8313 9542 8316
rect 9484 8307 9542 8313
rect 9766 8304 9772 8316
rect 9824 8304 9830 8356
rect 10686 8304 10692 8356
rect 10744 8344 10750 8356
rect 11333 8347 11391 8353
rect 11333 8344 11345 8347
rect 10744 8316 11345 8344
rect 10744 8304 10750 8316
rect 11333 8313 11345 8316
rect 11379 8344 11391 8347
rect 11974 8344 11980 8356
rect 11379 8316 11980 8344
rect 11379 8313 11391 8316
rect 11333 8307 11391 8313
rect 11974 8304 11980 8316
rect 12032 8304 12038 8356
rect 12802 8344 12808 8356
rect 12763 8316 12808 8344
rect 12802 8304 12808 8316
rect 12860 8304 12866 8356
rect 13722 8304 13728 8356
rect 13780 8344 13786 8356
rect 14274 8344 14280 8356
rect 13780 8316 14280 8344
rect 13780 8304 13786 8316
rect 14274 8304 14280 8316
rect 14332 8304 14338 8356
rect 16114 8344 16120 8356
rect 15488 8316 15976 8344
rect 16075 8316 16120 8344
rect 12894 8276 12900 8288
rect 12855 8248 12900 8276
rect 12894 8236 12900 8248
rect 12952 8236 12958 8288
rect 13814 8276 13820 8288
rect 13775 8248 13820 8276
rect 13814 8236 13820 8248
rect 13872 8236 13878 8288
rect 14185 8279 14243 8285
rect 14185 8245 14197 8279
rect 14231 8276 14243 8279
rect 15488 8276 15516 8316
rect 14231 8248 15516 8276
rect 14231 8245 14243 8248
rect 14185 8239 14243 8245
rect 15562 8236 15568 8288
rect 15620 8276 15626 8288
rect 15749 8279 15807 8285
rect 15749 8276 15761 8279
rect 15620 8248 15761 8276
rect 15620 8236 15626 8248
rect 15749 8245 15761 8248
rect 15795 8245 15807 8279
rect 15948 8276 15976 8316
rect 16114 8304 16120 8316
rect 16172 8304 16178 8356
rect 16209 8347 16267 8353
rect 16209 8313 16221 8347
rect 16255 8344 16267 8347
rect 16574 8344 16580 8356
rect 16255 8316 16580 8344
rect 16255 8313 16267 8316
rect 16209 8307 16267 8313
rect 16574 8304 16580 8316
rect 16632 8304 16638 8356
rect 16684 8344 16712 8384
rect 16758 8372 16764 8424
rect 16816 8412 16822 8424
rect 17221 8415 17279 8421
rect 17221 8412 17233 8415
rect 16816 8384 17233 8412
rect 16816 8372 16822 8384
rect 17221 8381 17233 8384
rect 17267 8381 17279 8415
rect 17221 8375 17279 8381
rect 19153 8415 19211 8421
rect 19153 8381 19165 8415
rect 19199 8381 19211 8415
rect 19521 8415 19579 8421
rect 19521 8412 19533 8415
rect 19153 8375 19211 8381
rect 19251 8384 19533 8412
rect 17129 8347 17187 8353
rect 17129 8344 17141 8347
rect 16684 8316 17141 8344
rect 17129 8313 17141 8316
rect 17175 8313 17187 8347
rect 17129 8307 17187 8313
rect 18598 8304 18604 8356
rect 18656 8344 18662 8356
rect 19061 8347 19119 8353
rect 19061 8344 19073 8347
rect 18656 8316 19073 8344
rect 18656 8304 18662 8316
rect 19061 8313 19073 8316
rect 19107 8313 19119 8347
rect 19168 8344 19196 8375
rect 19251 8344 19279 8384
rect 19521 8381 19533 8384
rect 19567 8381 19579 8415
rect 19521 8375 19579 8381
rect 20070 8372 20076 8424
rect 20128 8372 20134 8424
rect 19168 8316 19279 8344
rect 19061 8307 19119 8313
rect 20088 8288 20116 8372
rect 17494 8276 17500 8288
rect 15948 8248 17500 8276
rect 15749 8239 15807 8245
rect 17494 8236 17500 8248
rect 17552 8236 17558 8288
rect 20070 8276 20076 8288
rect 19983 8248 20076 8276
rect 20070 8236 20076 8248
rect 20128 8236 20134 8288
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 10045 8075 10103 8081
rect 10045 8041 10057 8075
rect 10091 8072 10103 8075
rect 11790 8072 11796 8084
rect 10091 8044 11796 8072
rect 10091 8041 10103 8044
rect 10045 8035 10103 8041
rect 11790 8032 11796 8044
rect 11848 8032 11854 8084
rect 12437 8075 12495 8081
rect 12437 8041 12449 8075
rect 12483 8072 12495 8075
rect 12526 8072 12532 8084
rect 12483 8044 12532 8072
rect 12483 8041 12495 8044
rect 12437 8035 12495 8041
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 12894 8072 12900 8084
rect 12855 8044 12900 8072
rect 12894 8032 12900 8044
rect 12952 8032 12958 8084
rect 13357 8075 13415 8081
rect 13357 8041 13369 8075
rect 13403 8072 13415 8075
rect 13814 8072 13820 8084
rect 13403 8044 13820 8072
rect 13403 8041 13415 8044
rect 13357 8035 13415 8041
rect 13814 8032 13820 8044
rect 13872 8032 13878 8084
rect 13909 8075 13967 8081
rect 13909 8041 13921 8075
rect 13955 8041 13967 8075
rect 13909 8035 13967 8041
rect 14277 8075 14335 8081
rect 14277 8041 14289 8075
rect 14323 8072 14335 8075
rect 14458 8072 14464 8084
rect 14323 8044 14464 8072
rect 14323 8041 14335 8044
rect 14277 8035 14335 8041
rect 9125 8007 9183 8013
rect 9125 7973 9137 8007
rect 9171 8004 9183 8007
rect 9950 8004 9956 8016
rect 9171 7976 9956 8004
rect 9171 7973 9183 7976
rect 9125 7967 9183 7973
rect 9950 7964 9956 7976
rect 10008 7964 10014 8016
rect 10870 7964 10876 8016
rect 10928 8004 10934 8016
rect 13265 8007 13323 8013
rect 10928 7976 13216 8004
rect 10928 7964 10934 7976
rect 8849 7939 8907 7945
rect 8849 7905 8861 7939
rect 8895 7936 8907 7939
rect 9674 7936 9680 7948
rect 8895 7908 9680 7936
rect 8895 7905 8907 7908
rect 8849 7899 8907 7905
rect 9674 7896 9680 7908
rect 9732 7896 9738 7948
rect 10318 7896 10324 7948
rect 10376 7936 10382 7948
rect 11330 7945 11336 7948
rect 10413 7939 10471 7945
rect 10413 7936 10425 7939
rect 10376 7908 10425 7936
rect 10376 7896 10382 7908
rect 10413 7905 10425 7908
rect 10459 7905 10471 7939
rect 10413 7899 10471 7905
rect 11313 7939 11336 7945
rect 11313 7905 11325 7939
rect 11313 7899 11336 7905
rect 11330 7896 11336 7899
rect 11388 7896 11394 7948
rect 13188 7936 13216 7976
rect 13265 7973 13277 8007
rect 13311 8004 13323 8007
rect 13924 8004 13952 8035
rect 14458 8032 14464 8044
rect 14516 8032 14522 8084
rect 15749 8075 15807 8081
rect 15749 8041 15761 8075
rect 15795 8072 15807 8075
rect 16114 8072 16120 8084
rect 15795 8044 16120 8072
rect 15795 8041 15807 8044
rect 15749 8035 15807 8041
rect 16114 8032 16120 8044
rect 16172 8032 16178 8084
rect 16209 8075 16267 8081
rect 16209 8041 16221 8075
rect 16255 8072 16267 8075
rect 17034 8072 17040 8084
rect 16255 8044 17040 8072
rect 16255 8041 16267 8044
rect 16209 8035 16267 8041
rect 17034 8032 17040 8044
rect 17092 8032 17098 8084
rect 18506 8032 18512 8084
rect 18564 8072 18570 8084
rect 18782 8072 18788 8084
rect 18564 8044 18788 8072
rect 18564 8032 18570 8044
rect 18782 8032 18788 8044
rect 18840 8032 18846 8084
rect 19978 8032 19984 8084
rect 20036 8072 20042 8084
rect 20349 8075 20407 8081
rect 20349 8072 20361 8075
rect 20036 8044 20361 8072
rect 20036 8032 20042 8044
rect 20349 8041 20361 8044
rect 20395 8041 20407 8075
rect 20898 8072 20904 8084
rect 20859 8044 20904 8072
rect 20349 8035 20407 8041
rect 20898 8032 20904 8044
rect 20956 8032 20962 8084
rect 13311 7976 13952 8004
rect 13311 7973 13323 7976
rect 13265 7967 13323 7973
rect 13998 7964 14004 8016
rect 14056 8004 14062 8016
rect 17954 8004 17960 8016
rect 14056 7976 17960 8004
rect 14056 7964 14062 7976
rect 17954 7964 17960 7976
rect 18012 7964 18018 8016
rect 19236 8007 19294 8013
rect 19236 7973 19248 8007
rect 19282 8004 19294 8007
rect 20622 8004 20628 8016
rect 19282 7976 20628 8004
rect 19282 7973 19294 7976
rect 19236 7967 19294 7973
rect 20622 7964 20628 7976
rect 20680 7964 20686 8016
rect 13906 7936 13912 7948
rect 13188 7908 13912 7936
rect 13906 7896 13912 7908
rect 13964 7896 13970 7948
rect 14369 7939 14427 7945
rect 14369 7905 14381 7939
rect 14415 7936 14427 7939
rect 15102 7936 15108 7948
rect 14415 7908 15108 7936
rect 14415 7905 14427 7908
rect 14369 7899 14427 7905
rect 15102 7896 15108 7908
rect 15160 7936 15166 7948
rect 15286 7936 15292 7948
rect 15160 7908 15292 7936
rect 15160 7896 15166 7908
rect 15286 7896 15292 7908
rect 15344 7896 15350 7948
rect 16117 7939 16175 7945
rect 16117 7905 16129 7939
rect 16163 7936 16175 7939
rect 16574 7936 16580 7948
rect 16163 7908 16580 7936
rect 16163 7905 16175 7908
rect 16117 7899 16175 7905
rect 16574 7896 16580 7908
rect 16632 7896 16638 7948
rect 16761 7939 16819 7945
rect 16761 7905 16773 7939
rect 16807 7936 16819 7939
rect 16850 7936 16856 7948
rect 16807 7908 16856 7936
rect 16807 7905 16819 7908
rect 16761 7899 16819 7905
rect 16850 7896 16856 7908
rect 16908 7896 16914 7948
rect 17028 7939 17086 7945
rect 17028 7905 17040 7939
rect 17074 7936 17086 7939
rect 17402 7936 17408 7948
rect 17074 7908 17408 7936
rect 17074 7905 17086 7908
rect 17028 7899 17086 7905
rect 17402 7896 17408 7908
rect 17460 7936 17466 7948
rect 18598 7936 18604 7948
rect 17460 7908 18604 7936
rect 17460 7896 17466 7908
rect 18598 7896 18604 7908
rect 18656 7896 18662 7948
rect 18969 7939 19027 7945
rect 18969 7905 18981 7939
rect 19015 7936 19027 7939
rect 19058 7936 19064 7948
rect 19015 7908 19064 7936
rect 19015 7905 19027 7908
rect 18969 7899 19027 7905
rect 19058 7896 19064 7908
rect 19116 7896 19122 7948
rect 10502 7868 10508 7880
rect 10463 7840 10508 7868
rect 10502 7828 10508 7840
rect 10560 7828 10566 7880
rect 10689 7871 10747 7877
rect 10689 7837 10701 7871
rect 10735 7868 10747 7871
rect 10962 7868 10968 7880
rect 10735 7840 10968 7868
rect 10735 7837 10747 7840
rect 10689 7831 10747 7837
rect 10962 7828 10968 7840
rect 11020 7828 11026 7880
rect 11057 7871 11115 7877
rect 11057 7837 11069 7871
rect 11103 7837 11115 7871
rect 11057 7831 11115 7837
rect 11072 7732 11100 7831
rect 13446 7828 13452 7880
rect 13504 7868 13510 7880
rect 13504 7840 13549 7868
rect 13504 7828 13510 7840
rect 14458 7828 14464 7880
rect 14516 7868 14522 7880
rect 16393 7871 16451 7877
rect 14516 7840 14561 7868
rect 14516 7828 14522 7840
rect 16393 7837 16405 7871
rect 16439 7868 16451 7871
rect 16439 7840 16712 7868
rect 16439 7837 16451 7840
rect 16393 7831 16451 7837
rect 12066 7760 12072 7812
rect 12124 7800 12130 7812
rect 16482 7800 16488 7812
rect 12124 7772 16488 7800
rect 12124 7760 12130 7772
rect 16482 7760 16488 7772
rect 16540 7760 16546 7812
rect 11790 7732 11796 7744
rect 11072 7704 11796 7732
rect 11790 7692 11796 7704
rect 11848 7692 11854 7744
rect 13446 7692 13452 7744
rect 13504 7732 13510 7744
rect 13998 7732 14004 7744
rect 13504 7704 14004 7732
rect 13504 7692 13510 7704
rect 13998 7692 14004 7704
rect 14056 7692 14062 7744
rect 16574 7692 16580 7744
rect 16632 7732 16638 7744
rect 16684 7732 16712 7840
rect 17494 7732 17500 7744
rect 16632 7704 17500 7732
rect 16632 7692 16638 7704
rect 17494 7692 17500 7704
rect 17552 7732 17558 7744
rect 18141 7735 18199 7741
rect 18141 7732 18153 7735
rect 17552 7704 18153 7732
rect 17552 7692 17558 7704
rect 18141 7701 18153 7704
rect 18187 7701 18199 7735
rect 18141 7695 18199 7701
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 9766 7528 9772 7540
rect 9727 7500 9772 7528
rect 9766 7488 9772 7500
rect 9824 7488 9830 7540
rect 10318 7528 10324 7540
rect 10279 7500 10324 7528
rect 10318 7488 10324 7500
rect 10376 7488 10382 7540
rect 10502 7488 10508 7540
rect 10560 7528 10566 7540
rect 11333 7531 11391 7537
rect 11333 7528 11345 7531
rect 10560 7500 11345 7528
rect 10560 7488 10566 7500
rect 11333 7497 11345 7500
rect 11379 7497 11391 7531
rect 12802 7528 12808 7540
rect 12763 7500 12808 7528
rect 11333 7491 11391 7497
rect 12802 7488 12808 7500
rect 12860 7488 12866 7540
rect 15197 7531 15255 7537
rect 15197 7528 15209 7531
rect 13372 7500 15209 7528
rect 10594 7352 10600 7404
rect 10652 7392 10658 7404
rect 10873 7395 10931 7401
rect 10873 7392 10885 7395
rect 10652 7364 10885 7392
rect 10652 7352 10658 7364
rect 10873 7361 10885 7364
rect 10919 7392 10931 7395
rect 11885 7395 11943 7401
rect 11885 7392 11897 7395
rect 10919 7364 11897 7392
rect 10919 7361 10931 7364
rect 10873 7355 10931 7361
rect 11885 7361 11897 7364
rect 11931 7361 11943 7395
rect 11885 7355 11943 7361
rect 13170 7352 13176 7404
rect 13228 7392 13234 7404
rect 13372 7401 13400 7500
rect 15197 7497 15209 7500
rect 15243 7497 15255 7531
rect 15197 7491 15255 7497
rect 16482 7488 16488 7540
rect 16540 7488 16546 7540
rect 16942 7528 16948 7540
rect 16903 7500 16948 7528
rect 16942 7488 16948 7500
rect 17000 7488 17006 7540
rect 16500 7460 16528 7488
rect 17402 7460 17408 7472
rect 16500 7432 17408 7460
rect 17402 7420 17408 7432
rect 17460 7460 17466 7472
rect 18230 7460 18236 7472
rect 17460 7432 18236 7460
rect 17460 7420 17466 7432
rect 18230 7420 18236 7432
rect 18288 7420 18294 7472
rect 13357 7395 13415 7401
rect 13357 7392 13369 7395
rect 13228 7364 13369 7392
rect 13228 7352 13234 7364
rect 13357 7361 13369 7364
rect 13403 7361 13415 7395
rect 13357 7355 13415 7361
rect 16666 7352 16672 7404
rect 16724 7392 16730 7404
rect 17221 7395 17279 7401
rect 17221 7392 17233 7395
rect 16724 7364 17233 7392
rect 16724 7352 16730 7364
rect 17221 7361 17233 7364
rect 17267 7361 17279 7395
rect 18598 7392 18604 7404
rect 18559 7364 18604 7392
rect 17221 7355 17279 7361
rect 18598 7352 18604 7364
rect 18656 7352 18662 7404
rect 20438 7392 20444 7404
rect 20399 7364 20444 7392
rect 20438 7352 20444 7364
rect 20496 7352 20502 7404
rect 8386 7324 8392 7336
rect 8347 7296 8392 7324
rect 8386 7284 8392 7296
rect 8444 7284 8450 7336
rect 10781 7327 10839 7333
rect 10781 7293 10793 7327
rect 10827 7324 10839 7327
rect 13722 7324 13728 7336
rect 10827 7296 13728 7324
rect 10827 7293 10839 7296
rect 10781 7287 10839 7293
rect 13722 7284 13728 7296
rect 13780 7284 13786 7336
rect 13817 7327 13875 7333
rect 13817 7293 13829 7327
rect 13863 7324 13875 7327
rect 14084 7327 14142 7333
rect 13863 7296 14044 7324
rect 13863 7293 13875 7296
rect 13817 7287 13875 7293
rect 8656 7259 8714 7265
rect 8656 7225 8668 7259
rect 8702 7256 8714 7259
rect 9858 7256 9864 7268
rect 8702 7228 9864 7256
rect 8702 7225 8714 7228
rect 8656 7219 8714 7225
rect 9858 7216 9864 7228
rect 9916 7216 9922 7268
rect 11701 7259 11759 7265
rect 11701 7225 11713 7259
rect 11747 7256 11759 7259
rect 13446 7256 13452 7268
rect 11747 7228 13452 7256
rect 11747 7225 11759 7228
rect 11701 7219 11759 7225
rect 13446 7216 13452 7228
rect 13504 7216 13510 7268
rect 9950 7148 9956 7200
rect 10008 7188 10014 7200
rect 10689 7191 10747 7197
rect 10689 7188 10701 7191
rect 10008 7160 10701 7188
rect 10008 7148 10014 7160
rect 10689 7157 10701 7160
rect 10735 7188 10747 7191
rect 10870 7188 10876 7200
rect 10735 7160 10876 7188
rect 10735 7157 10747 7160
rect 10689 7151 10747 7157
rect 10870 7148 10876 7160
rect 10928 7148 10934 7200
rect 11793 7191 11851 7197
rect 11793 7157 11805 7191
rect 11839 7188 11851 7191
rect 12894 7188 12900 7200
rect 11839 7160 12900 7188
rect 11839 7157 11851 7160
rect 11793 7151 11851 7157
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 13170 7188 13176 7200
rect 13131 7160 13176 7188
rect 13170 7148 13176 7160
rect 13228 7148 13234 7200
rect 13265 7191 13323 7197
rect 13265 7157 13277 7191
rect 13311 7188 13323 7191
rect 13906 7188 13912 7200
rect 13311 7160 13912 7188
rect 13311 7157 13323 7160
rect 13265 7151 13323 7157
rect 13906 7148 13912 7160
rect 13964 7148 13970 7200
rect 14016 7188 14044 7296
rect 14084 7293 14096 7327
rect 14130 7324 14142 7327
rect 14458 7324 14464 7336
rect 14130 7296 14464 7324
rect 14130 7293 14142 7296
rect 14084 7287 14142 7293
rect 14458 7284 14464 7296
rect 14516 7284 14522 7336
rect 15565 7327 15623 7333
rect 15565 7324 15577 7327
rect 15488 7296 15577 7324
rect 15378 7188 15384 7200
rect 14016 7160 15384 7188
rect 15378 7148 15384 7160
rect 15436 7188 15442 7200
rect 15488 7188 15516 7296
rect 15565 7293 15577 7296
rect 15611 7293 15623 7327
rect 15565 7287 15623 7293
rect 15832 7327 15890 7333
rect 15832 7293 15844 7327
rect 15878 7324 15890 7327
rect 16574 7324 16580 7336
rect 15878 7296 16580 7324
rect 15878 7293 15890 7296
rect 15832 7287 15890 7293
rect 16574 7284 16580 7296
rect 16632 7284 16638 7336
rect 18417 7327 18475 7333
rect 18417 7293 18429 7327
rect 18463 7324 18475 7327
rect 18966 7324 18972 7336
rect 18463 7296 18972 7324
rect 18463 7293 18475 7296
rect 18417 7287 18475 7293
rect 18966 7284 18972 7296
rect 19024 7284 19030 7336
rect 19886 7284 19892 7336
rect 19944 7324 19950 7336
rect 20349 7327 20407 7333
rect 20349 7324 20361 7327
rect 19944 7296 20361 7324
rect 19944 7284 19950 7296
rect 20349 7293 20361 7296
rect 20395 7293 20407 7327
rect 20349 7287 20407 7293
rect 15654 7216 15660 7268
rect 15712 7256 15718 7268
rect 18782 7256 18788 7268
rect 15712 7228 18788 7256
rect 15712 7216 15718 7228
rect 18782 7216 18788 7228
rect 18840 7216 18846 7268
rect 20257 7259 20315 7265
rect 20257 7225 20269 7259
rect 20303 7256 20315 7259
rect 20898 7256 20904 7268
rect 20303 7228 20904 7256
rect 20303 7225 20315 7228
rect 20257 7219 20315 7225
rect 20898 7216 20904 7228
rect 20956 7216 20962 7268
rect 16298 7188 16304 7200
rect 15436 7160 16304 7188
rect 15436 7148 15442 7160
rect 16298 7148 16304 7160
rect 16356 7148 16362 7200
rect 18046 7188 18052 7200
rect 18007 7160 18052 7188
rect 18046 7148 18052 7160
rect 18104 7148 18110 7200
rect 18506 7188 18512 7200
rect 18467 7160 18512 7188
rect 18506 7148 18512 7160
rect 18564 7148 18570 7200
rect 19150 7148 19156 7200
rect 19208 7188 19214 7200
rect 19889 7191 19947 7197
rect 19889 7188 19901 7191
rect 19208 7160 19901 7188
rect 19208 7148 19214 7160
rect 19889 7157 19901 7160
rect 19935 7157 19947 7191
rect 19889 7151 19947 7157
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 9674 6984 9680 6996
rect 9635 6956 9680 6984
rect 9674 6944 9680 6956
rect 9732 6944 9738 6996
rect 13170 6944 13176 6996
rect 13228 6984 13234 6996
rect 13449 6987 13507 6993
rect 13449 6984 13461 6987
rect 13228 6956 13461 6984
rect 13228 6944 13234 6956
rect 13449 6953 13461 6956
rect 13495 6953 13507 6987
rect 13906 6984 13912 6996
rect 13867 6956 13912 6984
rect 13449 6947 13507 6953
rect 13906 6944 13912 6956
rect 13964 6944 13970 6996
rect 15654 6984 15660 6996
rect 14200 6956 15240 6984
rect 15615 6956 15660 6984
rect 9766 6876 9772 6928
rect 9824 6916 9830 6928
rect 11057 6919 11115 6925
rect 9824 6888 10272 6916
rect 9824 6876 9830 6888
rect 10042 6848 10048 6860
rect 10003 6820 10048 6848
rect 10042 6808 10048 6820
rect 10100 6808 10106 6860
rect 9122 6780 9128 6792
rect 9083 6752 9128 6780
rect 9122 6740 9128 6752
rect 9180 6740 9186 6792
rect 9766 6740 9772 6792
rect 9824 6780 9830 6792
rect 10244 6789 10272 6888
rect 11057 6885 11069 6919
rect 11103 6916 11115 6919
rect 14200 6916 14228 6956
rect 11103 6888 14228 6916
rect 14277 6919 14335 6925
rect 11103 6885 11115 6888
rect 11057 6879 11115 6885
rect 14277 6885 14289 6919
rect 14323 6916 14335 6919
rect 14366 6916 14372 6928
rect 14323 6888 14372 6916
rect 14323 6885 14335 6888
rect 14277 6879 14335 6885
rect 14366 6876 14372 6888
rect 14424 6876 14430 6928
rect 15212 6916 15240 6956
rect 15654 6944 15660 6956
rect 15712 6944 15718 6996
rect 15930 6944 15936 6996
rect 15988 6984 15994 6996
rect 16114 6984 16120 6996
rect 15988 6956 16120 6984
rect 15988 6944 15994 6956
rect 16114 6944 16120 6956
rect 16172 6944 16178 6996
rect 16298 6984 16304 6996
rect 16259 6956 16304 6984
rect 16298 6944 16304 6956
rect 16356 6944 16362 6996
rect 17313 6987 17371 6993
rect 17313 6953 17325 6987
rect 17359 6984 17371 6987
rect 17865 6987 17923 6993
rect 17865 6984 17877 6987
rect 17359 6956 17877 6984
rect 17359 6953 17371 6956
rect 17313 6947 17371 6953
rect 17865 6953 17877 6956
rect 17911 6953 17923 6987
rect 18230 6984 18236 6996
rect 18191 6956 18236 6984
rect 17865 6947 17923 6953
rect 18230 6944 18236 6956
rect 18288 6944 18294 6996
rect 20533 6987 20591 6993
rect 20533 6953 20545 6987
rect 20579 6984 20591 6987
rect 20622 6984 20628 6996
rect 20579 6956 20628 6984
rect 20579 6953 20591 6956
rect 20533 6947 20591 6953
rect 20622 6944 20628 6956
rect 20680 6944 20686 6996
rect 17221 6919 17279 6925
rect 15212 6888 17172 6916
rect 10962 6808 10968 6860
rect 11020 6848 11026 6860
rect 12060 6851 12118 6857
rect 11020 6820 11284 6848
rect 11020 6808 11026 6820
rect 11256 6789 11284 6820
rect 12060 6817 12072 6851
rect 12106 6848 12118 6851
rect 12526 6848 12532 6860
rect 12106 6820 12532 6848
rect 12106 6817 12118 6820
rect 12060 6811 12118 6817
rect 12526 6808 12532 6820
rect 12584 6808 12590 6860
rect 13722 6808 13728 6860
rect 13780 6848 13786 6860
rect 14826 6848 14832 6860
rect 13780 6820 14832 6848
rect 13780 6808 13786 6820
rect 14826 6808 14832 6820
rect 14884 6808 14890 6860
rect 15749 6851 15807 6857
rect 15749 6817 15761 6851
rect 15795 6848 15807 6851
rect 15930 6848 15936 6860
rect 15795 6820 15936 6848
rect 15795 6817 15807 6820
rect 15749 6811 15807 6817
rect 15930 6808 15936 6820
rect 15988 6808 15994 6860
rect 16206 6808 16212 6860
rect 16264 6848 16270 6860
rect 16485 6851 16543 6857
rect 16485 6848 16497 6851
rect 16264 6820 16497 6848
rect 16264 6808 16270 6820
rect 16485 6817 16497 6820
rect 16531 6817 16543 6851
rect 17144 6848 17172 6888
rect 17221 6885 17233 6919
rect 17267 6916 17279 6919
rect 18046 6916 18052 6928
rect 17267 6888 18052 6916
rect 17267 6885 17279 6888
rect 17221 6879 17279 6885
rect 18046 6876 18052 6888
rect 18104 6876 18110 6928
rect 17586 6848 17592 6860
rect 17144 6820 17592 6848
rect 16485 6811 16543 6817
rect 17586 6808 17592 6820
rect 17644 6808 17650 6860
rect 19426 6857 19432 6860
rect 19420 6848 19432 6857
rect 19387 6820 19432 6848
rect 19420 6811 19432 6820
rect 19426 6808 19432 6811
rect 19484 6808 19490 6860
rect 10137 6783 10195 6789
rect 10137 6780 10149 6783
rect 9824 6752 10149 6780
rect 9824 6740 9830 6752
rect 10137 6749 10149 6752
rect 10183 6749 10195 6783
rect 10137 6743 10195 6749
rect 10229 6783 10287 6789
rect 10229 6749 10241 6783
rect 10275 6749 10287 6783
rect 10229 6743 10287 6749
rect 11149 6783 11207 6789
rect 11149 6749 11161 6783
rect 11195 6749 11207 6783
rect 11149 6743 11207 6749
rect 11241 6783 11299 6789
rect 11241 6749 11253 6783
rect 11287 6749 11299 6783
rect 11790 6780 11796 6792
rect 11751 6752 11796 6780
rect 11241 6743 11299 6749
rect 10502 6604 10508 6656
rect 10560 6644 10566 6656
rect 10689 6647 10747 6653
rect 10689 6644 10701 6647
rect 10560 6616 10701 6644
rect 10560 6604 10566 6616
rect 10689 6613 10701 6616
rect 10735 6613 10747 6647
rect 11164 6644 11192 6743
rect 11790 6740 11796 6752
rect 11848 6740 11854 6792
rect 13814 6740 13820 6792
rect 13872 6780 13878 6792
rect 14369 6783 14427 6789
rect 14369 6780 14381 6783
rect 13872 6752 14381 6780
rect 13872 6740 13878 6752
rect 14369 6749 14381 6752
rect 14415 6749 14427 6783
rect 14369 6743 14427 6749
rect 14458 6740 14464 6792
rect 14516 6780 14522 6792
rect 15838 6780 15844 6792
rect 14516 6752 14561 6780
rect 15799 6752 15844 6780
rect 14516 6740 14522 6752
rect 15838 6740 15844 6752
rect 15896 6740 15902 6792
rect 17494 6780 17500 6792
rect 17455 6752 17500 6780
rect 17494 6740 17500 6752
rect 17552 6740 17558 6792
rect 17770 6740 17776 6792
rect 17828 6780 17834 6792
rect 18325 6783 18383 6789
rect 18325 6780 18337 6783
rect 17828 6752 18337 6780
rect 17828 6740 17834 6752
rect 18325 6749 18337 6752
rect 18371 6749 18383 6783
rect 18325 6743 18383 6749
rect 18509 6783 18567 6789
rect 18509 6749 18521 6783
rect 18555 6780 18567 6783
rect 18598 6780 18604 6792
rect 18555 6752 18604 6780
rect 18555 6749 18567 6752
rect 18509 6743 18567 6749
rect 18598 6740 18604 6752
rect 18656 6740 18662 6792
rect 18966 6740 18972 6792
rect 19024 6780 19030 6792
rect 19153 6783 19211 6789
rect 19153 6780 19165 6783
rect 19024 6752 19165 6780
rect 19024 6740 19030 6752
rect 19153 6749 19165 6752
rect 19199 6749 19211 6783
rect 19153 6743 19211 6749
rect 15654 6712 15660 6724
rect 13004 6684 15660 6712
rect 13004 6644 13032 6684
rect 15654 6672 15660 6684
rect 15712 6672 15718 6724
rect 16758 6672 16764 6724
rect 16816 6712 16822 6724
rect 16853 6715 16911 6721
rect 16853 6712 16865 6715
rect 16816 6684 16865 6712
rect 16816 6672 16822 6684
rect 16853 6681 16865 6684
rect 16899 6681 16911 6715
rect 16853 6675 16911 6681
rect 13170 6644 13176 6656
rect 11164 6616 13032 6644
rect 13131 6616 13176 6644
rect 10689 6607 10747 6613
rect 13170 6604 13176 6616
rect 13228 6604 13234 6656
rect 14550 6604 14556 6656
rect 14608 6644 14614 6656
rect 15289 6647 15347 6653
rect 15289 6644 15301 6647
rect 14608 6616 15301 6644
rect 14608 6604 14614 6616
rect 15289 6613 15301 6616
rect 15335 6613 15347 6647
rect 15289 6607 15347 6613
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 9858 6440 9864 6452
rect 9819 6412 9864 6440
rect 9858 6400 9864 6412
rect 9916 6400 9922 6452
rect 10042 6400 10048 6452
rect 10100 6440 10106 6452
rect 10137 6443 10195 6449
rect 10137 6440 10149 6443
rect 10100 6412 10149 6440
rect 10100 6400 10106 6412
rect 10137 6409 10149 6412
rect 10183 6409 10195 6443
rect 14642 6440 14648 6452
rect 10137 6403 10195 6409
rect 11808 6412 14648 6440
rect 9876 6304 9904 6400
rect 10318 6304 10324 6316
rect 9876 6276 10324 6304
rect 10318 6264 10324 6276
rect 10376 6304 10382 6316
rect 10689 6307 10747 6313
rect 10689 6304 10701 6307
rect 10376 6276 10701 6304
rect 10376 6264 10382 6276
rect 10689 6273 10701 6276
rect 10735 6273 10747 6307
rect 10689 6267 10747 6273
rect 10962 6264 10968 6316
rect 11020 6304 11026 6316
rect 11701 6307 11759 6313
rect 11701 6304 11713 6307
rect 11020 6276 11713 6304
rect 11020 6264 11026 6276
rect 11701 6273 11713 6276
rect 11747 6273 11759 6307
rect 11701 6267 11759 6273
rect 6825 6239 6883 6245
rect 6825 6205 6837 6239
rect 6871 6236 6883 6239
rect 8386 6236 8392 6248
rect 6871 6208 8392 6236
rect 6871 6205 6883 6208
rect 6825 6199 6883 6205
rect 8386 6196 8392 6208
rect 8444 6236 8450 6248
rect 8481 6239 8539 6245
rect 8481 6236 8493 6239
rect 8444 6208 8493 6236
rect 8444 6196 8450 6208
rect 8481 6205 8493 6208
rect 8527 6205 8539 6239
rect 8481 6199 8539 6205
rect 9122 6196 9128 6248
rect 9180 6236 9186 6248
rect 10505 6239 10563 6245
rect 10505 6236 10517 6239
rect 9180 6208 10517 6236
rect 9180 6196 9186 6208
rect 10505 6205 10517 6208
rect 10551 6205 10563 6239
rect 10505 6199 10563 6205
rect 10594 6196 10600 6248
rect 10652 6236 10658 6248
rect 10652 6208 11100 6236
rect 10652 6196 10658 6208
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 7070 6171 7128 6177
rect 7070 6168 7082 6171
rect 4120 6140 7082 6168
rect 4120 6128 4126 6140
rect 7070 6137 7082 6140
rect 7116 6137 7128 6171
rect 8726 6171 8784 6177
rect 8726 6168 8738 6171
rect 7070 6131 7128 6137
rect 8220 6140 8738 6168
rect 8220 6109 8248 6140
rect 8726 6137 8738 6140
rect 8772 6168 8784 6171
rect 10962 6168 10968 6180
rect 8772 6140 10968 6168
rect 8772 6137 8784 6140
rect 8726 6131 8784 6137
rect 10962 6128 10968 6140
rect 11020 6128 11026 6180
rect 11072 6168 11100 6208
rect 11146 6196 11152 6248
rect 11204 6236 11210 6248
rect 11609 6239 11667 6245
rect 11609 6236 11621 6239
rect 11204 6208 11621 6236
rect 11204 6196 11210 6208
rect 11609 6205 11621 6208
rect 11655 6236 11667 6239
rect 11808 6236 11836 6412
rect 14642 6400 14648 6412
rect 14700 6400 14706 6452
rect 14918 6400 14924 6452
rect 14976 6440 14982 6452
rect 17310 6440 17316 6452
rect 14976 6412 17316 6440
rect 14976 6400 14982 6412
rect 17310 6400 17316 6412
rect 17368 6400 17374 6452
rect 18233 6443 18291 6449
rect 18233 6409 18245 6443
rect 18279 6440 18291 6443
rect 18690 6440 18696 6452
rect 18279 6412 18696 6440
rect 18279 6409 18291 6412
rect 18233 6403 18291 6409
rect 18690 6400 18696 6412
rect 18748 6400 18754 6452
rect 19426 6400 19432 6452
rect 19484 6440 19490 6452
rect 20625 6443 20683 6449
rect 20625 6440 20637 6443
rect 19484 6412 20637 6440
rect 19484 6400 19490 6412
rect 20625 6409 20637 6412
rect 20671 6409 20683 6443
rect 20625 6403 20683 6409
rect 13354 6372 13360 6384
rect 11655 6208 11836 6236
rect 11900 6344 13360 6372
rect 11655 6205 11667 6208
rect 11609 6199 11667 6205
rect 11517 6171 11575 6177
rect 11517 6168 11529 6171
rect 11072 6140 11529 6168
rect 11517 6137 11529 6140
rect 11563 6168 11575 6171
rect 11900 6168 11928 6344
rect 13354 6332 13360 6344
rect 13412 6332 13418 6384
rect 13814 6332 13820 6384
rect 13872 6372 13878 6384
rect 14182 6372 14188 6384
rect 13872 6344 14188 6372
rect 13872 6332 13878 6344
rect 14182 6332 14188 6344
rect 14240 6332 14246 6384
rect 14277 6375 14335 6381
rect 14277 6341 14289 6375
rect 14323 6372 14335 6375
rect 18782 6372 18788 6384
rect 14323 6344 18788 6372
rect 14323 6341 14335 6344
rect 14277 6335 14335 6341
rect 18782 6332 18788 6344
rect 18840 6332 18846 6384
rect 13078 6304 13084 6316
rect 13039 6276 13084 6304
rect 13078 6264 13084 6276
rect 13136 6264 13142 6316
rect 13170 6264 13176 6316
rect 13228 6304 13234 6316
rect 14093 6307 14151 6313
rect 14093 6304 14105 6307
rect 13228 6276 14105 6304
rect 13228 6264 13234 6276
rect 14093 6273 14105 6276
rect 14139 6304 14151 6307
rect 15013 6307 15071 6313
rect 15013 6304 15025 6307
rect 14139 6276 15025 6304
rect 14139 6273 14151 6276
rect 14093 6267 14151 6273
rect 15013 6273 15025 6276
rect 15059 6273 15071 6307
rect 15013 6267 15071 6273
rect 16301 6307 16359 6313
rect 16301 6273 16313 6307
rect 16347 6273 16359 6307
rect 16301 6267 16359 6273
rect 12894 6196 12900 6248
rect 12952 6236 12958 6248
rect 13817 6239 13875 6245
rect 12952 6208 13584 6236
rect 12952 6196 12958 6208
rect 11563 6140 11928 6168
rect 12805 6171 12863 6177
rect 11563 6137 11575 6140
rect 11517 6131 11575 6137
rect 12805 6137 12817 6171
rect 12851 6168 12863 6171
rect 13556 6168 13584 6208
rect 13817 6205 13829 6239
rect 13863 6236 13875 6239
rect 13998 6236 14004 6248
rect 13863 6208 14004 6236
rect 13863 6205 13875 6208
rect 13817 6199 13875 6205
rect 13998 6196 14004 6208
rect 14056 6196 14062 6248
rect 14182 6196 14188 6248
rect 14240 6236 14246 6248
rect 16117 6239 16175 6245
rect 16117 6236 16129 6239
rect 14240 6208 16129 6236
rect 14240 6196 14246 6208
rect 16117 6205 16129 6208
rect 16163 6205 16175 6239
rect 16316 6236 16344 6267
rect 16482 6264 16488 6316
rect 16540 6304 16546 6316
rect 17221 6307 17279 6313
rect 17221 6304 17233 6307
rect 16540 6276 17233 6304
rect 16540 6264 16546 6276
rect 17221 6273 17233 6276
rect 17267 6273 17279 6307
rect 17221 6267 17279 6273
rect 18877 6307 18935 6313
rect 18877 6273 18889 6307
rect 18923 6304 18935 6307
rect 18923 6276 19380 6304
rect 18923 6273 18935 6276
rect 18877 6267 18935 6273
rect 19352 6248 19380 6276
rect 16942 6236 16948 6248
rect 16316 6208 16948 6236
rect 16117 6199 16175 6205
rect 16942 6196 16948 6208
rect 17000 6196 17006 6248
rect 17129 6239 17187 6245
rect 17129 6205 17141 6239
rect 17175 6236 17187 6239
rect 17586 6236 17592 6248
rect 17175 6208 17592 6236
rect 17175 6205 17187 6208
rect 17129 6199 17187 6205
rect 17586 6196 17592 6208
rect 17644 6196 17650 6248
rect 18966 6196 18972 6248
rect 19024 6236 19030 6248
rect 19245 6239 19303 6245
rect 19245 6236 19257 6239
rect 19024 6208 19257 6236
rect 19024 6196 19030 6208
rect 19245 6205 19257 6208
rect 19291 6205 19303 6239
rect 19245 6199 19303 6205
rect 19334 6196 19340 6248
rect 19392 6196 19398 6248
rect 19512 6239 19570 6245
rect 19512 6205 19524 6239
rect 19558 6236 19570 6239
rect 19886 6236 19892 6248
rect 19558 6208 19892 6236
rect 19558 6205 19570 6208
rect 19512 6199 19570 6205
rect 19886 6196 19892 6208
rect 19944 6236 19950 6248
rect 20438 6236 20444 6248
rect 19944 6208 20444 6236
rect 19944 6196 19950 6208
rect 20438 6196 20444 6208
rect 20496 6196 20502 6248
rect 13909 6171 13967 6177
rect 13909 6168 13921 6171
rect 12851 6140 13492 6168
rect 13556 6140 13921 6168
rect 12851 6137 12863 6140
rect 12805 6131 12863 6137
rect 8205 6103 8263 6109
rect 8205 6069 8217 6103
rect 8251 6069 8263 6103
rect 8205 6063 8263 6069
rect 9858 6060 9864 6112
rect 9916 6100 9922 6112
rect 10226 6100 10232 6112
rect 9916 6072 10232 6100
rect 9916 6060 9922 6072
rect 10226 6060 10232 6072
rect 10284 6060 10290 6112
rect 10597 6103 10655 6109
rect 10597 6069 10609 6103
rect 10643 6100 10655 6103
rect 11149 6103 11207 6109
rect 11149 6100 11161 6103
rect 10643 6072 11161 6100
rect 10643 6069 10655 6072
rect 10597 6063 10655 6069
rect 11149 6069 11161 6072
rect 11195 6069 11207 6103
rect 11149 6063 11207 6069
rect 12434 6060 12440 6112
rect 12492 6100 12498 6112
rect 12894 6100 12900 6112
rect 12492 6072 12537 6100
rect 12855 6072 12900 6100
rect 12492 6060 12498 6072
rect 12894 6060 12900 6072
rect 12952 6060 12958 6112
rect 13464 6109 13492 6140
rect 13909 6137 13921 6140
rect 13955 6168 13967 6171
rect 14277 6171 14335 6177
rect 14277 6168 14289 6171
rect 13955 6140 14289 6168
rect 13955 6137 13967 6140
rect 13909 6131 13967 6137
rect 14277 6137 14289 6140
rect 14323 6137 14335 6171
rect 14277 6131 14335 6137
rect 14366 6128 14372 6180
rect 14424 6168 14430 6180
rect 14918 6168 14924 6180
rect 14424 6140 14596 6168
rect 14879 6140 14924 6168
rect 14424 6128 14430 6140
rect 13449 6103 13507 6109
rect 13449 6069 13461 6103
rect 13495 6069 13507 6103
rect 14458 6100 14464 6112
rect 14419 6072 14464 6100
rect 13449 6063 13507 6069
rect 14458 6060 14464 6072
rect 14516 6060 14522 6112
rect 14568 6100 14596 6140
rect 14918 6128 14924 6140
rect 14976 6128 14982 6180
rect 16025 6171 16083 6177
rect 16025 6137 16037 6171
rect 16071 6168 16083 6171
rect 18601 6171 18659 6177
rect 16071 6140 16712 6168
rect 16071 6137 16083 6140
rect 16025 6131 16083 6137
rect 14829 6103 14887 6109
rect 14829 6100 14841 6103
rect 14568 6072 14841 6100
rect 14829 6069 14841 6072
rect 14875 6069 14887 6103
rect 14829 6063 14887 6069
rect 15657 6103 15715 6109
rect 15657 6069 15669 6103
rect 15703 6100 15715 6103
rect 15746 6100 15752 6112
rect 15703 6072 15752 6100
rect 15703 6069 15715 6072
rect 15657 6063 15715 6069
rect 15746 6060 15752 6072
rect 15804 6060 15810 6112
rect 16684 6109 16712 6140
rect 18601 6137 18613 6171
rect 18647 6168 18659 6171
rect 18647 6140 19288 6168
rect 18647 6137 18659 6140
rect 18601 6131 18659 6137
rect 19260 6112 19288 6140
rect 16669 6103 16727 6109
rect 16669 6069 16681 6103
rect 16715 6069 16727 6103
rect 17034 6100 17040 6112
rect 16995 6072 17040 6100
rect 16669 6063 16727 6069
rect 17034 6060 17040 6072
rect 17092 6060 17098 6112
rect 18690 6100 18696 6112
rect 18651 6072 18696 6100
rect 18690 6060 18696 6072
rect 18748 6060 18754 6112
rect 19242 6060 19248 6112
rect 19300 6060 19306 6112
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 9766 5896 9772 5908
rect 9727 5868 9772 5896
rect 9766 5856 9772 5868
rect 9824 5856 9830 5908
rect 10137 5899 10195 5905
rect 10137 5865 10149 5899
rect 10183 5896 10195 5899
rect 10502 5896 10508 5908
rect 10183 5868 10508 5896
rect 10183 5865 10195 5868
rect 10137 5859 10195 5865
rect 10502 5856 10508 5868
rect 10560 5856 10566 5908
rect 12434 5856 12440 5908
rect 12492 5896 12498 5908
rect 12989 5899 13047 5905
rect 12989 5896 13001 5899
rect 12492 5868 13001 5896
rect 12492 5856 12498 5868
rect 12989 5865 13001 5868
rect 13035 5865 13047 5899
rect 14182 5896 14188 5908
rect 14143 5868 14188 5896
rect 12989 5859 13047 5865
rect 14182 5856 14188 5868
rect 14240 5856 14246 5908
rect 14550 5896 14556 5908
rect 14511 5868 14556 5896
rect 14550 5856 14556 5868
rect 14608 5856 14614 5908
rect 15013 5899 15071 5905
rect 15013 5865 15025 5899
rect 15059 5896 15071 5899
rect 16482 5896 16488 5908
rect 15059 5868 16488 5896
rect 15059 5865 15071 5868
rect 15013 5859 15071 5865
rect 16482 5856 16488 5868
rect 16540 5896 16546 5908
rect 16669 5899 16727 5905
rect 16669 5896 16681 5899
rect 16540 5868 16681 5896
rect 16540 5856 16546 5868
rect 16669 5865 16681 5868
rect 16715 5865 16727 5899
rect 18138 5896 18144 5908
rect 16669 5859 16727 5865
rect 16776 5868 18144 5896
rect 11140 5831 11198 5837
rect 11140 5797 11152 5831
rect 11186 5828 11198 5831
rect 13170 5828 13176 5840
rect 11186 5800 13176 5828
rect 11186 5797 11198 5800
rect 11140 5791 11198 5797
rect 13170 5788 13176 5800
rect 13228 5788 13234 5840
rect 15556 5831 15614 5837
rect 15556 5797 15568 5831
rect 15602 5828 15614 5831
rect 15838 5828 15844 5840
rect 15602 5800 15844 5828
rect 15602 5797 15614 5800
rect 15556 5791 15614 5797
rect 15838 5788 15844 5800
rect 15896 5788 15902 5840
rect 16390 5788 16396 5840
rect 16448 5828 16454 5840
rect 16776 5828 16804 5868
rect 18138 5856 18144 5868
rect 18196 5856 18202 5908
rect 18598 5896 18604 5908
rect 18559 5868 18604 5896
rect 18598 5856 18604 5868
rect 18656 5856 18662 5908
rect 20898 5896 20904 5908
rect 20859 5868 20904 5896
rect 20898 5856 20904 5868
rect 20956 5856 20962 5908
rect 16448 5800 16804 5828
rect 16448 5788 16454 5800
rect 16942 5788 16948 5840
rect 17000 5828 17006 5840
rect 19122 5831 19180 5837
rect 19122 5828 19134 5831
rect 17000 5800 19134 5828
rect 17000 5788 17006 5800
rect 19122 5797 19134 5800
rect 19168 5797 19180 5831
rect 19122 5791 19180 5797
rect 8386 5720 8392 5772
rect 8444 5760 8450 5772
rect 10870 5760 10876 5772
rect 8444 5732 10876 5760
rect 8444 5720 8450 5732
rect 10870 5720 10876 5732
rect 10928 5720 10934 5772
rect 12894 5760 12900 5772
rect 12855 5732 12900 5760
rect 12894 5720 12900 5732
rect 12952 5720 12958 5772
rect 14645 5763 14703 5769
rect 14645 5729 14657 5763
rect 14691 5760 14703 5763
rect 15194 5760 15200 5772
rect 14691 5732 15200 5760
rect 14691 5729 14703 5732
rect 14645 5723 14703 5729
rect 15194 5720 15200 5732
rect 15252 5720 15258 5772
rect 15289 5763 15347 5769
rect 15289 5729 15301 5763
rect 15335 5760 15347 5763
rect 15378 5760 15384 5772
rect 15335 5732 15384 5760
rect 15335 5729 15347 5732
rect 15289 5723 15347 5729
rect 15378 5720 15384 5732
rect 15436 5760 15442 5772
rect 17221 5763 17279 5769
rect 17221 5760 17233 5763
rect 15436 5732 17233 5760
rect 15436 5720 15442 5732
rect 17221 5729 17233 5732
rect 17267 5729 17279 5763
rect 17221 5723 17279 5729
rect 17488 5763 17546 5769
rect 17488 5729 17500 5763
rect 17534 5760 17546 5763
rect 17954 5760 17960 5772
rect 17534 5732 17960 5760
rect 17534 5729 17546 5732
rect 17488 5723 17546 5729
rect 10226 5692 10232 5704
rect 10187 5664 10232 5692
rect 10226 5652 10232 5664
rect 10284 5652 10290 5704
rect 10318 5652 10324 5704
rect 10376 5692 10382 5704
rect 13170 5692 13176 5704
rect 10376 5664 10421 5692
rect 13131 5664 13176 5692
rect 10376 5652 10382 5664
rect 13170 5652 13176 5664
rect 13228 5652 13234 5704
rect 14829 5695 14887 5701
rect 14829 5661 14841 5695
rect 14875 5692 14887 5695
rect 15013 5695 15071 5701
rect 15013 5692 15025 5695
rect 14875 5664 15025 5692
rect 14875 5661 14887 5664
rect 14829 5655 14887 5661
rect 15013 5661 15025 5664
rect 15059 5661 15071 5695
rect 15013 5655 15071 5661
rect 12253 5627 12311 5633
rect 12253 5593 12265 5627
rect 12299 5624 12311 5627
rect 13078 5624 13084 5636
rect 12299 5596 13084 5624
rect 12299 5593 12311 5596
rect 12253 5587 12311 5593
rect 13078 5584 13084 5596
rect 13136 5584 13142 5636
rect 12529 5559 12587 5565
rect 12529 5525 12541 5559
rect 12575 5556 12587 5559
rect 13446 5556 13452 5568
rect 12575 5528 13452 5556
rect 12575 5525 12587 5528
rect 12529 5519 12587 5525
rect 13446 5516 13452 5528
rect 13504 5516 13510 5568
rect 17236 5556 17264 5723
rect 17954 5720 17960 5732
rect 18012 5720 18018 5772
rect 18966 5760 18972 5772
rect 18892 5732 18972 5760
rect 18892 5701 18920 5732
rect 18966 5720 18972 5732
rect 19024 5720 19030 5772
rect 18877 5695 18935 5701
rect 18877 5692 18889 5695
rect 18524 5664 18889 5692
rect 18524 5568 18552 5664
rect 18877 5661 18889 5664
rect 18923 5661 18935 5695
rect 18877 5655 18935 5661
rect 18506 5556 18512 5568
rect 17236 5528 18512 5556
rect 18506 5516 18512 5528
rect 18564 5516 18570 5568
rect 20254 5556 20260 5568
rect 20215 5528 20260 5556
rect 20254 5516 20260 5528
rect 20312 5516 20318 5568
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 10226 5312 10232 5364
rect 10284 5352 10290 5364
rect 10321 5355 10379 5361
rect 10321 5352 10333 5355
rect 10284 5324 10333 5352
rect 10284 5312 10290 5324
rect 10321 5321 10333 5324
rect 10367 5321 10379 5355
rect 10321 5315 10379 5321
rect 10870 5312 10876 5364
rect 10928 5352 10934 5364
rect 11333 5355 11391 5361
rect 11333 5352 11345 5355
rect 10928 5324 11345 5352
rect 10928 5312 10934 5324
rect 11333 5321 11345 5324
rect 11379 5352 11391 5355
rect 11790 5352 11796 5364
rect 11379 5324 11796 5352
rect 11379 5321 11391 5324
rect 11333 5315 11391 5321
rect 11790 5312 11796 5324
rect 11848 5312 11854 5364
rect 12437 5355 12495 5361
rect 12437 5321 12449 5355
rect 12483 5352 12495 5355
rect 12894 5352 12900 5364
rect 12483 5324 12900 5352
rect 12483 5321 12495 5324
rect 12437 5315 12495 5321
rect 12894 5312 12900 5324
rect 12952 5312 12958 5364
rect 15013 5355 15071 5361
rect 15013 5321 15025 5355
rect 15059 5352 15071 5355
rect 15838 5352 15844 5364
rect 15059 5324 15844 5352
rect 15059 5321 15071 5324
rect 15013 5315 15071 5321
rect 15838 5312 15844 5324
rect 15896 5312 15902 5364
rect 16942 5312 16948 5364
rect 17000 5352 17006 5364
rect 17221 5355 17279 5361
rect 17221 5352 17233 5355
rect 17000 5324 17233 5352
rect 17000 5312 17006 5324
rect 17221 5321 17233 5324
rect 17267 5321 17279 5355
rect 17221 5315 17279 5321
rect 17310 5312 17316 5364
rect 17368 5352 17374 5364
rect 19886 5352 19892 5364
rect 17368 5324 19748 5352
rect 19847 5324 19892 5352
rect 17368 5312 17374 5324
rect 19720 5296 19748 5324
rect 19886 5312 19892 5324
rect 19944 5312 19950 5364
rect 19702 5244 19708 5296
rect 19760 5284 19766 5296
rect 20530 5284 20536 5296
rect 19760 5256 20536 5284
rect 19760 5244 19766 5256
rect 20530 5244 20536 5256
rect 20588 5244 20594 5296
rect 10778 5216 10784 5228
rect 10739 5188 10784 5216
rect 10778 5176 10784 5188
rect 10836 5176 10842 5228
rect 10962 5216 10968 5228
rect 10923 5188 10968 5216
rect 10962 5176 10968 5188
rect 11020 5176 11026 5228
rect 11882 5176 11888 5228
rect 11940 5176 11946 5228
rect 13078 5216 13084 5228
rect 13039 5188 13084 5216
rect 13078 5176 13084 5188
rect 13136 5176 13142 5228
rect 15378 5176 15384 5228
rect 15436 5216 15442 5228
rect 15654 5216 15660 5228
rect 15436 5188 15660 5216
rect 15436 5176 15442 5188
rect 15654 5176 15660 5188
rect 15712 5216 15718 5228
rect 15841 5219 15899 5225
rect 15841 5216 15853 5219
rect 15712 5188 15853 5216
rect 15712 5176 15718 5188
rect 15841 5185 15853 5188
rect 15887 5185 15899 5219
rect 18506 5216 18512 5228
rect 18467 5188 18512 5216
rect 15841 5179 15899 5185
rect 18506 5176 18512 5188
rect 18564 5176 18570 5228
rect 20717 5219 20775 5225
rect 20717 5216 20729 5219
rect 20272 5188 20729 5216
rect 10042 5108 10048 5160
rect 10100 5148 10106 5160
rect 10686 5148 10692 5160
rect 10100 5120 10692 5148
rect 10100 5108 10106 5120
rect 10686 5108 10692 5120
rect 10744 5108 10750 5160
rect 11517 5151 11575 5157
rect 11517 5117 11529 5151
rect 11563 5148 11575 5151
rect 11900 5148 11928 5176
rect 11563 5120 11928 5148
rect 13633 5151 13691 5157
rect 11563 5117 11575 5120
rect 11517 5111 11575 5117
rect 13633 5117 13645 5151
rect 13679 5148 13691 5151
rect 15396 5148 15424 5176
rect 20272 5160 20300 5188
rect 20717 5185 20729 5188
rect 20763 5185 20775 5219
rect 20717 5179 20775 5185
rect 13679 5120 15424 5148
rect 16108 5151 16166 5157
rect 13679 5117 13691 5120
rect 13633 5111 13691 5117
rect 16108 5117 16120 5151
rect 16154 5148 16166 5151
rect 16482 5148 16488 5160
rect 16154 5120 16488 5148
rect 16154 5117 16166 5120
rect 16108 5111 16166 5117
rect 16482 5108 16488 5120
rect 16540 5108 16546 5160
rect 18776 5151 18834 5157
rect 18776 5117 18788 5151
rect 18822 5148 18834 5151
rect 20254 5148 20260 5160
rect 18822 5120 20260 5148
rect 18822 5117 18834 5120
rect 18776 5111 18834 5117
rect 20254 5108 20260 5120
rect 20312 5108 20318 5160
rect 11885 5083 11943 5089
rect 11885 5049 11897 5083
rect 11931 5080 11943 5083
rect 12805 5083 12863 5089
rect 12805 5080 12817 5083
rect 11931 5052 12817 5080
rect 11931 5049 11943 5052
rect 11885 5043 11943 5049
rect 12805 5049 12817 5052
rect 12851 5049 12863 5083
rect 12805 5043 12863 5049
rect 13170 5040 13176 5092
rect 13228 5080 13234 5092
rect 13878 5083 13936 5089
rect 13878 5080 13890 5083
rect 13228 5052 13890 5080
rect 13228 5040 13234 5052
rect 13878 5049 13890 5052
rect 13924 5049 13936 5083
rect 13878 5043 13936 5049
rect 19794 5040 19800 5092
rect 19852 5080 19858 5092
rect 20533 5083 20591 5089
rect 20533 5080 20545 5083
rect 19852 5052 20545 5080
rect 19852 5040 19858 5052
rect 20533 5049 20545 5052
rect 20579 5080 20591 5083
rect 20714 5080 20720 5092
rect 20579 5052 20720 5080
rect 20579 5049 20591 5052
rect 20533 5043 20591 5049
rect 20714 5040 20720 5052
rect 20772 5040 20778 5092
rect 10686 5012 10692 5024
rect 10647 4984 10692 5012
rect 10686 4972 10692 4984
rect 10744 4972 10750 5024
rect 12897 5015 12955 5021
rect 12897 4981 12909 5015
rect 12943 5012 12955 5015
rect 14458 5012 14464 5024
rect 12943 4984 14464 5012
rect 12943 4981 12955 4984
rect 12897 4975 12955 4981
rect 14458 4972 14464 4984
rect 14516 4972 14522 5024
rect 15289 5015 15347 5021
rect 15289 4981 15301 5015
rect 15335 5012 15347 5015
rect 15378 5012 15384 5024
rect 15335 4984 15384 5012
rect 15335 4981 15347 4984
rect 15289 4975 15347 4981
rect 15378 4972 15384 4984
rect 15436 4972 15442 5024
rect 18049 5015 18107 5021
rect 18049 4981 18061 5015
rect 18095 5012 18107 5015
rect 18138 5012 18144 5024
rect 18095 4984 18144 5012
rect 18095 4981 18107 4984
rect 18049 4975 18107 4981
rect 18138 4972 18144 4984
rect 18196 4972 18202 5024
rect 20162 5012 20168 5024
rect 20123 4984 20168 5012
rect 20162 4972 20168 4984
rect 20220 4972 20226 5024
rect 20622 5012 20628 5024
rect 20583 4984 20628 5012
rect 20622 4972 20628 4984
rect 20680 4972 20686 5024
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 13170 4768 13176 4820
rect 13228 4808 13234 4820
rect 13449 4811 13507 4817
rect 13449 4808 13461 4811
rect 13228 4780 13461 4808
rect 13228 4768 13234 4780
rect 13449 4777 13461 4780
rect 13495 4777 13507 4811
rect 13449 4771 13507 4777
rect 15194 4768 15200 4820
rect 15252 4808 15258 4820
rect 15289 4811 15347 4817
rect 15289 4808 15301 4811
rect 15252 4780 15301 4808
rect 15252 4768 15258 4780
rect 15289 4777 15301 4780
rect 15335 4777 15347 4811
rect 15289 4771 15347 4777
rect 16301 4811 16359 4817
rect 16301 4777 16313 4811
rect 16347 4808 16359 4811
rect 17034 4808 17040 4820
rect 16347 4780 17040 4808
rect 16347 4777 16359 4780
rect 16301 4771 16359 4777
rect 17034 4768 17040 4780
rect 17092 4768 17098 4820
rect 17773 4811 17831 4817
rect 17773 4777 17785 4811
rect 17819 4808 17831 4811
rect 17862 4808 17868 4820
rect 17819 4780 17868 4808
rect 17819 4777 17831 4780
rect 17773 4771 17831 4777
rect 17862 4768 17868 4780
rect 17920 4768 17926 4820
rect 18138 4808 18144 4820
rect 18099 4780 18144 4808
rect 18138 4768 18144 4780
rect 18196 4768 18202 4820
rect 19150 4808 19156 4820
rect 19111 4780 19156 4808
rect 19150 4768 19156 4780
rect 19208 4768 19214 4820
rect 19242 4768 19248 4820
rect 19300 4808 19306 4820
rect 20165 4811 20223 4817
rect 20165 4808 20177 4811
rect 19300 4780 20177 4808
rect 19300 4768 19306 4780
rect 20165 4777 20177 4780
rect 20211 4777 20223 4811
rect 20165 4771 20223 4777
rect 17954 4700 17960 4752
rect 18012 4700 18018 4752
rect 18690 4700 18696 4752
rect 18748 4740 18754 4752
rect 18748 4712 20300 4740
rect 18748 4700 18754 4712
rect 11790 4632 11796 4684
rect 11848 4672 11854 4684
rect 12069 4675 12127 4681
rect 12069 4672 12081 4675
rect 11848 4644 12081 4672
rect 11848 4632 11854 4644
rect 12069 4641 12081 4644
rect 12115 4641 12127 4675
rect 12069 4635 12127 4641
rect 12336 4675 12394 4681
rect 12336 4641 12348 4675
rect 12382 4672 12394 4675
rect 13078 4672 13084 4684
rect 12382 4644 13084 4672
rect 12382 4641 12394 4644
rect 12336 4635 12394 4641
rect 13078 4632 13084 4644
rect 13136 4632 13142 4684
rect 13722 4672 13728 4684
rect 13683 4644 13728 4672
rect 13722 4632 13728 4644
rect 13780 4632 13786 4684
rect 14274 4632 14280 4684
rect 14332 4672 14338 4684
rect 14553 4675 14611 4681
rect 14553 4672 14565 4675
rect 14332 4644 14565 4672
rect 14332 4632 14338 4644
rect 14553 4641 14565 4644
rect 14599 4641 14611 4675
rect 14553 4635 14611 4641
rect 15657 4675 15715 4681
rect 15657 4641 15669 4675
rect 15703 4672 15715 4675
rect 17310 4672 17316 4684
rect 15703 4644 17316 4672
rect 15703 4641 15715 4644
rect 15657 4635 15715 4641
rect 17310 4632 17316 4644
rect 17368 4632 17374 4684
rect 17972 4672 18000 4700
rect 19245 4675 19303 4681
rect 17972 4644 18368 4672
rect 15286 4564 15292 4616
rect 15344 4604 15350 4616
rect 15749 4607 15807 4613
rect 15749 4604 15761 4607
rect 15344 4576 15761 4604
rect 15344 4564 15350 4576
rect 15749 4573 15761 4576
rect 15795 4573 15807 4607
rect 15749 4567 15807 4573
rect 13909 4471 13967 4477
rect 13909 4437 13921 4471
rect 13955 4468 13967 4471
rect 14182 4468 14188 4480
rect 13955 4440 14188 4468
rect 13955 4437 13967 4440
rect 13909 4431 13967 4437
rect 14182 4428 14188 4440
rect 14240 4428 14246 4480
rect 14737 4471 14795 4477
rect 14737 4437 14749 4471
rect 14783 4468 14795 4471
rect 15286 4468 15292 4480
rect 14783 4440 15292 4468
rect 14783 4437 14795 4440
rect 14737 4431 14795 4437
rect 15286 4428 15292 4440
rect 15344 4428 15350 4480
rect 15764 4468 15792 4567
rect 15838 4564 15844 4616
rect 15896 4604 15902 4616
rect 16942 4604 16948 4616
rect 15896 4576 15941 4604
rect 16903 4576 16948 4604
rect 15896 4564 15902 4576
rect 16942 4564 16948 4576
rect 17000 4564 17006 4616
rect 17954 4564 17960 4616
rect 18012 4604 18018 4616
rect 18340 4613 18368 4644
rect 19245 4641 19257 4675
rect 19291 4672 19303 4675
rect 19702 4672 19708 4684
rect 19291 4644 19708 4672
rect 19291 4641 19303 4644
rect 19245 4635 19303 4641
rect 19702 4632 19708 4644
rect 19760 4632 19766 4684
rect 20272 4616 20300 4712
rect 18233 4607 18291 4613
rect 18233 4604 18245 4607
rect 18012 4576 18245 4604
rect 18012 4564 18018 4576
rect 18233 4573 18245 4576
rect 18279 4573 18291 4607
rect 18233 4567 18291 4573
rect 18325 4607 18383 4613
rect 18325 4573 18337 4607
rect 18371 4604 18383 4607
rect 19150 4604 19156 4616
rect 18371 4576 19156 4604
rect 18371 4573 18383 4576
rect 18325 4567 18383 4573
rect 19150 4564 19156 4576
rect 19208 4564 19214 4616
rect 19426 4604 19432 4616
rect 19387 4576 19432 4604
rect 19426 4564 19432 4576
rect 19484 4564 19490 4616
rect 20254 4604 20260 4616
rect 20215 4576 20260 4604
rect 20254 4564 20260 4576
rect 20312 4564 20318 4616
rect 20346 4564 20352 4616
rect 20404 4604 20410 4616
rect 20404 4576 20449 4604
rect 20404 4564 20410 4576
rect 17310 4496 17316 4548
rect 17368 4536 17374 4548
rect 20622 4536 20628 4548
rect 17368 4508 20628 4536
rect 17368 4496 17374 4508
rect 20622 4496 20628 4508
rect 20680 4496 20686 4548
rect 15930 4468 15936 4480
rect 15764 4440 15936 4468
rect 15930 4428 15936 4440
rect 15988 4428 15994 4480
rect 18785 4471 18843 4477
rect 18785 4437 18797 4471
rect 18831 4468 18843 4471
rect 19058 4468 19064 4480
rect 18831 4440 19064 4468
rect 18831 4437 18843 4440
rect 18785 4431 18843 4437
rect 19058 4428 19064 4440
rect 19116 4428 19122 4480
rect 19794 4468 19800 4480
rect 19755 4440 19800 4468
rect 19794 4428 19800 4440
rect 19852 4428 19858 4480
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 7742 4224 7748 4276
rect 7800 4264 7806 4276
rect 17310 4264 17316 4276
rect 7800 4236 17316 4264
rect 7800 4224 7806 4236
rect 17310 4224 17316 4236
rect 17368 4224 17374 4276
rect 19702 4264 19708 4276
rect 19663 4236 19708 4264
rect 19702 4224 19708 4236
rect 19760 4224 19766 4276
rect 10686 4156 10692 4208
rect 10744 4196 10750 4208
rect 12618 4196 12624 4208
rect 10744 4168 12624 4196
rect 10744 4156 10750 4168
rect 12618 4156 12624 4168
rect 12676 4156 12682 4208
rect 13262 4156 13268 4208
rect 13320 4196 13326 4208
rect 13320 4168 13400 4196
rect 13320 4156 13326 4168
rect 8386 4088 8392 4140
rect 8444 4128 8450 4140
rect 9125 4131 9183 4137
rect 9125 4128 9137 4131
rect 8444 4100 9137 4128
rect 8444 4088 8450 4100
rect 9125 4097 9137 4100
rect 9171 4097 9183 4131
rect 11422 4128 11428 4140
rect 11383 4100 11428 4128
rect 9125 4091 9183 4097
rect 11422 4088 11428 4100
rect 11480 4088 11486 4140
rect 13372 4137 13400 4168
rect 14384 4168 14688 4196
rect 13357 4131 13415 4137
rect 13357 4097 13369 4131
rect 13403 4097 13415 4131
rect 13357 4091 13415 4097
rect 13630 4088 13636 4140
rect 13688 4128 13694 4140
rect 14384 4128 14412 4168
rect 14550 4128 14556 4140
rect 13688 4100 14412 4128
rect 14511 4100 14556 4128
rect 13688 4088 13694 4100
rect 14550 4088 14556 4100
rect 14608 4088 14614 4140
rect 14660 4128 14688 4168
rect 19886 4156 19892 4208
rect 19944 4196 19950 4208
rect 19944 4168 20300 4196
rect 19944 4156 19950 4168
rect 20162 4128 20168 4140
rect 14660 4100 16528 4128
rect 20123 4100 20168 4128
rect 9858 4060 9864 4072
rect 9039 4032 9864 4060
rect 842 3952 848 4004
rect 900 3992 906 4004
rect 9039 3992 9067 4032
rect 9858 4020 9864 4032
rect 9916 4020 9922 4072
rect 15010 4060 15016 4072
rect 14971 4032 15016 4060
rect 15010 4020 15016 4032
rect 15068 4020 15074 4072
rect 15746 4060 15752 4072
rect 15707 4032 15752 4060
rect 15746 4020 15752 4032
rect 15804 4020 15810 4072
rect 16500 4069 16528 4100
rect 20162 4088 20168 4100
rect 20220 4088 20226 4140
rect 20272 4137 20300 4168
rect 20257 4131 20315 4137
rect 20257 4097 20269 4131
rect 20303 4097 20315 4131
rect 20257 4091 20315 4097
rect 16485 4063 16543 4069
rect 16485 4029 16497 4063
rect 16531 4029 16543 4063
rect 16485 4023 16543 4029
rect 17218 4020 17224 4072
rect 17276 4060 17282 4072
rect 17405 4063 17463 4069
rect 17405 4060 17417 4063
rect 17276 4032 17417 4060
rect 17276 4020 17282 4032
rect 17405 4029 17417 4032
rect 17451 4029 17463 4063
rect 17405 4023 17463 4029
rect 18049 4063 18107 4069
rect 18049 4029 18061 4063
rect 18095 4060 18107 4063
rect 18598 4060 18604 4072
rect 18095 4032 18604 4060
rect 18095 4029 18107 4032
rect 18049 4023 18107 4029
rect 18598 4020 18604 4032
rect 18656 4020 18662 4072
rect 19794 4020 19800 4072
rect 19852 4060 19858 4072
rect 20073 4063 20131 4069
rect 20073 4060 20085 4063
rect 19852 4032 20085 4060
rect 19852 4020 19858 4032
rect 20073 4029 20085 4032
rect 20119 4029 20131 4063
rect 20714 4060 20720 4072
rect 20675 4032 20720 4060
rect 20073 4023 20131 4029
rect 20714 4020 20720 4032
rect 20772 4020 20778 4072
rect 900 3964 9067 3992
rect 9392 3995 9450 4001
rect 900 3952 906 3964
rect 9392 3961 9404 3995
rect 9438 3992 9450 3995
rect 9582 3992 9588 4004
rect 9438 3964 9588 3992
rect 9438 3961 9450 3964
rect 9392 3955 9450 3961
rect 9582 3952 9588 3964
rect 9640 3952 9646 4004
rect 10594 3992 10600 4004
rect 10244 3964 10600 3992
rect 7466 3884 7472 3936
rect 7524 3924 7530 3936
rect 10244 3924 10272 3964
rect 10594 3952 10600 3964
rect 10652 3952 10658 4004
rect 11149 3995 11207 4001
rect 11149 3961 11161 3995
rect 11195 3992 11207 3995
rect 11793 3995 11851 4001
rect 11793 3992 11805 3995
rect 11195 3964 11805 3992
rect 11195 3961 11207 3964
rect 11149 3955 11207 3961
rect 11793 3961 11805 3964
rect 11839 3961 11851 3995
rect 11793 3955 11851 3961
rect 13265 3995 13323 4001
rect 13265 3961 13277 3995
rect 13311 3992 13323 3995
rect 13354 3992 13360 4004
rect 13311 3964 13360 3992
rect 13311 3961 13323 3964
rect 13265 3955 13323 3961
rect 13354 3952 13360 3964
rect 13412 3992 13418 4004
rect 13630 3992 13636 4004
rect 13412 3964 13636 3992
rect 13412 3952 13418 3964
rect 13630 3952 13636 3964
rect 13688 3952 13694 4004
rect 14369 3995 14427 4001
rect 14369 3961 14381 3995
rect 14415 3992 14427 3995
rect 15378 3992 15384 4004
rect 14415 3964 15384 3992
rect 14415 3961 14427 3964
rect 14369 3955 14427 3961
rect 15378 3952 15384 3964
rect 15436 3952 15442 4004
rect 16025 3995 16083 4001
rect 16025 3961 16037 3995
rect 16071 3992 16083 3995
rect 16758 3992 16764 4004
rect 16071 3964 16764 3992
rect 16071 3961 16083 3964
rect 16025 3955 16083 3961
rect 16758 3952 16764 3964
rect 16816 3952 16822 4004
rect 16850 3952 16856 4004
rect 16908 3992 16914 4004
rect 17678 3992 17684 4004
rect 16908 3964 17684 3992
rect 16908 3952 16914 3964
rect 17678 3952 17684 3964
rect 17736 3952 17742 4004
rect 18316 3995 18374 4001
rect 18316 3961 18328 3995
rect 18362 3992 18374 3995
rect 18690 3992 18696 4004
rect 18362 3964 18696 3992
rect 18362 3961 18374 3964
rect 18316 3955 18374 3961
rect 18690 3952 18696 3964
rect 18748 3952 18754 4004
rect 7524 3896 10272 3924
rect 7524 3884 7530 3896
rect 10318 3884 10324 3936
rect 10376 3924 10382 3936
rect 10505 3927 10563 3933
rect 10505 3924 10517 3927
rect 10376 3896 10517 3924
rect 10376 3884 10382 3896
rect 10505 3893 10517 3896
rect 10551 3893 10563 3927
rect 10778 3924 10784 3936
rect 10739 3896 10784 3924
rect 10505 3887 10563 3893
rect 10778 3884 10784 3896
rect 10836 3884 10842 3936
rect 10870 3884 10876 3936
rect 10928 3924 10934 3936
rect 11241 3927 11299 3933
rect 11241 3924 11253 3927
rect 10928 3896 11253 3924
rect 10928 3884 10934 3896
rect 11241 3893 11253 3896
rect 11287 3893 11299 3927
rect 11241 3887 11299 3893
rect 11330 3884 11336 3936
rect 11388 3924 11394 3936
rect 12342 3924 12348 3936
rect 11388 3896 12348 3924
rect 11388 3884 11394 3896
rect 12342 3884 12348 3896
rect 12400 3884 12406 3936
rect 12802 3924 12808 3936
rect 12763 3896 12808 3924
rect 12802 3884 12808 3896
rect 12860 3884 12866 3936
rect 13173 3927 13231 3933
rect 13173 3893 13185 3927
rect 13219 3924 13231 3927
rect 13906 3924 13912 3936
rect 13219 3896 13912 3924
rect 13219 3893 13231 3896
rect 13173 3887 13231 3893
rect 13906 3884 13912 3896
rect 13964 3884 13970 3936
rect 14001 3927 14059 3933
rect 14001 3893 14013 3927
rect 14047 3924 14059 3927
rect 14090 3924 14096 3936
rect 14047 3896 14096 3924
rect 14047 3893 14059 3896
rect 14001 3887 14059 3893
rect 14090 3884 14096 3896
rect 14148 3884 14154 3936
rect 14274 3884 14280 3936
rect 14332 3924 14338 3936
rect 14461 3927 14519 3933
rect 14461 3924 14473 3927
rect 14332 3896 14473 3924
rect 14332 3884 14338 3896
rect 14461 3893 14473 3896
rect 14507 3893 14519 3927
rect 14461 3887 14519 3893
rect 15010 3884 15016 3936
rect 15068 3924 15074 3936
rect 15197 3927 15255 3933
rect 15197 3924 15209 3927
rect 15068 3896 15209 3924
rect 15068 3884 15074 3896
rect 15197 3893 15209 3896
rect 15243 3893 15255 3927
rect 15197 3887 15255 3893
rect 15838 3884 15844 3936
rect 15896 3924 15902 3936
rect 16669 3927 16727 3933
rect 16669 3924 16681 3927
rect 15896 3896 16681 3924
rect 15896 3884 15902 3896
rect 16669 3893 16681 3896
rect 16715 3893 16727 3927
rect 16669 3887 16727 3893
rect 17589 3927 17647 3933
rect 17589 3893 17601 3927
rect 17635 3924 17647 3927
rect 17862 3924 17868 3936
rect 17635 3896 17868 3924
rect 17635 3893 17647 3896
rect 17589 3887 17647 3893
rect 17862 3884 17868 3896
rect 17920 3884 17926 3936
rect 19150 3884 19156 3936
rect 19208 3924 19214 3936
rect 19429 3927 19487 3933
rect 19429 3924 19441 3927
rect 19208 3896 19441 3924
rect 19208 3884 19214 3896
rect 19429 3893 19441 3896
rect 19475 3893 19487 3927
rect 19429 3887 19487 3893
rect 20901 3927 20959 3933
rect 20901 3893 20913 3927
rect 20947 3924 20959 3927
rect 22462 3924 22468 3936
rect 20947 3896 22468 3924
rect 20947 3893 20959 3896
rect 20901 3887 20959 3893
rect 22462 3884 22468 3896
rect 22520 3884 22526 3936
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 9582 3680 9588 3732
rect 9640 3720 9646 3732
rect 11146 3720 11152 3732
rect 9640 3692 11152 3720
rect 9640 3680 9646 3692
rect 11146 3680 11152 3692
rect 11204 3680 11210 3732
rect 11422 3720 11428 3732
rect 11383 3692 11428 3720
rect 11422 3680 11428 3692
rect 11480 3680 11486 3732
rect 11698 3680 11704 3732
rect 11756 3720 11762 3732
rect 11756 3692 13400 3720
rect 11756 3680 11762 3692
rect 3602 3612 3608 3664
rect 3660 3652 3666 3664
rect 3660 3624 10456 3652
rect 3660 3612 3666 3624
rect 290 3544 296 3596
rect 348 3584 354 3596
rect 7190 3584 7196 3596
rect 348 3556 7196 3584
rect 348 3544 354 3556
rect 7190 3544 7196 3556
rect 7248 3544 7254 3596
rect 8386 3544 8392 3596
rect 8444 3584 8450 3596
rect 10318 3593 10324 3596
rect 10045 3587 10103 3593
rect 10045 3584 10057 3587
rect 8444 3556 10057 3584
rect 8444 3544 8450 3556
rect 10045 3553 10057 3556
rect 10091 3553 10103 3587
rect 10312 3584 10324 3593
rect 10279 3556 10324 3584
rect 10045 3547 10103 3553
rect 10312 3547 10324 3556
rect 10318 3544 10324 3547
rect 10376 3544 10382 3596
rect 10428 3584 10456 3624
rect 10502 3612 10508 3664
rect 10560 3652 10566 3664
rect 11330 3652 11336 3664
rect 10560 3624 11336 3652
rect 10560 3612 10566 3624
rect 11330 3612 11336 3624
rect 11388 3612 11394 3664
rect 11440 3652 11468 3680
rect 11946 3655 12004 3661
rect 11946 3652 11958 3655
rect 11440 3624 11958 3652
rect 11946 3621 11958 3624
rect 11992 3621 12004 3655
rect 11946 3615 12004 3621
rect 12710 3584 12716 3596
rect 10428 3556 12716 3584
rect 12710 3544 12716 3556
rect 12768 3544 12774 3596
rect 13372 3593 13400 3692
rect 13906 3680 13912 3732
rect 13964 3680 13970 3732
rect 14550 3680 14556 3732
rect 14608 3720 14614 3732
rect 14737 3723 14795 3729
rect 14737 3720 14749 3723
rect 14608 3692 14749 3720
rect 14608 3680 14614 3692
rect 14737 3689 14749 3692
rect 14783 3689 14795 3723
rect 16850 3720 16856 3732
rect 14737 3683 14795 3689
rect 14844 3692 16856 3720
rect 13924 3652 13952 3680
rect 14844 3652 14872 3692
rect 16850 3680 16856 3692
rect 16908 3680 16914 3732
rect 17037 3723 17095 3729
rect 17037 3689 17049 3723
rect 17083 3689 17095 3723
rect 18690 3720 18696 3732
rect 18651 3692 18696 3720
rect 17037 3683 17095 3689
rect 13924 3624 14872 3652
rect 15924 3655 15982 3661
rect 15924 3621 15936 3655
rect 15970 3652 15982 3655
rect 16114 3652 16120 3664
rect 15970 3624 16120 3652
rect 15970 3621 15982 3624
rect 15924 3615 15982 3621
rect 16114 3612 16120 3624
rect 16172 3612 16178 3664
rect 17052 3652 17080 3683
rect 18690 3680 18696 3692
rect 18748 3680 18754 3732
rect 17218 3652 17224 3664
rect 17052 3624 17224 3652
rect 17218 3612 17224 3624
rect 17276 3652 17282 3664
rect 17558 3655 17616 3661
rect 17558 3652 17570 3655
rect 17276 3624 17570 3652
rect 17276 3612 17282 3624
rect 17558 3621 17570 3624
rect 17604 3621 17616 3655
rect 17558 3615 17616 3621
rect 13357 3587 13415 3593
rect 13357 3553 13369 3587
rect 13403 3553 13415 3587
rect 13613 3587 13671 3593
rect 13613 3584 13625 3587
rect 13357 3547 13415 3553
rect 13464 3556 13625 3584
rect 3050 3476 3056 3528
rect 3108 3516 3114 3528
rect 9950 3516 9956 3528
rect 3108 3488 9956 3516
rect 3108 3476 3114 3488
rect 9950 3476 9956 3488
rect 10008 3476 10014 3528
rect 11698 3516 11704 3528
rect 11659 3488 11704 3516
rect 11698 3476 11704 3488
rect 11756 3476 11762 3528
rect 13464 3516 13492 3556
rect 13613 3553 13625 3556
rect 13659 3584 13671 3587
rect 13906 3584 13912 3596
rect 13659 3556 13912 3584
rect 13659 3553 13671 3556
rect 13613 3547 13671 3553
rect 13906 3544 13912 3556
rect 13964 3544 13970 3596
rect 15654 3584 15660 3596
rect 15615 3556 15660 3584
rect 15654 3544 15660 3556
rect 15712 3584 15718 3596
rect 17313 3587 17371 3593
rect 17313 3584 17325 3587
rect 15712 3556 17325 3584
rect 15712 3544 15718 3556
rect 17313 3553 17325 3556
rect 17359 3553 17371 3587
rect 19058 3584 19064 3596
rect 19019 3556 19064 3584
rect 17313 3547 17371 3553
rect 19058 3544 19064 3556
rect 19116 3544 19122 3596
rect 19610 3544 19616 3596
rect 19668 3584 19674 3596
rect 19797 3587 19855 3593
rect 19797 3584 19809 3587
rect 19668 3556 19809 3584
rect 19668 3544 19674 3556
rect 19797 3553 19809 3556
rect 19843 3553 19855 3587
rect 19797 3547 19855 3553
rect 13096 3488 13492 3516
rect 19337 3519 19395 3525
rect 8202 3408 8208 3460
rect 8260 3448 8266 3460
rect 10042 3448 10048 3460
rect 8260 3420 10048 3448
rect 8260 3408 8266 3420
rect 10042 3408 10048 3420
rect 10100 3408 10106 3460
rect 13096 3457 13124 3488
rect 19337 3485 19349 3519
rect 19383 3516 19395 3519
rect 19518 3516 19524 3528
rect 19383 3488 19524 3516
rect 19383 3485 19395 3488
rect 19337 3479 19395 3485
rect 19518 3476 19524 3488
rect 19576 3476 19582 3528
rect 20073 3519 20131 3525
rect 20073 3485 20085 3519
rect 20119 3516 20131 3519
rect 20346 3516 20352 3528
rect 20119 3488 20352 3516
rect 20119 3485 20131 3488
rect 20073 3479 20131 3485
rect 20346 3476 20352 3488
rect 20404 3476 20410 3528
rect 13081 3451 13139 3457
rect 13081 3417 13093 3451
rect 13127 3417 13139 3451
rect 13081 3411 13139 3417
rect 5810 3340 5816 3392
rect 5868 3380 5874 3392
rect 9306 3380 9312 3392
rect 5868 3352 9312 3380
rect 5868 3340 5874 3352
rect 9306 3340 9312 3352
rect 9364 3340 9370 3392
rect 9674 3340 9680 3392
rect 9732 3380 9738 3392
rect 12342 3380 12348 3392
rect 9732 3352 12348 3380
rect 9732 3340 9738 3352
rect 12342 3340 12348 3352
rect 12400 3340 12406 3392
rect 13998 3340 14004 3392
rect 14056 3380 14062 3392
rect 16298 3380 16304 3392
rect 14056 3352 16304 3380
rect 14056 3340 14062 3352
rect 16298 3340 16304 3352
rect 16356 3340 16362 3392
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 6362 3136 6368 3188
rect 6420 3176 6426 3188
rect 10226 3176 10232 3188
rect 6420 3148 10232 3176
rect 6420 3136 6426 3148
rect 10226 3136 10232 3148
rect 10284 3136 10290 3188
rect 10413 3179 10471 3185
rect 10413 3145 10425 3179
rect 10459 3176 10471 3179
rect 10870 3176 10876 3188
rect 10459 3148 10876 3176
rect 10459 3145 10471 3148
rect 10413 3139 10471 3145
rect 10870 3136 10876 3148
rect 10928 3136 10934 3188
rect 13357 3179 13415 3185
rect 13357 3145 13369 3179
rect 13403 3176 13415 3179
rect 14274 3176 14280 3188
rect 13403 3148 14280 3176
rect 13403 3145 13415 3148
rect 13357 3139 13415 3145
rect 14274 3136 14280 3148
rect 14332 3136 14338 3188
rect 15654 3176 15660 3188
rect 14384 3148 15660 3176
rect 7190 3068 7196 3120
rect 7248 3108 7254 3120
rect 7248 3080 14320 3108
rect 7248 3068 7254 3080
rect 14292 3052 14320 3080
rect 4154 3000 4160 3052
rect 4212 3040 4218 3052
rect 10226 3040 10232 3052
rect 4212 3012 10232 3040
rect 4212 3000 4218 3012
rect 10226 3000 10232 3012
rect 10284 3000 10290 3052
rect 10318 3000 10324 3052
rect 10376 3040 10382 3052
rect 10965 3043 11023 3049
rect 10965 3040 10977 3043
rect 10376 3012 10977 3040
rect 10376 3000 10382 3012
rect 10965 3009 10977 3012
rect 11011 3009 11023 3043
rect 13906 3040 13912 3052
rect 13867 3012 13912 3040
rect 10965 3003 11023 3009
rect 13906 3000 13912 3012
rect 13964 3000 13970 3052
rect 14274 3000 14280 3052
rect 14332 3000 14338 3052
rect 14384 3049 14412 3148
rect 15654 3136 15660 3148
rect 15712 3136 15718 3188
rect 16577 3179 16635 3185
rect 16577 3145 16589 3179
rect 16623 3176 16635 3179
rect 17126 3176 17132 3188
rect 16623 3148 17132 3176
rect 16623 3145 16635 3148
rect 16577 3139 16635 3145
rect 17126 3136 17132 3148
rect 17184 3136 17190 3188
rect 17954 3136 17960 3188
rect 18012 3176 18018 3188
rect 18049 3179 18107 3185
rect 18049 3176 18061 3179
rect 18012 3148 18061 3176
rect 18012 3136 18018 3148
rect 18049 3145 18061 3148
rect 18095 3145 18107 3179
rect 18049 3139 18107 3145
rect 16209 3111 16267 3117
rect 16209 3077 16221 3111
rect 16255 3108 16267 3111
rect 16850 3108 16856 3120
rect 16255 3080 16856 3108
rect 16255 3077 16267 3080
rect 16209 3071 16267 3077
rect 16850 3068 16856 3080
rect 16908 3068 16914 3120
rect 17678 3068 17684 3120
rect 17736 3108 17742 3120
rect 19613 3111 19671 3117
rect 17736 3080 19564 3108
rect 17736 3068 17742 3080
rect 14369 3043 14427 3049
rect 14369 3009 14381 3043
rect 14415 3009 14427 3043
rect 17218 3040 17224 3052
rect 17179 3012 17224 3040
rect 14369 3003 14427 3009
rect 17218 3000 17224 3012
rect 17276 3000 17282 3052
rect 18506 3040 18512 3052
rect 18467 3012 18512 3040
rect 18506 3000 18512 3012
rect 18564 3000 18570 3052
rect 18690 3040 18696 3052
rect 18651 3012 18696 3040
rect 18690 3000 18696 3012
rect 18748 3000 18754 3052
rect 8570 2932 8576 2984
rect 8628 2972 8634 2984
rect 10686 2972 10692 2984
rect 8628 2944 10692 2972
rect 8628 2932 8634 2944
rect 10686 2932 10692 2944
rect 10744 2932 10750 2984
rect 11606 2972 11612 2984
rect 11567 2944 11612 2972
rect 11606 2932 11612 2944
rect 11664 2932 11670 2984
rect 12437 2975 12495 2981
rect 12437 2941 12449 2975
rect 12483 2972 12495 2975
rect 13817 2975 13875 2981
rect 12483 2944 12940 2972
rect 12483 2941 12495 2944
rect 12437 2935 12495 2941
rect 2498 2864 2504 2916
rect 2556 2904 2562 2916
rect 2556 2876 11284 2904
rect 2556 2864 2562 2876
rect 4706 2796 4712 2848
rect 4764 2836 4770 2848
rect 10781 2839 10839 2845
rect 10781 2836 10793 2839
rect 4764 2808 10793 2836
rect 4764 2796 4770 2808
rect 10781 2805 10793 2808
rect 10827 2805 10839 2839
rect 10781 2799 10839 2805
rect 10873 2839 10931 2845
rect 10873 2805 10885 2839
rect 10919 2836 10931 2839
rect 11146 2836 11152 2848
rect 10919 2808 11152 2836
rect 10919 2805 10931 2808
rect 10873 2799 10931 2805
rect 11146 2796 11152 2808
rect 11204 2796 11210 2848
rect 11256 2836 11284 2876
rect 11330 2864 11336 2916
rect 11388 2904 11394 2916
rect 11885 2907 11943 2913
rect 11885 2904 11897 2907
rect 11388 2876 11897 2904
rect 11388 2864 11394 2876
rect 11885 2873 11897 2876
rect 11931 2873 11943 2907
rect 11885 2867 11943 2873
rect 12526 2864 12532 2916
rect 12584 2904 12590 2916
rect 12713 2907 12771 2913
rect 12713 2904 12725 2907
rect 12584 2876 12725 2904
rect 12584 2864 12590 2876
rect 12713 2873 12725 2876
rect 12759 2873 12771 2907
rect 12912 2904 12940 2944
rect 13817 2941 13829 2975
rect 13863 2972 13875 2975
rect 13998 2972 14004 2984
rect 13863 2944 14004 2972
rect 13863 2941 13875 2944
rect 13817 2935 13875 2941
rect 13998 2932 14004 2944
rect 14056 2932 14062 2984
rect 15930 2932 15936 2984
rect 15988 2972 15994 2984
rect 16025 2975 16083 2981
rect 16025 2972 16037 2975
rect 15988 2944 16037 2972
rect 15988 2932 15994 2944
rect 16025 2941 16037 2944
rect 16071 2941 16083 2975
rect 16942 2972 16948 2984
rect 16903 2944 16948 2972
rect 16025 2935 16083 2941
rect 16942 2932 16948 2944
rect 17000 2932 17006 2984
rect 18414 2972 18420 2984
rect 18375 2944 18420 2972
rect 18414 2932 18420 2944
rect 18472 2972 18478 2984
rect 18877 2975 18935 2981
rect 18877 2972 18889 2975
rect 18472 2944 18889 2972
rect 18472 2932 18478 2944
rect 18877 2941 18889 2944
rect 18923 2941 18935 2975
rect 19426 2972 19432 2984
rect 19387 2944 19432 2972
rect 18877 2935 18935 2941
rect 19426 2932 19432 2944
rect 19484 2932 19490 2984
rect 19536 2972 19564 3080
rect 19613 3077 19625 3111
rect 19659 3108 19671 3111
rect 20254 3108 20260 3120
rect 19659 3080 20260 3108
rect 19659 3077 19671 3080
rect 19613 3071 19671 3077
rect 20254 3068 20260 3080
rect 20312 3068 20318 3120
rect 19981 2975 20039 2981
rect 19981 2972 19993 2975
rect 19536 2944 19993 2972
rect 19981 2941 19993 2944
rect 20027 2941 20039 2975
rect 20530 2972 20536 2984
rect 20491 2944 20536 2972
rect 19981 2935 20039 2941
rect 20530 2932 20536 2944
rect 20588 2932 20594 2984
rect 12912 2876 13952 2904
rect 12713 2867 12771 2873
rect 13725 2839 13783 2845
rect 13725 2836 13737 2839
rect 11256 2808 13737 2836
rect 13725 2805 13737 2808
rect 13771 2805 13783 2839
rect 13924 2836 13952 2876
rect 14550 2864 14556 2916
rect 14608 2913 14614 2916
rect 14608 2907 14672 2913
rect 14608 2873 14626 2907
rect 14660 2873 14672 2907
rect 21358 2904 21364 2916
rect 14608 2867 14672 2873
rect 20180 2876 21364 2904
rect 14608 2864 14614 2867
rect 15562 2836 15568 2848
rect 13924 2808 15568 2836
rect 13725 2799 13783 2805
rect 15562 2796 15568 2808
rect 15620 2796 15626 2848
rect 15749 2839 15807 2845
rect 15749 2805 15761 2839
rect 15795 2836 15807 2839
rect 16114 2836 16120 2848
rect 15795 2808 16120 2836
rect 15795 2805 15807 2808
rect 15749 2799 15807 2805
rect 16114 2796 16120 2808
rect 16172 2796 16178 2848
rect 17034 2836 17040 2848
rect 16995 2808 17040 2836
rect 17034 2796 17040 2808
rect 17092 2796 17098 2848
rect 20180 2845 20208 2876
rect 21358 2864 21364 2876
rect 21416 2864 21422 2916
rect 20165 2839 20223 2845
rect 20165 2805 20177 2839
rect 20211 2805 20223 2839
rect 20165 2799 20223 2805
rect 20717 2839 20775 2845
rect 20717 2805 20729 2839
rect 20763 2836 20775 2839
rect 21910 2836 21916 2848
rect 20763 2808 21916 2836
rect 20763 2805 20775 2808
rect 20717 2799 20775 2805
rect 21910 2796 21916 2808
rect 21968 2796 21974 2848
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 9766 2592 9772 2644
rect 9824 2632 9830 2644
rect 10226 2632 10232 2644
rect 9824 2604 10232 2632
rect 9824 2592 9830 2604
rect 10226 2592 10232 2604
rect 10284 2592 10290 2644
rect 10778 2592 10784 2644
rect 10836 2632 10842 2644
rect 12250 2632 12256 2644
rect 10836 2604 12256 2632
rect 10836 2592 10842 2604
rect 12250 2592 12256 2604
rect 12308 2592 12314 2644
rect 16022 2592 16028 2644
rect 16080 2632 16086 2644
rect 18138 2632 18144 2644
rect 16080 2604 18144 2632
rect 16080 2592 16086 2604
rect 18138 2592 18144 2604
rect 18196 2592 18202 2644
rect 13722 2564 13728 2576
rect 7576 2536 13584 2564
rect 13683 2536 13728 2564
rect 1394 2388 1400 2440
rect 1452 2428 1458 2440
rect 7576 2428 7604 2536
rect 11330 2496 11336 2508
rect 11291 2468 11336 2496
rect 11330 2456 11336 2468
rect 11388 2456 11394 2508
rect 11885 2499 11943 2505
rect 11885 2465 11897 2499
rect 11931 2496 11943 2499
rect 12526 2496 12532 2508
rect 11931 2468 12532 2496
rect 11931 2465 11943 2468
rect 11885 2459 11943 2465
rect 12526 2456 12532 2468
rect 12584 2456 12590 2508
rect 12713 2499 12771 2505
rect 12713 2465 12725 2499
rect 12759 2496 12771 2499
rect 12986 2496 12992 2508
rect 12759 2468 12992 2496
rect 12759 2465 12771 2468
rect 12713 2459 12771 2465
rect 12986 2456 12992 2468
rect 13044 2456 13050 2508
rect 13446 2496 13452 2508
rect 13407 2468 13452 2496
rect 13446 2456 13452 2468
rect 13504 2456 13510 2508
rect 13556 2496 13584 2536
rect 13722 2524 13728 2536
rect 13780 2524 13786 2576
rect 17770 2564 17776 2576
rect 13832 2536 14320 2564
rect 13832 2496 13860 2536
rect 13556 2468 13860 2496
rect 14185 2499 14243 2505
rect 14185 2465 14197 2499
rect 14231 2465 14243 2499
rect 14185 2459 14243 2465
rect 1452 2400 7604 2428
rect 12897 2431 12955 2437
rect 1452 2388 1458 2400
rect 12897 2397 12909 2431
rect 12943 2428 12955 2431
rect 14200 2428 14228 2459
rect 12943 2400 14228 2428
rect 14292 2428 14320 2536
rect 14752 2536 17776 2564
rect 14752 2505 14780 2536
rect 17770 2524 17776 2536
rect 17828 2524 17834 2576
rect 14737 2499 14795 2505
rect 14737 2465 14749 2499
rect 14783 2465 14795 2499
rect 14737 2459 14795 2465
rect 15933 2499 15991 2505
rect 15933 2465 15945 2499
rect 15979 2465 15991 2499
rect 15933 2459 15991 2465
rect 16577 2499 16635 2505
rect 16577 2465 16589 2499
rect 16623 2496 16635 2499
rect 16758 2496 16764 2508
rect 16623 2468 16764 2496
rect 16623 2465 16635 2468
rect 16577 2459 16635 2465
rect 15948 2428 15976 2459
rect 16758 2456 16764 2468
rect 16816 2456 16822 2508
rect 17310 2496 17316 2508
rect 17271 2468 17316 2496
rect 17310 2456 17316 2468
rect 17368 2456 17374 2508
rect 17402 2456 17408 2508
rect 17460 2496 17466 2508
rect 18417 2499 18475 2505
rect 18417 2496 18429 2499
rect 17460 2468 18429 2496
rect 17460 2456 17466 2468
rect 18417 2465 18429 2468
rect 18463 2465 18475 2499
rect 18966 2496 18972 2508
rect 18927 2468 18972 2496
rect 18417 2459 18475 2465
rect 18966 2456 18972 2468
rect 19024 2456 19030 2508
rect 19518 2496 19524 2508
rect 19479 2468 19524 2496
rect 19518 2456 19524 2468
rect 19576 2456 19582 2508
rect 20346 2496 20352 2508
rect 20307 2468 20352 2496
rect 20346 2456 20352 2468
rect 20404 2456 20410 2508
rect 14292 2400 15976 2428
rect 12943 2397 12955 2400
rect 12897 2391 12955 2397
rect 16114 2388 16120 2440
rect 16172 2428 16178 2440
rect 16172 2400 16217 2428
rect 16172 2388 16178 2400
rect 16298 2388 16304 2440
rect 16356 2428 16362 2440
rect 19242 2428 19248 2440
rect 16356 2400 19248 2428
rect 16356 2388 16362 2400
rect 19242 2388 19248 2400
rect 19300 2388 19306 2440
rect 11517 2363 11575 2369
rect 11517 2329 11529 2363
rect 11563 2360 11575 2363
rect 13078 2360 13084 2372
rect 11563 2332 13084 2360
rect 11563 2329 11575 2332
rect 11517 2323 11575 2329
rect 13078 2320 13084 2332
rect 13136 2320 13142 2372
rect 13630 2320 13636 2372
rect 13688 2360 13694 2372
rect 14921 2363 14979 2369
rect 14921 2360 14933 2363
rect 13688 2332 14933 2360
rect 13688 2320 13694 2332
rect 14921 2329 14933 2332
rect 14967 2329 14979 2363
rect 14921 2323 14979 2329
rect 15565 2363 15623 2369
rect 15565 2329 15577 2363
rect 15611 2360 15623 2363
rect 17034 2360 17040 2372
rect 15611 2332 17040 2360
rect 15611 2329 15623 2332
rect 15565 2323 15623 2329
rect 17034 2320 17040 2332
rect 17092 2320 17098 2372
rect 18690 2320 18696 2372
rect 18748 2360 18754 2372
rect 19705 2363 19763 2369
rect 19705 2360 19717 2363
rect 18748 2332 19717 2360
rect 18748 2320 18754 2332
rect 19705 2329 19717 2332
rect 19751 2329 19763 2363
rect 19705 2323 19763 2329
rect 11974 2252 11980 2304
rect 12032 2292 12038 2304
rect 12069 2295 12127 2301
rect 12069 2292 12081 2295
rect 12032 2264 12081 2292
rect 12032 2252 12038 2264
rect 12069 2261 12081 2264
rect 12115 2261 12127 2295
rect 12069 2255 12127 2261
rect 12526 2252 12532 2304
rect 12584 2292 12590 2304
rect 14369 2295 14427 2301
rect 14369 2292 14381 2295
rect 12584 2264 14381 2292
rect 12584 2252 12590 2264
rect 14369 2261 14381 2264
rect 14415 2261 14427 2295
rect 14369 2255 14427 2261
rect 16390 2252 16396 2304
rect 16448 2292 16454 2304
rect 16761 2295 16819 2301
rect 16761 2292 16773 2295
rect 16448 2264 16773 2292
rect 16448 2252 16454 2264
rect 16761 2261 16773 2264
rect 16807 2261 16819 2295
rect 17494 2292 17500 2304
rect 17455 2264 17500 2292
rect 16761 2255 16819 2261
rect 17494 2252 17500 2264
rect 17552 2252 17558 2304
rect 18601 2295 18659 2301
rect 18601 2261 18613 2295
rect 18647 2292 18659 2295
rect 19058 2292 19064 2304
rect 18647 2264 19064 2292
rect 18647 2261 18659 2264
rect 18601 2255 18659 2261
rect 19058 2252 19064 2264
rect 19116 2252 19122 2304
rect 19153 2295 19211 2301
rect 19153 2261 19165 2295
rect 19199 2292 19211 2295
rect 19610 2292 19616 2304
rect 19199 2264 19616 2292
rect 19199 2261 19211 2264
rect 19153 2255 19211 2261
rect 19610 2252 19616 2264
rect 19668 2252 19674 2304
rect 20533 2295 20591 2301
rect 20533 2261 20545 2295
rect 20579 2292 20591 2295
rect 20806 2292 20812 2304
rect 20579 2264 20812 2292
rect 20579 2261 20591 2264
rect 20533 2255 20591 2261
rect 20806 2252 20812 2264
rect 20864 2252 20870 2304
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 11146 2048 11152 2100
rect 11204 2088 11210 2100
rect 13538 2088 13544 2100
rect 11204 2060 13544 2088
rect 11204 2048 11210 2060
rect 13538 2048 13544 2060
rect 13596 2088 13602 2100
rect 18506 2088 18512 2100
rect 13596 2060 18512 2088
rect 13596 2048 13602 2060
rect 18506 2048 18512 2060
rect 18564 2048 18570 2100
rect 5258 1980 5264 2032
rect 5316 2020 5322 2032
rect 8938 2020 8944 2032
rect 5316 1992 8944 2020
rect 5316 1980 5322 1992
rect 8938 1980 8944 1992
rect 8996 1980 9002 2032
rect 1946 1096 1952 1148
rect 2004 1136 2010 1148
rect 9582 1136 9588 1148
rect 2004 1108 9588 1136
rect 2004 1096 2010 1108
rect 9582 1096 9588 1108
rect 9640 1096 9646 1148
<< via1 >>
rect 7472 20204 7524 20256
rect 12072 20204 12124 20256
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 11152 20000 11204 20052
rect 11336 20000 11388 20052
rect 12072 20000 12124 20052
rect 12348 20000 12400 20052
rect 13084 20000 13136 20052
rect 10784 19932 10836 19984
rect 14188 20000 14240 20052
rect 14556 20000 14608 20052
rect 15292 20000 15344 20052
rect 16580 20000 16632 20052
rect 17500 20000 17552 20052
rect 18052 20000 18104 20052
rect 19156 20000 19208 20052
rect 19708 20000 19760 20052
rect 20168 20043 20220 20052
rect 20168 20009 20177 20043
rect 20177 20009 20211 20043
rect 20211 20009 20220 20043
rect 20168 20000 20220 20009
rect 20628 20000 20680 20052
rect 10876 19864 10928 19916
rect 12624 19907 12676 19916
rect 12624 19873 12633 19907
rect 12633 19873 12667 19907
rect 12667 19873 12676 19907
rect 12624 19864 12676 19873
rect 10692 19796 10744 19848
rect 12072 19839 12124 19848
rect 12072 19805 12081 19839
rect 12081 19805 12115 19839
rect 12115 19805 12124 19839
rect 12072 19796 12124 19805
rect 11888 19728 11940 19780
rect 20260 19932 20312 19984
rect 13084 19864 13136 19916
rect 14096 19907 14148 19916
rect 14096 19873 14105 19907
rect 14105 19873 14139 19907
rect 14139 19873 14148 19907
rect 14096 19864 14148 19873
rect 13912 19796 13964 19848
rect 15016 19864 15068 19916
rect 15384 19796 15436 19848
rect 17132 19864 17184 19916
rect 17408 19796 17460 19848
rect 18696 19864 18748 19916
rect 19432 19907 19484 19916
rect 19432 19873 19441 19907
rect 19441 19873 19475 19907
rect 19475 19873 19484 19907
rect 19432 19864 19484 19873
rect 19984 19907 20036 19916
rect 19984 19873 19993 19907
rect 19993 19873 20027 19907
rect 20027 19873 20036 19907
rect 19984 19864 20036 19873
rect 20168 19864 20220 19916
rect 10324 19660 10376 19712
rect 12164 19660 12216 19712
rect 17960 19660 18012 19712
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 8484 19456 8536 19508
rect 10508 19456 10560 19508
rect 7748 19252 7800 19304
rect 8484 19295 8536 19304
rect 8484 19261 8493 19295
rect 8493 19261 8527 19295
rect 8527 19261 8536 19295
rect 8484 19252 8536 19261
rect 11796 19295 11848 19304
rect 8208 19184 8260 19236
rect 8944 19184 8996 19236
rect 11796 19261 11805 19295
rect 11805 19261 11839 19295
rect 11839 19261 11848 19295
rect 11796 19252 11848 19261
rect 6368 19116 6420 19168
rect 9312 19116 9364 19168
rect 11888 19184 11940 19236
rect 12072 19184 12124 19236
rect 10692 19116 10744 19168
rect 11520 19159 11572 19168
rect 11520 19125 11529 19159
rect 11529 19125 11563 19159
rect 11563 19125 11572 19159
rect 11520 19116 11572 19125
rect 12532 19116 12584 19168
rect 12808 19116 12860 19168
rect 14188 19252 14240 19304
rect 14280 19252 14332 19304
rect 15016 19295 15068 19304
rect 15016 19261 15025 19295
rect 15025 19261 15059 19295
rect 15059 19261 15068 19295
rect 15016 19252 15068 19261
rect 16672 19320 16724 19372
rect 16856 19252 16908 19304
rect 13636 19184 13688 19236
rect 13820 19159 13872 19168
rect 13820 19125 13829 19159
rect 13829 19125 13863 19159
rect 13863 19125 13872 19159
rect 13820 19116 13872 19125
rect 16120 19159 16172 19168
rect 16120 19125 16129 19159
rect 16129 19125 16163 19159
rect 16163 19125 16172 19159
rect 16120 19116 16172 19125
rect 16212 19159 16264 19168
rect 16212 19125 16221 19159
rect 16221 19125 16255 19159
rect 16255 19125 16264 19159
rect 17316 19227 17368 19236
rect 17316 19193 17325 19227
rect 17325 19193 17359 19227
rect 17359 19193 17368 19227
rect 17868 19252 17920 19304
rect 19156 19252 19208 19304
rect 17316 19184 17368 19193
rect 20076 19184 20128 19236
rect 20536 19227 20588 19236
rect 20536 19193 20545 19227
rect 20545 19193 20579 19227
rect 20579 19193 20588 19227
rect 20536 19184 20588 19193
rect 16212 19116 16264 19125
rect 19064 19116 19116 19168
rect 19248 19159 19300 19168
rect 19248 19125 19257 19159
rect 19257 19125 19291 19159
rect 19291 19125 19300 19159
rect 19248 19116 19300 19125
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 296 18912 348 18964
rect 8944 18912 8996 18964
rect 12072 18912 12124 18964
rect 9864 18844 9916 18896
rect 10600 18844 10652 18896
rect 11520 18844 11572 18896
rect 13544 18912 13596 18964
rect 13820 18912 13872 18964
rect 16672 18955 16724 18964
rect 16672 18921 16681 18955
rect 16681 18921 16715 18955
rect 16715 18921 16724 18955
rect 16672 18912 16724 18921
rect 16948 18912 17000 18964
rect 18512 18912 18564 18964
rect 18604 18912 18656 18964
rect 18880 18912 18932 18964
rect 21916 18912 21968 18964
rect 7748 18819 7800 18828
rect 7748 18785 7757 18819
rect 7757 18785 7791 18819
rect 7791 18785 7800 18819
rect 7748 18776 7800 18785
rect 8852 18776 8904 18828
rect 10232 18776 10284 18828
rect 10508 18819 10560 18828
rect 10508 18785 10517 18819
rect 10517 18785 10551 18819
rect 10551 18785 10560 18819
rect 10508 18776 10560 18785
rect 12072 18776 12124 18828
rect 13636 18844 13688 18896
rect 15292 18844 15344 18896
rect 15476 18844 15528 18896
rect 19984 18887 20036 18896
rect 19984 18853 19993 18887
rect 19993 18853 20027 18887
rect 20027 18853 20036 18887
rect 19984 18844 20036 18853
rect 13268 18776 13320 18828
rect 9680 18708 9732 18760
rect 10416 18708 10468 18760
rect 14188 18708 14240 18760
rect 15108 18708 15160 18760
rect 15292 18751 15344 18760
rect 15292 18717 15301 18751
rect 15301 18717 15335 18751
rect 15335 18717 15344 18751
rect 15292 18708 15344 18717
rect 16580 18776 16632 18828
rect 17316 18776 17368 18828
rect 18788 18776 18840 18828
rect 19524 18776 19576 18828
rect 19708 18819 19760 18828
rect 19708 18785 19717 18819
rect 19717 18785 19751 18819
rect 19751 18785 19760 18819
rect 19708 18776 19760 18785
rect 16764 18708 16816 18760
rect 17040 18708 17092 18760
rect 21364 18708 21416 18760
rect 3056 18640 3108 18692
rect 4712 18572 4764 18624
rect 6184 18572 6236 18624
rect 9772 18640 9824 18692
rect 12256 18572 12308 18624
rect 14188 18572 14240 18624
rect 20812 18640 20864 18692
rect 19248 18572 19300 18624
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 9588 18368 9640 18420
rect 11980 18368 12032 18420
rect 13268 18368 13320 18420
rect 9956 18343 10008 18352
rect 3608 18232 3660 18284
rect 8208 18232 8260 18284
rect 8944 18232 8996 18284
rect 9956 18309 9965 18343
rect 9965 18309 9999 18343
rect 9999 18309 10008 18343
rect 9956 18300 10008 18309
rect 10508 18300 10560 18352
rect 10692 18300 10744 18352
rect 15844 18368 15896 18420
rect 17040 18368 17092 18420
rect 19156 18368 19208 18420
rect 10140 18232 10192 18284
rect 10416 18275 10468 18284
rect 10416 18241 10425 18275
rect 10425 18241 10459 18275
rect 10459 18241 10468 18275
rect 10416 18232 10468 18241
rect 10600 18275 10652 18284
rect 10600 18241 10609 18275
rect 10609 18241 10643 18275
rect 10643 18241 10652 18275
rect 10600 18232 10652 18241
rect 11152 18232 11204 18284
rect 9128 18164 9180 18216
rect 9312 18207 9364 18216
rect 9312 18173 9321 18207
rect 9321 18173 9355 18207
rect 9355 18173 9364 18207
rect 9312 18164 9364 18173
rect 4160 18096 4212 18148
rect 9496 18096 9548 18148
rect 10324 18139 10376 18148
rect 10324 18105 10333 18139
rect 10333 18105 10367 18139
rect 10367 18105 10376 18139
rect 10324 18096 10376 18105
rect 5816 18028 5868 18080
rect 7472 18028 7524 18080
rect 10600 18028 10652 18080
rect 13176 18164 13228 18216
rect 13636 18164 13688 18216
rect 15292 18232 15344 18284
rect 16304 18275 16356 18284
rect 16304 18241 16313 18275
rect 16313 18241 16347 18275
rect 16347 18241 16356 18275
rect 16304 18232 16356 18241
rect 17960 18300 18012 18352
rect 18880 18232 18932 18284
rect 19064 18232 19116 18284
rect 14188 18207 14240 18216
rect 14188 18173 14222 18207
rect 14222 18173 14240 18207
rect 14188 18164 14240 18173
rect 15752 18164 15804 18216
rect 16672 18096 16724 18148
rect 19984 18096 20036 18148
rect 13268 18071 13320 18080
rect 13268 18037 13277 18071
rect 13277 18037 13311 18071
rect 13311 18037 13320 18071
rect 13268 18028 13320 18037
rect 13360 18071 13412 18080
rect 13360 18037 13369 18071
rect 13369 18037 13403 18071
rect 13403 18037 13412 18071
rect 13360 18028 13412 18037
rect 15476 18028 15528 18080
rect 16304 18028 16356 18080
rect 18144 18071 18196 18080
rect 18144 18037 18153 18071
rect 18153 18037 18187 18071
rect 18187 18037 18196 18071
rect 18144 18028 18196 18037
rect 18604 18071 18656 18080
rect 18604 18037 18613 18071
rect 18613 18037 18647 18071
rect 18647 18037 18656 18071
rect 18604 18028 18656 18037
rect 18696 18028 18748 18080
rect 20812 18139 20864 18148
rect 20812 18105 20821 18139
rect 20821 18105 20855 18139
rect 20855 18105 20864 18139
rect 20812 18096 20864 18105
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 7748 17824 7800 17876
rect 8668 17824 8720 17876
rect 8852 17824 8904 17876
rect 9680 17867 9732 17876
rect 9680 17833 9689 17867
rect 9689 17833 9723 17867
rect 9723 17833 9732 17867
rect 9680 17824 9732 17833
rect 12900 17824 12952 17876
rect 13268 17824 13320 17876
rect 16120 17824 16172 17876
rect 16396 17824 16448 17876
rect 848 17756 900 17808
rect 8484 17756 8536 17808
rect 9956 17756 10008 17808
rect 18144 17824 18196 17876
rect 19984 17824 20036 17876
rect 7656 17688 7708 17740
rect 8392 17688 8444 17740
rect 10140 17731 10192 17740
rect 10140 17697 10149 17731
rect 10149 17697 10183 17731
rect 10183 17697 10192 17731
rect 10140 17688 10192 17697
rect 11888 17731 11940 17740
rect 11888 17697 11897 17731
rect 11897 17697 11931 17731
rect 11931 17697 11940 17731
rect 11888 17688 11940 17697
rect 10324 17663 10376 17672
rect 10324 17629 10333 17663
rect 10333 17629 10367 17663
rect 10367 17629 10376 17663
rect 10324 17620 10376 17629
rect 11612 17620 11664 17672
rect 14556 17731 14608 17740
rect 14556 17697 14565 17731
rect 14565 17697 14599 17731
rect 14599 17697 14608 17731
rect 14556 17688 14608 17697
rect 12992 17620 13044 17672
rect 13452 17663 13504 17672
rect 13452 17629 13461 17663
rect 13461 17629 13495 17663
rect 13495 17629 13504 17663
rect 13452 17620 13504 17629
rect 13544 17663 13596 17672
rect 13544 17629 13553 17663
rect 13553 17629 13587 17663
rect 13587 17629 13596 17663
rect 13544 17620 13596 17629
rect 14004 17620 14056 17672
rect 15016 17620 15068 17672
rect 15936 17620 15988 17672
rect 16304 17663 16356 17672
rect 16304 17629 16313 17663
rect 16313 17629 16347 17663
rect 16347 17629 16356 17663
rect 16672 17688 16724 17740
rect 18880 17756 18932 17808
rect 19156 17688 19208 17740
rect 16304 17620 16356 17629
rect 16948 17552 17000 17604
rect 11060 17484 11112 17536
rect 15568 17484 15620 17536
rect 16488 17484 16540 17536
rect 18512 17595 18564 17604
rect 18512 17561 18521 17595
rect 18521 17561 18555 17595
rect 18555 17561 18564 17595
rect 19616 17620 19668 17672
rect 18512 17552 18564 17561
rect 19432 17484 19484 17536
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 8392 17323 8444 17332
rect 8392 17289 8401 17323
rect 8401 17289 8435 17323
rect 8435 17289 8444 17323
rect 8392 17280 8444 17289
rect 8484 17280 8536 17332
rect 8852 17212 8904 17264
rect 8760 17144 8812 17196
rect 10692 17144 10744 17196
rect 11704 17144 11756 17196
rect 8668 17076 8720 17128
rect 9312 17076 9364 17128
rect 7656 17008 7708 17060
rect 10600 17076 10652 17128
rect 11520 17076 11572 17128
rect 11612 17076 11664 17128
rect 13360 17280 13412 17332
rect 14004 17212 14056 17264
rect 14556 17280 14608 17332
rect 16212 17280 16264 17332
rect 22468 17280 22520 17332
rect 18052 17212 18104 17264
rect 12164 17144 12216 17196
rect 13544 17144 13596 17196
rect 14464 17144 14516 17196
rect 16304 17187 16356 17196
rect 16304 17153 16313 17187
rect 16313 17153 16347 17187
rect 16347 17153 16356 17187
rect 16304 17144 16356 17153
rect 20720 17144 20772 17196
rect 16396 17076 16448 17128
rect 16764 17076 16816 17128
rect 17960 17076 18012 17128
rect 9036 16983 9088 16992
rect 9036 16949 9045 16983
rect 9045 16949 9079 16983
rect 9079 16949 9088 16983
rect 9036 16940 9088 16949
rect 9312 16940 9364 16992
rect 9772 16940 9824 16992
rect 9864 16940 9916 16992
rect 10784 16983 10836 16992
rect 10784 16949 10793 16983
rect 10793 16949 10827 16983
rect 10827 16949 10836 16983
rect 10784 16940 10836 16949
rect 11244 16983 11296 16992
rect 11244 16949 11253 16983
rect 11253 16949 11287 16983
rect 11287 16949 11296 16983
rect 11244 16940 11296 16949
rect 15660 17008 15712 17060
rect 13452 16940 13504 16992
rect 13820 16940 13872 16992
rect 14188 16940 14240 16992
rect 14372 16940 14424 16992
rect 15476 16940 15528 16992
rect 17776 17008 17828 17060
rect 19432 17076 19484 17128
rect 20444 17119 20496 17128
rect 20444 17085 20453 17119
rect 20453 17085 20487 17119
rect 20487 17085 20496 17119
rect 20444 17076 20496 17085
rect 18512 17008 18564 17060
rect 19524 17008 19576 17060
rect 16304 16940 16356 16992
rect 17960 16940 18012 16992
rect 19340 16940 19392 16992
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 6920 16736 6972 16788
rect 7472 16779 7524 16788
rect 7472 16745 7481 16779
rect 7481 16745 7515 16779
rect 7515 16745 7524 16779
rect 7472 16736 7524 16745
rect 7748 16736 7800 16788
rect 9864 16736 9916 16788
rect 11520 16736 11572 16788
rect 11888 16736 11940 16788
rect 16212 16736 16264 16788
rect 14464 16668 14516 16720
rect 17040 16668 17092 16720
rect 9220 16600 9272 16652
rect 9496 16643 9548 16652
rect 9496 16609 9505 16643
rect 9505 16609 9539 16643
rect 9539 16609 9548 16643
rect 9496 16600 9548 16609
rect 9680 16643 9732 16652
rect 9680 16609 9689 16643
rect 9689 16609 9723 16643
rect 9723 16609 9732 16643
rect 9680 16600 9732 16609
rect 10692 16643 10744 16652
rect 10692 16609 10726 16643
rect 10726 16609 10744 16643
rect 10692 16600 10744 16609
rect 13636 16600 13688 16652
rect 16120 16643 16172 16652
rect 7656 16575 7708 16584
rect 7656 16541 7665 16575
rect 7665 16541 7699 16575
rect 7699 16541 7708 16575
rect 7656 16532 7708 16541
rect 8208 16532 8260 16584
rect 8760 16575 8812 16584
rect 8760 16541 8769 16575
rect 8769 16541 8803 16575
rect 8803 16541 8812 16575
rect 8760 16532 8812 16541
rect 10324 16532 10376 16584
rect 8668 16464 8720 16516
rect 9404 16464 9456 16516
rect 12256 16532 12308 16584
rect 16120 16609 16129 16643
rect 16129 16609 16163 16643
rect 16163 16609 16172 16643
rect 16120 16600 16172 16609
rect 12348 16464 12400 16516
rect 12440 16396 12492 16448
rect 13728 16396 13780 16448
rect 15200 16532 15252 16584
rect 16028 16532 16080 16584
rect 16488 16600 16540 16652
rect 16948 16643 17000 16652
rect 16948 16609 16957 16643
rect 16957 16609 16991 16643
rect 16991 16609 17000 16643
rect 16948 16600 17000 16609
rect 18972 16779 19024 16788
rect 18972 16745 18981 16779
rect 18981 16745 19015 16779
rect 19015 16745 19024 16779
rect 18972 16736 19024 16745
rect 17960 16600 18012 16652
rect 16396 16575 16448 16584
rect 16396 16541 16405 16575
rect 16405 16541 16439 16575
rect 16439 16541 16448 16575
rect 16396 16532 16448 16541
rect 18604 16600 18656 16652
rect 18696 16532 18748 16584
rect 15016 16396 15068 16448
rect 15752 16439 15804 16448
rect 15752 16405 15761 16439
rect 15761 16405 15795 16439
rect 15795 16405 15804 16439
rect 15752 16396 15804 16405
rect 16948 16396 17000 16448
rect 19064 16600 19116 16652
rect 19892 16643 19944 16652
rect 19892 16609 19901 16643
rect 19901 16609 19935 16643
rect 19935 16609 19944 16643
rect 19892 16600 19944 16609
rect 19340 16532 19392 16584
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 8208 16235 8260 16244
rect 8208 16201 8217 16235
rect 8217 16201 8251 16235
rect 8251 16201 8260 16235
rect 8208 16192 8260 16201
rect 8668 16056 8720 16108
rect 7564 15988 7616 16040
rect 9772 16192 9824 16244
rect 11704 16192 11756 16244
rect 12348 16192 12400 16244
rect 13544 16192 13596 16244
rect 15016 16192 15068 16244
rect 15844 16124 15896 16176
rect 9404 16056 9456 16108
rect 10692 16056 10744 16108
rect 10968 16056 11020 16108
rect 11704 16099 11756 16108
rect 11704 16065 11713 16099
rect 11713 16065 11747 16099
rect 11747 16065 11756 16099
rect 11704 16056 11756 16065
rect 12440 16099 12492 16108
rect 12440 16065 12449 16099
rect 12449 16065 12483 16099
rect 12483 16065 12492 16099
rect 12440 16056 12492 16065
rect 13636 16056 13688 16108
rect 15752 16056 15804 16108
rect 16488 16192 16540 16244
rect 17776 16192 17828 16244
rect 16396 16056 16448 16108
rect 17776 16056 17828 16108
rect 18052 16099 18104 16108
rect 18052 16065 18061 16099
rect 18061 16065 18095 16099
rect 18095 16065 18104 16099
rect 18052 16056 18104 16065
rect 20352 16099 20404 16108
rect 20352 16065 20361 16099
rect 20361 16065 20395 16099
rect 20395 16065 20404 16099
rect 20352 16056 20404 16065
rect 8668 15920 8720 15972
rect 10600 15920 10652 15972
rect 10048 15852 10100 15904
rect 12716 15963 12768 15972
rect 12716 15929 12750 15963
rect 12750 15929 12768 15963
rect 12716 15920 12768 15929
rect 14004 15988 14056 16040
rect 15016 15920 15068 15972
rect 10968 15852 11020 15904
rect 11152 15895 11204 15904
rect 11152 15861 11161 15895
rect 11161 15861 11195 15895
rect 11195 15861 11204 15895
rect 11152 15852 11204 15861
rect 12532 15852 12584 15904
rect 13268 15852 13320 15904
rect 13820 15852 13872 15904
rect 15660 15852 15712 15904
rect 17040 15988 17092 16040
rect 19340 15920 19392 15972
rect 19616 15920 19668 15972
rect 20168 15963 20220 15972
rect 18696 15852 18748 15904
rect 19800 15895 19852 15904
rect 19800 15861 19809 15895
rect 19809 15861 19843 15895
rect 19843 15861 19852 15895
rect 19800 15852 19852 15861
rect 20168 15929 20177 15963
rect 20177 15929 20211 15963
rect 20211 15929 20220 15963
rect 20168 15920 20220 15929
rect 20904 15920 20956 15972
rect 20076 15852 20128 15904
rect 20996 15895 21048 15904
rect 20996 15861 21005 15895
rect 21005 15861 21039 15895
rect 21039 15861 21048 15895
rect 20996 15852 21048 15861
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 9036 15648 9088 15700
rect 9680 15648 9732 15700
rect 11060 15648 11112 15700
rect 12992 15691 13044 15700
rect 12992 15657 13001 15691
rect 13001 15657 13035 15691
rect 13035 15657 13044 15691
rect 12992 15648 13044 15657
rect 15200 15648 15252 15700
rect 15660 15691 15712 15700
rect 15660 15657 15669 15691
rect 15669 15657 15703 15691
rect 15703 15657 15712 15691
rect 15660 15648 15712 15657
rect 17776 15691 17828 15700
rect 17776 15657 17785 15691
rect 17785 15657 17819 15691
rect 17819 15657 17828 15691
rect 17776 15648 17828 15657
rect 10968 15580 11020 15632
rect 12440 15580 12492 15632
rect 13728 15580 13780 15632
rect 14004 15580 14056 15632
rect 7564 15512 7616 15564
rect 9680 15555 9732 15564
rect 8116 15444 8168 15496
rect 9036 15487 9088 15496
rect 9036 15453 9045 15487
rect 9045 15453 9079 15487
rect 9079 15453 9088 15487
rect 9036 15444 9088 15453
rect 7472 15351 7524 15360
rect 7472 15317 7481 15351
rect 7481 15317 7515 15351
rect 7515 15317 7524 15351
rect 7472 15308 7524 15317
rect 8852 15308 8904 15360
rect 9680 15521 9689 15555
rect 9689 15521 9723 15555
rect 9723 15521 9732 15555
rect 9680 15512 9732 15521
rect 14556 15555 14608 15564
rect 10968 15487 11020 15496
rect 10968 15453 10977 15487
rect 10977 15453 11011 15487
rect 11011 15453 11020 15487
rect 10968 15444 11020 15453
rect 14556 15521 14565 15555
rect 14565 15521 14599 15555
rect 14599 15521 14608 15555
rect 14556 15512 14608 15521
rect 15568 15580 15620 15632
rect 16120 15580 16172 15632
rect 18696 15580 18748 15632
rect 19248 15648 19300 15700
rect 20168 15580 20220 15632
rect 12348 15487 12400 15496
rect 12348 15453 12357 15487
rect 12357 15453 12391 15487
rect 12391 15453 12400 15487
rect 12348 15444 12400 15453
rect 13084 15444 13136 15496
rect 13544 15487 13596 15496
rect 13544 15453 13553 15487
rect 13553 15453 13587 15487
rect 13587 15453 13596 15487
rect 13544 15444 13596 15453
rect 15016 15444 15068 15496
rect 16488 15512 16540 15564
rect 17500 15512 17552 15564
rect 19892 15512 19944 15564
rect 20812 15512 20864 15564
rect 15568 15444 15620 15496
rect 15844 15487 15896 15496
rect 15844 15453 15853 15487
rect 15853 15453 15887 15487
rect 15887 15453 15896 15487
rect 15844 15444 15896 15453
rect 18144 15444 18196 15496
rect 11704 15308 11756 15360
rect 12808 15308 12860 15360
rect 13912 15308 13964 15360
rect 15292 15351 15344 15360
rect 15292 15317 15301 15351
rect 15301 15317 15335 15351
rect 15335 15317 15344 15351
rect 15292 15308 15344 15317
rect 19156 15308 19208 15360
rect 19432 15308 19484 15360
rect 20352 15308 20404 15360
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 8116 15104 8168 15156
rect 8208 15104 8260 15156
rect 6184 15011 6236 15020
rect 6184 14977 6193 15011
rect 6193 14977 6227 15011
rect 6227 14977 6236 15011
rect 6184 14968 6236 14977
rect 7472 15036 7524 15088
rect 8668 15104 8720 15156
rect 10968 15104 11020 15156
rect 12348 15104 12400 15156
rect 12716 15104 12768 15156
rect 13636 15104 13688 15156
rect 15016 15104 15068 15156
rect 15476 15104 15528 15156
rect 15936 15104 15988 15156
rect 19524 15104 19576 15156
rect 21180 15104 21232 15156
rect 9036 14968 9088 15020
rect 10600 14968 10652 15020
rect 5540 14900 5592 14952
rect 6092 14943 6144 14952
rect 6092 14909 6101 14943
rect 6101 14909 6135 14943
rect 6135 14909 6144 14943
rect 6092 14900 6144 14909
rect 7564 14900 7616 14952
rect 10784 14900 10836 14952
rect 17960 15036 18012 15088
rect 11888 14968 11940 15020
rect 11980 15011 12032 15020
rect 11980 14977 11989 15011
rect 11989 14977 12023 15011
rect 12023 14977 12032 15011
rect 11980 14968 12032 14977
rect 14004 14900 14056 14952
rect 17316 15011 17368 15020
rect 17316 14977 17325 15011
rect 17325 14977 17359 15011
rect 17359 14977 17368 15011
rect 17316 14968 17368 14977
rect 18604 14968 18656 15020
rect 18972 14968 19024 15020
rect 8760 14832 8812 14884
rect 11888 14832 11940 14884
rect 13084 14832 13136 14884
rect 15844 14900 15896 14952
rect 16212 14943 16264 14952
rect 16212 14909 16221 14943
rect 16221 14909 16255 14943
rect 16255 14909 16264 14943
rect 16212 14900 16264 14909
rect 9128 14807 9180 14816
rect 9128 14773 9137 14807
rect 9137 14773 9171 14807
rect 9171 14773 9180 14807
rect 9128 14764 9180 14773
rect 9588 14807 9640 14816
rect 9588 14773 9597 14807
rect 9597 14773 9631 14807
rect 9631 14773 9640 14807
rect 9588 14764 9640 14773
rect 11152 14764 11204 14816
rect 12624 14764 12676 14816
rect 15660 14832 15712 14884
rect 18880 14832 18932 14884
rect 16764 14807 16816 14816
rect 16764 14773 16773 14807
rect 16773 14773 16807 14807
rect 16807 14773 16816 14807
rect 16764 14764 16816 14773
rect 17224 14807 17276 14816
rect 17224 14773 17233 14807
rect 17233 14773 17267 14807
rect 17267 14773 17276 14807
rect 17224 14764 17276 14773
rect 18696 14764 18748 14816
rect 20720 14900 20772 14952
rect 19432 14875 19484 14884
rect 19432 14841 19466 14875
rect 19466 14841 19484 14875
rect 19432 14832 19484 14841
rect 19892 14764 19944 14816
rect 20168 14764 20220 14816
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 9128 14560 9180 14612
rect 9496 14560 9548 14612
rect 7472 14492 7524 14544
rect 8852 14535 8904 14544
rect 8852 14501 8861 14535
rect 8861 14501 8895 14535
rect 8895 14501 8904 14535
rect 8852 14492 8904 14501
rect 9404 14424 9456 14476
rect 12624 14560 12676 14612
rect 12808 14560 12860 14612
rect 19248 14603 19300 14612
rect 8668 14356 8720 14408
rect 14096 14492 14148 14544
rect 15660 14492 15712 14544
rect 11980 14467 12032 14476
rect 11980 14433 12014 14467
rect 12014 14433 12032 14467
rect 11980 14424 12032 14433
rect 13452 14424 13504 14476
rect 14372 14467 14424 14476
rect 14372 14433 14381 14467
rect 14381 14433 14415 14467
rect 14415 14433 14424 14467
rect 14372 14424 14424 14433
rect 15292 14467 15344 14476
rect 15292 14433 15301 14467
rect 15301 14433 15335 14467
rect 15335 14433 15344 14467
rect 15292 14424 15344 14433
rect 16212 14424 16264 14476
rect 17316 14492 17368 14544
rect 19248 14569 19257 14603
rect 19257 14569 19291 14603
rect 19291 14569 19300 14603
rect 19248 14560 19300 14569
rect 19800 14560 19852 14612
rect 16672 14424 16724 14476
rect 17960 14424 18012 14476
rect 18512 14424 18564 14476
rect 9036 14288 9088 14340
rect 13636 14356 13688 14408
rect 14096 14356 14148 14408
rect 14280 14356 14332 14408
rect 16028 14356 16080 14408
rect 17316 14356 17368 14408
rect 19156 14424 19208 14476
rect 19800 14424 19852 14476
rect 20168 14399 20220 14408
rect 20168 14365 20177 14399
rect 20177 14365 20211 14399
rect 20211 14365 20220 14399
rect 20168 14356 20220 14365
rect 20352 14356 20404 14408
rect 17684 14288 17736 14340
rect 19340 14288 19392 14340
rect 20444 14288 20496 14340
rect 9680 14220 9732 14272
rect 11060 14263 11112 14272
rect 11060 14229 11069 14263
rect 11069 14229 11103 14263
rect 11103 14229 11112 14263
rect 11060 14220 11112 14229
rect 13084 14263 13136 14272
rect 13084 14229 13093 14263
rect 13093 14229 13127 14263
rect 13127 14229 13136 14263
rect 13084 14220 13136 14229
rect 13176 14220 13228 14272
rect 14004 14220 14056 14272
rect 15384 14220 15436 14272
rect 17500 14263 17552 14272
rect 17500 14229 17509 14263
rect 17509 14229 17543 14263
rect 17543 14229 17552 14263
rect 17500 14220 17552 14229
rect 17776 14263 17828 14272
rect 17776 14229 17785 14263
rect 17785 14229 17819 14263
rect 17819 14229 17828 14263
rect 17776 14220 17828 14229
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 6092 14016 6144 14068
rect 12440 14059 12492 14068
rect 12440 14025 12449 14059
rect 12449 14025 12483 14059
rect 12483 14025 12492 14059
rect 12440 14016 12492 14025
rect 15292 14016 15344 14068
rect 13084 13948 13136 14000
rect 8760 13923 8812 13932
rect 8760 13889 8769 13923
rect 8769 13889 8803 13923
rect 8803 13889 8812 13923
rect 8760 13880 8812 13889
rect 9404 13880 9456 13932
rect 10692 13880 10744 13932
rect 11520 13880 11572 13932
rect 11060 13812 11112 13864
rect 11980 13880 12032 13932
rect 13912 13923 13964 13932
rect 12532 13812 12584 13864
rect 12900 13812 12952 13864
rect 13912 13889 13921 13923
rect 13921 13889 13955 13923
rect 13955 13889 13964 13923
rect 13912 13880 13964 13889
rect 15384 13948 15436 14000
rect 16212 13948 16264 14000
rect 17316 14016 17368 14068
rect 17960 14016 18012 14068
rect 18604 14016 18656 14068
rect 19800 14059 19852 14068
rect 19800 14025 19809 14059
rect 19809 14025 19843 14059
rect 19843 14025 19852 14059
rect 19800 14016 19852 14025
rect 20628 14016 20680 14068
rect 17592 13948 17644 14000
rect 15016 13923 15068 13932
rect 15016 13889 15025 13923
rect 15025 13889 15059 13923
rect 15059 13889 15068 13923
rect 15016 13880 15068 13889
rect 15660 13855 15712 13864
rect 15660 13821 15669 13855
rect 15669 13821 15703 13855
rect 15703 13821 15712 13855
rect 15660 13812 15712 13821
rect 16212 13812 16264 13864
rect 17316 13880 17368 13932
rect 18052 13880 18104 13932
rect 18420 13880 18472 13932
rect 19432 13880 19484 13932
rect 19064 13855 19116 13864
rect 19064 13821 19073 13855
rect 19073 13821 19107 13855
rect 19107 13821 19116 13855
rect 19064 13812 19116 13821
rect 19340 13812 19392 13864
rect 19800 13812 19852 13864
rect 20812 13855 20864 13864
rect 20812 13821 20821 13855
rect 20821 13821 20855 13855
rect 20855 13821 20864 13855
rect 20812 13812 20864 13821
rect 1400 13744 1452 13796
rect 10876 13719 10928 13728
rect 10876 13685 10885 13719
rect 10885 13685 10919 13719
rect 10919 13685 10928 13719
rect 10876 13676 10928 13685
rect 11152 13719 11204 13728
rect 11152 13685 11161 13719
rect 11161 13685 11195 13719
rect 11195 13685 11204 13719
rect 11152 13676 11204 13685
rect 11704 13676 11756 13728
rect 13084 13676 13136 13728
rect 13452 13719 13504 13728
rect 13452 13685 13461 13719
rect 13461 13685 13495 13719
rect 13495 13685 13504 13719
rect 13452 13676 13504 13685
rect 14556 13676 14608 13728
rect 18328 13744 18380 13796
rect 18604 13744 18656 13796
rect 20352 13744 20404 13796
rect 17684 13676 17736 13728
rect 19248 13676 19300 13728
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 9404 13472 9456 13524
rect 11152 13472 11204 13524
rect 12624 13472 12676 13524
rect 14372 13472 14424 13524
rect 16396 13472 16448 13524
rect 10508 13404 10560 13456
rect 12716 13404 12768 13456
rect 9496 13379 9548 13388
rect 9496 13345 9505 13379
rect 9505 13345 9539 13379
rect 9539 13345 9548 13379
rect 9496 13336 9548 13345
rect 10232 13379 10284 13388
rect 10232 13345 10241 13379
rect 10241 13345 10275 13379
rect 10275 13345 10284 13379
rect 10232 13336 10284 13345
rect 11612 13336 11664 13388
rect 9496 13200 9548 13252
rect 10876 13268 10928 13320
rect 12440 13336 12492 13388
rect 15568 13404 15620 13456
rect 15752 13447 15804 13456
rect 15752 13413 15761 13447
rect 15761 13413 15795 13447
rect 15795 13413 15804 13447
rect 15752 13404 15804 13413
rect 16764 13472 16816 13524
rect 17776 13472 17828 13524
rect 18512 13472 18564 13524
rect 18604 13472 18656 13524
rect 18880 13515 18932 13524
rect 18880 13481 18889 13515
rect 18889 13481 18923 13515
rect 18923 13481 18932 13515
rect 18880 13472 18932 13481
rect 19524 13472 19576 13524
rect 17960 13404 18012 13456
rect 13176 13379 13228 13388
rect 13176 13345 13185 13379
rect 13185 13345 13219 13379
rect 13219 13345 13228 13379
rect 13176 13336 13228 13345
rect 14188 13336 14240 13388
rect 14924 13336 14976 13388
rect 15200 13336 15252 13388
rect 16028 13336 16080 13388
rect 17776 13336 17828 13388
rect 18604 13336 18656 13388
rect 12256 13268 12308 13320
rect 14464 13268 14516 13320
rect 12532 13132 12584 13184
rect 13728 13132 13780 13184
rect 14372 13132 14424 13184
rect 16764 13268 16816 13320
rect 17224 13268 17276 13320
rect 17500 13268 17552 13320
rect 17684 13311 17736 13320
rect 17684 13277 17693 13311
rect 17693 13277 17727 13311
rect 17727 13277 17736 13311
rect 17684 13268 17736 13277
rect 18512 13311 18564 13320
rect 18512 13277 18521 13311
rect 18521 13277 18555 13311
rect 18555 13277 18564 13311
rect 18512 13268 18564 13277
rect 19984 13311 20036 13320
rect 19984 13277 19993 13311
rect 19993 13277 20027 13311
rect 20027 13277 20036 13311
rect 19984 13268 20036 13277
rect 19064 13200 19116 13252
rect 15844 13132 15896 13184
rect 15936 13132 15988 13184
rect 20444 13132 20496 13184
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 9404 12928 9456 12980
rect 10232 12928 10284 12980
rect 12440 12971 12492 12980
rect 12440 12937 12449 12971
rect 12449 12937 12483 12971
rect 12483 12937 12492 12971
rect 12440 12928 12492 12937
rect 12072 12860 12124 12912
rect 16120 12928 16172 12980
rect 16396 12928 16448 12980
rect 16764 12971 16816 12980
rect 16764 12937 16773 12971
rect 16773 12937 16807 12971
rect 16807 12937 16816 12971
rect 16764 12928 16816 12937
rect 8760 12835 8812 12844
rect 8760 12801 8769 12835
rect 8769 12801 8803 12835
rect 8803 12801 8812 12835
rect 8760 12792 8812 12801
rect 12992 12835 13044 12844
rect 10876 12724 10928 12776
rect 12992 12801 13001 12835
rect 13001 12801 13035 12835
rect 13035 12801 13044 12835
rect 12992 12792 13044 12801
rect 16764 12792 16816 12844
rect 17132 12792 17184 12844
rect 18788 12860 18840 12912
rect 13084 12724 13136 12776
rect 15200 12724 15252 12776
rect 12440 12656 12492 12708
rect 14372 12656 14424 12708
rect 9496 12588 9548 12640
rect 11060 12588 11112 12640
rect 12900 12631 12952 12640
rect 12900 12597 12909 12631
rect 12909 12597 12943 12631
rect 12943 12597 12952 12631
rect 12900 12588 12952 12597
rect 16212 12724 16264 12776
rect 16948 12724 17000 12776
rect 17592 12724 17644 12776
rect 15016 12588 15068 12640
rect 16672 12588 16724 12640
rect 17224 12588 17276 12640
rect 18420 12724 18472 12776
rect 18880 12724 18932 12776
rect 19984 12724 20036 12776
rect 20444 12767 20496 12776
rect 20444 12733 20453 12767
rect 20453 12733 20487 12767
rect 20487 12733 20496 12767
rect 20444 12724 20496 12733
rect 18512 12588 18564 12640
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 9496 12316 9548 12368
rect 9588 12316 9640 12368
rect 12992 12384 13044 12436
rect 14372 12427 14424 12436
rect 14372 12393 14381 12427
rect 14381 12393 14415 12427
rect 14415 12393 14424 12427
rect 14372 12384 14424 12393
rect 14556 12384 14608 12436
rect 9680 12291 9732 12300
rect 9680 12257 9689 12291
rect 9689 12257 9723 12291
rect 9723 12257 9732 12291
rect 9680 12248 9732 12257
rect 8760 12180 8812 12232
rect 12072 12248 12124 12300
rect 9128 12087 9180 12096
rect 9128 12053 9137 12087
rect 9137 12053 9171 12087
rect 9171 12053 9180 12087
rect 9128 12044 9180 12053
rect 10968 12180 11020 12232
rect 14740 12316 14792 12368
rect 17408 12384 17460 12436
rect 18512 12384 18564 12436
rect 16120 12359 16172 12368
rect 16120 12325 16154 12359
rect 16154 12325 16172 12359
rect 16120 12316 16172 12325
rect 12992 12291 13044 12300
rect 12992 12257 13001 12291
rect 13001 12257 13035 12291
rect 13035 12257 13044 12291
rect 12992 12248 13044 12257
rect 16580 12316 16632 12368
rect 18880 12384 18932 12436
rect 19984 12427 20036 12436
rect 19984 12393 19993 12427
rect 19993 12393 20027 12427
rect 20027 12393 20036 12427
rect 19984 12384 20036 12393
rect 20352 12384 20404 12436
rect 15292 12223 15344 12232
rect 15292 12189 15301 12223
rect 15301 12189 15335 12223
rect 15335 12189 15344 12223
rect 15292 12180 15344 12189
rect 15752 12180 15804 12232
rect 18052 12223 18104 12232
rect 18052 12189 18061 12223
rect 18061 12189 18095 12223
rect 18095 12189 18104 12223
rect 18052 12180 18104 12189
rect 18880 12291 18932 12300
rect 18880 12257 18914 12291
rect 18914 12257 18932 12291
rect 18880 12248 18932 12257
rect 19432 12248 19484 12300
rect 17960 12112 18012 12164
rect 15752 12044 15804 12096
rect 17224 12087 17276 12096
rect 17224 12053 17233 12087
rect 17233 12053 17267 12087
rect 17267 12053 17276 12087
rect 17224 12044 17276 12053
rect 18880 12044 18932 12096
rect 19708 12044 19760 12096
rect 20352 12044 20404 12096
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 12440 11840 12492 11892
rect 12900 11840 12952 11892
rect 14924 11840 14976 11892
rect 15568 11883 15620 11892
rect 15568 11849 15577 11883
rect 15577 11849 15611 11883
rect 15611 11849 15620 11883
rect 15568 11840 15620 11849
rect 15752 11840 15804 11892
rect 12072 11747 12124 11756
rect 12072 11713 12081 11747
rect 12081 11713 12115 11747
rect 12115 11713 12124 11747
rect 12072 11704 12124 11713
rect 14372 11704 14424 11756
rect 15660 11704 15712 11756
rect 15936 11704 15988 11756
rect 17224 11772 17276 11824
rect 16212 11747 16264 11756
rect 16212 11713 16221 11747
rect 16221 11713 16255 11747
rect 16255 11713 16264 11747
rect 16212 11704 16264 11713
rect 17684 11704 17736 11756
rect 19156 11840 19208 11892
rect 18880 11772 18932 11824
rect 8760 11636 8812 11688
rect 8944 11636 8996 11688
rect 9588 11636 9640 11688
rect 9956 11636 10008 11688
rect 10876 11636 10928 11688
rect 14464 11636 14516 11688
rect 19616 11636 19668 11688
rect 20812 11636 20864 11688
rect 9128 11568 9180 11620
rect 12716 11568 12768 11620
rect 14924 11568 14976 11620
rect 16580 11568 16632 11620
rect 17500 11568 17552 11620
rect 18972 11568 19024 11620
rect 19984 11611 20036 11620
rect 19984 11577 20018 11611
rect 20018 11577 20036 11611
rect 19984 11568 20036 11577
rect 9496 11500 9548 11552
rect 10048 11500 10100 11552
rect 12440 11500 12492 11552
rect 12992 11543 13044 11552
rect 12992 11509 13001 11543
rect 13001 11509 13035 11543
rect 13035 11509 13044 11543
rect 12992 11500 13044 11509
rect 14464 11500 14516 11552
rect 14556 11500 14608 11552
rect 15476 11500 15528 11552
rect 15752 11500 15804 11552
rect 16488 11500 16540 11552
rect 16948 11543 17000 11552
rect 16948 11509 16957 11543
rect 16957 11509 16991 11543
rect 16991 11509 17000 11543
rect 16948 11500 17000 11509
rect 17316 11543 17368 11552
rect 17316 11509 17325 11543
rect 17325 11509 17359 11543
rect 17359 11509 17368 11543
rect 17316 11500 17368 11509
rect 18788 11500 18840 11552
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 9680 11339 9732 11348
rect 9680 11305 9689 11339
rect 9689 11305 9723 11339
rect 9723 11305 9732 11339
rect 9680 11296 9732 11305
rect 10048 11339 10100 11348
rect 10048 11305 10057 11339
rect 10057 11305 10091 11339
rect 10091 11305 10100 11339
rect 10048 11296 10100 11305
rect 12072 11296 12124 11348
rect 14188 11339 14240 11348
rect 14188 11305 14197 11339
rect 14197 11305 14231 11339
rect 14231 11305 14240 11339
rect 14188 11296 14240 11305
rect 17316 11296 17368 11348
rect 9036 11228 9088 11280
rect 9220 11160 9272 11212
rect 12164 11228 12216 11280
rect 9496 11160 9548 11212
rect 10968 11203 11020 11212
rect 9128 11135 9180 11144
rect 9128 11101 9137 11135
rect 9137 11101 9171 11135
rect 9171 11101 9180 11135
rect 10968 11169 10977 11203
rect 10977 11169 11011 11203
rect 11011 11169 11020 11203
rect 10968 11160 11020 11169
rect 11796 11160 11848 11212
rect 9128 11092 9180 11101
rect 15752 11160 15804 11212
rect 17224 11228 17276 11280
rect 18420 11228 18472 11280
rect 19248 11296 19300 11348
rect 19064 11228 19116 11280
rect 17408 11160 17460 11212
rect 17960 11160 18012 11212
rect 18604 11203 18656 11212
rect 18604 11169 18613 11203
rect 18613 11169 18647 11203
rect 18647 11169 18656 11203
rect 18604 11160 18656 11169
rect 20904 11160 20956 11212
rect 14464 11024 14516 11076
rect 15752 11024 15804 11076
rect 13728 10956 13780 11008
rect 14372 10956 14424 11008
rect 16396 11092 16448 11144
rect 16488 11024 16540 11076
rect 17684 11024 17736 11076
rect 20076 11135 20128 11144
rect 20076 11101 20085 11135
rect 20085 11101 20119 11135
rect 20119 11101 20128 11135
rect 20076 11092 20128 11101
rect 18052 11024 18104 11076
rect 20536 11024 20588 11076
rect 19340 10956 19392 11008
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 12440 10795 12492 10804
rect 12440 10761 12449 10795
rect 12449 10761 12483 10795
rect 12483 10761 12492 10795
rect 12440 10752 12492 10761
rect 12992 10752 13044 10804
rect 12716 10684 12768 10736
rect 11796 10616 11848 10668
rect 9496 10548 9548 10600
rect 9680 10591 9732 10600
rect 9680 10557 9689 10591
rect 9689 10557 9723 10591
rect 9723 10557 9732 10591
rect 9680 10548 9732 10557
rect 11612 10548 11664 10600
rect 12440 10548 12492 10600
rect 12716 10548 12768 10600
rect 14004 10684 14056 10736
rect 14372 10752 14424 10804
rect 15108 10752 15160 10804
rect 15384 10795 15436 10804
rect 15384 10761 15393 10795
rect 15393 10761 15427 10795
rect 15427 10761 15436 10795
rect 15384 10752 15436 10761
rect 15108 10659 15160 10668
rect 15108 10625 15117 10659
rect 15117 10625 15151 10659
rect 15151 10625 15160 10659
rect 15108 10616 15160 10625
rect 15844 10659 15896 10668
rect 15844 10625 15853 10659
rect 15853 10625 15887 10659
rect 15887 10625 15896 10659
rect 15844 10616 15896 10625
rect 16212 10616 16264 10668
rect 13728 10548 13780 10600
rect 14464 10548 14516 10600
rect 14556 10548 14608 10600
rect 15292 10548 15344 10600
rect 16120 10548 16172 10600
rect 16488 10752 16540 10804
rect 18512 10752 18564 10804
rect 17592 10684 17644 10736
rect 18328 10684 18380 10736
rect 17684 10616 17736 10668
rect 18604 10616 18656 10668
rect 19340 10548 19392 10600
rect 8208 10480 8260 10532
rect 9220 10412 9272 10464
rect 10692 10412 10744 10464
rect 10876 10412 10928 10464
rect 12624 10412 12676 10464
rect 12808 10455 12860 10464
rect 12808 10421 12817 10455
rect 12817 10421 12851 10455
rect 12851 10421 12860 10455
rect 12808 10412 12860 10421
rect 14004 10412 14056 10464
rect 16396 10480 16448 10532
rect 19432 10480 19484 10532
rect 19616 10591 19668 10600
rect 19616 10557 19625 10591
rect 19625 10557 19659 10591
rect 19659 10557 19668 10591
rect 19616 10548 19668 10557
rect 20444 10480 20496 10532
rect 18052 10412 18104 10464
rect 19064 10455 19116 10464
rect 19064 10421 19073 10455
rect 19073 10421 19107 10455
rect 19107 10421 19116 10455
rect 19064 10412 19116 10421
rect 19340 10412 19392 10464
rect 19984 10412 20036 10464
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 9680 10251 9732 10260
rect 9680 10217 9689 10251
rect 9689 10217 9723 10251
rect 9723 10217 9732 10251
rect 9680 10208 9732 10217
rect 11796 10208 11848 10260
rect 9956 10140 10008 10192
rect 10784 10140 10836 10192
rect 11152 10140 11204 10192
rect 11888 10140 11940 10192
rect 14004 10140 14056 10192
rect 14280 10140 14332 10192
rect 15016 10140 15068 10192
rect 12348 10115 12400 10124
rect 12348 10081 12357 10115
rect 12357 10081 12391 10115
rect 12391 10081 12400 10115
rect 12348 10072 12400 10081
rect 15568 10072 15620 10124
rect 16948 10208 17000 10260
rect 19064 10208 19116 10260
rect 20444 10251 20496 10260
rect 20444 10217 20453 10251
rect 20453 10217 20487 10251
rect 20487 10217 20496 10251
rect 20444 10208 20496 10217
rect 20904 10251 20956 10260
rect 20904 10217 20913 10251
rect 20913 10217 20947 10251
rect 20947 10217 20956 10251
rect 20904 10208 20956 10217
rect 17040 10140 17092 10192
rect 17960 10140 18012 10192
rect 10140 10047 10192 10056
rect 10140 10013 10149 10047
rect 10149 10013 10183 10047
rect 10183 10013 10192 10047
rect 10140 10004 10192 10013
rect 10692 10047 10744 10056
rect 9588 9936 9640 9988
rect 10692 10013 10701 10047
rect 10701 10013 10735 10047
rect 10735 10013 10744 10047
rect 10692 10004 10744 10013
rect 13728 10047 13780 10056
rect 13728 10013 13737 10047
rect 13737 10013 13771 10047
rect 13771 10013 13780 10047
rect 13728 10004 13780 10013
rect 14004 10004 14056 10056
rect 15108 10004 15160 10056
rect 12440 9936 12492 9988
rect 14924 9936 14976 9988
rect 16764 10072 16816 10124
rect 16212 10004 16264 10056
rect 16488 10004 16540 10056
rect 17960 10004 18012 10056
rect 18512 10047 18564 10056
rect 18512 10013 18521 10047
rect 18521 10013 18555 10047
rect 18555 10013 18564 10047
rect 18512 10004 18564 10013
rect 20076 10140 20128 10192
rect 19616 10072 19668 10124
rect 19064 10047 19116 10056
rect 19064 10013 19073 10047
rect 19073 10013 19107 10047
rect 19107 10013 19116 10047
rect 19064 10004 19116 10013
rect 16304 9936 16356 9988
rect 18604 9936 18656 9988
rect 12992 9868 13044 9920
rect 14372 9868 14424 9920
rect 17592 9868 17644 9920
rect 19248 9868 19300 9920
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 9312 9664 9364 9716
rect 14372 9664 14424 9716
rect 11152 9596 11204 9648
rect 11888 9596 11940 9648
rect 15752 9664 15804 9716
rect 16764 9664 16816 9716
rect 15568 9596 15620 9648
rect 16212 9596 16264 9648
rect 15844 9528 15896 9580
rect 8208 9503 8260 9512
rect 8208 9469 8217 9503
rect 8217 9469 8251 9503
rect 8251 9469 8260 9503
rect 8208 9460 8260 9469
rect 9220 9460 9272 9512
rect 9680 9460 9732 9512
rect 10692 9460 10744 9512
rect 12440 9503 12492 9512
rect 12440 9469 12449 9503
rect 12449 9469 12483 9503
rect 12483 9469 12492 9503
rect 12440 9460 12492 9469
rect 14004 9460 14056 9512
rect 14188 9460 14240 9512
rect 16120 9460 16172 9512
rect 16488 9528 16540 9580
rect 19064 9664 19116 9716
rect 20168 9664 20220 9716
rect 20812 9664 20864 9716
rect 20536 9571 20588 9580
rect 20536 9537 20545 9571
rect 20545 9537 20579 9571
rect 20579 9537 20588 9571
rect 20536 9528 20588 9537
rect 20628 9571 20680 9580
rect 20628 9537 20637 9571
rect 20637 9537 20671 9571
rect 20671 9537 20680 9571
rect 20628 9528 20680 9537
rect 18144 9460 18196 9512
rect 10324 9435 10376 9444
rect 10324 9401 10358 9435
rect 10358 9401 10376 9435
rect 10324 9392 10376 9401
rect 14924 9392 14976 9444
rect 15292 9392 15344 9444
rect 15476 9392 15528 9444
rect 16396 9392 16448 9444
rect 17960 9392 18012 9444
rect 20904 9392 20956 9444
rect 9588 9367 9640 9376
rect 9588 9333 9597 9367
rect 9597 9333 9631 9367
rect 9631 9333 9640 9367
rect 9588 9324 9640 9333
rect 11704 9367 11756 9376
rect 11704 9333 11713 9367
rect 11713 9333 11747 9367
rect 11747 9333 11756 9367
rect 11704 9324 11756 9333
rect 13728 9324 13780 9376
rect 14004 9324 14056 9376
rect 15108 9324 15160 9376
rect 16304 9324 16356 9376
rect 19432 9367 19484 9376
rect 19432 9333 19441 9367
rect 19441 9333 19475 9367
rect 19475 9333 19484 9367
rect 19432 9324 19484 9333
rect 19524 9324 19576 9376
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 10140 9120 10192 9172
rect 10324 9120 10376 9172
rect 10968 9120 11020 9172
rect 12348 9120 12400 9172
rect 16488 9120 16540 9172
rect 18512 9120 18564 9172
rect 19984 9163 20036 9172
rect 19984 9129 19993 9163
rect 19993 9129 20027 9163
rect 20027 9129 20036 9163
rect 19984 9120 20036 9129
rect 12532 9052 12584 9104
rect 13728 9052 13780 9104
rect 16304 9052 16356 9104
rect 6920 8984 6972 9036
rect 9680 9027 9732 9036
rect 9680 8993 9689 9027
rect 9689 8993 9723 9027
rect 9723 8993 9732 9027
rect 9680 8984 9732 8993
rect 10508 8984 10560 9036
rect 10876 8984 10928 9036
rect 11980 8984 12032 9036
rect 12348 8984 12400 9036
rect 12440 8984 12492 9036
rect 15752 9027 15804 9036
rect 15752 8993 15761 9027
rect 15761 8993 15795 9027
rect 15795 8993 15804 9027
rect 15752 8984 15804 8993
rect 16948 8984 17000 9036
rect 18144 9052 18196 9104
rect 18328 8984 18380 9036
rect 9220 8959 9272 8968
rect 9220 8925 9229 8959
rect 9229 8925 9263 8959
rect 9263 8925 9272 8959
rect 9220 8916 9272 8925
rect 11796 8959 11848 8968
rect 11796 8925 11805 8959
rect 11805 8925 11839 8959
rect 11839 8925 11848 8959
rect 11796 8916 11848 8925
rect 11888 8959 11940 8968
rect 11888 8925 11897 8959
rect 11897 8925 11931 8959
rect 11931 8925 11940 8959
rect 11888 8916 11940 8925
rect 19432 9052 19484 9104
rect 19156 8984 19208 9036
rect 8852 8780 8904 8832
rect 12900 8848 12952 8900
rect 11612 8780 11664 8832
rect 11888 8780 11940 8832
rect 11980 8780 12032 8832
rect 15660 8848 15712 8900
rect 18512 8848 18564 8900
rect 14372 8823 14424 8832
rect 14372 8789 14381 8823
rect 14381 8789 14415 8823
rect 14415 8789 14424 8823
rect 14372 8780 14424 8789
rect 14464 8780 14516 8832
rect 17960 8780 18012 8832
rect 18604 8780 18656 8832
rect 19984 8780 20036 8832
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 3424 8576 3476 8628
rect 10324 8576 10376 8628
rect 10508 8576 10560 8628
rect 10876 8619 10928 8628
rect 10876 8585 10885 8619
rect 10885 8585 10919 8619
rect 10919 8585 10928 8619
rect 10876 8576 10928 8585
rect 11888 8619 11940 8628
rect 11888 8585 11897 8619
rect 11897 8585 11931 8619
rect 11931 8585 11940 8619
rect 11888 8576 11940 8585
rect 16212 8576 16264 8628
rect 11612 8508 11664 8560
rect 12900 8508 12952 8560
rect 17224 8576 17276 8628
rect 18604 8576 18656 8628
rect 19616 8576 19668 8628
rect 19984 8576 20036 8628
rect 17040 8508 17092 8560
rect 18328 8508 18380 8560
rect 10968 8440 11020 8492
rect 12532 8440 12584 8492
rect 14372 8483 14424 8492
rect 14372 8449 14381 8483
rect 14381 8449 14415 8483
rect 14415 8449 14424 8483
rect 14372 8440 14424 8449
rect 15844 8440 15896 8492
rect 16304 8440 16356 8492
rect 16580 8440 16632 8492
rect 17408 8483 17460 8492
rect 17408 8449 17417 8483
rect 17417 8449 17451 8483
rect 17451 8449 17460 8483
rect 17408 8440 17460 8449
rect 19984 8440 20036 8492
rect 20628 8440 20680 8492
rect 9864 8372 9916 8424
rect 11704 8372 11756 8424
rect 14004 8372 14056 8424
rect 16488 8372 16540 8424
rect 9772 8304 9824 8356
rect 10692 8304 10744 8356
rect 11980 8304 12032 8356
rect 12808 8347 12860 8356
rect 12808 8313 12817 8347
rect 12817 8313 12851 8347
rect 12851 8313 12860 8347
rect 12808 8304 12860 8313
rect 13728 8304 13780 8356
rect 14280 8347 14332 8356
rect 14280 8313 14289 8347
rect 14289 8313 14323 8347
rect 14323 8313 14332 8347
rect 14280 8304 14332 8313
rect 16120 8347 16172 8356
rect 12900 8279 12952 8288
rect 12900 8245 12909 8279
rect 12909 8245 12943 8279
rect 12943 8245 12952 8279
rect 12900 8236 12952 8245
rect 13820 8279 13872 8288
rect 13820 8245 13829 8279
rect 13829 8245 13863 8279
rect 13863 8245 13872 8279
rect 13820 8236 13872 8245
rect 15568 8236 15620 8288
rect 16120 8313 16129 8347
rect 16129 8313 16163 8347
rect 16163 8313 16172 8347
rect 16120 8304 16172 8313
rect 16580 8304 16632 8356
rect 16764 8372 16816 8424
rect 18604 8304 18656 8356
rect 20076 8372 20128 8424
rect 17500 8236 17552 8288
rect 20076 8279 20128 8288
rect 20076 8245 20085 8279
rect 20085 8245 20119 8279
rect 20119 8245 20128 8279
rect 20076 8236 20128 8245
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 11796 8032 11848 8084
rect 12532 8032 12584 8084
rect 12900 8075 12952 8084
rect 12900 8041 12909 8075
rect 12909 8041 12943 8075
rect 12943 8041 12952 8075
rect 12900 8032 12952 8041
rect 13820 8032 13872 8084
rect 9956 7964 10008 8016
rect 10876 7964 10928 8016
rect 9680 7896 9732 7948
rect 10324 7896 10376 7948
rect 11336 7939 11388 7948
rect 11336 7905 11359 7939
rect 11359 7905 11388 7939
rect 11336 7896 11388 7905
rect 14464 8032 14516 8084
rect 16120 8032 16172 8084
rect 17040 8032 17092 8084
rect 18512 8032 18564 8084
rect 18788 8032 18840 8084
rect 19984 8032 20036 8084
rect 20904 8075 20956 8084
rect 20904 8041 20913 8075
rect 20913 8041 20947 8075
rect 20947 8041 20956 8075
rect 20904 8032 20956 8041
rect 14004 7964 14056 8016
rect 17960 7964 18012 8016
rect 20628 7964 20680 8016
rect 13912 7896 13964 7948
rect 15108 7896 15160 7948
rect 15292 7896 15344 7948
rect 16580 7896 16632 7948
rect 16856 7896 16908 7948
rect 17408 7896 17460 7948
rect 18604 7896 18656 7948
rect 19064 7896 19116 7948
rect 10508 7871 10560 7880
rect 10508 7837 10517 7871
rect 10517 7837 10551 7871
rect 10551 7837 10560 7871
rect 10508 7828 10560 7837
rect 10968 7828 11020 7880
rect 13452 7871 13504 7880
rect 13452 7837 13461 7871
rect 13461 7837 13495 7871
rect 13495 7837 13504 7871
rect 13452 7828 13504 7837
rect 14464 7871 14516 7880
rect 14464 7837 14473 7871
rect 14473 7837 14507 7871
rect 14507 7837 14516 7871
rect 14464 7828 14516 7837
rect 12072 7760 12124 7812
rect 16488 7760 16540 7812
rect 11796 7692 11848 7744
rect 13452 7692 13504 7744
rect 14004 7692 14056 7744
rect 16580 7692 16632 7744
rect 17500 7692 17552 7744
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 9772 7531 9824 7540
rect 9772 7497 9781 7531
rect 9781 7497 9815 7531
rect 9815 7497 9824 7531
rect 9772 7488 9824 7497
rect 10324 7531 10376 7540
rect 10324 7497 10333 7531
rect 10333 7497 10367 7531
rect 10367 7497 10376 7531
rect 10324 7488 10376 7497
rect 10508 7488 10560 7540
rect 12808 7531 12860 7540
rect 12808 7497 12817 7531
rect 12817 7497 12851 7531
rect 12851 7497 12860 7531
rect 12808 7488 12860 7497
rect 10600 7352 10652 7404
rect 13176 7352 13228 7404
rect 16488 7488 16540 7540
rect 16948 7531 17000 7540
rect 16948 7497 16957 7531
rect 16957 7497 16991 7531
rect 16991 7497 17000 7531
rect 16948 7488 17000 7497
rect 17408 7420 17460 7472
rect 18236 7420 18288 7472
rect 16672 7352 16724 7404
rect 18604 7395 18656 7404
rect 18604 7361 18613 7395
rect 18613 7361 18647 7395
rect 18647 7361 18656 7395
rect 18604 7352 18656 7361
rect 20444 7395 20496 7404
rect 20444 7361 20453 7395
rect 20453 7361 20487 7395
rect 20487 7361 20496 7395
rect 20444 7352 20496 7361
rect 8392 7327 8444 7336
rect 8392 7293 8401 7327
rect 8401 7293 8435 7327
rect 8435 7293 8444 7327
rect 8392 7284 8444 7293
rect 13728 7284 13780 7336
rect 9864 7216 9916 7268
rect 13452 7216 13504 7268
rect 9956 7148 10008 7200
rect 10876 7148 10928 7200
rect 12900 7148 12952 7200
rect 13176 7191 13228 7200
rect 13176 7157 13185 7191
rect 13185 7157 13219 7191
rect 13219 7157 13228 7191
rect 13176 7148 13228 7157
rect 13912 7148 13964 7200
rect 14464 7284 14516 7336
rect 15384 7148 15436 7200
rect 16580 7284 16632 7336
rect 18972 7284 19024 7336
rect 19892 7284 19944 7336
rect 15660 7216 15712 7268
rect 18788 7216 18840 7268
rect 20904 7216 20956 7268
rect 16304 7148 16356 7200
rect 18052 7191 18104 7200
rect 18052 7157 18061 7191
rect 18061 7157 18095 7191
rect 18095 7157 18104 7191
rect 18052 7148 18104 7157
rect 18512 7191 18564 7200
rect 18512 7157 18521 7191
rect 18521 7157 18555 7191
rect 18555 7157 18564 7191
rect 18512 7148 18564 7157
rect 19156 7148 19208 7200
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 9680 6987 9732 6996
rect 9680 6953 9689 6987
rect 9689 6953 9723 6987
rect 9723 6953 9732 6987
rect 9680 6944 9732 6953
rect 13176 6944 13228 6996
rect 13912 6987 13964 6996
rect 13912 6953 13921 6987
rect 13921 6953 13955 6987
rect 13955 6953 13964 6987
rect 13912 6944 13964 6953
rect 15660 6987 15712 6996
rect 9772 6876 9824 6928
rect 10048 6851 10100 6860
rect 10048 6817 10057 6851
rect 10057 6817 10091 6851
rect 10091 6817 10100 6851
rect 10048 6808 10100 6817
rect 9128 6783 9180 6792
rect 9128 6749 9137 6783
rect 9137 6749 9171 6783
rect 9171 6749 9180 6783
rect 9128 6740 9180 6749
rect 9772 6740 9824 6792
rect 14372 6876 14424 6928
rect 15660 6953 15669 6987
rect 15669 6953 15703 6987
rect 15703 6953 15712 6987
rect 15660 6944 15712 6953
rect 15936 6944 15988 6996
rect 16120 6944 16172 6996
rect 16304 6987 16356 6996
rect 16304 6953 16313 6987
rect 16313 6953 16347 6987
rect 16347 6953 16356 6987
rect 16304 6944 16356 6953
rect 18236 6987 18288 6996
rect 18236 6953 18245 6987
rect 18245 6953 18279 6987
rect 18279 6953 18288 6987
rect 18236 6944 18288 6953
rect 20628 6944 20680 6996
rect 10968 6808 11020 6860
rect 12532 6808 12584 6860
rect 13728 6808 13780 6860
rect 14832 6808 14884 6860
rect 15936 6808 15988 6860
rect 16212 6808 16264 6860
rect 18052 6876 18104 6928
rect 17592 6808 17644 6860
rect 19432 6851 19484 6860
rect 19432 6817 19466 6851
rect 19466 6817 19484 6851
rect 19432 6808 19484 6817
rect 11796 6783 11848 6792
rect 10508 6604 10560 6656
rect 11796 6749 11805 6783
rect 11805 6749 11839 6783
rect 11839 6749 11848 6783
rect 11796 6740 11848 6749
rect 13820 6740 13872 6792
rect 14464 6783 14516 6792
rect 14464 6749 14473 6783
rect 14473 6749 14507 6783
rect 14507 6749 14516 6783
rect 15844 6783 15896 6792
rect 14464 6740 14516 6749
rect 15844 6749 15853 6783
rect 15853 6749 15887 6783
rect 15887 6749 15896 6783
rect 15844 6740 15896 6749
rect 17500 6783 17552 6792
rect 17500 6749 17509 6783
rect 17509 6749 17543 6783
rect 17543 6749 17552 6783
rect 17500 6740 17552 6749
rect 17776 6740 17828 6792
rect 18604 6740 18656 6792
rect 18972 6740 19024 6792
rect 15660 6672 15712 6724
rect 16764 6672 16816 6724
rect 13176 6647 13228 6656
rect 13176 6613 13185 6647
rect 13185 6613 13219 6647
rect 13219 6613 13228 6647
rect 13176 6604 13228 6613
rect 14556 6604 14608 6656
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 9864 6443 9916 6452
rect 9864 6409 9873 6443
rect 9873 6409 9907 6443
rect 9907 6409 9916 6443
rect 9864 6400 9916 6409
rect 10048 6400 10100 6452
rect 10324 6264 10376 6316
rect 10968 6264 11020 6316
rect 8392 6196 8444 6248
rect 9128 6196 9180 6248
rect 10600 6196 10652 6248
rect 4068 6128 4120 6180
rect 10968 6128 11020 6180
rect 11152 6196 11204 6248
rect 14648 6400 14700 6452
rect 14924 6400 14976 6452
rect 17316 6400 17368 6452
rect 18696 6400 18748 6452
rect 19432 6400 19484 6452
rect 13360 6332 13412 6384
rect 13820 6332 13872 6384
rect 14188 6332 14240 6384
rect 18788 6332 18840 6384
rect 13084 6307 13136 6316
rect 13084 6273 13093 6307
rect 13093 6273 13127 6307
rect 13127 6273 13136 6307
rect 13084 6264 13136 6273
rect 13176 6264 13228 6316
rect 12900 6196 12952 6248
rect 14004 6196 14056 6248
rect 14188 6196 14240 6248
rect 16488 6264 16540 6316
rect 16948 6196 17000 6248
rect 17592 6196 17644 6248
rect 18972 6196 19024 6248
rect 19340 6196 19392 6248
rect 19892 6196 19944 6248
rect 20444 6196 20496 6248
rect 9864 6060 9916 6112
rect 10232 6060 10284 6112
rect 12440 6103 12492 6112
rect 12440 6069 12449 6103
rect 12449 6069 12483 6103
rect 12483 6069 12492 6103
rect 12900 6103 12952 6112
rect 12440 6060 12492 6069
rect 12900 6069 12909 6103
rect 12909 6069 12943 6103
rect 12943 6069 12952 6103
rect 12900 6060 12952 6069
rect 14372 6128 14424 6180
rect 14924 6171 14976 6180
rect 14464 6103 14516 6112
rect 14464 6069 14473 6103
rect 14473 6069 14507 6103
rect 14507 6069 14516 6103
rect 14464 6060 14516 6069
rect 14924 6137 14933 6171
rect 14933 6137 14967 6171
rect 14967 6137 14976 6171
rect 14924 6128 14976 6137
rect 15752 6060 15804 6112
rect 17040 6103 17092 6112
rect 17040 6069 17049 6103
rect 17049 6069 17083 6103
rect 17083 6069 17092 6103
rect 17040 6060 17092 6069
rect 18696 6103 18748 6112
rect 18696 6069 18705 6103
rect 18705 6069 18739 6103
rect 18739 6069 18748 6103
rect 18696 6060 18748 6069
rect 19248 6060 19300 6112
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 9772 5899 9824 5908
rect 9772 5865 9781 5899
rect 9781 5865 9815 5899
rect 9815 5865 9824 5899
rect 9772 5856 9824 5865
rect 10508 5856 10560 5908
rect 12440 5856 12492 5908
rect 14188 5899 14240 5908
rect 14188 5865 14197 5899
rect 14197 5865 14231 5899
rect 14231 5865 14240 5899
rect 14188 5856 14240 5865
rect 14556 5899 14608 5908
rect 14556 5865 14565 5899
rect 14565 5865 14599 5899
rect 14599 5865 14608 5899
rect 14556 5856 14608 5865
rect 16488 5856 16540 5908
rect 13176 5788 13228 5840
rect 15844 5788 15896 5840
rect 16396 5788 16448 5840
rect 18144 5856 18196 5908
rect 18604 5899 18656 5908
rect 18604 5865 18613 5899
rect 18613 5865 18647 5899
rect 18647 5865 18656 5899
rect 18604 5856 18656 5865
rect 20904 5899 20956 5908
rect 20904 5865 20913 5899
rect 20913 5865 20947 5899
rect 20947 5865 20956 5899
rect 20904 5856 20956 5865
rect 16948 5788 17000 5840
rect 8392 5720 8444 5772
rect 10876 5763 10928 5772
rect 10876 5729 10885 5763
rect 10885 5729 10919 5763
rect 10919 5729 10928 5763
rect 10876 5720 10928 5729
rect 12900 5763 12952 5772
rect 12900 5729 12909 5763
rect 12909 5729 12943 5763
rect 12943 5729 12952 5763
rect 12900 5720 12952 5729
rect 15200 5720 15252 5772
rect 15384 5720 15436 5772
rect 10232 5695 10284 5704
rect 10232 5661 10241 5695
rect 10241 5661 10275 5695
rect 10275 5661 10284 5695
rect 10232 5652 10284 5661
rect 10324 5695 10376 5704
rect 10324 5661 10333 5695
rect 10333 5661 10367 5695
rect 10367 5661 10376 5695
rect 13176 5695 13228 5704
rect 10324 5652 10376 5661
rect 13176 5661 13185 5695
rect 13185 5661 13219 5695
rect 13219 5661 13228 5695
rect 13176 5652 13228 5661
rect 13084 5584 13136 5636
rect 13452 5516 13504 5568
rect 17960 5720 18012 5772
rect 18972 5720 19024 5772
rect 18512 5516 18564 5568
rect 20260 5559 20312 5568
rect 20260 5525 20269 5559
rect 20269 5525 20303 5559
rect 20303 5525 20312 5559
rect 20260 5516 20312 5525
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 10232 5312 10284 5364
rect 10876 5312 10928 5364
rect 11796 5312 11848 5364
rect 12900 5312 12952 5364
rect 15844 5312 15896 5364
rect 16948 5312 17000 5364
rect 17316 5312 17368 5364
rect 19892 5355 19944 5364
rect 19892 5321 19901 5355
rect 19901 5321 19935 5355
rect 19935 5321 19944 5355
rect 19892 5312 19944 5321
rect 19708 5244 19760 5296
rect 20536 5244 20588 5296
rect 10784 5219 10836 5228
rect 10784 5185 10793 5219
rect 10793 5185 10827 5219
rect 10827 5185 10836 5219
rect 10784 5176 10836 5185
rect 10968 5219 11020 5228
rect 10968 5185 10977 5219
rect 10977 5185 11011 5219
rect 11011 5185 11020 5219
rect 10968 5176 11020 5185
rect 11888 5176 11940 5228
rect 13084 5219 13136 5228
rect 13084 5185 13093 5219
rect 13093 5185 13127 5219
rect 13127 5185 13136 5219
rect 13084 5176 13136 5185
rect 15384 5176 15436 5228
rect 15660 5176 15712 5228
rect 18512 5219 18564 5228
rect 18512 5185 18521 5219
rect 18521 5185 18555 5219
rect 18555 5185 18564 5219
rect 18512 5176 18564 5185
rect 10048 5108 10100 5160
rect 10692 5108 10744 5160
rect 16488 5108 16540 5160
rect 20260 5108 20312 5160
rect 13176 5040 13228 5092
rect 19800 5040 19852 5092
rect 20720 5040 20772 5092
rect 10692 5015 10744 5024
rect 10692 4981 10701 5015
rect 10701 4981 10735 5015
rect 10735 4981 10744 5015
rect 10692 4972 10744 4981
rect 14464 4972 14516 5024
rect 15384 4972 15436 5024
rect 18144 4972 18196 5024
rect 20168 5015 20220 5024
rect 20168 4981 20177 5015
rect 20177 4981 20211 5015
rect 20211 4981 20220 5015
rect 20168 4972 20220 4981
rect 20628 5015 20680 5024
rect 20628 4981 20637 5015
rect 20637 4981 20671 5015
rect 20671 4981 20680 5015
rect 20628 4972 20680 4981
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 13176 4768 13228 4820
rect 15200 4768 15252 4820
rect 17040 4768 17092 4820
rect 17868 4768 17920 4820
rect 18144 4811 18196 4820
rect 18144 4777 18153 4811
rect 18153 4777 18187 4811
rect 18187 4777 18196 4811
rect 18144 4768 18196 4777
rect 19156 4811 19208 4820
rect 19156 4777 19165 4811
rect 19165 4777 19199 4811
rect 19199 4777 19208 4811
rect 19156 4768 19208 4777
rect 19248 4768 19300 4820
rect 17960 4700 18012 4752
rect 18696 4700 18748 4752
rect 11796 4632 11848 4684
rect 13084 4632 13136 4684
rect 13728 4675 13780 4684
rect 13728 4641 13737 4675
rect 13737 4641 13771 4675
rect 13771 4641 13780 4675
rect 13728 4632 13780 4641
rect 14280 4632 14332 4684
rect 17316 4632 17368 4684
rect 15292 4564 15344 4616
rect 14188 4428 14240 4480
rect 15292 4428 15344 4480
rect 15844 4607 15896 4616
rect 15844 4573 15853 4607
rect 15853 4573 15887 4607
rect 15887 4573 15896 4607
rect 16948 4607 17000 4616
rect 15844 4564 15896 4573
rect 16948 4573 16957 4607
rect 16957 4573 16991 4607
rect 16991 4573 17000 4607
rect 16948 4564 17000 4573
rect 17960 4564 18012 4616
rect 19708 4632 19760 4684
rect 19156 4564 19208 4616
rect 19432 4607 19484 4616
rect 19432 4573 19441 4607
rect 19441 4573 19475 4607
rect 19475 4573 19484 4607
rect 19432 4564 19484 4573
rect 20260 4607 20312 4616
rect 20260 4573 20269 4607
rect 20269 4573 20303 4607
rect 20303 4573 20312 4607
rect 20260 4564 20312 4573
rect 20352 4607 20404 4616
rect 20352 4573 20361 4607
rect 20361 4573 20395 4607
rect 20395 4573 20404 4607
rect 20352 4564 20404 4573
rect 17316 4496 17368 4548
rect 20628 4496 20680 4548
rect 15936 4428 15988 4480
rect 19064 4428 19116 4480
rect 19800 4471 19852 4480
rect 19800 4437 19809 4471
rect 19809 4437 19843 4471
rect 19843 4437 19852 4471
rect 19800 4428 19852 4437
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 7748 4224 7800 4276
rect 17316 4224 17368 4276
rect 19708 4267 19760 4276
rect 19708 4233 19717 4267
rect 19717 4233 19751 4267
rect 19751 4233 19760 4267
rect 19708 4224 19760 4233
rect 10692 4156 10744 4208
rect 12624 4156 12676 4208
rect 13268 4156 13320 4208
rect 8392 4088 8444 4140
rect 11428 4131 11480 4140
rect 11428 4097 11437 4131
rect 11437 4097 11471 4131
rect 11471 4097 11480 4131
rect 11428 4088 11480 4097
rect 13636 4088 13688 4140
rect 14556 4131 14608 4140
rect 14556 4097 14565 4131
rect 14565 4097 14599 4131
rect 14599 4097 14608 4131
rect 14556 4088 14608 4097
rect 19892 4156 19944 4208
rect 20168 4131 20220 4140
rect 848 3952 900 4004
rect 9864 4020 9916 4072
rect 15016 4063 15068 4072
rect 15016 4029 15025 4063
rect 15025 4029 15059 4063
rect 15059 4029 15068 4063
rect 15016 4020 15068 4029
rect 15752 4063 15804 4072
rect 15752 4029 15761 4063
rect 15761 4029 15795 4063
rect 15795 4029 15804 4063
rect 15752 4020 15804 4029
rect 20168 4097 20177 4131
rect 20177 4097 20211 4131
rect 20211 4097 20220 4131
rect 20168 4088 20220 4097
rect 17224 4020 17276 4072
rect 18604 4020 18656 4072
rect 19800 4020 19852 4072
rect 20720 4063 20772 4072
rect 20720 4029 20729 4063
rect 20729 4029 20763 4063
rect 20763 4029 20772 4063
rect 20720 4020 20772 4029
rect 9588 3952 9640 4004
rect 7472 3884 7524 3936
rect 10600 3952 10652 4004
rect 13360 3952 13412 4004
rect 13636 3952 13688 4004
rect 15384 3952 15436 4004
rect 16764 3952 16816 4004
rect 16856 3952 16908 4004
rect 17684 3952 17736 4004
rect 18696 3952 18748 4004
rect 10324 3884 10376 3936
rect 10784 3927 10836 3936
rect 10784 3893 10793 3927
rect 10793 3893 10827 3927
rect 10827 3893 10836 3927
rect 10784 3884 10836 3893
rect 10876 3884 10928 3936
rect 11336 3884 11388 3936
rect 12348 3884 12400 3936
rect 12808 3927 12860 3936
rect 12808 3893 12817 3927
rect 12817 3893 12851 3927
rect 12851 3893 12860 3927
rect 12808 3884 12860 3893
rect 13912 3884 13964 3936
rect 14096 3884 14148 3936
rect 14280 3884 14332 3936
rect 15016 3884 15068 3936
rect 15844 3884 15896 3936
rect 17868 3884 17920 3936
rect 19156 3884 19208 3936
rect 22468 3884 22520 3936
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 9588 3680 9640 3732
rect 11152 3680 11204 3732
rect 11428 3723 11480 3732
rect 11428 3689 11437 3723
rect 11437 3689 11471 3723
rect 11471 3689 11480 3723
rect 11428 3680 11480 3689
rect 11704 3680 11756 3732
rect 3608 3612 3660 3664
rect 296 3544 348 3596
rect 7196 3544 7248 3596
rect 8392 3544 8444 3596
rect 10324 3587 10376 3596
rect 10324 3553 10358 3587
rect 10358 3553 10376 3587
rect 10324 3544 10376 3553
rect 10508 3612 10560 3664
rect 11336 3612 11388 3664
rect 12716 3544 12768 3596
rect 13912 3680 13964 3732
rect 14556 3680 14608 3732
rect 16856 3680 16908 3732
rect 18696 3723 18748 3732
rect 16120 3612 16172 3664
rect 18696 3689 18705 3723
rect 18705 3689 18739 3723
rect 18739 3689 18748 3723
rect 18696 3680 18748 3689
rect 17224 3612 17276 3664
rect 3056 3476 3108 3528
rect 9956 3476 10008 3528
rect 11704 3519 11756 3528
rect 11704 3485 11713 3519
rect 11713 3485 11747 3519
rect 11747 3485 11756 3519
rect 11704 3476 11756 3485
rect 13912 3544 13964 3596
rect 15660 3587 15712 3596
rect 15660 3553 15669 3587
rect 15669 3553 15703 3587
rect 15703 3553 15712 3587
rect 15660 3544 15712 3553
rect 19064 3587 19116 3596
rect 19064 3553 19073 3587
rect 19073 3553 19107 3587
rect 19107 3553 19116 3587
rect 19064 3544 19116 3553
rect 19616 3544 19668 3596
rect 8208 3408 8260 3460
rect 10048 3408 10100 3460
rect 19524 3476 19576 3528
rect 20352 3476 20404 3528
rect 5816 3340 5868 3392
rect 9312 3340 9364 3392
rect 9680 3340 9732 3392
rect 12348 3340 12400 3392
rect 14004 3340 14056 3392
rect 16304 3340 16356 3392
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 6368 3136 6420 3188
rect 10232 3136 10284 3188
rect 10876 3136 10928 3188
rect 14280 3136 14332 3188
rect 7196 3068 7248 3120
rect 4160 3000 4212 3052
rect 10232 3000 10284 3052
rect 10324 3000 10376 3052
rect 13912 3043 13964 3052
rect 13912 3009 13921 3043
rect 13921 3009 13955 3043
rect 13955 3009 13964 3043
rect 13912 3000 13964 3009
rect 14280 3000 14332 3052
rect 15660 3136 15712 3188
rect 17132 3136 17184 3188
rect 17960 3136 18012 3188
rect 16856 3068 16908 3120
rect 17684 3068 17736 3120
rect 17224 3043 17276 3052
rect 17224 3009 17233 3043
rect 17233 3009 17267 3043
rect 17267 3009 17276 3043
rect 17224 3000 17276 3009
rect 18512 3043 18564 3052
rect 18512 3009 18521 3043
rect 18521 3009 18555 3043
rect 18555 3009 18564 3043
rect 18512 3000 18564 3009
rect 18696 3043 18748 3052
rect 18696 3009 18705 3043
rect 18705 3009 18739 3043
rect 18739 3009 18748 3043
rect 18696 3000 18748 3009
rect 8576 2932 8628 2984
rect 10692 2932 10744 2984
rect 11612 2975 11664 2984
rect 11612 2941 11621 2975
rect 11621 2941 11655 2975
rect 11655 2941 11664 2975
rect 11612 2932 11664 2941
rect 2504 2864 2556 2916
rect 4712 2796 4764 2848
rect 11152 2796 11204 2848
rect 11336 2864 11388 2916
rect 12532 2864 12584 2916
rect 14004 2932 14056 2984
rect 15936 2932 15988 2984
rect 16948 2975 17000 2984
rect 16948 2941 16957 2975
rect 16957 2941 16991 2975
rect 16991 2941 17000 2975
rect 16948 2932 17000 2941
rect 18420 2975 18472 2984
rect 18420 2941 18429 2975
rect 18429 2941 18463 2975
rect 18463 2941 18472 2975
rect 18420 2932 18472 2941
rect 19432 2975 19484 2984
rect 19432 2941 19441 2975
rect 19441 2941 19475 2975
rect 19475 2941 19484 2975
rect 19432 2932 19484 2941
rect 20260 3068 20312 3120
rect 20536 2975 20588 2984
rect 20536 2941 20545 2975
rect 20545 2941 20579 2975
rect 20579 2941 20588 2975
rect 20536 2932 20588 2941
rect 14556 2864 14608 2916
rect 15568 2796 15620 2848
rect 16120 2796 16172 2848
rect 17040 2839 17092 2848
rect 17040 2805 17049 2839
rect 17049 2805 17083 2839
rect 17083 2805 17092 2839
rect 17040 2796 17092 2805
rect 21364 2864 21416 2916
rect 21916 2796 21968 2848
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 9772 2592 9824 2644
rect 10232 2592 10284 2644
rect 10784 2592 10836 2644
rect 12256 2592 12308 2644
rect 16028 2635 16080 2644
rect 16028 2601 16037 2635
rect 16037 2601 16071 2635
rect 16071 2601 16080 2635
rect 16028 2592 16080 2601
rect 18144 2592 18196 2644
rect 13728 2567 13780 2576
rect 1400 2388 1452 2440
rect 11336 2499 11388 2508
rect 11336 2465 11345 2499
rect 11345 2465 11379 2499
rect 11379 2465 11388 2499
rect 11336 2456 11388 2465
rect 12532 2456 12584 2508
rect 12992 2456 13044 2508
rect 13452 2499 13504 2508
rect 13452 2465 13461 2499
rect 13461 2465 13495 2499
rect 13495 2465 13504 2499
rect 13452 2456 13504 2465
rect 13728 2533 13737 2567
rect 13737 2533 13771 2567
rect 13771 2533 13780 2567
rect 13728 2524 13780 2533
rect 17776 2524 17828 2576
rect 16764 2456 16816 2508
rect 17316 2499 17368 2508
rect 17316 2465 17325 2499
rect 17325 2465 17359 2499
rect 17359 2465 17368 2499
rect 17316 2456 17368 2465
rect 17408 2456 17460 2508
rect 18972 2499 19024 2508
rect 18972 2465 18981 2499
rect 18981 2465 19015 2499
rect 19015 2465 19024 2499
rect 18972 2456 19024 2465
rect 19524 2499 19576 2508
rect 19524 2465 19533 2499
rect 19533 2465 19567 2499
rect 19567 2465 19576 2499
rect 19524 2456 19576 2465
rect 20352 2499 20404 2508
rect 20352 2465 20361 2499
rect 20361 2465 20395 2499
rect 20395 2465 20404 2499
rect 20352 2456 20404 2465
rect 16120 2431 16172 2440
rect 16120 2397 16129 2431
rect 16129 2397 16163 2431
rect 16163 2397 16172 2431
rect 16120 2388 16172 2397
rect 16304 2388 16356 2440
rect 19248 2388 19300 2440
rect 13084 2320 13136 2372
rect 13636 2320 13688 2372
rect 17040 2320 17092 2372
rect 18696 2320 18748 2372
rect 11980 2252 12032 2304
rect 12532 2252 12584 2304
rect 16396 2252 16448 2304
rect 17500 2295 17552 2304
rect 17500 2261 17509 2295
rect 17509 2261 17543 2295
rect 17543 2261 17552 2295
rect 17500 2252 17552 2261
rect 19064 2252 19116 2304
rect 19616 2252 19668 2304
rect 20812 2252 20864 2304
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 11152 2048 11204 2100
rect 13544 2048 13596 2100
rect 18512 2048 18564 2100
rect 5264 1980 5316 2032
rect 8944 1980 8996 2032
rect 1952 1096 2004 1148
rect 9588 1096 9640 1148
<< metal2 >>
rect 294 22320 350 22800
rect 846 22320 902 22800
rect 1398 22320 1454 22800
rect 1950 22320 2006 22800
rect 2502 22320 2558 22800
rect 3054 22320 3110 22800
rect 3606 22320 3662 22800
rect 4158 22320 4214 22800
rect 4710 22320 4766 22800
rect 5262 22320 5318 22800
rect 5814 22320 5870 22800
rect 6366 22320 6422 22800
rect 6918 22320 6974 22800
rect 7470 22320 7526 22800
rect 8022 22320 8078 22800
rect 8574 22320 8630 22800
rect 9126 22320 9182 22800
rect 9678 22320 9734 22800
rect 10230 22320 10286 22800
rect 10782 22320 10838 22800
rect 11334 22320 11390 22800
rect 11978 22320 12034 22800
rect 12530 22320 12586 22800
rect 13082 22320 13138 22800
rect 13634 22320 13690 22800
rect 14186 22320 14242 22800
rect 14738 22320 14794 22800
rect 15290 22320 15346 22800
rect 15842 22320 15898 22800
rect 16394 22320 16450 22800
rect 16946 22320 17002 22800
rect 17498 22320 17554 22800
rect 18050 22320 18106 22800
rect 18602 22320 18658 22800
rect 19062 22536 19118 22545
rect 19062 22471 19118 22480
rect 308 18970 336 22320
rect 296 18964 348 18970
rect 296 18906 348 18912
rect 860 17814 888 22320
rect 1412 18329 1440 22320
rect 1964 22250 1992 22320
rect 1504 22222 1992 22250
rect 1398 18320 1454 18329
rect 1398 18255 1454 18264
rect 1504 18170 1532 22222
rect 2516 19281 2544 22320
rect 2502 19272 2558 19281
rect 2502 19207 2558 19216
rect 3068 18698 3096 22320
rect 3056 18692 3108 18698
rect 3056 18634 3108 18640
rect 3620 18290 3648 22320
rect 3608 18284 3660 18290
rect 3608 18226 3660 18232
rect 1412 18142 1532 18170
rect 4172 18154 4200 22320
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 4724 18630 4752 22320
rect 4712 18624 4764 18630
rect 4712 18566 4764 18572
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4160 18148 4212 18154
rect 848 17808 900 17814
rect 848 17750 900 17756
rect 1412 13802 1440 18142
rect 4160 18090 4212 18096
rect 5276 18034 5304 22320
rect 5828 18086 5856 22320
rect 6380 19174 6408 22320
rect 6368 19168 6420 19174
rect 6368 19110 6420 19116
rect 6184 18624 6236 18630
rect 6184 18566 6236 18572
rect 5816 18080 5868 18086
rect 5276 18006 5580 18034
rect 5816 18022 5868 18028
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 3422 17232 3478 17241
rect 3422 17167 3478 17176
rect 1400 13796 1452 13802
rect 1400 13738 1452 13744
rect 3436 8634 3464 17167
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 5552 14958 5580 18006
rect 6196 15026 6224 18566
rect 6932 16794 6960 22320
rect 7484 20262 7512 22320
rect 8036 20890 8064 22320
rect 8036 20862 8248 20890
rect 7472 20256 7524 20262
rect 7472 20198 7524 20204
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 7748 19304 7800 19310
rect 7748 19246 7800 19252
rect 7760 18834 7788 19246
rect 8220 19242 8248 20862
rect 8484 19508 8536 19514
rect 8484 19450 8536 19456
rect 8496 19310 8524 19450
rect 8484 19304 8536 19310
rect 8484 19246 8536 19252
rect 8208 19236 8260 19242
rect 8208 19178 8260 19184
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 7748 18828 7800 18834
rect 7748 18770 7800 18776
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 7484 16794 7512 18022
rect 7760 17882 7788 18770
rect 8588 18737 8616 22320
rect 8944 19236 8996 19242
rect 8944 19178 8996 19184
rect 8956 18970 8984 19178
rect 8944 18964 8996 18970
rect 8944 18906 8996 18912
rect 8852 18828 8904 18834
rect 8852 18770 8904 18776
rect 8574 18728 8630 18737
rect 8574 18663 8630 18672
rect 8208 18284 8260 18290
rect 8208 18226 8260 18232
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 7748 17876 7800 17882
rect 7748 17818 7800 17824
rect 7760 17762 7788 17818
rect 7668 17746 7788 17762
rect 7656 17740 7788 17746
rect 7708 17734 7788 17740
rect 7656 17682 7708 17688
rect 7656 17060 7708 17066
rect 7656 17002 7708 17008
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 7472 16788 7524 16794
rect 7472 16730 7524 16736
rect 7668 16590 7696 17002
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 7748 16788 7800 16794
rect 7748 16730 7800 16736
rect 7656 16584 7708 16590
rect 7656 16526 7708 16532
rect 7564 16040 7616 16046
rect 7564 15982 7616 15988
rect 7576 15570 7604 15982
rect 7564 15564 7616 15570
rect 7564 15506 7616 15512
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7484 15094 7512 15302
rect 7472 15088 7524 15094
rect 7472 15030 7524 15036
rect 6184 15020 6236 15026
rect 6184 14962 6236 14968
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 6092 14952 6144 14958
rect 6092 14894 6144 14900
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 6104 14074 6132 14894
rect 7484 14550 7512 15030
rect 7576 14958 7604 15506
rect 7564 14952 7616 14958
rect 7564 14894 7616 14900
rect 7472 14544 7524 14550
rect 7472 14486 7524 14492
rect 6092 14068 6144 14074
rect 6092 14010 6144 14016
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 4080 5817 4108 6122
rect 4066 5808 4122 5817
rect 4066 5743 4122 5752
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 848 4004 900 4010
rect 848 3946 900 3952
rect 296 3596 348 3602
rect 296 3538 348 3544
rect 308 480 336 3538
rect 860 480 888 3946
rect 3608 3664 3660 3670
rect 3608 3606 3660 3612
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 2504 2916 2556 2922
rect 2504 2858 2556 2864
rect 1400 2440 1452 2446
rect 1400 2382 1452 2388
rect 1412 480 1440 2382
rect 1952 1148 2004 1154
rect 1952 1090 2004 1096
rect 1964 480 1992 1090
rect 2516 480 2544 2858
rect 3068 480 3096 3470
rect 3620 480 3648 3606
rect 5816 3392 5868 3398
rect 5816 3334 5868 3340
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 4172 480 4200 2994
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4724 480 4752 2790
rect 5264 2032 5316 2038
rect 5264 1974 5316 1980
rect 5276 480 5304 1974
rect 5828 480 5856 3334
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 6380 480 6408 3130
rect 6932 480 6960 8978
rect 7760 4282 7788 16730
rect 8220 16674 8248 18226
rect 8864 17882 8892 18770
rect 8956 18290 8984 18906
rect 8944 18284 8996 18290
rect 8944 18226 8996 18232
rect 9140 18222 9168 22320
rect 9692 19802 9720 22320
rect 9692 19774 10088 19802
rect 10060 19281 10088 19774
rect 9862 19272 9918 19281
rect 9862 19207 9918 19216
rect 10046 19272 10102 19281
rect 10046 19207 10102 19216
rect 9312 19168 9364 19174
rect 9312 19110 9364 19116
rect 9876 19122 9904 19207
rect 10244 19145 10272 22320
rect 10796 20074 10824 22320
rect 10796 20046 11008 20074
rect 11348 20058 11376 22320
rect 10784 19984 10836 19990
rect 10784 19926 10836 19932
rect 10692 19848 10744 19854
rect 10692 19790 10744 19796
rect 10324 19712 10376 19718
rect 10324 19654 10376 19660
rect 10230 19136 10286 19145
rect 9324 18222 9352 19110
rect 9876 19094 10088 19122
rect 9770 19000 9826 19009
rect 9770 18935 9826 18944
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9494 18456 9550 18465
rect 9494 18391 9550 18400
rect 9588 18420 9640 18426
rect 9128 18216 9180 18222
rect 9128 18158 9180 18164
rect 9312 18216 9364 18222
rect 9312 18158 9364 18164
rect 8668 17876 8720 17882
rect 8668 17818 8720 17824
rect 8852 17876 8904 17882
rect 8852 17818 8904 17824
rect 8484 17808 8536 17814
rect 8484 17750 8536 17756
rect 8392 17740 8444 17746
rect 8392 17682 8444 17688
rect 8404 17338 8432 17682
rect 8496 17338 8524 17750
rect 8392 17332 8444 17338
rect 8392 17274 8444 17280
rect 8484 17332 8536 17338
rect 8484 17274 8536 17280
rect 8680 17134 8708 17818
rect 8864 17270 8892 17818
rect 8852 17264 8904 17270
rect 9324 17218 9352 18158
rect 9508 18154 9536 18391
rect 9588 18362 9640 18368
rect 9600 18329 9628 18362
rect 9586 18320 9642 18329
rect 9586 18255 9642 18264
rect 9496 18148 9548 18154
rect 9496 18090 9548 18096
rect 9692 17882 9720 18702
rect 9784 18698 9812 18935
rect 9864 18896 9916 18902
rect 9864 18838 9916 18844
rect 9772 18692 9824 18698
rect 9772 18634 9824 18640
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9876 17626 9904 18838
rect 9956 18352 10008 18358
rect 9956 18294 10008 18300
rect 9968 17814 9996 18294
rect 9956 17808 10008 17814
rect 9956 17750 10008 17756
rect 9876 17598 9996 17626
rect 8852 17206 8904 17212
rect 8760 17196 8812 17202
rect 8760 17138 8812 17144
rect 8956 17190 9352 17218
rect 8668 17128 8720 17134
rect 8668 17070 8720 17076
rect 8128 16646 8248 16674
rect 8128 15960 8156 16646
rect 8208 16584 8260 16590
rect 8208 16526 8260 16532
rect 8220 16250 8248 16526
rect 8680 16522 8708 17070
rect 8772 16590 8800 17138
rect 8760 16584 8812 16590
rect 8760 16526 8812 16532
rect 8668 16516 8720 16522
rect 8668 16458 8720 16464
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 8680 16114 8708 16458
rect 8668 16108 8720 16114
rect 8668 16050 8720 16056
rect 8668 15972 8720 15978
rect 8128 15932 8248 15960
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 8128 15162 8156 15438
rect 8220 15162 8248 15932
rect 8668 15914 8720 15920
rect 8680 15162 8708 15914
rect 8852 15360 8904 15366
rect 8852 15302 8904 15308
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8668 15156 8720 15162
rect 8668 15098 8720 15104
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 8680 14414 8708 15098
rect 8760 14884 8812 14890
rect 8760 14826 8812 14832
rect 8668 14408 8720 14414
rect 8668 14350 8720 14356
rect 8772 13938 8800 14826
rect 8864 14550 8892 15302
rect 8852 14544 8904 14550
rect 8852 14486 8904 14492
rect 8956 14362 8984 17190
rect 9312 17128 9364 17134
rect 9232 17076 9312 17082
rect 9232 17070 9364 17076
rect 9232 17054 9352 17070
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 9048 15706 9076 16934
rect 9232 16658 9260 17054
rect 9312 16992 9364 16998
rect 9312 16934 9364 16940
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 9220 16652 9272 16658
rect 9220 16594 9272 16600
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 9036 15496 9088 15502
rect 9036 15438 9088 15444
rect 9048 15026 9076 15438
rect 9036 15020 9088 15026
rect 9036 14962 9088 14968
rect 8864 14334 8984 14362
rect 9048 14346 9076 14962
rect 9128 14816 9180 14822
rect 9128 14758 9180 14764
rect 9140 14618 9168 14758
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 9036 14340 9088 14346
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 8772 12238 8800 12786
rect 8760 12232 8812 12238
rect 8760 12174 8812 12180
rect 8772 11694 8800 12174
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 8208 10532 8260 10538
rect 8208 10474 8260 10480
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 8220 9518 8248 10474
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 8864 8838 8892 14334
rect 9036 14282 9088 14288
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 8944 11688 8996 11694
rect 8944 11630 8996 11636
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 8392 7336 8444 7342
rect 8392 7278 8444 7284
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 8404 6254 8432 7278
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 8404 5778 8432 6190
rect 8392 5772 8444 5778
rect 8392 5714 8444 5720
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 8404 4146 8432 5714
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 7208 3126 7236 3538
rect 7196 3120 7248 3126
rect 7196 3062 7248 3068
rect 7484 480 7512 3878
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 8404 3602 8432 4082
rect 8392 3596 8444 3602
rect 8392 3538 8444 3544
rect 8208 3460 8260 3466
rect 8208 3402 8260 3408
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 8220 1442 8248 3402
rect 8576 2984 8628 2990
rect 8576 2926 8628 2932
rect 8036 1414 8248 1442
rect 8036 480 8064 1414
rect 8588 480 8616 2926
rect 8956 2038 8984 11630
rect 9140 11626 9168 12038
rect 9128 11620 9180 11626
rect 9128 11562 9180 11568
rect 9036 11280 9088 11286
rect 9036 11222 9088 11228
rect 9048 2836 9076 11222
rect 9140 11150 9168 11562
rect 9232 11218 9260 16594
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 9232 9518 9260 10406
rect 9324 9722 9352 16934
rect 9402 16688 9458 16697
rect 9402 16623 9458 16632
rect 9496 16652 9548 16658
rect 9416 16522 9444 16623
rect 9496 16594 9548 16600
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9404 16516 9456 16522
rect 9404 16458 9456 16464
rect 9416 16114 9444 16458
rect 9404 16108 9456 16114
rect 9404 16050 9456 16056
rect 9508 14618 9536 16594
rect 9692 15706 9720 16594
rect 9784 16250 9812 16934
rect 9876 16794 9904 16934
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9588 14816 9640 14822
rect 9588 14758 9640 14764
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 9404 14476 9456 14482
rect 9404 14418 9456 14424
rect 9416 13938 9444 14418
rect 9404 13932 9456 13938
rect 9404 13874 9456 13880
rect 9416 13530 9444 13874
rect 9404 13524 9456 13530
rect 9404 13466 9456 13472
rect 9416 12986 9444 13466
rect 9508 13394 9536 14554
rect 9496 13388 9548 13394
rect 9496 13330 9548 13336
rect 9496 13252 9548 13258
rect 9496 13194 9548 13200
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9508 12646 9536 13194
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9508 12374 9536 12582
rect 9600 12374 9628 14758
rect 9692 14278 9720 15506
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9496 12368 9548 12374
rect 9496 12310 9548 12316
rect 9588 12368 9640 12374
rect 9588 12310 9640 12316
rect 9600 11694 9628 12310
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 9588 11688 9640 11694
rect 9588 11630 9640 11636
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9508 11218 9536 11494
rect 9692 11354 9720 12242
rect 9968 11694 9996 17598
rect 10060 15910 10088 19094
rect 10230 19071 10286 19080
rect 10232 18828 10284 18834
rect 10232 18770 10284 18776
rect 10140 18284 10192 18290
rect 10140 18226 10192 18232
rect 10152 17746 10180 18226
rect 10140 17740 10192 17746
rect 10140 17682 10192 17688
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 10244 13569 10272 18770
rect 10336 18154 10364 19654
rect 10508 19508 10560 19514
rect 10508 19450 10560 19456
rect 10520 18834 10548 19450
rect 10704 19174 10732 19790
rect 10692 19168 10744 19174
rect 10692 19110 10744 19116
rect 10600 18896 10652 18902
rect 10600 18838 10652 18844
rect 10508 18828 10560 18834
rect 10508 18770 10560 18776
rect 10416 18760 10468 18766
rect 10416 18702 10468 18708
rect 10428 18290 10456 18702
rect 10508 18352 10560 18358
rect 10508 18294 10560 18300
rect 10416 18284 10468 18290
rect 10416 18226 10468 18232
rect 10324 18148 10376 18154
rect 10520 18136 10548 18294
rect 10612 18290 10640 18838
rect 10704 18358 10732 19110
rect 10692 18352 10744 18358
rect 10692 18294 10744 18300
rect 10600 18284 10652 18290
rect 10600 18226 10652 18232
rect 10324 18090 10376 18096
rect 10428 18108 10548 18136
rect 10428 18034 10456 18108
rect 10600 18080 10652 18086
rect 10336 18006 10456 18034
rect 10520 18040 10600 18068
rect 10336 17678 10364 18006
rect 10324 17672 10376 17678
rect 10324 17614 10376 17620
rect 10322 16688 10378 16697
rect 10322 16623 10378 16632
rect 10336 16590 10364 16623
rect 10324 16584 10376 16590
rect 10324 16526 10376 16532
rect 10230 13560 10286 13569
rect 10230 13495 10286 13504
rect 10520 13462 10548 18040
rect 10796 18057 10824 19926
rect 10876 19916 10928 19922
rect 10876 19858 10928 19864
rect 10600 18022 10652 18028
rect 10782 18048 10838 18057
rect 10782 17983 10838 17992
rect 10692 17196 10744 17202
rect 10692 17138 10744 17144
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10612 15978 10640 17070
rect 10704 16658 10732 17138
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 10692 16652 10744 16658
rect 10692 16594 10744 16600
rect 10692 16108 10744 16114
rect 10692 16050 10744 16056
rect 10600 15972 10652 15978
rect 10600 15914 10652 15920
rect 10612 15026 10640 15914
rect 10600 15020 10652 15026
rect 10600 14962 10652 14968
rect 10704 13938 10732 16050
rect 10796 14958 10824 16934
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 10888 14804 10916 19858
rect 10980 16114 11008 20046
rect 11152 20052 11204 20058
rect 11152 19994 11204 20000
rect 11336 20052 11388 20058
rect 11336 19994 11388 20000
rect 11164 18290 11192 19994
rect 11992 19802 12020 22320
rect 12072 20256 12124 20262
rect 12072 20198 12124 20204
rect 12084 20058 12112 20198
rect 12072 20052 12124 20058
rect 12072 19994 12124 20000
rect 12348 20052 12400 20058
rect 12348 19994 12400 20000
rect 11900 19786 12020 19802
rect 12072 19848 12124 19854
rect 12072 19790 12124 19796
rect 11888 19780 12020 19786
rect 11940 19774 12020 19780
rect 11888 19722 11940 19728
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 11796 19304 11848 19310
rect 11796 19246 11848 19252
rect 11520 19168 11572 19174
rect 11520 19110 11572 19116
rect 11532 18902 11560 19110
rect 11520 18896 11572 18902
rect 11520 18838 11572 18844
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 11152 18284 11204 18290
rect 11152 18226 11204 18232
rect 11612 17672 11664 17678
rect 11612 17614 11664 17620
rect 11060 17536 11112 17542
rect 11060 17478 11112 17484
rect 10968 16108 11020 16114
rect 10968 16050 11020 16056
rect 10968 15904 11020 15910
rect 10968 15846 11020 15852
rect 10980 15638 11008 15846
rect 11072 15706 11100 17478
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 11624 17218 11652 17614
rect 11532 17190 11652 17218
rect 11704 17196 11756 17202
rect 11532 17134 11560 17190
rect 11704 17138 11756 17144
rect 11520 17128 11572 17134
rect 11520 17070 11572 17076
rect 11612 17128 11664 17134
rect 11612 17070 11664 17076
rect 11244 16992 11296 16998
rect 11242 16960 11244 16969
rect 11296 16960 11298 16969
rect 11242 16895 11298 16904
rect 11532 16794 11560 17070
rect 11520 16788 11572 16794
rect 11520 16730 11572 16736
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 10968 15632 11020 15638
rect 10968 15574 11020 15580
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 10980 15162 11008 15438
rect 10968 15156 11020 15162
rect 10968 15098 11020 15104
rect 11164 14822 11192 15846
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 10796 14776 10916 14804
rect 11152 14816 11204 14822
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 10508 13456 10560 13462
rect 10508 13398 10560 13404
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 10244 12986 10272 13330
rect 10232 12980 10284 12986
rect 10232 12922 10284 12928
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 10060 11354 10088 11494
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 9508 10606 9536 11154
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9692 10266 9720 10542
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9956 10192 10008 10198
rect 9956 10134 10008 10140
rect 9588 9988 9640 9994
rect 9588 9930 9640 9936
rect 9312 9716 9364 9722
rect 9312 9658 9364 9664
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 9232 8974 9260 9454
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9140 6254 9168 6734
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 9324 3398 9352 9658
rect 9600 9382 9628 9930
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9600 4010 9628 9318
rect 9692 9042 9720 9454
rect 9680 9036 9732 9042
rect 9732 8996 9904 9024
rect 9680 8978 9732 8984
rect 9876 8430 9904 8996
rect 9864 8424 9916 8430
rect 9864 8366 9916 8372
rect 9772 8356 9824 8362
rect 9772 8298 9824 8304
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9692 7002 9720 7890
rect 9784 7546 9812 8298
rect 9968 8022 9996 10134
rect 10704 10062 10732 10406
rect 10796 10198 10824 14776
rect 11152 14758 11204 14764
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 11072 13870 11100 14214
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11518 13968 11574 13977
rect 11518 13903 11520 13912
rect 11572 13903 11574 13912
rect 11520 13874 11572 13880
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 10888 13326 10916 13670
rect 11164 13530 11192 13670
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 11624 13394 11652 17070
rect 11716 16250 11744 17138
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 11716 16114 11744 16186
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11704 15360 11756 15366
rect 11704 15302 11756 15308
rect 11716 13734 11744 15302
rect 11808 14090 11836 19246
rect 12084 19242 12112 19790
rect 12164 19712 12216 19718
rect 12164 19654 12216 19660
rect 11888 19236 11940 19242
rect 11888 19178 11940 19184
rect 12072 19236 12124 19242
rect 12072 19178 12124 19184
rect 11900 18601 11928 19178
rect 12084 18970 12112 19178
rect 12072 18964 12124 18970
rect 12072 18906 12124 18912
rect 12072 18828 12124 18834
rect 12072 18770 12124 18776
rect 11886 18592 11942 18601
rect 11886 18527 11942 18536
rect 11980 18420 12032 18426
rect 11980 18362 12032 18368
rect 11888 17740 11940 17746
rect 11888 17682 11940 17688
rect 11900 16794 11928 17682
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11992 16674 12020 18362
rect 11900 16646 12020 16674
rect 11900 15026 11928 16646
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 11888 14884 11940 14890
rect 11888 14826 11940 14832
rect 11900 14249 11928 14826
rect 11992 14482 12020 14962
rect 11980 14476 12032 14482
rect 11980 14418 12032 14424
rect 11886 14240 11942 14249
rect 11886 14175 11942 14184
rect 11808 14062 11928 14090
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10888 12782 10916 13262
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10888 10470 10916 11630
rect 10980 11218 11008 12174
rect 10968 11212 11020 11218
rect 10968 11154 11020 11160
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 10784 10192 10836 10198
rect 10784 10134 10836 10140
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10152 9178 10180 9998
rect 10414 9616 10470 9625
rect 10414 9551 10470 9560
rect 10324 9444 10376 9450
rect 10324 9386 10376 9392
rect 10336 9178 10364 9386
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10324 9172 10376 9178
rect 10324 9114 10376 9120
rect 10138 9072 10194 9081
rect 10138 9007 10194 9016
rect 10152 8344 10180 9007
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10336 8401 10364 8570
rect 10322 8392 10378 8401
rect 10152 8316 10272 8344
rect 10322 8327 10378 8336
rect 9956 8016 10008 8022
rect 9956 7958 10008 7964
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9784 6934 9812 7482
rect 9864 7268 9916 7274
rect 9864 7210 9916 7216
rect 9772 6928 9824 6934
rect 9772 6870 9824 6876
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9784 5914 9812 6734
rect 9876 6458 9904 7210
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9876 4162 9904 6054
rect 9784 4134 9904 4162
rect 9588 4004 9640 4010
rect 9588 3946 9640 3952
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9039 2808 9076 2836
rect 9039 2666 9067 2808
rect 9039 2638 9168 2666
rect 8944 2032 8996 2038
rect 8944 1974 8996 1980
rect 9140 480 9168 2638
rect 9600 1154 9628 3674
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9588 1148 9640 1154
rect 9588 1090 9640 1096
rect 9692 480 9720 3334
rect 9784 2650 9812 4134
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 9876 3097 9904 4014
rect 9968 3534 9996 7142
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10060 6458 10088 6802
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10244 6118 10272 8316
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 10336 7546 10364 7890
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10336 5710 10364 6258
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10244 5370 10272 5646
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 10428 5250 10456 9551
rect 10704 9518 10732 9998
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10888 9194 10916 10406
rect 10796 9166 10916 9194
rect 10968 9172 11020 9178
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10520 8634 10548 8978
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10520 7970 10548 8570
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10520 7942 10640 7970
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10520 7546 10548 7822
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 10612 7410 10640 7942
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10508 6656 10560 6662
rect 10508 6598 10560 6604
rect 10520 5914 10548 6598
rect 10600 6248 10652 6254
rect 10600 6190 10652 6196
rect 10508 5908 10560 5914
rect 10508 5850 10560 5856
rect 10244 5222 10456 5250
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10060 3466 10088 5102
rect 10048 3460 10100 3466
rect 10048 3402 10100 3408
rect 10244 3194 10272 5222
rect 10612 4010 10640 6190
rect 10704 5166 10732 8298
rect 10796 5234 10824 9166
rect 10968 9114 11020 9120
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 10888 8634 10916 8978
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10980 8498 11008 9114
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10876 8016 10928 8022
rect 10876 7958 10928 7964
rect 10888 7206 10916 7958
rect 10980 7886 11008 8434
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10980 6322 11008 6802
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 10980 6186 11008 6258
rect 10968 6180 11020 6186
rect 10968 6122 11020 6128
rect 10876 5772 10928 5778
rect 10876 5714 10928 5720
rect 10888 5370 10916 5714
rect 10876 5364 10928 5370
rect 10876 5306 10928 5312
rect 10980 5234 11008 6122
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10704 4593 10732 4966
rect 10690 4584 10746 4593
rect 10690 4519 10746 4528
rect 10692 4208 10744 4214
rect 10692 4150 10744 4156
rect 10600 4004 10652 4010
rect 10600 3946 10652 3952
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10336 3602 10364 3878
rect 10508 3664 10560 3670
rect 10508 3606 10560 3612
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 9862 3088 9918 3097
rect 10336 3058 10364 3538
rect 9862 3023 9918 3032
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10244 2938 10272 2994
rect 10520 2938 10548 3606
rect 10704 2990 10732 4150
rect 10782 4040 10838 4049
rect 10782 3975 10838 3984
rect 10796 3942 10824 3975
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 10876 3936 10928 3942
rect 10876 3878 10928 3884
rect 10888 3194 10916 3878
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10244 2910 10548 2938
rect 10692 2984 10744 2990
rect 10692 2926 10744 2932
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 10244 480 10272 2586
rect 10796 480 10824 2586
rect 11072 1442 11100 12582
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11796 11212 11848 11218
rect 11796 11154 11848 11160
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11808 10674 11836 11154
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11612 10600 11664 10606
rect 11612 10542 11664 10548
rect 11152 10192 11204 10198
rect 11152 10134 11204 10140
rect 11164 9654 11192 10134
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11152 9648 11204 9654
rect 11152 9590 11204 9596
rect 11624 8838 11652 10542
rect 11808 10266 11836 10610
rect 11796 10260 11848 10266
rect 11796 10202 11848 10208
rect 11900 10198 11928 14062
rect 11992 13938 12020 14418
rect 11980 13932 12032 13938
rect 11980 13874 12032 13880
rect 11978 13424 12034 13433
rect 11978 13359 12034 13368
rect 11888 10192 11940 10198
rect 11888 10134 11940 10140
rect 11888 9648 11940 9654
rect 11888 9590 11940 9596
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 11612 8832 11664 8838
rect 11612 8774 11664 8780
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11612 8560 11664 8566
rect 11612 8502 11664 8508
rect 11336 7948 11388 7954
rect 11336 7890 11388 7896
rect 11348 7857 11376 7890
rect 11334 7848 11390 7857
rect 11334 7783 11390 7792
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 11164 3738 11192 6190
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 11428 4140 11480 4146
rect 11428 4082 11480 4088
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 11348 3670 11376 3878
rect 11440 3738 11468 4082
rect 11428 3732 11480 3738
rect 11428 3674 11480 3680
rect 11336 3664 11388 3670
rect 11336 3606 11388 3612
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11624 2990 11652 8502
rect 11716 8430 11744 9318
rect 11900 8974 11928 9590
rect 11992 9042 12020 13359
rect 12084 12918 12112 18770
rect 12176 17202 12204 19654
rect 12254 18864 12310 18873
rect 12254 18799 12310 18808
rect 12268 18630 12296 18799
rect 12256 18624 12308 18630
rect 12256 18566 12308 18572
rect 12164 17196 12216 17202
rect 12164 17138 12216 17144
rect 12360 16697 12388 19994
rect 12544 19174 12572 22320
rect 13096 20058 13124 22320
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 12624 19916 12676 19922
rect 12624 19858 12676 19864
rect 13084 19916 13136 19922
rect 13084 19858 13136 19864
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12530 18320 12586 18329
rect 12530 18255 12586 18264
rect 12346 16688 12402 16697
rect 12346 16623 12402 16632
rect 12256 16584 12308 16590
rect 12256 16526 12308 16532
rect 12268 13433 12296 16526
rect 12348 16516 12400 16522
rect 12348 16458 12400 16464
rect 12360 16250 12388 16458
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12348 16244 12400 16250
rect 12348 16186 12400 16192
rect 12452 16114 12480 16390
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 12544 15910 12572 18255
rect 12532 15904 12584 15910
rect 12532 15846 12584 15852
rect 12440 15632 12492 15638
rect 12440 15574 12492 15580
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 12360 15162 12388 15438
rect 12348 15156 12400 15162
rect 12348 15098 12400 15104
rect 12452 14074 12480 15574
rect 12636 14906 12664 19858
rect 12808 19168 12860 19174
rect 12806 19136 12808 19145
rect 12860 19136 12862 19145
rect 12806 19071 12862 19080
rect 13096 18193 13124 19858
rect 13648 19242 13676 22320
rect 14200 20058 14228 22320
rect 14752 20346 14780 22320
rect 14568 20318 14780 20346
rect 14568 20058 14596 20318
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 15304 20058 15332 22320
rect 14188 20052 14240 20058
rect 14188 19994 14240 20000
rect 14556 20052 14608 20058
rect 14556 19994 14608 20000
rect 15292 20052 15344 20058
rect 15292 19994 15344 20000
rect 14096 19916 14148 19922
rect 14096 19858 14148 19864
rect 15016 19916 15068 19922
rect 15016 19858 15068 19864
rect 13912 19848 13964 19854
rect 13912 19790 13964 19796
rect 13636 19236 13688 19242
rect 13636 19178 13688 19184
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13832 18970 13860 19110
rect 13544 18964 13596 18970
rect 13544 18906 13596 18912
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 13268 18828 13320 18834
rect 13268 18770 13320 18776
rect 13280 18426 13308 18770
rect 13268 18420 13320 18426
rect 13268 18362 13320 18368
rect 13450 18320 13506 18329
rect 13450 18255 13506 18264
rect 13176 18216 13228 18222
rect 13082 18184 13138 18193
rect 13176 18158 13228 18164
rect 13082 18119 13138 18128
rect 12900 17876 12952 17882
rect 12900 17818 12952 17824
rect 12716 15972 12768 15978
rect 12716 15914 12768 15920
rect 12728 15162 12756 15914
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 12636 14878 12756 14906
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12636 14618 12664 14758
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 12254 13424 12310 13433
rect 12254 13359 12310 13368
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12256 13320 12308 13326
rect 12256 13262 12308 13268
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 12084 11762 12112 12242
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 12084 11354 12112 11698
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 12164 11280 12216 11286
rect 12070 11248 12126 11257
rect 12164 11222 12216 11228
rect 12070 11183 12126 11192
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 11796 8968 11848 8974
rect 11796 8910 11848 8916
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 11808 8090 11836 8910
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 11900 8634 11928 8774
rect 11888 8628 11940 8634
rect 11888 8570 11940 8576
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11808 6798 11836 7686
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11808 5370 11836 6734
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11808 4690 11836 5306
rect 11900 5234 11928 8570
rect 11992 8362 12020 8774
rect 11980 8356 12032 8362
rect 11980 8298 12032 8304
rect 12084 7818 12112 11183
rect 12072 7812 12124 7818
rect 12072 7754 12124 7760
rect 12176 7698 12204 11222
rect 12268 10713 12296 13262
rect 12452 12986 12480 13330
rect 12544 13190 12572 13806
rect 12636 13530 12664 14554
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12728 13462 12756 14878
rect 12820 14618 12848 15302
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 12912 13870 12940 17818
rect 12992 17672 13044 17678
rect 12992 17614 13044 17620
rect 13004 15706 13032 17614
rect 12992 15700 13044 15706
rect 12992 15642 13044 15648
rect 13096 15586 13124 18119
rect 13004 15558 13124 15586
rect 12900 13864 12952 13870
rect 12900 13806 12952 13812
rect 13004 13716 13032 15558
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 13096 14890 13124 15438
rect 13084 14884 13136 14890
rect 13084 14826 13136 14832
rect 13096 14278 13124 14826
rect 13188 14385 13216 18158
rect 13268 18080 13320 18086
rect 13268 18022 13320 18028
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13280 17882 13308 18022
rect 13268 17876 13320 17882
rect 13268 17818 13320 17824
rect 13372 17338 13400 18022
rect 13464 17678 13492 18255
rect 13556 17678 13584 18906
rect 13636 18896 13688 18902
rect 13636 18838 13688 18844
rect 13818 18864 13874 18873
rect 13648 18222 13676 18838
rect 13818 18799 13874 18808
rect 13636 18216 13688 18222
rect 13636 18158 13688 18164
rect 13452 17672 13504 17678
rect 13452 17614 13504 17620
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13360 17332 13412 17338
rect 13360 17274 13412 17280
rect 13464 17082 13492 17614
rect 13556 17202 13584 17614
rect 13544 17196 13596 17202
rect 13544 17138 13596 17144
rect 13372 17054 13492 17082
rect 13268 15904 13320 15910
rect 13268 15846 13320 15852
rect 13174 14376 13230 14385
rect 13174 14311 13230 14320
rect 13084 14272 13136 14278
rect 13084 14214 13136 14220
rect 13176 14272 13228 14278
rect 13176 14214 13228 14220
rect 13096 14006 13124 14214
rect 13084 14000 13136 14006
rect 13084 13942 13136 13948
rect 12820 13688 13032 13716
rect 13084 13728 13136 13734
rect 12716 13456 12768 13462
rect 12716 13398 12768 13404
rect 12532 13184 12584 13190
rect 12532 13126 12584 13132
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12440 12708 12492 12714
rect 12440 12650 12492 12656
rect 12452 11898 12480 12650
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 12452 10810 12480 11494
rect 12440 10804 12492 10810
rect 12440 10746 12492 10752
rect 12254 10704 12310 10713
rect 12254 10639 12310 10648
rect 11992 7670 12204 7698
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 11796 4684 11848 4690
rect 11796 4626 11848 4632
rect 11808 4026 11836 4626
rect 11716 3998 11836 4026
rect 11716 3738 11744 3998
rect 11704 3732 11756 3738
rect 11704 3674 11756 3680
rect 11716 3534 11744 3674
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 11992 3074 12020 7670
rect 11992 3046 12112 3074
rect 11612 2984 11664 2990
rect 11612 2926 11664 2932
rect 11336 2916 11388 2922
rect 11336 2858 11388 2864
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 11164 2106 11192 2790
rect 11348 2514 11376 2858
rect 11336 2508 11388 2514
rect 11336 2450 11388 2456
rect 11980 2304 12032 2310
rect 11980 2246 12032 2252
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11152 2100 11204 2106
rect 11152 2042 11204 2048
rect 11072 1414 11376 1442
rect 11348 480 11376 1414
rect 11992 480 12020 2246
rect 12084 649 12112 3046
rect 12268 2650 12296 10639
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 12360 9178 12388 10066
rect 12452 9994 12480 10542
rect 12440 9988 12492 9994
rect 12440 9930 12492 9936
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 12452 9042 12480 9454
rect 12544 9110 12572 13126
rect 12716 11620 12768 11626
rect 12716 11562 12768 11568
rect 12728 10742 12756 11562
rect 12716 10736 12768 10742
rect 12716 10678 12768 10684
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 12624 10464 12676 10470
rect 12624 10406 12676 10412
rect 12532 9104 12584 9110
rect 12532 9046 12584 9052
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 12360 3942 12388 8978
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12544 8090 12572 8434
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12544 6866 12572 8026
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12452 5914 12480 6054
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12636 4214 12664 10406
rect 12624 4208 12676 4214
rect 12624 4150 12676 4156
rect 12348 3936 12400 3942
rect 12348 3878 12400 3884
rect 12728 3602 12756 10542
rect 12820 10470 12848 13688
rect 13084 13670 13136 13676
rect 13096 13161 13124 13670
rect 13188 13394 13216 14214
rect 13176 13388 13228 13394
rect 13176 13330 13228 13336
rect 13082 13152 13138 13161
rect 13082 13087 13138 13096
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 12900 12640 12952 12646
rect 12900 12582 12952 12588
rect 12912 11898 12940 12582
rect 13004 12442 13032 12786
rect 13084 12776 13136 12782
rect 13084 12718 13136 12724
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 12992 12300 13044 12306
rect 13096 12288 13124 12718
rect 13044 12260 13124 12288
rect 12992 12242 13044 12248
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 13004 10810 13032 11494
rect 12992 10804 13044 10810
rect 12992 10746 13044 10752
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12992 9920 13044 9926
rect 12992 9862 13044 9868
rect 12900 8900 12952 8906
rect 12900 8842 12952 8848
rect 12912 8566 12940 8842
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 12808 8356 12860 8362
rect 12808 8298 12860 8304
rect 12820 7546 12848 8298
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12912 8090 12940 8230
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12912 6254 12940 7142
rect 12900 6248 12952 6254
rect 12900 6190 12952 6196
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 12912 5930 12940 6054
rect 12820 5902 12940 5930
rect 12820 3942 12848 5902
rect 12900 5772 12952 5778
rect 12900 5714 12952 5720
rect 12912 5370 12940 5714
rect 12900 5364 12952 5370
rect 12900 5306 12952 5312
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12346 3496 12402 3505
rect 12346 3431 12402 3440
rect 12360 3398 12388 3431
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 12532 2916 12584 2922
rect 12532 2858 12584 2864
rect 12256 2644 12308 2650
rect 12256 2586 12308 2592
rect 12544 2514 12572 2858
rect 13004 2514 13032 9862
rect 13174 7848 13230 7857
rect 13174 7783 13230 7792
rect 13188 7410 13216 7783
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13188 7002 13216 7142
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 13188 6322 13216 6598
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 13096 5642 13124 6258
rect 13188 5846 13216 6258
rect 13280 5930 13308 15846
rect 13372 6390 13400 17054
rect 13452 16992 13504 16998
rect 13452 16934 13504 16940
rect 13464 15314 13492 16934
rect 13648 16658 13676 18158
rect 13832 16998 13860 18799
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13924 16810 13952 19790
rect 14004 17672 14056 17678
rect 14004 17614 14056 17620
rect 14016 17270 14044 17614
rect 14004 17264 14056 17270
rect 14004 17206 14056 17212
rect 13832 16782 13952 16810
rect 13636 16652 13688 16658
rect 13636 16594 13688 16600
rect 13544 16244 13596 16250
rect 13544 16186 13596 16192
rect 13556 15502 13584 16186
rect 13648 16114 13676 16594
rect 13728 16448 13780 16454
rect 13728 16390 13780 16396
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 13740 15638 13768 16390
rect 13832 15910 13860 16782
rect 14004 16040 14056 16046
rect 14004 15982 14056 15988
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 13728 15632 13780 15638
rect 13728 15574 13780 15580
rect 13544 15496 13596 15502
rect 13544 15438 13596 15444
rect 13464 15286 13584 15314
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13464 13734 13492 14418
rect 13452 13728 13504 13734
rect 13452 13670 13504 13676
rect 13452 7880 13504 7886
rect 13450 7848 13452 7857
rect 13504 7848 13506 7857
rect 13450 7783 13506 7792
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13464 7274 13492 7686
rect 13452 7268 13504 7274
rect 13452 7210 13504 7216
rect 13360 6384 13412 6390
rect 13360 6326 13412 6332
rect 13280 5902 13400 5930
rect 13176 5840 13228 5846
rect 13228 5788 13308 5794
rect 13176 5782 13308 5788
rect 13188 5766 13308 5782
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 13084 5636 13136 5642
rect 13084 5578 13136 5584
rect 13096 5234 13124 5578
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 13096 4690 13124 5170
rect 13188 5098 13216 5646
rect 13176 5092 13228 5098
rect 13176 5034 13228 5040
rect 13188 4826 13216 5034
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 13280 4214 13308 5766
rect 13268 4208 13320 4214
rect 13268 4150 13320 4156
rect 13372 4010 13400 5902
rect 13452 5568 13504 5574
rect 13452 5510 13504 5516
rect 13360 4004 13412 4010
rect 13360 3946 13412 3952
rect 13464 2514 13492 5510
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 12992 2508 13044 2514
rect 12992 2450 13044 2456
rect 13452 2508 13504 2514
rect 13452 2450 13504 2456
rect 13084 2372 13136 2378
rect 13084 2314 13136 2320
rect 12532 2304 12584 2310
rect 12532 2246 12584 2252
rect 12070 640 12126 649
rect 12070 575 12126 584
rect 12544 480 12572 2246
rect 13096 480 13124 2314
rect 13556 2106 13584 15286
rect 13636 15156 13688 15162
rect 13636 15098 13688 15104
rect 13648 14414 13676 15098
rect 13636 14408 13688 14414
rect 13832 14362 13860 15846
rect 14016 15638 14044 15982
rect 14004 15632 14056 15638
rect 14004 15574 14056 15580
rect 13912 15360 13964 15366
rect 13912 15302 13964 15308
rect 13636 14350 13688 14356
rect 13740 14334 13860 14362
rect 13634 14240 13690 14249
rect 13634 14175 13690 14184
rect 13648 13682 13676 14175
rect 13740 13818 13768 14334
rect 13924 13938 13952 15302
rect 14016 14958 14044 15574
rect 14004 14952 14056 14958
rect 14004 14894 14056 14900
rect 14108 14550 14136 19858
rect 15028 19310 15056 19858
rect 15384 19848 15436 19854
rect 15384 19790 15436 19796
rect 14188 19304 14240 19310
rect 14188 19246 14240 19252
rect 14280 19304 14332 19310
rect 14280 19246 14332 19252
rect 15016 19304 15068 19310
rect 15016 19246 15068 19252
rect 14200 18766 14228 19246
rect 14188 18760 14240 18766
rect 14188 18702 14240 18708
rect 14188 18624 14240 18630
rect 14188 18566 14240 18572
rect 14200 18222 14228 18566
rect 14188 18216 14240 18222
rect 14188 18158 14240 18164
rect 14188 16992 14240 16998
rect 14188 16934 14240 16940
rect 14096 14544 14148 14550
rect 14096 14486 14148 14492
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 14004 14272 14056 14278
rect 14004 14214 14056 14220
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 13740 13790 13952 13818
rect 13648 13654 13860 13682
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13740 12753 13768 13126
rect 13726 12744 13782 12753
rect 13726 12679 13782 12688
rect 13728 11008 13780 11014
rect 13728 10950 13780 10956
rect 13740 10606 13768 10950
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13740 10146 13768 10542
rect 13648 10118 13768 10146
rect 13648 7970 13676 10118
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13740 9382 13768 9998
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13740 9110 13768 9318
rect 13728 9104 13780 9110
rect 13728 9046 13780 9052
rect 13832 8378 13860 13654
rect 13740 8362 13860 8378
rect 13728 8356 13860 8362
rect 13780 8350 13860 8356
rect 13728 8298 13780 8304
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13832 8090 13860 8230
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13648 7942 13860 7970
rect 13924 7954 13952 13790
rect 14016 10742 14044 14214
rect 14004 10736 14056 10742
rect 14004 10678 14056 10684
rect 14004 10464 14056 10470
rect 14004 10406 14056 10412
rect 14016 10198 14044 10406
rect 14004 10192 14056 10198
rect 14004 10134 14056 10140
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 14016 9518 14044 9998
rect 14004 9512 14056 9518
rect 14004 9454 14056 9460
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 14016 8430 14044 9318
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 14004 8016 14056 8022
rect 14004 7958 14056 7964
rect 13728 7336 13780 7342
rect 13728 7278 13780 7284
rect 13740 6866 13768 7278
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13832 6798 13860 7942
rect 13912 7948 13964 7954
rect 13912 7890 13964 7896
rect 14016 7750 14044 7958
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 13912 7200 13964 7206
rect 13912 7142 13964 7148
rect 13924 7002 13952 7142
rect 13912 6996 13964 7002
rect 13912 6938 13964 6944
rect 13820 6792 13872 6798
rect 13820 6734 13872 6740
rect 13820 6384 13872 6390
rect 13820 6326 13872 6332
rect 13728 4684 13780 4690
rect 13728 4626 13780 4632
rect 13636 4140 13688 4146
rect 13636 4082 13688 4088
rect 13648 4010 13676 4082
rect 13636 4004 13688 4010
rect 13636 3946 13688 3952
rect 13740 2582 13768 4626
rect 13832 3505 13860 6326
rect 14016 6254 14044 7686
rect 14004 6248 14056 6254
rect 14004 6190 14056 6196
rect 14108 3942 14136 14350
rect 14200 14226 14228 16934
rect 14292 14414 14320 19246
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 15292 18896 15344 18902
rect 15292 18838 15344 18844
rect 15304 18766 15332 18838
rect 15108 18760 15160 18766
rect 15108 18702 15160 18708
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 14556 17740 14608 17746
rect 14556 17682 14608 17688
rect 14568 17338 14596 17682
rect 15016 17672 15068 17678
rect 15016 17614 15068 17620
rect 14556 17332 14608 17338
rect 14556 17274 14608 17280
rect 14464 17196 14516 17202
rect 14464 17138 14516 17144
rect 14372 16992 14424 16998
rect 14370 16960 14372 16969
rect 14424 16960 14426 16969
rect 14370 16895 14426 16904
rect 14476 16726 14504 17138
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 14464 16720 14516 16726
rect 14464 16662 14516 16668
rect 15028 16454 15056 17614
rect 15016 16448 15068 16454
rect 15016 16390 15068 16396
rect 15028 16250 15056 16390
rect 15016 16244 15068 16250
rect 15016 16186 15068 16192
rect 15028 15978 15056 16186
rect 15016 15972 15068 15978
rect 15016 15914 15068 15920
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 14554 15600 14610 15609
rect 14554 15535 14556 15544
rect 14608 15535 14610 15544
rect 14556 15506 14608 15512
rect 15016 15496 15068 15502
rect 15016 15438 15068 15444
rect 15028 15162 15056 15438
rect 15016 15156 15068 15162
rect 15016 15098 15068 15104
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14200 14198 14320 14226
rect 14188 13388 14240 13394
rect 14188 13330 14240 13336
rect 14200 11354 14228 13330
rect 14188 11348 14240 11354
rect 14188 11290 14240 11296
rect 14200 9518 14228 11290
rect 14292 10198 14320 14198
rect 14384 13530 14412 14418
rect 15028 13938 15056 15098
rect 15016 13932 15068 13938
rect 15016 13874 15068 13880
rect 14556 13728 14608 13734
rect 14556 13670 14608 13676
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14372 13184 14424 13190
rect 14372 13126 14424 13132
rect 14384 12714 14412 13126
rect 14372 12708 14424 12714
rect 14372 12650 14424 12656
rect 14384 12442 14412 12650
rect 14372 12436 14424 12442
rect 14372 12378 14424 12384
rect 14384 11762 14412 12378
rect 14372 11756 14424 11762
rect 14372 11698 14424 11704
rect 14476 11694 14504 13262
rect 14568 12442 14596 13670
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 15120 13444 15148 18702
rect 15304 18290 15332 18702
rect 15292 18284 15344 18290
rect 15292 18226 15344 18232
rect 15200 16584 15252 16590
rect 15200 16526 15252 16532
rect 15212 15706 15240 16526
rect 15200 15700 15252 15706
rect 15200 15642 15252 15648
rect 15292 15360 15344 15366
rect 15292 15302 15344 15308
rect 15304 14482 15332 15302
rect 15292 14476 15344 14482
rect 15292 14418 15344 14424
rect 15198 14376 15254 14385
rect 15198 14311 15254 14320
rect 15028 13416 15148 13444
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 14936 13297 14964 13330
rect 14922 13288 14978 13297
rect 14922 13223 14978 13232
rect 15028 12646 15056 13416
rect 15212 13394 15240 14311
rect 15396 14278 15424 19790
rect 15476 18896 15528 18902
rect 15476 18838 15528 18844
rect 15488 18086 15516 18838
rect 15658 18592 15714 18601
rect 15658 18527 15714 18536
rect 15476 18080 15528 18086
rect 15476 18022 15528 18028
rect 15568 17536 15620 17542
rect 15568 17478 15620 17484
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 15488 15484 15516 16934
rect 15580 15638 15608 17478
rect 15672 17066 15700 18527
rect 15856 18426 15884 22320
rect 16408 20074 16436 22320
rect 16408 20058 16620 20074
rect 16408 20052 16632 20058
rect 16408 20046 16580 20052
rect 16580 19994 16632 20000
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16120 19168 16172 19174
rect 16120 19110 16172 19116
rect 16212 19168 16264 19174
rect 16212 19110 16264 19116
rect 15844 18420 15896 18426
rect 15844 18362 15896 18368
rect 15752 18216 15804 18222
rect 15752 18158 15804 18164
rect 15660 17060 15712 17066
rect 15660 17002 15712 17008
rect 15764 16946 15792 18158
rect 16132 17882 16160 19110
rect 16120 17876 16172 17882
rect 16120 17818 16172 17824
rect 15936 17672 15988 17678
rect 15936 17614 15988 17620
rect 15672 16918 15792 16946
rect 15672 15994 15700 16918
rect 15752 16448 15804 16454
rect 15752 16390 15804 16396
rect 15764 16114 15792 16390
rect 15844 16176 15896 16182
rect 15844 16118 15896 16124
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 15672 15966 15792 15994
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15672 15706 15700 15846
rect 15660 15700 15712 15706
rect 15660 15642 15712 15648
rect 15568 15632 15620 15638
rect 15568 15574 15620 15580
rect 15568 15496 15620 15502
rect 15488 15456 15568 15484
rect 15568 15438 15620 15444
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 15200 13388 15252 13394
rect 15120 13348 15200 13376
rect 15016 12640 15068 12646
rect 15016 12582 15068 12588
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 14556 12436 14608 12442
rect 14556 12378 14608 12384
rect 14740 12368 14792 12374
rect 14740 12310 14792 12316
rect 14752 11744 14780 12310
rect 14924 11892 14976 11898
rect 14924 11834 14976 11840
rect 14568 11716 14780 11744
rect 14464 11688 14516 11694
rect 14370 11656 14426 11665
rect 14464 11630 14516 11636
rect 14370 11591 14426 11600
rect 14384 11014 14412 11591
rect 14568 11558 14596 11716
rect 14936 11626 14964 11834
rect 14924 11620 14976 11626
rect 14924 11562 14976 11568
rect 14464 11552 14516 11558
rect 14464 11494 14516 11500
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 14476 11082 14504 11494
rect 14464 11076 14516 11082
rect 14464 11018 14516 11024
rect 14372 11008 14424 11014
rect 14372 10950 14424 10956
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14280 10192 14332 10198
rect 14280 10134 14332 10140
rect 14384 10044 14412 10746
rect 14568 10606 14596 11494
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14292 10016 14412 10044
rect 14188 9512 14240 9518
rect 14188 9454 14240 9460
rect 14292 8514 14320 10016
rect 14372 9920 14424 9926
rect 14372 9862 14424 9868
rect 14384 9722 14412 9862
rect 14372 9716 14424 9722
rect 14372 9658 14424 9664
rect 14476 8838 14504 10542
rect 15028 10452 15056 12582
rect 15120 10810 15148 13348
rect 15200 13330 15252 13336
rect 15198 12880 15254 12889
rect 15198 12815 15254 12824
rect 15212 12782 15240 12815
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15304 12628 15332 14010
rect 15396 14006 15424 14214
rect 15384 14000 15436 14006
rect 15384 13942 15436 13948
rect 15382 13288 15438 13297
rect 15382 13223 15438 13232
rect 15212 12600 15332 12628
rect 15108 10804 15160 10810
rect 15108 10746 15160 10752
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 14568 10424 15056 10452
rect 14372 8832 14424 8838
rect 14372 8774 14424 8780
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14200 8486 14320 8514
rect 14384 8498 14412 8774
rect 14372 8492 14424 8498
rect 14200 6390 14228 8486
rect 14372 8434 14424 8440
rect 14280 8356 14332 8362
rect 14280 8298 14332 8304
rect 14188 6384 14240 6390
rect 14188 6326 14240 6332
rect 14188 6248 14240 6254
rect 14188 6190 14240 6196
rect 14200 5914 14228 6190
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 14292 4690 14320 8298
rect 14384 7970 14412 8434
rect 14476 8090 14504 8774
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 14384 7942 14504 7970
rect 14476 7886 14504 7942
rect 14464 7880 14516 7886
rect 14370 7848 14426 7857
rect 14464 7822 14516 7828
rect 14370 7783 14426 7792
rect 14384 6934 14412 7783
rect 14476 7342 14504 7822
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 14372 6928 14424 6934
rect 14372 6870 14424 6876
rect 14384 6186 14412 6870
rect 14476 6798 14504 7278
rect 14568 6882 14596 10424
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 15016 10192 15068 10198
rect 15016 10134 15068 10140
rect 14924 9988 14976 9994
rect 14924 9930 14976 9936
rect 14936 9450 14964 9930
rect 14924 9444 14976 9450
rect 14924 9386 14976 9392
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 14568 6854 14688 6882
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14372 6180 14424 6186
rect 14372 6122 14424 6128
rect 14280 4684 14332 4690
rect 14280 4626 14332 4632
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 13912 3936 13964 3942
rect 13912 3878 13964 3884
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 13924 3738 13952 3878
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 13818 3496 13874 3505
rect 13818 3431 13874 3440
rect 13924 3058 13952 3538
rect 14004 3392 14056 3398
rect 14004 3334 14056 3340
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 14016 2990 14044 3334
rect 14004 2984 14056 2990
rect 14004 2926 14056 2932
rect 13728 2576 13780 2582
rect 13728 2518 13780 2524
rect 13636 2372 13688 2378
rect 13636 2314 13688 2320
rect 13544 2100 13596 2106
rect 13544 2042 13596 2048
rect 13648 480 13676 2314
rect 14200 480 14228 4422
rect 14280 3936 14332 3942
rect 14280 3878 14332 3884
rect 14292 3194 14320 3878
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14280 3052 14332 3058
rect 14384 3040 14412 6122
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14476 5030 14504 6054
rect 14568 5914 14596 6598
rect 14660 6458 14688 6854
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 14844 6610 14872 6802
rect 14844 6582 14964 6610
rect 14936 6458 14964 6582
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 14924 6452 14976 6458
rect 14924 6394 14976 6400
rect 14936 6186 14964 6394
rect 14924 6180 14976 6186
rect 14924 6122 14976 6128
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 14556 5908 14608 5914
rect 14556 5850 14608 5856
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 14568 3738 14596 4082
rect 15028 4078 15056 10134
rect 15120 10062 15148 10610
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 15120 9382 15148 9998
rect 15108 9376 15160 9382
rect 15108 9318 15160 9324
rect 15108 7948 15160 7954
rect 15108 7890 15160 7896
rect 15120 5273 15148 7890
rect 15212 6100 15240 12600
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 15304 10606 15332 12174
rect 15396 10810 15424 13223
rect 15488 11642 15516 15098
rect 15580 13682 15608 15438
rect 15660 14884 15712 14890
rect 15660 14826 15712 14832
rect 15672 14550 15700 14826
rect 15660 14544 15712 14550
rect 15660 14486 15712 14492
rect 15672 13870 15700 14486
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 15580 13654 15700 13682
rect 15568 13456 15620 13462
rect 15568 13398 15620 13404
rect 15580 11898 15608 13398
rect 15672 13274 15700 13654
rect 15764 13462 15792 15966
rect 15856 15502 15884 16118
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15856 14958 15884 15438
rect 15948 15162 15976 17614
rect 16224 17338 16252 19110
rect 16684 18970 16712 19314
rect 16856 19304 16908 19310
rect 16856 19246 16908 19252
rect 16672 18964 16724 18970
rect 16672 18906 16724 18912
rect 16580 18828 16632 18834
rect 16580 18770 16632 18776
rect 16304 18284 16356 18290
rect 16356 18244 16436 18272
rect 16304 18226 16356 18232
rect 16304 18080 16356 18086
rect 16304 18022 16356 18028
rect 16316 17678 16344 18022
rect 16408 17882 16436 18244
rect 16396 17876 16448 17882
rect 16396 17818 16448 17824
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 16316 17202 16344 17614
rect 16488 17536 16540 17542
rect 16488 17478 16540 17484
rect 16304 17196 16356 17202
rect 16304 17138 16356 17144
rect 16396 17128 16448 17134
rect 16396 17070 16448 17076
rect 16304 16992 16356 16998
rect 16304 16934 16356 16940
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16120 16652 16172 16658
rect 16120 16594 16172 16600
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 15936 15156 15988 15162
rect 15936 15098 15988 15104
rect 15844 14952 15896 14958
rect 15844 14894 15896 14900
rect 16040 14498 16068 16526
rect 16132 15638 16160 16594
rect 16120 15632 16172 15638
rect 16120 15574 16172 15580
rect 16224 14958 16252 16730
rect 16212 14952 16264 14958
rect 16212 14894 16264 14900
rect 16040 14470 16160 14498
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 15752 13456 15804 13462
rect 15750 13424 15752 13433
rect 15804 13424 15806 13433
rect 16040 13394 16068 14350
rect 15750 13359 15806 13368
rect 16028 13388 16080 13394
rect 16028 13330 16080 13336
rect 16132 13274 16160 14470
rect 16212 14476 16264 14482
rect 16212 14418 16264 14424
rect 16224 14006 16252 14418
rect 16212 14000 16264 14006
rect 16212 13942 16264 13948
rect 16224 13870 16252 13942
rect 16212 13864 16264 13870
rect 16210 13832 16212 13841
rect 16264 13832 16266 13841
rect 16210 13767 16266 13776
rect 15672 13246 15976 13274
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15672 11762 15700 13246
rect 15948 13190 15976 13246
rect 16040 13246 16160 13274
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 15750 12880 15806 12889
rect 15750 12815 15806 12824
rect 15764 12238 15792 12815
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15764 11898 15792 12038
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15488 11614 15700 11642
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15488 9450 15516 11494
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 15580 9654 15608 10066
rect 15568 9648 15620 9654
rect 15568 9590 15620 9596
rect 15292 9444 15344 9450
rect 15292 9386 15344 9392
rect 15476 9444 15528 9450
rect 15476 9386 15528 9392
rect 15304 7954 15332 9386
rect 15672 8906 15700 11614
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 15764 11218 15792 11494
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 15752 11076 15804 11082
rect 15752 11018 15804 11024
rect 15764 10554 15792 11018
rect 15856 10674 15884 13126
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 15844 10668 15896 10674
rect 15844 10610 15896 10616
rect 15764 10526 15884 10554
rect 15750 10432 15806 10441
rect 15750 10367 15806 10376
rect 15764 9722 15792 10367
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 15764 9042 15792 9658
rect 15856 9586 15884 10526
rect 15844 9580 15896 9586
rect 15844 9522 15896 9528
rect 15752 9036 15804 9042
rect 15752 8978 15804 8984
rect 15660 8900 15712 8906
rect 15660 8842 15712 8848
rect 15856 8498 15884 9522
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 15568 8288 15620 8294
rect 15568 8230 15620 8236
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 15212 6072 15332 6100
rect 15200 5772 15252 5778
rect 15200 5714 15252 5720
rect 15106 5264 15162 5273
rect 15106 5199 15162 5208
rect 15212 4826 15240 5714
rect 15200 4820 15252 4826
rect 15200 4762 15252 4768
rect 15304 4622 15332 6072
rect 15396 5778 15424 7142
rect 15384 5772 15436 5778
rect 15384 5714 15436 5720
rect 15396 5234 15424 5714
rect 15384 5228 15436 5234
rect 15384 5170 15436 5176
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15292 4616 15344 4622
rect 15292 4558 15344 4564
rect 15292 4480 15344 4486
rect 15292 4422 15344 4428
rect 15016 4072 15068 4078
rect 15016 4014 15068 4020
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 14556 3732 14608 3738
rect 14556 3674 14608 3680
rect 14332 3012 14412 3040
rect 14280 2994 14332 3000
rect 14568 2922 14596 3674
rect 14556 2916 14608 2922
rect 14556 2858 14608 2864
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 15028 1034 15056 3878
rect 14752 1006 15056 1034
rect 14752 480 14780 1006
rect 15304 480 15332 4422
rect 15396 4010 15424 4966
rect 15384 4004 15436 4010
rect 15384 3946 15436 3952
rect 15580 2854 15608 8230
rect 15660 7268 15712 7274
rect 15660 7210 15712 7216
rect 15672 7002 15700 7210
rect 15948 7002 15976 11698
rect 15660 6996 15712 7002
rect 15660 6938 15712 6944
rect 15936 6996 15988 7002
rect 15936 6938 15988 6944
rect 15672 6730 15700 6938
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 15844 6792 15896 6798
rect 15844 6734 15896 6740
rect 15660 6724 15712 6730
rect 15660 6666 15712 6672
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 15672 3602 15700 5170
rect 15764 4078 15792 6054
rect 15856 5846 15884 6734
rect 15844 5840 15896 5846
rect 15844 5782 15896 5788
rect 15856 5370 15884 5782
rect 15844 5364 15896 5370
rect 15844 5306 15896 5312
rect 15856 4622 15884 5306
rect 15844 4616 15896 4622
rect 15948 4593 15976 6802
rect 15844 4558 15896 4564
rect 15934 4584 15990 4593
rect 15934 4519 15990 4528
rect 15936 4480 15988 4486
rect 15936 4422 15988 4428
rect 15752 4072 15804 4078
rect 15752 4014 15804 4020
rect 15844 3936 15896 3942
rect 15844 3878 15896 3884
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 15672 3194 15700 3538
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 15568 2848 15620 2854
rect 15568 2790 15620 2796
rect 15856 480 15884 3878
rect 15948 2990 15976 4422
rect 15936 2984 15988 2990
rect 15936 2926 15988 2932
rect 16040 2650 16068 13246
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 16132 12374 16160 12922
rect 16224 12889 16252 13767
rect 16210 12880 16266 12889
rect 16210 12815 16266 12824
rect 16212 12776 16264 12782
rect 16212 12718 16264 12724
rect 16120 12368 16172 12374
rect 16120 12310 16172 12316
rect 16224 11762 16252 12718
rect 16212 11756 16264 11762
rect 16212 11698 16264 11704
rect 16224 10674 16252 11698
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16120 10600 16172 10606
rect 16120 10542 16172 10548
rect 16132 10441 16160 10542
rect 16118 10432 16174 10441
rect 16118 10367 16174 10376
rect 16212 10056 16264 10062
rect 16212 9998 16264 10004
rect 16224 9738 16252 9998
rect 16316 9994 16344 16934
rect 16408 16590 16436 17070
rect 16500 16658 16528 17478
rect 16488 16652 16540 16658
rect 16488 16594 16540 16600
rect 16396 16584 16448 16590
rect 16396 16526 16448 16532
rect 16408 16114 16436 16526
rect 16488 16244 16540 16250
rect 16488 16186 16540 16192
rect 16396 16108 16448 16114
rect 16396 16050 16448 16056
rect 16500 15570 16528 16186
rect 16488 15564 16540 15570
rect 16488 15506 16540 15512
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 16408 12986 16436 13466
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16592 12374 16620 18770
rect 16684 18154 16712 18906
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 16672 18148 16724 18154
rect 16672 18090 16724 18096
rect 16672 17740 16724 17746
rect 16672 17682 16724 17688
rect 16684 14482 16712 17682
rect 16776 17134 16804 18702
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 16764 14816 16816 14822
rect 16764 14758 16816 14764
rect 16672 14476 16724 14482
rect 16672 14418 16724 14424
rect 16670 14376 16726 14385
rect 16670 14311 16726 14320
rect 16684 12646 16712 14311
rect 16776 13530 16804 14758
rect 16764 13524 16816 13530
rect 16764 13466 16816 13472
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16776 12986 16804 13262
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 16764 12844 16816 12850
rect 16764 12786 16816 12792
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 16580 12368 16632 12374
rect 16580 12310 16632 12316
rect 16592 11744 16620 12310
rect 16500 11716 16620 11744
rect 16500 11558 16528 11716
rect 16580 11620 16632 11626
rect 16580 11562 16632 11568
rect 16488 11552 16540 11558
rect 16488 11494 16540 11500
rect 16396 11144 16448 11150
rect 16396 11086 16448 11092
rect 16408 10792 16436 11086
rect 16488 11076 16540 11082
rect 16488 11018 16540 11024
rect 16500 10962 16528 11018
rect 16592 10962 16620 11562
rect 16670 11248 16726 11257
rect 16670 11183 16726 11192
rect 16500 10934 16620 10962
rect 16488 10804 16540 10810
rect 16408 10764 16488 10792
rect 16488 10746 16540 10752
rect 16396 10532 16448 10538
rect 16396 10474 16448 10480
rect 16304 9988 16356 9994
rect 16304 9930 16356 9936
rect 16132 9710 16252 9738
rect 16132 9518 16160 9710
rect 16212 9648 16264 9654
rect 16212 9590 16264 9596
rect 16120 9512 16172 9518
rect 16120 9454 16172 9460
rect 16224 8634 16252 9590
rect 16408 9450 16436 10474
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16500 9586 16528 9998
rect 16488 9580 16540 9586
rect 16488 9522 16540 9528
rect 16396 9444 16448 9450
rect 16396 9386 16448 9392
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16316 9110 16344 9318
rect 16500 9178 16528 9522
rect 16488 9172 16540 9178
rect 16488 9114 16540 9120
rect 16304 9104 16356 9110
rect 16304 9046 16356 9052
rect 16592 8922 16620 10934
rect 16684 9081 16712 11183
rect 16776 10130 16804 12786
rect 16764 10124 16816 10130
rect 16764 10066 16816 10072
rect 16764 9716 16816 9722
rect 16764 9658 16816 9664
rect 16670 9072 16726 9081
rect 16670 9007 16726 9016
rect 16776 9024 16804 9658
rect 16868 9160 16896 19246
rect 16960 18970 16988 22320
rect 17512 20058 17540 22320
rect 17958 20632 18014 20641
rect 17958 20567 18014 20576
rect 17500 20052 17552 20058
rect 17500 19994 17552 20000
rect 17132 19916 17184 19922
rect 17132 19858 17184 19864
rect 16948 18964 17000 18970
rect 16948 18906 17000 18912
rect 17040 18760 17092 18766
rect 17040 18702 17092 18708
rect 17052 18426 17080 18702
rect 17040 18420 17092 18426
rect 17040 18362 17092 18368
rect 16948 17604 17000 17610
rect 16948 17546 17000 17552
rect 16960 16658 16988 17546
rect 17040 16720 17092 16726
rect 17040 16662 17092 16668
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 16948 16448 17000 16454
rect 16948 16390 17000 16396
rect 16960 15609 16988 16390
rect 17052 16046 17080 16662
rect 17040 16040 17092 16046
rect 17040 15982 17092 15988
rect 16946 15600 17002 15609
rect 16946 15535 17002 15544
rect 16960 12782 16988 15535
rect 17144 12850 17172 19858
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 17316 19236 17368 19242
rect 17316 19178 17368 19184
rect 17328 18834 17356 19178
rect 17316 18828 17368 18834
rect 17316 18770 17368 18776
rect 17316 15020 17368 15026
rect 17316 14962 17368 14968
rect 17224 14816 17276 14822
rect 17224 14758 17276 14764
rect 17236 13326 17264 14758
rect 17328 14550 17356 14962
rect 17316 14544 17368 14550
rect 17316 14486 17368 14492
rect 17328 14414 17356 14486
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 17328 14074 17356 14350
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 17328 12889 17356 13874
rect 17314 12880 17370 12889
rect 17132 12844 17184 12850
rect 17314 12815 17370 12824
rect 17132 12786 17184 12792
rect 16948 12776 17000 12782
rect 17420 12730 17448 19790
rect 17972 19718 18000 20567
rect 18064 20058 18092 22320
rect 18510 21176 18566 21185
rect 18510 21111 18566 21120
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 17960 19712 18012 19718
rect 17960 19654 18012 19660
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 17868 19304 17920 19310
rect 17868 19246 17920 19252
rect 17590 18728 17646 18737
rect 17590 18663 17646 18672
rect 17500 15564 17552 15570
rect 17500 15506 17552 15512
rect 17512 14278 17540 15506
rect 17604 14385 17632 18663
rect 17776 17060 17828 17066
rect 17776 17002 17828 17008
rect 17788 16250 17816 17002
rect 17776 16244 17828 16250
rect 17776 16186 17828 16192
rect 17776 16108 17828 16114
rect 17776 16050 17828 16056
rect 17788 15706 17816 16050
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 17590 14376 17646 14385
rect 17590 14311 17646 14320
rect 17684 14340 17736 14346
rect 17684 14282 17736 14288
rect 17500 14272 17552 14278
rect 17500 14214 17552 14220
rect 17512 13326 17540 14214
rect 17592 14000 17644 14006
rect 17696 13977 17724 14282
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 17592 13942 17644 13948
rect 17682 13968 17738 13977
rect 17500 13320 17552 13326
rect 17604 13297 17632 13942
rect 17682 13903 17738 13912
rect 17684 13728 17736 13734
rect 17684 13670 17736 13676
rect 17696 13326 17724 13670
rect 17788 13530 17816 14214
rect 17776 13524 17828 13530
rect 17776 13466 17828 13472
rect 17776 13388 17828 13394
rect 17776 13330 17828 13336
rect 17684 13320 17736 13326
rect 17500 13262 17552 13268
rect 17590 13288 17646 13297
rect 17684 13262 17736 13268
rect 17590 13223 17646 13232
rect 17592 12776 17644 12782
rect 16948 12718 17000 12724
rect 17144 12702 17448 12730
rect 17498 12744 17554 12753
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16960 10266 16988 11494
rect 16948 10260 17000 10266
rect 16948 10202 17000 10208
rect 17040 10192 17092 10198
rect 17144 10180 17172 12702
rect 17592 12718 17644 12724
rect 17498 12679 17554 12688
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 17236 12186 17264 12582
rect 17408 12436 17460 12442
rect 17408 12378 17460 12384
rect 17420 12345 17448 12378
rect 17406 12336 17462 12345
rect 17406 12271 17462 12280
rect 17236 12158 17448 12186
rect 17224 12096 17276 12102
rect 17224 12038 17276 12044
rect 17236 11830 17264 12038
rect 17224 11824 17276 11830
rect 17224 11766 17276 11772
rect 17236 11286 17264 11766
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 17420 11506 17448 12158
rect 17512 11626 17540 12679
rect 17500 11620 17552 11626
rect 17500 11562 17552 11568
rect 17328 11354 17356 11494
rect 17420 11478 17540 11506
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17224 11280 17276 11286
rect 17224 11222 17276 11228
rect 17408 11212 17460 11218
rect 17408 11154 17460 11160
rect 17420 11098 17448 11154
rect 17092 10152 17172 10180
rect 17328 11070 17448 11098
rect 17040 10134 17092 10140
rect 16868 9132 17172 9160
rect 16948 9036 17000 9042
rect 16776 8996 16896 9024
rect 16592 8894 16804 8922
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16120 8356 16172 8362
rect 16120 8298 16172 8304
rect 16132 8090 16160 8298
rect 16120 8084 16172 8090
rect 16120 8026 16172 8032
rect 16120 6996 16172 7002
rect 16120 6938 16172 6944
rect 16132 6066 16160 6938
rect 16224 6866 16252 8570
rect 16578 8528 16634 8537
rect 16304 8492 16356 8498
rect 16578 8463 16580 8472
rect 16304 8434 16356 8440
rect 16632 8463 16634 8472
rect 16580 8434 16632 8440
rect 16316 8378 16344 8434
rect 16776 8430 16804 8894
rect 16488 8424 16540 8430
rect 16316 8350 16436 8378
rect 16488 8366 16540 8372
rect 16764 8424 16816 8430
rect 16764 8366 16816 8372
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16316 7002 16344 7142
rect 16304 6996 16356 7002
rect 16304 6938 16356 6944
rect 16212 6860 16264 6866
rect 16212 6802 16264 6808
rect 16132 6038 16344 6066
rect 16120 3664 16172 3670
rect 16120 3606 16172 3612
rect 16132 2854 16160 3606
rect 16316 3398 16344 6038
rect 16408 5846 16436 8350
rect 16500 7993 16528 8366
rect 16580 8356 16632 8362
rect 16632 8316 16712 8344
rect 16580 8298 16632 8304
rect 16486 7984 16542 7993
rect 16684 7970 16712 8316
rect 16486 7919 16542 7928
rect 16580 7948 16632 7954
rect 16684 7942 16804 7970
rect 16868 7954 16896 8996
rect 16948 8978 17000 8984
rect 16960 8537 16988 8978
rect 17040 8560 17092 8566
rect 16946 8528 17002 8537
rect 17040 8502 17092 8508
rect 16946 8463 17002 8472
rect 16580 7890 16632 7896
rect 16592 7834 16620 7890
rect 16488 7812 16540 7818
rect 16592 7806 16712 7834
rect 16488 7754 16540 7760
rect 16500 7546 16528 7754
rect 16580 7744 16632 7750
rect 16580 7686 16632 7692
rect 16488 7540 16540 7546
rect 16488 7482 16540 7488
rect 16592 7342 16620 7686
rect 16684 7410 16712 7806
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16580 7336 16632 7342
rect 16580 7278 16632 7284
rect 16776 6730 16804 7942
rect 16856 7948 16908 7954
rect 16856 7890 16908 7896
rect 16960 7546 16988 8463
rect 17052 8090 17080 8502
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 16764 6724 16816 6730
rect 16764 6666 16816 6672
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16500 5914 16528 6258
rect 16948 6248 17000 6254
rect 16948 6190 17000 6196
rect 16488 5908 16540 5914
rect 16488 5850 16540 5856
rect 16396 5840 16448 5846
rect 16396 5782 16448 5788
rect 16500 5166 16528 5850
rect 16960 5846 16988 6190
rect 17040 6112 17092 6118
rect 17040 6054 17092 6060
rect 16948 5840 17000 5846
rect 16948 5782 17000 5788
rect 16960 5370 16988 5782
rect 16948 5364 17000 5370
rect 16948 5306 17000 5312
rect 16488 5160 16540 5166
rect 16488 5102 16540 5108
rect 17052 4826 17080 6054
rect 17040 4820 17092 4826
rect 17040 4762 17092 4768
rect 16948 4616 17000 4622
rect 16948 4558 17000 4564
rect 16764 4004 16816 4010
rect 16764 3946 16816 3952
rect 16856 4004 16908 4010
rect 16856 3946 16908 3952
rect 16304 3392 16356 3398
rect 16304 3334 16356 3340
rect 16120 2848 16172 2854
rect 16120 2790 16172 2796
rect 16028 2644 16080 2650
rect 16028 2586 16080 2592
rect 16132 2446 16160 2790
rect 16316 2446 16344 3334
rect 16776 2514 16804 3946
rect 16868 3738 16896 3946
rect 16856 3732 16908 3738
rect 16856 3674 16908 3680
rect 16856 3120 16908 3126
rect 16856 3062 16908 3068
rect 16764 2508 16816 2514
rect 16764 2450 16816 2456
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 16396 2304 16448 2310
rect 16396 2246 16448 2252
rect 16408 480 16436 2246
rect 16868 626 16896 3062
rect 16960 2990 16988 4558
rect 17144 3194 17172 9132
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 17236 4078 17264 8570
rect 17328 6458 17356 11070
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 17420 7954 17448 8434
rect 17512 8294 17540 11478
rect 17604 10742 17632 12718
rect 17696 11914 17724 13262
rect 17788 13161 17816 13330
rect 17774 13152 17830 13161
rect 17774 13087 17830 13096
rect 17788 12617 17816 13087
rect 17774 12608 17830 12617
rect 17774 12543 17830 12552
rect 17696 11886 17816 11914
rect 17684 11756 17736 11762
rect 17684 11698 17736 11704
rect 17696 11082 17724 11698
rect 17684 11076 17736 11082
rect 17684 11018 17736 11024
rect 17592 10736 17644 10742
rect 17592 10678 17644 10684
rect 17696 10674 17724 11018
rect 17684 10668 17736 10674
rect 17684 10610 17736 10616
rect 17682 10568 17738 10577
rect 17682 10503 17738 10512
rect 17592 9920 17644 9926
rect 17592 9862 17644 9868
rect 17500 8288 17552 8294
rect 17498 8256 17500 8265
rect 17552 8256 17554 8265
rect 17498 8191 17554 8200
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 17500 7744 17552 7750
rect 17500 7686 17552 7692
rect 17408 7472 17460 7478
rect 17408 7414 17460 7420
rect 17316 6452 17368 6458
rect 17316 6394 17368 6400
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 17328 4690 17356 5306
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17316 4548 17368 4554
rect 17316 4490 17368 4496
rect 17328 4282 17356 4490
rect 17316 4276 17368 4282
rect 17316 4218 17368 4224
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 17224 3664 17276 3670
rect 17224 3606 17276 3612
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 17236 3058 17264 3606
rect 17224 3052 17276 3058
rect 17224 2994 17276 3000
rect 16948 2984 17000 2990
rect 16948 2926 17000 2932
rect 17040 2848 17092 2854
rect 17040 2790 17092 2796
rect 17052 2378 17080 2790
rect 17328 2514 17356 4218
rect 17420 2514 17448 7414
rect 17512 6798 17540 7686
rect 17604 6866 17632 9862
rect 17592 6860 17644 6866
rect 17592 6802 17644 6808
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17604 6254 17632 6802
rect 17592 6248 17644 6254
rect 17592 6190 17644 6196
rect 17696 4010 17724 10503
rect 17788 6798 17816 11886
rect 17776 6792 17828 6798
rect 17776 6734 17828 6740
rect 17684 4004 17736 4010
rect 17684 3946 17736 3952
rect 17696 3126 17724 3946
rect 17684 3120 17736 3126
rect 17684 3062 17736 3068
rect 17788 2582 17816 6734
rect 17880 4826 17908 19246
rect 18524 18970 18552 21111
rect 18616 18970 18644 22320
rect 18696 19916 18748 19922
rect 18696 19858 18748 19864
rect 18512 18964 18564 18970
rect 18512 18906 18564 18912
rect 18604 18964 18656 18970
rect 18604 18906 18656 18912
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 17960 18352 18012 18358
rect 18708 18329 18736 19858
rect 19076 19292 19104 22471
rect 19154 22320 19210 22800
rect 19706 22320 19762 22800
rect 20258 22320 20314 22800
rect 20810 22320 20866 22800
rect 21362 22320 21418 22800
rect 21914 22320 21970 22800
rect 22466 22320 22522 22800
rect 19168 20058 19196 22320
rect 19246 21584 19302 21593
rect 19246 21519 19302 21528
rect 19156 20052 19208 20058
rect 19156 19994 19208 20000
rect 19156 19304 19208 19310
rect 18970 19272 19026 19281
rect 19076 19264 19156 19292
rect 19156 19246 19208 19252
rect 18970 19207 19026 19216
rect 18880 18964 18932 18970
rect 18880 18906 18932 18912
rect 18892 18873 18920 18906
rect 18878 18864 18934 18873
rect 18788 18828 18840 18834
rect 18878 18799 18934 18808
rect 18788 18770 18840 18776
rect 17960 18294 18012 18300
rect 18694 18320 18750 18329
rect 17972 17134 18000 18294
rect 18694 18255 18750 18264
rect 18602 18184 18658 18193
rect 18602 18119 18658 18128
rect 18616 18086 18644 18119
rect 18144 18080 18196 18086
rect 18144 18022 18196 18028
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 18696 18080 18748 18086
rect 18696 18022 18748 18028
rect 18156 17882 18184 18022
rect 18144 17876 18196 17882
rect 18144 17818 18196 17824
rect 18512 17604 18564 17610
rect 18512 17546 18564 17552
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 18052 17264 18104 17270
rect 18052 17206 18104 17212
rect 17960 17128 18012 17134
rect 17960 17070 18012 17076
rect 17960 16992 18012 16998
rect 17958 16960 17960 16969
rect 18012 16960 18014 16969
rect 17958 16895 18014 16904
rect 17960 16652 18012 16658
rect 17960 16594 18012 16600
rect 17972 16017 18000 16594
rect 18064 16561 18092 17206
rect 18524 17066 18552 17546
rect 18512 17060 18564 17066
rect 18512 17002 18564 17008
rect 18708 16674 18736 18022
rect 18616 16658 18736 16674
rect 18604 16652 18736 16658
rect 18656 16646 18736 16652
rect 18604 16594 18656 16600
rect 18696 16584 18748 16590
rect 18050 16552 18106 16561
rect 18696 16526 18748 16532
rect 18050 16487 18106 16496
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 18052 16108 18104 16114
rect 18052 16050 18104 16056
rect 17958 16008 18014 16017
rect 17958 15943 18014 15952
rect 18064 15484 18092 16050
rect 18708 15910 18736 16526
rect 18696 15904 18748 15910
rect 18696 15846 18748 15852
rect 18708 15638 18736 15846
rect 18696 15632 18748 15638
rect 18696 15574 18748 15580
rect 18144 15496 18196 15502
rect 18064 15456 18144 15484
rect 18144 15438 18196 15444
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 17960 15088 18012 15094
rect 17960 15030 18012 15036
rect 17972 14657 18000 15030
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 17958 14648 18014 14657
rect 17958 14583 18014 14592
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 18512 14476 18564 14482
rect 18512 14418 18564 14424
rect 17972 14074 18000 14418
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 18052 13932 18104 13938
rect 18052 13874 18104 13880
rect 18420 13932 18472 13938
rect 18420 13874 18472 13880
rect 17958 13696 18014 13705
rect 17958 13631 18014 13640
rect 17972 13462 18000 13631
rect 17960 13456 18012 13462
rect 17960 13398 18012 13404
rect 18064 13274 18092 13874
rect 18432 13818 18460 13874
rect 18340 13802 18460 13818
rect 18328 13796 18460 13802
rect 18380 13790 18460 13796
rect 18328 13738 18380 13744
rect 18432 13410 18460 13790
rect 18524 13530 18552 14418
rect 18616 14074 18644 14962
rect 18696 14816 18748 14822
rect 18696 14758 18748 14764
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18604 13796 18656 13802
rect 18604 13738 18656 13744
rect 18616 13530 18644 13738
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18604 13524 18656 13530
rect 18604 13466 18656 13472
rect 18432 13382 18552 13410
rect 18524 13326 18552 13382
rect 18604 13388 18656 13394
rect 18604 13330 18656 13336
rect 17972 13246 18092 13274
rect 18512 13320 18564 13326
rect 18512 13262 18564 13268
rect 17972 12170 18000 13246
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 18052 12232 18104 12238
rect 18050 12200 18052 12209
rect 18104 12200 18106 12209
rect 17960 12164 18012 12170
rect 18050 12135 18106 12144
rect 17960 12106 18012 12112
rect 18432 12084 18460 12718
rect 18524 12646 18552 13262
rect 18512 12640 18564 12646
rect 18512 12582 18564 12588
rect 18512 12436 18564 12442
rect 18616 12424 18644 13330
rect 18564 12396 18644 12424
rect 18512 12378 18564 12384
rect 18432 12056 18552 12084
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 17958 11384 18014 11393
rect 17958 11319 18014 11328
rect 17972 11218 18000 11319
rect 18420 11280 18472 11286
rect 18420 11222 18472 11228
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 18432 11121 18460 11222
rect 18418 11112 18474 11121
rect 17972 11082 18092 11098
rect 17972 11076 18104 11082
rect 17972 11070 18052 11076
rect 17972 10198 18000 11070
rect 18418 11047 18474 11056
rect 18052 11018 18104 11024
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 18524 10810 18552 12056
rect 18604 11212 18656 11218
rect 18604 11154 18656 11160
rect 18512 10804 18564 10810
rect 18512 10746 18564 10752
rect 18328 10736 18380 10742
rect 18328 10678 18380 10684
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 17960 10192 18012 10198
rect 17960 10134 18012 10140
rect 17960 10056 18012 10062
rect 18064 10010 18092 10406
rect 18340 10033 18368 10678
rect 18616 10674 18644 11154
rect 18604 10668 18656 10674
rect 18604 10610 18656 10616
rect 18512 10056 18564 10062
rect 18012 10004 18092 10010
rect 17960 9998 18092 10004
rect 17972 9982 18092 9998
rect 18326 10024 18382 10033
rect 17972 9450 18000 9982
rect 18512 9998 18564 10004
rect 18326 9959 18382 9968
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 18144 9512 18196 9518
rect 18144 9454 18196 9460
rect 17960 9444 18012 9450
rect 17960 9386 18012 9392
rect 18156 9110 18184 9454
rect 18524 9178 18552 9998
rect 18604 9988 18656 9994
rect 18604 9930 18656 9936
rect 18512 9172 18564 9178
rect 18512 9114 18564 9120
rect 18144 9104 18196 9110
rect 18144 9046 18196 9052
rect 18326 9072 18382 9081
rect 18326 9007 18328 9016
rect 18380 9007 18382 9016
rect 18328 8978 18380 8984
rect 18616 8945 18644 9930
rect 18602 8936 18658 8945
rect 18512 8900 18564 8906
rect 18602 8871 18658 8880
rect 18512 8842 18564 8848
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 17972 8537 18000 8774
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 18524 8673 18552 8842
rect 18604 8832 18656 8838
rect 18604 8774 18656 8780
rect 18510 8664 18566 8673
rect 18616 8634 18644 8774
rect 18510 8599 18566 8608
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18328 8560 18380 8566
rect 17958 8528 18014 8537
rect 18328 8502 18380 8508
rect 17958 8463 18014 8472
rect 18340 8401 18368 8502
rect 18326 8392 18382 8401
rect 18326 8327 18382 8336
rect 18602 8392 18658 8401
rect 18602 8327 18604 8336
rect 18656 8327 18658 8336
rect 18604 8298 18656 8304
rect 17958 8120 18014 8129
rect 17958 8055 18014 8064
rect 18512 8084 18564 8090
rect 17972 8022 18000 8055
rect 18512 8026 18564 8032
rect 17960 8016 18012 8022
rect 17960 7958 18012 7964
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 18236 7472 18288 7478
rect 18236 7414 18288 7420
rect 18052 7200 18104 7206
rect 18052 7142 18104 7148
rect 18064 6934 18092 7142
rect 18248 7002 18276 7414
rect 18524 7206 18552 8026
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 18616 7410 18644 7890
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18512 7200 18564 7206
rect 18512 7142 18564 7148
rect 18236 6996 18288 7002
rect 18236 6938 18288 6944
rect 18052 6928 18104 6934
rect 18052 6870 18104 6876
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 18524 6225 18552 7142
rect 18616 6798 18644 7346
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 18510 6216 18566 6225
rect 18510 6151 18566 6160
rect 18616 5914 18644 6734
rect 18708 6458 18736 14758
rect 18800 12918 18828 18770
rect 18880 18284 18932 18290
rect 18880 18226 18932 18232
rect 18892 17814 18920 18226
rect 18880 17808 18932 17814
rect 18880 17750 18932 17756
rect 18984 16794 19012 19207
rect 19260 19174 19288 21519
rect 19720 20058 19748 22320
rect 20166 20224 20222 20233
rect 20166 20159 20222 20168
rect 20180 20058 20208 20159
rect 19708 20052 19760 20058
rect 19708 19994 19760 20000
rect 20168 20052 20220 20058
rect 20168 19994 20220 20000
rect 20272 19990 20300 22320
rect 20626 22128 20682 22137
rect 20626 22063 20682 22072
rect 20640 20058 20668 22063
rect 20628 20052 20680 20058
rect 20628 19994 20680 20000
rect 20260 19984 20312 19990
rect 20260 19926 20312 19932
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19984 19916 20036 19922
rect 19984 19858 20036 19864
rect 20168 19916 20220 19922
rect 20168 19858 20220 19864
rect 19064 19168 19116 19174
rect 19064 19110 19116 19116
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 19076 18290 19104 19110
rect 19154 18864 19210 18873
rect 19154 18799 19210 18808
rect 19168 18426 19196 18799
rect 19248 18624 19300 18630
rect 19248 18566 19300 18572
rect 19156 18420 19208 18426
rect 19156 18362 19208 18368
rect 19260 18329 19288 18566
rect 19246 18320 19302 18329
rect 19064 18284 19116 18290
rect 19246 18255 19302 18264
rect 19064 18226 19116 18232
rect 19444 18034 19472 19858
rect 19996 18902 20024 19858
rect 20076 19236 20128 19242
rect 20076 19178 20128 19184
rect 19984 18896 20036 18902
rect 19984 18838 20036 18844
rect 19524 18828 19576 18834
rect 19524 18770 19576 18776
rect 19708 18828 19760 18834
rect 19708 18770 19760 18776
rect 19168 18006 19472 18034
rect 19168 17746 19196 18006
rect 19246 17912 19302 17921
rect 19246 17847 19302 17856
rect 19156 17740 19208 17746
rect 19156 17682 19208 17688
rect 18972 16788 19024 16794
rect 18972 16730 19024 16736
rect 18984 15473 19012 16730
rect 19064 16652 19116 16658
rect 19064 16594 19116 16600
rect 18970 15464 19026 15473
rect 18970 15399 19026 15408
rect 18972 15020 19024 15026
rect 18972 14962 19024 14968
rect 18880 14884 18932 14890
rect 18880 14826 18932 14832
rect 18892 13530 18920 14826
rect 18984 13841 19012 14962
rect 19076 14521 19104 16594
rect 19260 15706 19288 17847
rect 19432 17536 19484 17542
rect 19432 17478 19484 17484
rect 19444 17134 19472 17478
rect 19432 17128 19484 17134
rect 19432 17070 19484 17076
rect 19536 17066 19564 18770
rect 19614 18728 19670 18737
rect 19614 18663 19670 18672
rect 19628 17678 19656 18663
rect 19616 17672 19668 17678
rect 19616 17614 19668 17620
rect 19524 17060 19576 17066
rect 19524 17002 19576 17008
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19352 16590 19380 16934
rect 19340 16584 19392 16590
rect 19340 16526 19392 16532
rect 19352 15978 19380 16526
rect 19340 15972 19392 15978
rect 19340 15914 19392 15920
rect 19616 15972 19668 15978
rect 19616 15914 19668 15920
rect 19248 15700 19300 15706
rect 19248 15642 19300 15648
rect 19156 15360 19208 15366
rect 19156 15302 19208 15308
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 19062 14512 19118 14521
rect 19168 14482 19196 15302
rect 19246 15056 19302 15065
rect 19246 14991 19302 15000
rect 19260 14618 19288 14991
rect 19444 14890 19472 15302
rect 19524 15156 19576 15162
rect 19524 15098 19576 15104
rect 19432 14884 19484 14890
rect 19432 14826 19484 14832
rect 19248 14612 19300 14618
rect 19248 14554 19300 14560
rect 19062 14447 19118 14456
rect 19156 14476 19208 14482
rect 19156 14418 19208 14424
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19154 14104 19210 14113
rect 19154 14039 19210 14048
rect 19064 13864 19116 13870
rect 18970 13832 19026 13841
rect 19064 13806 19116 13812
rect 18970 13767 19026 13776
rect 18880 13524 18932 13530
rect 18880 13466 18932 13472
rect 18788 12912 18840 12918
rect 18788 12854 18840 12860
rect 18880 12776 18932 12782
rect 18984 12764 19012 13767
rect 19076 13258 19104 13806
rect 19064 13252 19116 13258
rect 19064 13194 19116 13200
rect 18932 12736 19012 12764
rect 18880 12718 18932 12724
rect 18786 12608 18842 12617
rect 18786 12543 18842 12552
rect 18800 11676 18828 12543
rect 18892 12442 18920 12718
rect 18880 12436 18932 12442
rect 18880 12378 18932 12384
rect 18880 12300 18932 12306
rect 18880 12242 18932 12248
rect 18892 12102 18920 12242
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18892 11830 18920 12038
rect 19168 11898 19196 14039
rect 19352 13870 19380 14282
rect 19444 13938 19472 14826
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19248 13728 19300 13734
rect 19248 13670 19300 13676
rect 19156 11892 19208 11898
rect 19156 11834 19208 11840
rect 18880 11824 18932 11830
rect 18880 11766 18932 11772
rect 18800 11648 18920 11676
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18800 8090 18828 11494
rect 18788 8084 18840 8090
rect 18788 8026 18840 8032
rect 18786 7576 18842 7585
rect 18786 7511 18842 7520
rect 18800 7274 18828 7511
rect 18788 7268 18840 7274
rect 18788 7210 18840 7216
rect 18696 6452 18748 6458
rect 18696 6394 18748 6400
rect 18788 6384 18840 6390
rect 18788 6326 18840 6332
rect 18696 6112 18748 6118
rect 18696 6054 18748 6060
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 18156 5817 18184 5850
rect 18142 5808 18198 5817
rect 17960 5772 18012 5778
rect 18142 5743 18198 5752
rect 17960 5714 18012 5720
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 17972 4758 18000 5714
rect 18512 5568 18564 5574
rect 18512 5510 18564 5516
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 18524 5234 18552 5510
rect 18512 5228 18564 5234
rect 18564 5188 18644 5216
rect 18512 5170 18564 5176
rect 18144 5024 18196 5030
rect 18144 4966 18196 4972
rect 18156 4826 18184 4966
rect 18144 4820 18196 4826
rect 18144 4762 18196 4768
rect 17960 4752 18012 4758
rect 17960 4694 18012 4700
rect 17960 4616 18012 4622
rect 17960 4558 18012 4564
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 17880 3074 17908 3878
rect 17972 3194 18000 4558
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 18616 4078 18644 5188
rect 18708 4758 18736 6054
rect 18800 4865 18828 6326
rect 18786 4856 18842 4865
rect 18786 4791 18842 4800
rect 18696 4752 18748 4758
rect 18696 4694 18748 4700
rect 18604 4072 18656 4078
rect 18604 4014 18656 4020
rect 18696 4004 18748 4010
rect 18696 3946 18748 3952
rect 18708 3738 18736 3946
rect 18696 3732 18748 3738
rect 18696 3674 18748 3680
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 18510 3224 18566 3233
rect 17960 3188 18012 3194
rect 18510 3159 18566 3168
rect 17960 3130 18012 3136
rect 18418 3088 18474 3097
rect 17880 3046 18000 3074
rect 17776 2576 17828 2582
rect 17776 2518 17828 2524
rect 17316 2508 17368 2514
rect 17316 2450 17368 2456
rect 17408 2508 17460 2514
rect 17408 2450 17460 2456
rect 17040 2372 17092 2378
rect 17040 2314 17092 2320
rect 17500 2304 17552 2310
rect 17500 2246 17552 2252
rect 16868 598 16988 626
rect 16960 480 16988 598
rect 17512 480 17540 2246
rect 17972 1306 18000 3046
rect 18524 3058 18552 3159
rect 18708 3058 18736 3674
rect 18418 3023 18474 3032
rect 18512 3052 18564 3058
rect 18432 2990 18460 3023
rect 18512 2994 18564 3000
rect 18696 3052 18748 3058
rect 18696 2994 18748 3000
rect 18420 2984 18472 2990
rect 18524 2961 18552 2994
rect 18420 2926 18472 2932
rect 18510 2952 18566 2961
rect 18510 2887 18566 2896
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 18156 2553 18184 2586
rect 18142 2544 18198 2553
rect 18142 2479 18198 2488
rect 18696 2372 18748 2378
rect 18696 2314 18748 2320
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 18512 2100 18564 2106
rect 18512 2042 18564 2048
rect 18524 1601 18552 2042
rect 18510 1592 18566 1601
rect 18510 1527 18566 1536
rect 17972 1278 18092 1306
rect 18064 480 18092 1278
rect 18708 1170 18736 2314
rect 18616 1142 18736 1170
rect 18616 480 18644 1142
rect 294 0 350 480
rect 846 0 902 480
rect 1398 0 1454 480
rect 1950 0 2006 480
rect 2502 0 2558 480
rect 3054 0 3110 480
rect 3606 0 3662 480
rect 4158 0 4214 480
rect 4710 0 4766 480
rect 5262 0 5318 480
rect 5814 0 5870 480
rect 6366 0 6422 480
rect 6918 0 6974 480
rect 7470 0 7526 480
rect 8022 0 8078 480
rect 8574 0 8630 480
rect 9126 0 9182 480
rect 9678 0 9734 480
rect 10230 0 10286 480
rect 10782 0 10838 480
rect 11334 0 11390 480
rect 11978 0 12034 480
rect 12530 0 12586 480
rect 13082 0 13138 480
rect 13634 0 13690 480
rect 14186 0 14242 480
rect 14738 0 14794 480
rect 15290 0 15346 480
rect 15842 0 15898 480
rect 16394 0 16450 480
rect 16946 0 17002 480
rect 17498 0 17554 480
rect 18050 0 18106 480
rect 18602 0 18658 480
rect 18892 241 18920 11648
rect 18972 11620 19024 11626
rect 18972 11562 19024 11568
rect 18984 9489 19012 11562
rect 19260 11354 19288 13670
rect 19536 13530 19564 15098
rect 19524 13524 19576 13530
rect 19524 13466 19576 13472
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19064 11280 19116 11286
rect 19064 11222 19116 11228
rect 19076 10713 19104 11222
rect 19340 11008 19392 11014
rect 19340 10950 19392 10956
rect 19246 10840 19302 10849
rect 19246 10775 19302 10784
rect 19062 10704 19118 10713
rect 19062 10639 19118 10648
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 19076 10266 19104 10406
rect 19064 10260 19116 10266
rect 19064 10202 19116 10208
rect 19064 10056 19116 10062
rect 19064 9998 19116 10004
rect 19076 9722 19104 9998
rect 19260 9926 19288 10775
rect 19352 10606 19380 10950
rect 19340 10600 19392 10606
rect 19340 10542 19392 10548
rect 19444 10538 19472 12242
rect 19628 11778 19656 15914
rect 19720 12102 19748 18770
rect 19984 18148 20036 18154
rect 19984 18090 20036 18096
rect 19996 17882 20024 18090
rect 19984 17876 20036 17882
rect 19984 17818 20036 17824
rect 19892 16652 19944 16658
rect 19892 16594 19944 16600
rect 19800 15904 19852 15910
rect 19800 15846 19852 15852
rect 19812 14618 19840 15846
rect 19904 15570 19932 16594
rect 20088 15910 20116 19178
rect 20180 15978 20208 19858
rect 20258 19816 20314 19825
rect 20258 19751 20314 19760
rect 20168 15972 20220 15978
rect 20168 15914 20220 15920
rect 20076 15904 20128 15910
rect 20076 15846 20128 15852
rect 20180 15638 20208 15914
rect 20168 15632 20220 15638
rect 20168 15574 20220 15580
rect 19892 15564 19944 15570
rect 19892 15506 19944 15512
rect 19892 14816 19944 14822
rect 19892 14758 19944 14764
rect 20168 14816 20220 14822
rect 20168 14758 20220 14764
rect 19800 14612 19852 14618
rect 19800 14554 19852 14560
rect 19800 14476 19852 14482
rect 19800 14418 19852 14424
rect 19812 14074 19840 14418
rect 19800 14068 19852 14074
rect 19800 14010 19852 14016
rect 19800 13864 19852 13870
rect 19800 13806 19852 13812
rect 19708 12096 19760 12102
rect 19708 12038 19760 12044
rect 19628 11750 19748 11778
rect 19616 11688 19668 11694
rect 19616 11630 19668 11636
rect 19628 10606 19656 11630
rect 19616 10600 19668 10606
rect 19616 10542 19668 10548
rect 19432 10532 19484 10538
rect 19432 10474 19484 10480
rect 19340 10464 19392 10470
rect 19340 10406 19392 10412
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 19064 9716 19116 9722
rect 19116 9676 19196 9704
rect 19064 9658 19116 9664
rect 18970 9480 19026 9489
rect 18970 9415 19026 9424
rect 18984 7342 19012 9415
rect 19168 9042 19196 9676
rect 19156 9036 19208 9042
rect 19076 8996 19156 9024
rect 19076 7954 19104 8996
rect 19156 8978 19208 8984
rect 19352 8548 19380 10406
rect 19628 10130 19656 10542
rect 19616 10124 19668 10130
rect 19616 10066 19668 10072
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19524 9376 19576 9382
rect 19524 9318 19576 9324
rect 19444 9110 19472 9318
rect 19432 9104 19484 9110
rect 19432 9046 19484 9052
rect 19352 8520 19463 8548
rect 19435 8344 19463 8520
rect 19536 8401 19564 9318
rect 19616 8628 19668 8634
rect 19616 8570 19668 8576
rect 19352 8316 19463 8344
rect 19522 8392 19578 8401
rect 19522 8327 19578 8336
rect 19352 8276 19380 8316
rect 19352 8248 19463 8276
rect 19435 8106 19463 8248
rect 19522 8256 19578 8265
rect 19522 8191 19578 8200
rect 19352 8078 19463 8106
rect 19064 7948 19116 7954
rect 19064 7890 19116 7896
rect 18972 7336 19024 7342
rect 18972 7278 19024 7284
rect 19156 7200 19208 7206
rect 19156 7142 19208 7148
rect 19246 7168 19302 7177
rect 18972 6792 19024 6798
rect 18972 6734 19024 6740
rect 18984 6254 19012 6734
rect 18972 6248 19024 6254
rect 18972 6190 19024 6196
rect 18984 5778 19012 6190
rect 18972 5772 19024 5778
rect 18972 5714 19024 5720
rect 18970 5672 19026 5681
rect 18970 5607 19026 5616
rect 18984 2514 19012 5607
rect 19168 4826 19196 7142
rect 19246 7103 19302 7112
rect 19260 6118 19288 7103
rect 19352 6254 19380 8078
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 19444 6458 19472 6802
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 19340 6248 19392 6254
rect 19340 6190 19392 6196
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 19260 4826 19288 6054
rect 19156 4820 19208 4826
rect 19156 4762 19208 4768
rect 19248 4820 19300 4826
rect 19248 4762 19300 4768
rect 19444 4622 19472 6394
rect 19156 4616 19208 4622
rect 19156 4558 19208 4564
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19064 4480 19116 4486
rect 19064 4422 19116 4428
rect 19076 3602 19104 4422
rect 19168 3942 19196 4558
rect 19536 4468 19564 8191
rect 19444 4440 19564 4468
rect 19156 3936 19208 3942
rect 19156 3878 19208 3884
rect 19064 3596 19116 3602
rect 19064 3538 19116 3544
rect 19444 2990 19472 4440
rect 19628 3602 19656 8570
rect 19720 5302 19748 11750
rect 19708 5296 19760 5302
rect 19708 5238 19760 5244
rect 19812 5098 19840 13806
rect 19904 10441 19932 14758
rect 20180 14414 20208 14758
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 20272 13682 20300 19751
rect 20626 19272 20682 19281
rect 20536 19236 20588 19242
rect 20626 19207 20682 19216
rect 20536 19178 20588 19184
rect 20444 17128 20496 17134
rect 20444 17070 20496 17076
rect 20352 16108 20404 16114
rect 20352 16050 20404 16056
rect 20364 15366 20392 16050
rect 20352 15360 20404 15366
rect 20352 15302 20404 15308
rect 20352 14408 20404 14414
rect 20352 14350 20404 14356
rect 20364 13802 20392 14350
rect 20456 14346 20484 17070
rect 20444 14340 20496 14346
rect 20444 14282 20496 14288
rect 20352 13796 20404 13802
rect 20352 13738 20404 13744
rect 20272 13654 20392 13682
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 19996 12782 20024 13262
rect 19984 12776 20036 12782
rect 19984 12718 20036 12724
rect 19996 12442 20024 12718
rect 20364 12442 20392 13654
rect 20444 13184 20496 13190
rect 20444 13126 20496 13132
rect 20456 12782 20484 13126
rect 20444 12776 20496 12782
rect 20444 12718 20496 12724
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 20352 12436 20404 12442
rect 20352 12378 20404 12384
rect 20352 12096 20404 12102
rect 20352 12038 20404 12044
rect 19984 11620 20036 11626
rect 19984 11562 20036 11568
rect 19996 10470 20024 11562
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 19984 10464 20036 10470
rect 19890 10432 19946 10441
rect 19984 10406 20036 10412
rect 19890 10367 19946 10376
rect 19904 7342 19932 10367
rect 20088 10198 20116 11086
rect 20076 10192 20128 10198
rect 19996 10152 20076 10180
rect 19996 9178 20024 10152
rect 20076 10134 20128 10140
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 19984 9172 20036 9178
rect 19984 9114 20036 9120
rect 19984 8832 20036 8838
rect 19984 8774 20036 8780
rect 19996 8634 20024 8774
rect 20074 8664 20130 8673
rect 19984 8628 20036 8634
rect 20074 8599 20130 8608
rect 19984 8570 20036 8576
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 19996 8090 20024 8434
rect 20088 8430 20116 8599
rect 20076 8424 20128 8430
rect 20076 8366 20128 8372
rect 20076 8288 20128 8294
rect 20076 8230 20128 8236
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 19892 7336 19944 7342
rect 19892 7278 19944 7284
rect 20088 6769 20116 8230
rect 20074 6760 20130 6769
rect 20074 6695 20130 6704
rect 20180 6610 20208 9658
rect 20364 8922 20392 12038
rect 20548 11082 20576 19178
rect 20640 14074 20668 19207
rect 20824 18698 20852 22320
rect 21376 18766 21404 22320
rect 21928 18970 21956 22320
rect 21916 18964 21968 18970
rect 21916 18906 21968 18912
rect 21364 18760 21416 18766
rect 21364 18702 21416 18708
rect 20812 18692 20864 18698
rect 20812 18634 20864 18640
rect 20812 18148 20864 18154
rect 20812 18090 20864 18096
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 20732 14958 20760 17138
rect 20824 15570 20852 18090
rect 21178 17368 21234 17377
rect 22480 17338 22508 22320
rect 21178 17303 21234 17312
rect 22468 17332 22520 17338
rect 20904 15972 20956 15978
rect 20904 15914 20956 15920
rect 20812 15564 20864 15570
rect 20812 15506 20864 15512
rect 20720 14952 20772 14958
rect 20720 14894 20772 14900
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 20824 11694 20852 13806
rect 20812 11688 20864 11694
rect 20812 11630 20864 11636
rect 20916 11506 20944 15914
rect 20996 15904 21048 15910
rect 20996 15846 21048 15852
rect 21008 15609 21036 15846
rect 20994 15600 21050 15609
rect 20994 15535 21050 15544
rect 21192 15162 21220 17303
rect 22468 17274 22520 17280
rect 21180 15156 21232 15162
rect 21180 15098 21232 15104
rect 20824 11478 20944 11506
rect 20536 11076 20588 11082
rect 20536 11018 20588 11024
rect 20444 10532 20496 10538
rect 20444 10474 20496 10480
rect 20456 10266 20484 10474
rect 20444 10260 20496 10266
rect 20444 10202 20496 10208
rect 20534 10024 20590 10033
rect 20534 9959 20590 9968
rect 20548 9586 20576 9959
rect 20824 9722 20852 11478
rect 20904 11212 20956 11218
rect 20904 11154 20956 11160
rect 20916 10266 20944 11154
rect 20904 10260 20956 10266
rect 20904 10202 20956 10208
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 20536 9580 20588 9586
rect 20536 9522 20588 9528
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 20364 8894 20576 8922
rect 20444 7404 20496 7410
rect 20444 7346 20496 7352
rect 20088 6582 20208 6610
rect 19892 6248 19944 6254
rect 19892 6190 19944 6196
rect 19904 5370 19932 6190
rect 19892 5364 19944 5370
rect 19892 5306 19944 5312
rect 19800 5092 19852 5098
rect 19800 5034 19852 5040
rect 19708 4684 19760 4690
rect 19708 4626 19760 4632
rect 19720 4282 19748 4626
rect 19800 4480 19852 4486
rect 19800 4422 19852 4428
rect 19708 4276 19760 4282
rect 19708 4218 19760 4224
rect 19812 4078 19840 4422
rect 19904 4214 19932 5306
rect 19892 4208 19944 4214
rect 19892 4150 19944 4156
rect 19800 4072 19852 4078
rect 19800 4014 19852 4020
rect 19616 3596 19668 3602
rect 19616 3538 19668 3544
rect 19524 3528 19576 3534
rect 20088 3505 20116 6582
rect 20456 6254 20484 7346
rect 20444 6248 20496 6254
rect 20444 6190 20496 6196
rect 20260 5568 20312 5574
rect 20260 5510 20312 5516
rect 20272 5166 20300 5510
rect 20548 5386 20576 8894
rect 20640 8498 20668 9522
rect 20904 9444 20956 9450
rect 20904 9386 20956 9392
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20640 8022 20668 8434
rect 20916 8090 20944 9386
rect 20904 8084 20956 8090
rect 20904 8026 20956 8032
rect 20628 8016 20680 8022
rect 20628 7958 20680 7964
rect 20640 7002 20668 7958
rect 20904 7268 20956 7274
rect 20904 7210 20956 7216
rect 20628 6996 20680 7002
rect 20628 6938 20680 6944
rect 20916 5914 20944 7210
rect 20904 5908 20956 5914
rect 20904 5850 20956 5856
rect 20456 5358 20576 5386
rect 20260 5160 20312 5166
rect 20312 5108 20392 5114
rect 20260 5102 20392 5108
rect 20272 5086 20392 5102
rect 20168 5024 20220 5030
rect 20168 4966 20220 4972
rect 20180 4146 20208 4966
rect 20364 4622 20392 5086
rect 20260 4616 20312 4622
rect 20260 4558 20312 4564
rect 20352 4616 20404 4622
rect 20352 4558 20404 4564
rect 20168 4140 20220 4146
rect 20168 4082 20220 4088
rect 20272 3913 20300 4558
rect 20456 4049 20484 5358
rect 20536 5296 20588 5302
rect 20536 5238 20588 5244
rect 20442 4040 20498 4049
rect 20442 3975 20498 3984
rect 20258 3904 20314 3913
rect 20258 3839 20314 3848
rect 20352 3528 20404 3534
rect 19524 3470 19576 3476
rect 20074 3496 20130 3505
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 19536 2514 19564 3470
rect 20352 3470 20404 3476
rect 20074 3431 20130 3440
rect 20260 3120 20312 3126
rect 20260 3062 20312 3068
rect 18972 2508 19024 2514
rect 18972 2450 19024 2456
rect 19524 2508 19576 2514
rect 19524 2450 19576 2456
rect 19248 2440 19300 2446
rect 19248 2382 19300 2388
rect 19064 2304 19116 2310
rect 19116 2264 19196 2292
rect 19064 2246 19116 2252
rect 19168 480 19196 2264
rect 19260 2009 19288 2382
rect 19616 2304 19668 2310
rect 19668 2264 19748 2292
rect 19616 2246 19668 2252
rect 19246 2000 19302 2009
rect 19246 1935 19302 1944
rect 19720 480 19748 2264
rect 20272 480 20300 3062
rect 20364 2514 20392 3470
rect 20548 2990 20576 5238
rect 20720 5092 20772 5098
rect 20720 5034 20772 5040
rect 20628 5024 20680 5030
rect 20628 4966 20680 4972
rect 20640 4554 20668 4966
rect 20628 4548 20680 4554
rect 20628 4490 20680 4496
rect 20732 4078 20760 5034
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 22468 3936 22520 3942
rect 22468 3878 22520 3884
rect 20536 2984 20588 2990
rect 20536 2926 20588 2932
rect 21364 2916 21416 2922
rect 21364 2858 21416 2864
rect 20352 2508 20404 2514
rect 20352 2450 20404 2456
rect 20812 2304 20864 2310
rect 20812 2246 20864 2252
rect 20824 480 20852 2246
rect 21376 480 21404 2858
rect 21916 2848 21968 2854
rect 21916 2790 21968 2796
rect 21928 480 21956 2790
rect 22480 480 22508 3878
rect 18878 232 18934 241
rect 18878 167 18934 176
rect 19154 0 19210 480
rect 19706 0 19762 480
rect 20258 0 20314 480
rect 20810 0 20866 480
rect 21362 0 21418 480
rect 21914 0 21970 480
rect 22466 0 22522 480
<< via2 >>
rect 19062 22480 19118 22536
rect 1398 18264 1454 18320
rect 2502 19216 2558 19272
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 3422 17176 3478 17232
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 8574 18672 8630 18728
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4066 5752 4122 5808
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 9862 19216 9918 19272
rect 10046 19216 10102 19272
rect 9770 18944 9826 19000
rect 9494 18400 9550 18456
rect 9586 18264 9642 18320
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 9402 16632 9458 16688
rect 10230 19080 10286 19136
rect 10322 16632 10378 16688
rect 10230 13504 10286 13560
rect 10782 17992 10838 18048
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 11242 16940 11244 16960
rect 11244 16940 11296 16960
rect 11296 16940 11298 16960
rect 11242 16904 11298 16940
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11518 13932 11574 13968
rect 11518 13912 11520 13932
rect 11520 13912 11572 13932
rect 11572 13912 11574 13932
rect 11886 18536 11942 18592
rect 11886 14184 11942 14240
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 10414 9560 10470 9616
rect 10138 9016 10194 9072
rect 10322 8336 10378 8392
rect 10690 4528 10746 4584
rect 9862 3032 9918 3088
rect 10782 3984 10838 4040
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11978 13368 12034 13424
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11334 7792 11390 7848
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 12254 18808 12310 18864
rect 12530 18264 12586 18320
rect 12346 16632 12402 16688
rect 12806 19116 12808 19136
rect 12808 19116 12860 19136
rect 12860 19116 12862 19136
rect 12806 19080 12862 19116
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 13450 18264 13506 18320
rect 13082 18128 13138 18184
rect 12254 13368 12310 13424
rect 12070 11192 12126 11248
rect 13818 18808 13874 18864
rect 13174 14320 13230 14376
rect 12254 10648 12310 10704
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 13082 13096 13138 13152
rect 12346 3440 12402 3496
rect 13174 7792 13230 7848
rect 13450 7828 13452 7848
rect 13452 7828 13504 7848
rect 13504 7828 13506 7848
rect 13450 7792 13506 7828
rect 12070 584 12126 640
rect 13634 14184 13690 14240
rect 13726 12688 13782 12744
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 14370 16940 14372 16960
rect 14372 16940 14424 16960
rect 14424 16940 14426 16960
rect 14370 16904 14426 16940
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 14554 15564 14610 15600
rect 14554 15544 14556 15564
rect 14556 15544 14608 15564
rect 14608 15544 14610 15564
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 15198 14320 15254 14376
rect 14922 13232 14978 13288
rect 15658 18536 15714 18592
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 14370 11600 14426 11656
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 15198 12824 15254 12880
rect 15382 13232 15438 13288
rect 14370 7792 14426 7848
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 13818 3440 13874 3496
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 15750 13404 15752 13424
rect 15752 13404 15804 13424
rect 15804 13404 15806 13424
rect 15750 13368 15806 13404
rect 16210 13812 16212 13832
rect 16212 13812 16264 13832
rect 16264 13812 16266 13832
rect 16210 13776 16266 13812
rect 15750 12824 15806 12880
rect 15750 10376 15806 10432
rect 15106 5208 15162 5264
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 15934 4528 15990 4584
rect 16210 12824 16266 12880
rect 16118 10376 16174 10432
rect 16670 14320 16726 14376
rect 16670 11192 16726 11248
rect 16670 9016 16726 9072
rect 17958 20576 18014 20632
rect 16946 15544 17002 15600
rect 17314 12824 17370 12880
rect 18510 21120 18566 21176
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 17590 18672 17646 18728
rect 17590 14320 17646 14376
rect 17682 13912 17738 13968
rect 17590 13232 17646 13288
rect 17498 12688 17554 12744
rect 17406 12280 17462 12336
rect 16578 8492 16634 8528
rect 16578 8472 16580 8492
rect 16580 8472 16632 8492
rect 16632 8472 16634 8492
rect 16486 7928 16542 7984
rect 16946 8472 17002 8528
rect 17774 13096 17830 13152
rect 17774 12552 17830 12608
rect 17682 10512 17738 10568
rect 17498 8236 17500 8256
rect 17500 8236 17552 8256
rect 17552 8236 17554 8256
rect 17498 8200 17554 8236
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 19246 21528 19302 21584
rect 18970 19216 19026 19272
rect 18878 18808 18934 18864
rect 18694 18264 18750 18320
rect 18602 18128 18658 18184
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 17958 16940 17960 16960
rect 17960 16940 18012 16960
rect 18012 16940 18014 16960
rect 17958 16904 18014 16940
rect 18050 16496 18106 16552
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 17958 15952 18014 16008
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 17958 14592 18014 14648
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 17958 13640 18014 13696
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 18050 12180 18052 12200
rect 18052 12180 18104 12200
rect 18104 12180 18106 12200
rect 18050 12144 18106 12180
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 17958 11328 18014 11384
rect 18418 11056 18474 11112
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18326 9968 18382 10024
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 18326 9036 18382 9072
rect 18326 9016 18328 9036
rect 18328 9016 18380 9036
rect 18380 9016 18382 9036
rect 18602 8880 18658 8936
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 18510 8608 18566 8664
rect 17958 8472 18014 8528
rect 18326 8336 18382 8392
rect 18602 8356 18658 8392
rect 18602 8336 18604 8356
rect 18604 8336 18656 8356
rect 18656 8336 18658 8356
rect 17958 8064 18014 8120
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 18510 6160 18566 6216
rect 20166 20168 20222 20224
rect 20626 22072 20682 22128
rect 19154 18808 19210 18864
rect 19246 18264 19302 18320
rect 19246 17856 19302 17912
rect 18970 15408 19026 15464
rect 19614 18672 19670 18728
rect 19062 14456 19118 14512
rect 19246 15000 19302 15056
rect 19154 14048 19210 14104
rect 18970 13776 19026 13832
rect 18786 12552 18842 12608
rect 18786 7520 18842 7576
rect 18142 5752 18198 5808
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 18786 4800 18842 4856
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 18510 3168 18566 3224
rect 18418 3032 18474 3088
rect 18510 2896 18566 2952
rect 18142 2488 18198 2544
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 18510 1536 18566 1592
rect 19246 10784 19302 10840
rect 19062 10648 19118 10704
rect 20258 19760 20314 19816
rect 18970 9424 19026 9480
rect 19522 8336 19578 8392
rect 19522 8200 19578 8256
rect 18970 5616 19026 5672
rect 19246 7112 19302 7168
rect 20626 19216 20682 19272
rect 19890 10376 19946 10432
rect 20074 8608 20130 8664
rect 20074 6704 20130 6760
rect 21178 17312 21234 17368
rect 20994 15544 21050 15600
rect 20534 9968 20590 10024
rect 20442 3984 20498 4040
rect 20258 3848 20314 3904
rect 20074 3440 20130 3496
rect 19246 1944 19302 2000
rect 18878 176 18934 232
<< metal3 >>
rect 19057 22538 19123 22541
rect 22320 22538 22800 22568
rect 19057 22536 22800 22538
rect 19057 22480 19062 22536
rect 19118 22480 22800 22536
rect 19057 22478 22800 22480
rect 19057 22475 19123 22478
rect 22320 22448 22800 22478
rect 20621 22130 20687 22133
rect 22320 22130 22800 22160
rect 20621 22128 22800 22130
rect 20621 22072 20626 22128
rect 20682 22072 22800 22128
rect 20621 22070 22800 22072
rect 20621 22067 20687 22070
rect 22320 22040 22800 22070
rect 19241 21586 19307 21589
rect 22320 21586 22800 21616
rect 19241 21584 22800 21586
rect 19241 21528 19246 21584
rect 19302 21528 22800 21584
rect 19241 21526 22800 21528
rect 19241 21523 19307 21526
rect 22320 21496 22800 21526
rect 18505 21178 18571 21181
rect 22320 21178 22800 21208
rect 18505 21176 22800 21178
rect 18505 21120 18510 21176
rect 18566 21120 22800 21176
rect 18505 21118 22800 21120
rect 18505 21115 18571 21118
rect 22320 21088 22800 21118
rect 17953 20634 18019 20637
rect 22320 20634 22800 20664
rect 17953 20632 22800 20634
rect 17953 20576 17958 20632
rect 18014 20576 22800 20632
rect 17953 20574 22800 20576
rect 17953 20571 18019 20574
rect 22320 20544 22800 20574
rect 20161 20226 20227 20229
rect 22320 20226 22800 20256
rect 20161 20224 22800 20226
rect 20161 20168 20166 20224
rect 20222 20168 22800 20224
rect 20161 20166 22800 20168
rect 20161 20163 20227 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 22320 20136 22800 20166
rect 14672 20095 14992 20096
rect 20253 19818 20319 19821
rect 22320 19818 22800 19848
rect 20253 19816 22800 19818
rect 20253 19760 20258 19816
rect 20314 19760 22800 19816
rect 20253 19758 22800 19760
rect 20253 19755 20319 19758
rect 22320 19728 22800 19758
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 2497 19274 2563 19277
rect 9857 19274 9923 19277
rect 2497 19272 9923 19274
rect 2497 19216 2502 19272
rect 2558 19216 9862 19272
rect 9918 19216 9923 19272
rect 2497 19214 9923 19216
rect 2497 19211 2563 19214
rect 9857 19211 9923 19214
rect 10041 19274 10107 19277
rect 18965 19274 19031 19277
rect 10041 19272 19031 19274
rect 10041 19216 10046 19272
rect 10102 19216 18970 19272
rect 19026 19216 19031 19272
rect 10041 19214 19031 19216
rect 10041 19211 10107 19214
rect 18965 19211 19031 19214
rect 20621 19274 20687 19277
rect 22320 19274 22800 19304
rect 20621 19272 22800 19274
rect 20621 19216 20626 19272
rect 20682 19216 22800 19272
rect 20621 19214 22800 19216
rect 20621 19211 20687 19214
rect 22320 19184 22800 19214
rect 10225 19138 10291 19141
rect 12801 19138 12867 19141
rect 10225 19136 12867 19138
rect 10225 19080 10230 19136
rect 10286 19080 12806 19136
rect 12862 19080 12867 19136
rect 10225 19078 12867 19080
rect 10225 19075 10291 19078
rect 12801 19075 12867 19078
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 9765 19002 9831 19005
rect 9765 19000 14106 19002
rect 9765 18944 9770 19000
rect 9826 18944 14106 19000
rect 9765 18942 14106 18944
rect 9765 18939 9831 18942
rect 12249 18866 12315 18869
rect 13813 18866 13879 18869
rect 12249 18864 13879 18866
rect 12249 18808 12254 18864
rect 12310 18808 13818 18864
rect 13874 18808 13879 18864
rect 12249 18806 13879 18808
rect 14046 18866 14106 18942
rect 18873 18866 18939 18869
rect 14046 18864 18939 18866
rect 14046 18808 18878 18864
rect 18934 18808 18939 18864
rect 14046 18806 18939 18808
rect 12249 18803 12315 18806
rect 13813 18803 13879 18806
rect 18873 18803 18939 18806
rect 19149 18866 19215 18869
rect 22320 18866 22800 18896
rect 19149 18864 22800 18866
rect 19149 18808 19154 18864
rect 19210 18808 22800 18864
rect 19149 18806 22800 18808
rect 19149 18803 19215 18806
rect 22320 18776 22800 18806
rect 8569 18730 8635 18733
rect 17585 18730 17651 18733
rect 19609 18730 19675 18733
rect 8569 18728 19675 18730
rect 8569 18672 8574 18728
rect 8630 18672 17590 18728
rect 17646 18672 19614 18728
rect 19670 18672 19675 18728
rect 8569 18670 19675 18672
rect 8569 18667 8635 18670
rect 17585 18667 17651 18670
rect 19609 18667 19675 18670
rect 11881 18594 11947 18597
rect 15653 18594 15719 18597
rect 11881 18592 15719 18594
rect 11881 18536 11886 18592
rect 11942 18536 15658 18592
rect 15714 18536 15719 18592
rect 11881 18534 15719 18536
rect 11881 18531 11947 18534
rect 15653 18531 15719 18534
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 9489 18458 9555 18461
rect 9489 18456 10426 18458
rect 9489 18400 9494 18456
rect 9550 18400 10426 18456
rect 9489 18398 10426 18400
rect 9489 18395 9555 18398
rect 1393 18322 1459 18325
rect 9581 18322 9647 18325
rect 1393 18320 9647 18322
rect 1393 18264 1398 18320
rect 1454 18264 9586 18320
rect 9642 18264 9647 18320
rect 1393 18262 9647 18264
rect 10366 18322 10426 18398
rect 12525 18322 12591 18325
rect 10366 18320 12591 18322
rect 10366 18264 12530 18320
rect 12586 18264 12591 18320
rect 10366 18262 12591 18264
rect 1393 18259 1459 18262
rect 9581 18259 9647 18262
rect 12525 18259 12591 18262
rect 13445 18322 13511 18325
rect 18689 18322 18755 18325
rect 13445 18320 18755 18322
rect 13445 18264 13450 18320
rect 13506 18264 18694 18320
rect 18750 18264 18755 18320
rect 13445 18262 18755 18264
rect 13445 18259 13511 18262
rect 18689 18259 18755 18262
rect 19241 18322 19307 18325
rect 22320 18322 22800 18352
rect 19241 18320 22800 18322
rect 19241 18264 19246 18320
rect 19302 18264 22800 18320
rect 19241 18262 22800 18264
rect 19241 18259 19307 18262
rect 22320 18232 22800 18262
rect 13077 18186 13143 18189
rect 18597 18186 18663 18189
rect 13077 18184 18663 18186
rect 13077 18128 13082 18184
rect 13138 18128 18602 18184
rect 18658 18128 18663 18184
rect 13077 18126 18663 18128
rect 13077 18123 13143 18126
rect 18597 18123 18663 18126
rect 10777 18050 10843 18053
rect 10550 18048 10843 18050
rect 10550 17992 10782 18048
rect 10838 17992 10843 18048
rect 10550 17990 10843 17992
rect 7808 17984 8128 17985
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 10550 17916 10610 17990
rect 10777 17987 10843 17990
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 10542 17852 10548 17916
rect 10612 17852 10618 17916
rect 19241 17914 19307 17917
rect 22320 17914 22800 17944
rect 19241 17912 22800 17914
rect 19241 17856 19246 17912
rect 19302 17856 22800 17912
rect 19241 17854 22800 17856
rect 19241 17851 19307 17854
rect 22320 17824 22800 17854
rect 4376 17440 4696 17441
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 21173 17370 21239 17373
rect 22320 17370 22800 17400
rect 21173 17368 22800 17370
rect 21173 17312 21178 17368
rect 21234 17312 22800 17368
rect 21173 17310 22800 17312
rect 21173 17307 21239 17310
rect 22320 17280 22800 17310
rect 0 17234 480 17264
rect 3417 17234 3483 17237
rect 0 17232 3483 17234
rect 0 17176 3422 17232
rect 3478 17176 3483 17232
rect 0 17174 3483 17176
rect 0 17144 480 17174
rect 3417 17171 3483 17174
rect 11237 16962 11303 16965
rect 14365 16962 14431 16965
rect 11237 16960 14431 16962
rect 11237 16904 11242 16960
rect 11298 16904 14370 16960
rect 14426 16904 14431 16960
rect 11237 16902 14431 16904
rect 11237 16899 11303 16902
rect 14365 16899 14431 16902
rect 17953 16962 18019 16965
rect 22320 16962 22800 16992
rect 17953 16960 22800 16962
rect 17953 16904 17958 16960
rect 18014 16904 22800 16960
rect 17953 16902 22800 16904
rect 17953 16899 18019 16902
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 22320 16872 22800 16902
rect 14672 16831 14992 16832
rect 9397 16690 9463 16693
rect 10317 16690 10383 16693
rect 9397 16688 10383 16690
rect 9397 16632 9402 16688
rect 9458 16632 10322 16688
rect 10378 16632 10383 16688
rect 9397 16630 10383 16632
rect 9397 16627 9463 16630
rect 10317 16627 10383 16630
rect 12198 16628 12204 16692
rect 12268 16690 12274 16692
rect 12341 16690 12407 16693
rect 12268 16688 12407 16690
rect 12268 16632 12346 16688
rect 12402 16632 12407 16688
rect 12268 16630 12407 16632
rect 12268 16628 12274 16630
rect 12341 16627 12407 16630
rect 18045 16554 18111 16557
rect 22320 16554 22800 16584
rect 18045 16552 22800 16554
rect 18045 16496 18050 16552
rect 18106 16496 22800 16552
rect 18045 16494 22800 16496
rect 18045 16491 18111 16494
rect 22320 16464 22800 16494
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 17953 16010 18019 16013
rect 22320 16010 22800 16040
rect 17953 16008 22800 16010
rect 17953 15952 17958 16008
rect 18014 15952 22800 16008
rect 17953 15950 22800 15952
rect 17953 15947 18019 15950
rect 22320 15920 22800 15950
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 14549 15602 14615 15605
rect 16941 15602 17007 15605
rect 14549 15600 17007 15602
rect 14549 15544 14554 15600
rect 14610 15544 16946 15600
rect 17002 15544 17007 15600
rect 14549 15542 17007 15544
rect 14549 15539 14615 15542
rect 16941 15539 17007 15542
rect 20989 15602 21055 15605
rect 22320 15602 22800 15632
rect 20989 15600 22800 15602
rect 20989 15544 20994 15600
rect 21050 15544 22800 15600
rect 20989 15542 22800 15544
rect 20989 15539 21055 15542
rect 22320 15512 22800 15542
rect 17718 15404 17724 15468
rect 17788 15466 17794 15468
rect 18965 15466 19031 15469
rect 17788 15464 19031 15466
rect 17788 15408 18970 15464
rect 19026 15408 19031 15464
rect 17788 15406 19031 15408
rect 17788 15404 17794 15406
rect 18965 15403 19031 15406
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 19241 15058 19307 15061
rect 22320 15058 22800 15088
rect 19241 15056 22800 15058
rect 19241 15000 19246 15056
rect 19302 15000 22800 15056
rect 19241 14998 22800 15000
rect 19241 14995 19307 14998
rect 22320 14968 22800 14998
rect 7808 14720 8128 14721
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 17953 14650 18019 14653
rect 22320 14650 22800 14680
rect 17953 14648 22800 14650
rect 17953 14592 17958 14648
rect 18014 14592 22800 14648
rect 17953 14590 22800 14592
rect 17953 14587 18019 14590
rect 22320 14560 22800 14590
rect 19057 14514 19123 14517
rect 16438 14512 19123 14514
rect 16438 14456 19062 14512
rect 19118 14456 19123 14512
rect 16438 14454 19123 14456
rect 13169 14378 13235 14381
rect 15193 14378 15259 14381
rect 16438 14378 16498 14454
rect 19057 14451 19123 14454
rect 13169 14376 16498 14378
rect 13169 14320 13174 14376
rect 13230 14320 15198 14376
rect 15254 14320 16498 14376
rect 13169 14318 16498 14320
rect 16665 14378 16731 14381
rect 17585 14378 17651 14381
rect 16665 14376 17651 14378
rect 16665 14320 16670 14376
rect 16726 14320 17590 14376
rect 17646 14320 17651 14376
rect 16665 14318 17651 14320
rect 13169 14315 13235 14318
rect 15193 14315 15259 14318
rect 16665 14315 16731 14318
rect 17585 14315 17651 14318
rect 11881 14242 11947 14245
rect 13629 14242 13695 14245
rect 11881 14240 13695 14242
rect 11881 14184 11886 14240
rect 11942 14184 13634 14240
rect 13690 14184 13695 14240
rect 11881 14182 13695 14184
rect 11881 14179 11947 14182
rect 13629 14179 13695 14182
rect 4376 14176 4696 14177
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 19149 14106 19215 14109
rect 22320 14106 22800 14136
rect 19149 14104 22800 14106
rect 19149 14048 19154 14104
rect 19210 14048 22800 14104
rect 19149 14046 22800 14048
rect 19149 14043 19215 14046
rect 22320 14016 22800 14046
rect 11513 13970 11579 13973
rect 17677 13970 17743 13973
rect 11513 13968 17743 13970
rect 11513 13912 11518 13968
rect 11574 13912 17682 13968
rect 17738 13912 17743 13968
rect 11513 13910 17743 13912
rect 11513 13907 11579 13910
rect 17677 13907 17743 13910
rect 16205 13834 16271 13837
rect 18965 13834 19031 13837
rect 16205 13832 19031 13834
rect 16205 13776 16210 13832
rect 16266 13776 18970 13832
rect 19026 13776 19031 13832
rect 16205 13774 19031 13776
rect 16205 13771 16271 13774
rect 18965 13771 19031 13774
rect 17953 13698 18019 13701
rect 22320 13698 22800 13728
rect 17953 13696 22800 13698
rect 17953 13640 17958 13696
rect 18014 13640 22800 13696
rect 17953 13638 22800 13640
rect 17953 13635 18019 13638
rect 7808 13632 8128 13633
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 22320 13608 22800 13638
rect 14672 13567 14992 13568
rect 10225 13564 10291 13565
rect 10174 13562 10180 13564
rect 10134 13502 10180 13562
rect 10244 13560 10291 13564
rect 10286 13504 10291 13560
rect 10174 13500 10180 13502
rect 10244 13500 10291 13504
rect 10225 13499 10291 13500
rect 11973 13426 12039 13429
rect 12249 13426 12315 13429
rect 15745 13426 15811 13429
rect 11973 13424 15811 13426
rect 11973 13368 11978 13424
rect 12034 13368 12254 13424
rect 12310 13368 15750 13424
rect 15806 13368 15811 13424
rect 11973 13366 15811 13368
rect 11973 13363 12039 13366
rect 12249 13363 12315 13366
rect 15745 13363 15811 13366
rect 14917 13290 14983 13293
rect 15377 13290 15443 13293
rect 14917 13288 15443 13290
rect 14917 13232 14922 13288
rect 14978 13232 15382 13288
rect 15438 13232 15443 13288
rect 14917 13230 15443 13232
rect 14917 13227 14983 13230
rect 15377 13227 15443 13230
rect 17585 13290 17651 13293
rect 22320 13290 22800 13320
rect 17585 13288 22800 13290
rect 17585 13232 17590 13288
rect 17646 13232 22800 13288
rect 17585 13230 22800 13232
rect 17585 13227 17651 13230
rect 22320 13200 22800 13230
rect 13077 13154 13143 13157
rect 17769 13154 17835 13157
rect 13077 13152 17835 13154
rect 13077 13096 13082 13152
rect 13138 13096 17774 13152
rect 17830 13096 17835 13152
rect 13077 13094 17835 13096
rect 13077 13091 13143 13094
rect 17769 13091 17835 13094
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 15193 12882 15259 12885
rect 15745 12882 15811 12885
rect 16205 12882 16271 12885
rect 17309 12882 17375 12885
rect 15193 12880 16271 12882
rect 15193 12824 15198 12880
rect 15254 12824 15750 12880
rect 15806 12824 16210 12880
rect 16266 12824 16271 12880
rect 15193 12822 16271 12824
rect 15193 12819 15259 12822
rect 15745 12819 15811 12822
rect 16205 12819 16271 12822
rect 16438 12880 17375 12882
rect 16438 12824 17314 12880
rect 17370 12824 17375 12880
rect 16438 12822 17375 12824
rect 13721 12746 13787 12749
rect 16438 12748 16498 12822
rect 17309 12819 17375 12822
rect 16430 12746 16436 12748
rect 13721 12744 16436 12746
rect 13721 12688 13726 12744
rect 13782 12688 16436 12744
rect 13721 12686 16436 12688
rect 13721 12683 13787 12686
rect 16430 12684 16436 12686
rect 16500 12684 16506 12748
rect 17493 12746 17559 12749
rect 22320 12746 22800 12776
rect 17493 12744 22800 12746
rect 17493 12688 17498 12744
rect 17554 12688 22800 12744
rect 17493 12686 22800 12688
rect 17493 12683 17559 12686
rect 22320 12656 22800 12686
rect 17769 12610 17835 12613
rect 18781 12610 18847 12613
rect 17769 12608 18847 12610
rect 17769 12552 17774 12608
rect 17830 12552 18786 12608
rect 18842 12552 18847 12608
rect 17769 12550 18847 12552
rect 17769 12547 17835 12550
rect 18781 12547 18847 12550
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 17401 12338 17467 12341
rect 22320 12338 22800 12368
rect 17401 12336 22800 12338
rect 17401 12280 17406 12336
rect 17462 12280 22800 12336
rect 17401 12278 22800 12280
rect 17401 12275 17467 12278
rect 22320 12248 22800 12278
rect 10542 12140 10548 12204
rect 10612 12202 10618 12204
rect 18045 12202 18111 12205
rect 10612 12200 18111 12202
rect 10612 12144 18050 12200
rect 18106 12144 18111 12200
rect 10612 12142 18111 12144
rect 10612 12140 10618 12142
rect 18045 12139 18111 12142
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 22320 11794 22800 11824
rect 18094 11734 22800 11794
rect 14365 11658 14431 11661
rect 18094 11658 18154 11734
rect 22320 11704 22800 11734
rect 14365 11656 18154 11658
rect 14365 11600 14370 11656
rect 14426 11600 18154 11656
rect 14365 11598 18154 11600
rect 14365 11595 14431 11598
rect 7808 11456 8128 11457
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 17953 11386 18019 11389
rect 22320 11386 22800 11416
rect 17953 11384 22800 11386
rect 17953 11328 17958 11384
rect 18014 11328 22800 11384
rect 17953 11326 22800 11328
rect 17953 11323 18019 11326
rect 22320 11296 22800 11326
rect 12065 11250 12131 11253
rect 12198 11250 12204 11252
rect 12065 11248 12204 11250
rect 12065 11192 12070 11248
rect 12126 11192 12204 11248
rect 12065 11190 12204 11192
rect 12065 11187 12131 11190
rect 12198 11188 12204 11190
rect 12268 11188 12274 11252
rect 16430 11188 16436 11252
rect 16500 11250 16506 11252
rect 16665 11250 16731 11253
rect 16500 11248 16731 11250
rect 16500 11192 16670 11248
rect 16726 11192 16731 11248
rect 16500 11190 16731 11192
rect 16500 11188 16506 11190
rect 16665 11187 16731 11190
rect 10174 11052 10180 11116
rect 10244 11114 10250 11116
rect 18413 11114 18479 11117
rect 10244 11112 18479 11114
rect 10244 11056 18418 11112
rect 18474 11056 18479 11112
rect 10244 11054 18479 11056
rect 10244 11052 10250 11054
rect 18413 11051 18479 11054
rect 4376 10912 4696 10913
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 19241 10842 19307 10845
rect 22320 10842 22800 10872
rect 19241 10840 22800 10842
rect 19241 10784 19246 10840
rect 19302 10784 22800 10840
rect 19241 10782 22800 10784
rect 19241 10779 19307 10782
rect 22320 10752 22800 10782
rect 12249 10706 12315 10709
rect 19057 10706 19123 10709
rect 12249 10704 19123 10706
rect 12249 10648 12254 10704
rect 12310 10648 19062 10704
rect 19118 10648 19123 10704
rect 12249 10646 19123 10648
rect 12249 10643 12315 10646
rect 19057 10643 19123 10646
rect 17677 10572 17743 10573
rect 17677 10570 17724 10572
rect 17632 10568 17724 10570
rect 17632 10512 17682 10568
rect 17632 10510 17724 10512
rect 17677 10508 17724 10510
rect 17788 10508 17794 10572
rect 17677 10507 17743 10508
rect 15745 10434 15811 10437
rect 16113 10434 16179 10437
rect 15745 10432 16179 10434
rect 15745 10376 15750 10432
rect 15806 10376 16118 10432
rect 16174 10376 16179 10432
rect 15745 10374 16179 10376
rect 15745 10371 15811 10374
rect 16113 10371 16179 10374
rect 19885 10434 19951 10437
rect 22320 10434 22800 10464
rect 19885 10432 22800 10434
rect 19885 10376 19890 10432
rect 19946 10376 22800 10432
rect 19885 10374 22800 10376
rect 19885 10371 19951 10374
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 22320 10344 22800 10374
rect 14672 10303 14992 10304
rect 18321 10026 18387 10029
rect 18638 10026 18644 10028
rect 18321 10024 18644 10026
rect 18321 9968 18326 10024
rect 18382 9968 18644 10024
rect 18321 9966 18644 9968
rect 18321 9963 18387 9966
rect 18638 9964 18644 9966
rect 18708 9964 18714 10028
rect 20529 10026 20595 10029
rect 22320 10026 22800 10056
rect 20529 10024 22800 10026
rect 20529 9968 20534 10024
rect 20590 9968 22800 10024
rect 20529 9966 22800 9968
rect 20529 9963 20595 9966
rect 22320 9936 22800 9966
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 10409 9618 10475 9621
rect 10542 9618 10548 9620
rect 10409 9616 10548 9618
rect 10409 9560 10414 9616
rect 10470 9560 10548 9616
rect 10409 9558 10548 9560
rect 10409 9555 10475 9558
rect 10542 9556 10548 9558
rect 10612 9556 10618 9620
rect 18965 9482 19031 9485
rect 22320 9482 22800 9512
rect 18965 9480 22800 9482
rect 18965 9424 18970 9480
rect 19026 9424 22800 9480
rect 18965 9422 22800 9424
rect 18965 9419 19031 9422
rect 22320 9392 22800 9422
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 10133 9076 10199 9077
rect 10133 9074 10180 9076
rect 10088 9072 10180 9074
rect 10088 9016 10138 9072
rect 10088 9014 10180 9016
rect 10133 9012 10180 9014
rect 10244 9012 10250 9076
rect 16665 9074 16731 9077
rect 17902 9074 17908 9076
rect 16665 9072 17908 9074
rect 16665 9016 16670 9072
rect 16726 9016 17908 9072
rect 16665 9014 17908 9016
rect 10133 9011 10199 9012
rect 16665 9011 16731 9014
rect 17902 9012 17908 9014
rect 17972 9012 17978 9076
rect 18321 9074 18387 9077
rect 22320 9074 22800 9104
rect 18321 9072 22800 9074
rect 18321 9016 18326 9072
rect 18382 9016 22800 9072
rect 18321 9014 22800 9016
rect 18321 9011 18387 9014
rect 22320 8984 22800 9014
rect 18597 8938 18663 8941
rect 18822 8938 18828 8940
rect 18597 8936 18828 8938
rect 18597 8880 18602 8936
rect 18658 8880 18828 8936
rect 18597 8878 18828 8880
rect 18597 8875 18663 8878
rect 18822 8876 18828 8878
rect 18892 8876 18898 8940
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 8671 18424 8672
rect 18505 8666 18571 8669
rect 20069 8666 20135 8669
rect 18505 8664 20135 8666
rect 18505 8608 18510 8664
rect 18566 8608 20074 8664
rect 20130 8608 20135 8664
rect 18505 8606 20135 8608
rect 18505 8603 18571 8606
rect 20069 8603 20135 8606
rect 16573 8530 16639 8533
rect 16941 8530 17007 8533
rect 16573 8528 17007 8530
rect 16573 8472 16578 8528
rect 16634 8472 16946 8528
rect 17002 8472 17007 8528
rect 16573 8470 17007 8472
rect 16573 8467 16639 8470
rect 16941 8467 17007 8470
rect 17953 8530 18019 8533
rect 22320 8530 22800 8560
rect 17953 8528 22800 8530
rect 17953 8472 17958 8528
rect 18014 8472 22800 8528
rect 17953 8470 22800 8472
rect 17953 8467 18019 8470
rect 22320 8440 22800 8470
rect 10317 8394 10383 8397
rect 18321 8394 18387 8397
rect 10317 8392 18387 8394
rect 10317 8336 10322 8392
rect 10378 8336 18326 8392
rect 18382 8336 18387 8392
rect 10317 8334 18387 8336
rect 10317 8331 10383 8334
rect 18321 8331 18387 8334
rect 18597 8394 18663 8397
rect 19517 8394 19583 8397
rect 18597 8392 19583 8394
rect 18597 8336 18602 8392
rect 18658 8336 19522 8392
rect 19578 8336 19583 8392
rect 18597 8334 19583 8336
rect 18597 8331 18663 8334
rect 19517 8331 19583 8334
rect 17493 8258 17559 8261
rect 19517 8258 19583 8261
rect 17493 8256 19583 8258
rect 17493 8200 17498 8256
rect 17554 8200 19522 8256
rect 19578 8200 19583 8256
rect 17493 8198 19583 8200
rect 17493 8195 17559 8198
rect 19517 8195 19583 8198
rect 7808 8192 8128 8193
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 17953 8122 18019 8125
rect 22320 8122 22800 8152
rect 17953 8120 22800 8122
rect 17953 8064 17958 8120
rect 18014 8064 22800 8120
rect 17953 8062 22800 8064
rect 17953 8059 18019 8062
rect 22320 8032 22800 8062
rect 16481 7986 16547 7989
rect 16438 7984 16547 7986
rect 16438 7928 16486 7984
rect 16542 7928 16547 7984
rect 16438 7923 16547 7928
rect 11329 7850 11395 7853
rect 13169 7850 13235 7853
rect 13445 7850 13511 7853
rect 11329 7848 13511 7850
rect 11329 7792 11334 7848
rect 11390 7792 13174 7848
rect 13230 7792 13450 7848
rect 13506 7792 13511 7848
rect 11329 7790 13511 7792
rect 11329 7787 11395 7790
rect 13169 7787 13235 7790
rect 13445 7787 13511 7790
rect 14365 7850 14431 7853
rect 16438 7850 16498 7923
rect 14365 7848 16498 7850
rect 14365 7792 14370 7848
rect 14426 7792 16498 7848
rect 14365 7790 16498 7792
rect 14365 7787 14431 7790
rect 4376 7648 4696 7649
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 18781 7578 18847 7581
rect 22320 7578 22800 7608
rect 18781 7576 22800 7578
rect 18781 7520 18786 7576
rect 18842 7520 22800 7576
rect 18781 7518 22800 7520
rect 18781 7515 18847 7518
rect 22320 7488 22800 7518
rect 19241 7170 19307 7173
rect 22320 7170 22800 7200
rect 19241 7168 22800 7170
rect 19241 7112 19246 7168
rect 19302 7112 22800 7168
rect 19241 7110 22800 7112
rect 19241 7107 19307 7110
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 22320 7080 22800 7110
rect 14672 7039 14992 7040
rect 20069 6762 20135 6765
rect 22320 6762 22800 6792
rect 20069 6760 22800 6762
rect 20069 6704 20074 6760
rect 20130 6704 22800 6760
rect 20069 6702 22800 6704
rect 20069 6699 20135 6702
rect 22320 6672 22800 6702
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 18505 6218 18571 6221
rect 22320 6218 22800 6248
rect 18505 6216 22800 6218
rect 18505 6160 18510 6216
rect 18566 6160 22800 6216
rect 18505 6158 22800 6160
rect 18505 6155 18571 6158
rect 22320 6128 22800 6158
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 0 5810 480 5840
rect 4061 5810 4127 5813
rect 0 5808 4127 5810
rect 0 5752 4066 5808
rect 4122 5752 4127 5808
rect 0 5750 4127 5752
rect 0 5720 480 5750
rect 4061 5747 4127 5750
rect 18137 5810 18203 5813
rect 22320 5810 22800 5840
rect 18137 5808 22800 5810
rect 18137 5752 18142 5808
rect 18198 5752 22800 5808
rect 18137 5750 22800 5752
rect 18137 5747 18203 5750
rect 22320 5720 22800 5750
rect 18822 5612 18828 5676
rect 18892 5674 18898 5676
rect 18965 5674 19031 5677
rect 18892 5672 19031 5674
rect 18892 5616 18970 5672
rect 19026 5616 19031 5672
rect 18892 5614 19031 5616
rect 18892 5612 18898 5614
rect 18965 5611 19031 5614
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 15101 5266 15167 5269
rect 22320 5266 22800 5296
rect 15101 5264 22800 5266
rect 15101 5208 15106 5264
rect 15162 5208 22800 5264
rect 15101 5206 22800 5208
rect 15101 5203 15167 5206
rect 22320 5176 22800 5206
rect 7808 4928 8128 4929
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 18781 4858 18847 4861
rect 22320 4858 22800 4888
rect 18781 4856 22800 4858
rect 18781 4800 18786 4856
rect 18842 4800 22800 4856
rect 18781 4798 22800 4800
rect 18781 4795 18847 4798
rect 22320 4768 22800 4798
rect 10685 4586 10751 4589
rect 15929 4586 15995 4589
rect 10685 4584 18568 4586
rect 10685 4528 10690 4584
rect 10746 4528 15934 4584
rect 15990 4528 18568 4584
rect 10685 4526 18568 4528
rect 10685 4523 10751 4526
rect 15929 4523 15995 4526
rect 4376 4384 4696 4385
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 18508 4314 18568 4526
rect 22320 4314 22800 4344
rect 18508 4254 22800 4314
rect 22320 4224 22800 4254
rect 10777 4042 10843 4045
rect 20437 4042 20503 4045
rect 10777 4040 20503 4042
rect 10777 3984 10782 4040
rect 10838 3984 20442 4040
rect 20498 3984 20503 4040
rect 10777 3982 20503 3984
rect 10777 3979 10843 3982
rect 20437 3979 20503 3982
rect 20253 3906 20319 3909
rect 22320 3906 22800 3936
rect 20253 3904 22800 3906
rect 20253 3848 20258 3904
rect 20314 3848 22800 3904
rect 20253 3846 22800 3848
rect 20253 3843 20319 3846
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 22320 3816 22800 3846
rect 14672 3775 14992 3776
rect 12341 3498 12407 3501
rect 13813 3498 13879 3501
rect 12341 3496 13879 3498
rect 12341 3440 12346 3496
rect 12402 3440 13818 3496
rect 13874 3440 13879 3496
rect 12341 3438 13879 3440
rect 12341 3435 12407 3438
rect 13813 3435 13879 3438
rect 20069 3498 20135 3501
rect 22320 3498 22800 3528
rect 20069 3496 22800 3498
rect 20069 3440 20074 3496
rect 20130 3440 22800 3496
rect 20069 3438 22800 3440
rect 20069 3435 20135 3438
rect 22320 3408 22800 3438
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 18505 3226 18571 3229
rect 18638 3226 18644 3228
rect 18505 3224 18644 3226
rect 18505 3168 18510 3224
rect 18566 3168 18644 3224
rect 18505 3166 18644 3168
rect 18505 3163 18571 3166
rect 18638 3164 18644 3166
rect 18708 3164 18714 3228
rect 9857 3090 9923 3093
rect 18413 3090 18479 3093
rect 9857 3088 18479 3090
rect 9857 3032 9862 3088
rect 9918 3032 18418 3088
rect 18474 3032 18479 3088
rect 9857 3030 18479 3032
rect 9857 3027 9923 3030
rect 18413 3027 18479 3030
rect 18505 2954 18571 2957
rect 22320 2954 22800 2984
rect 18505 2952 22800 2954
rect 18505 2896 18510 2952
rect 18566 2896 22800 2952
rect 18505 2894 22800 2896
rect 18505 2891 18571 2894
rect 22320 2864 22800 2894
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 18137 2546 18203 2549
rect 22320 2546 22800 2576
rect 18137 2544 22800 2546
rect 18137 2488 18142 2544
rect 18198 2488 22800 2544
rect 18137 2486 22800 2488
rect 18137 2483 18203 2486
rect 22320 2456 22800 2486
rect 4376 2208 4696 2209
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 19241 2002 19307 2005
rect 22320 2002 22800 2032
rect 19241 2000 22800 2002
rect 19241 1944 19246 2000
rect 19302 1944 22800 2000
rect 19241 1942 22800 1944
rect 19241 1939 19307 1942
rect 22320 1912 22800 1942
rect 18505 1594 18571 1597
rect 22320 1594 22800 1624
rect 18505 1592 22800 1594
rect 18505 1536 18510 1592
rect 18566 1536 22800 1592
rect 18505 1534 22800 1536
rect 18505 1531 18571 1534
rect 22320 1504 22800 1534
rect 17902 988 17908 1052
rect 17972 1050 17978 1052
rect 22320 1050 22800 1080
rect 17972 990 22800 1050
rect 17972 988 17978 990
rect 22320 960 22800 990
rect 12065 642 12131 645
rect 22320 642 22800 672
rect 12065 640 22800 642
rect 12065 584 12070 640
rect 12126 584 22800 640
rect 12065 582 22800 584
rect 12065 579 12131 582
rect 22320 552 22800 582
rect 18873 234 18939 237
rect 22320 234 22800 264
rect 18873 232 22800 234
rect 18873 176 18878 232
rect 18934 176 22800 232
rect 18873 174 22800 176
rect 18873 171 18939 174
rect 22320 144 22800 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 10548 17852 10612 17916
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 12204 16628 12268 16692
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 17724 15404 17788 15468
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 10180 13560 10244 13564
rect 10180 13504 10230 13560
rect 10230 13504 10244 13560
rect 10180 13500 10244 13504
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 16436 12684 16500 12748
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 10548 12140 10612 12204
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 12204 11188 12268 11252
rect 16436 11188 16500 11252
rect 10180 11052 10244 11116
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 17724 10568 17788 10572
rect 17724 10512 17738 10568
rect 17738 10512 17788 10568
rect 17724 10508 17788 10512
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 18644 9964 18708 10028
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 10548 9556 10612 9620
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 10180 9072 10244 9076
rect 10180 9016 10194 9072
rect 10194 9016 10244 9072
rect 10180 9012 10244 9016
rect 17908 9012 17972 9076
rect 18828 8876 18892 8940
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 18828 5612 18892 5676
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 18644 3164 18708 3228
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
rect 17908 988 17972 1052
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 10547 17916 10613 17917
rect 10547 17852 10548 17916
rect 10612 17852 10613 17916
rect 10547 17851 10613 17852
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 10179 13564 10245 13565
rect 10179 13500 10180 13564
rect 10244 13500 10245 13564
rect 10179 13499 10245 13500
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 10182 11117 10242 13499
rect 10550 12205 10610 17851
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 12203 16692 12269 16693
rect 12203 16628 12204 16692
rect 12268 16628 12269 16692
rect 12203 16627 12269 16628
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 10547 12204 10613 12205
rect 10547 12140 10548 12204
rect 10612 12140 10613 12204
rect 10547 12139 10613 12140
rect 10179 11116 10245 11117
rect 10179 11052 10180 11116
rect 10244 11052 10245 11116
rect 10179 11051 10245 11052
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 10182 9077 10242 11051
rect 10550 9621 10610 12139
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 12206 11253 12266 16627
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 17723 15468 17789 15469
rect 17723 15404 17724 15468
rect 17788 15404 17789 15468
rect 17723 15403 17789 15404
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 16435 12748 16501 12749
rect 16435 12684 16436 12748
rect 16500 12684 16501 12748
rect 16435 12683 16501 12684
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 12203 11252 12269 11253
rect 12203 11188 12204 11252
rect 12268 11188 12269 11252
rect 12203 11187 12269 11188
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 10547 9620 10613 9621
rect 10547 9556 10548 9620
rect 10612 9556 10613 9620
rect 10547 9555 10613 9556
rect 10179 9076 10245 9077
rect 10179 9012 10180 9076
rect 10244 9012 10245 9076
rect 10179 9011 10245 9012
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 10368 14992 11392
rect 16438 11253 16498 12683
rect 16435 11252 16501 11253
rect 16435 11188 16436 11252
rect 16500 11188 16501 11252
rect 16435 11187 16501 11188
rect 17726 10573 17786 15403
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 17723 10572 17789 10573
rect 17723 10508 17724 10572
rect 17788 10508 17789 10572
rect 17723 10507 17789 10508
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 18104 9824 18424 10848
rect 18643 10028 18709 10029
rect 18643 9964 18644 10028
rect 18708 9964 18709 10028
rect 18643 9963 18709 9964
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 17907 9076 17973 9077
rect 17907 9012 17908 9076
rect 17972 9012 17973 9076
rect 17907 9011 17973 9012
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 17910 1053 17970 9011
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18646 3229 18706 9963
rect 18827 8940 18893 8941
rect 18827 8876 18828 8940
rect 18892 8876 18893 8940
rect 18827 8875 18893 8876
rect 18830 5677 18890 8875
rect 18827 5676 18893 5677
rect 18827 5612 18828 5676
rect 18892 5612 18893 5676
rect 18827 5611 18893 5612
rect 18643 3228 18709 3229
rect 18643 3164 18644 3228
rect 18708 3164 18709 3228
rect 18643 3163 18709 3164
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
rect 17907 1052 17973 1053
rect 17907 988 17908 1052
rect 17972 988 17973 1052
rect 17907 987 17973 988
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606821651
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1606821651
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1606821651
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1606821651
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1606821651
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1606821651
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1606821651
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606821651
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606821651
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1606821651
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1606821651
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1606821651
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1606821651
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1606821651
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 10396 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606821651
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1606821651
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1606821651
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1606821651
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_98
timestamp 1606821651
transform 1 0 10120 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_110
timestamp 1606821651
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 11224 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_106
timestamp 1606821651
transform 1 0 10856 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 11316 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_115
timestamp 1606821651
transform 1 0 11684 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 11592 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1606821651
transform 1 0 11868 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1606821651
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_121
timestamp 1606821651
transform 1 0 12236 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606821651
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606821651
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 12420 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_125
timestamp 1606821651
transform 1 0 12604 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1606821651
transform 1 0 14168 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 14352 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 12696 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 13432 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13340 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_132
timestamp 1606821651
transform 1 0 13248 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_140
timestamp 1606821651
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_129
timestamp 1606821651
transform 1 0 12972 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_142
timestamp 1606821651
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_152
timestamp 1606821651
transform 1 0 15088 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_146
timestamp 1606821651
transform 1 0 14536 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606821651
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1606821651
transform 1 0 14720 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_160
timestamp 1606821651
transform 1 0 15824 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156
timestamp 1606821651
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1606821651
transform 1 0 15548 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1606821651
transform 1 0 16008 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1606821651
transform 1 0 16376 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1606821651
transform 1 0 16376 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_172
timestamp 1606821651
transform 1 0 16928 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16560 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1606821651
transform 1 0 16560 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1606821651
transform 1 0 17296 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_177
timestamp 1606821651
transform 1 0 17388 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1606821651
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606821651
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606821651
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1606821651
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_0_187
timestamp 1606821651
transform 1 0 18308 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_192
timestamp 1606821651
transform 1 0 18768 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1606821651
transform 1 0 18400 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_195
timestamp 1606821651
transform 1 0 19044 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1606821651
transform 1 0 18952 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_198
timestamp 1606821651
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1606821651
transform 1 0 19504 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1606821651
transform 1 0 19412 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_203
timestamp 1606821651
transform 1 0 19780 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_204
timestamp 1606821651
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1606821651
transform 1 0 19964 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_208
timestamp 1606821651
transform 1 0 20240 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_209
timestamp 1606821651
transform 1 0 20332 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_213
timestamp 1606821651
transform 1 0 20700 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1606821651
transform 1 0 20332 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1606821651
transform 1 0 20516 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1606821651
transform 1 0 20884 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1606821651
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606821651
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_219
timestamp 1606821651
transform 1 0 21252 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606821651
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606821651
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606821651
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1606821651
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1606821651
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606821651
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1606821651
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1606821651
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1606821651
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1606821651
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1606821651
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1606821651
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10028 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606821651
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_93
timestamp 1606821651
transform 1 0 9660 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 11684 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_113
timestamp 1606821651
transform 1 0 11500 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 13340 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_131
timestamp 1606821651
transform 1 0 13156 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15640 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606821651
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_149
timestamp 1606821651
transform 1 0 14812 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_154
timestamp 1606821651
transform 1 0 15272 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 17296 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_174
timestamp 1606821651
transform 1 0 17112 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19044 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19780 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_2_192
timestamp 1606821651
transform 1 0 18768 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_201
timestamp 1606821651
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606821651
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606821651
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1606821651
transform 1 0 20332 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1606821651
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1606821651
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1606821651
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606821651
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1606821651
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1606821651
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1606821651
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1606821651
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606821651
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1606821651
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1606821651
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1606821651
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1606821651
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 9108 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_3_86
timestamp 1606821651
transform 1 0 9016 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_103
timestamp 1606821651
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _040_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 11776 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10764 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606821651
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_114
timestamp 1606821651
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_119
timestamp 1606821651
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_123
timestamp 1606821651
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12788 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1606821651
transform 1 0 13984 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_136
timestamp 1606821651
transform 1 0 13616 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1606821651
transform 1 0 14996 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 15732 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_149
timestamp 1606821651
transform 1 0 14812 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_155
timestamp 1606821651
transform 1 0 15364 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_165
timestamp 1606821651
transform 1 0 16284 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1606821651
transform 1 0 17388 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1606821651
transform 1 0 16468 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 18032 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606821651
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_171
timestamp 1606821651
transform 1 0 16836 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1606821651
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1606821651
transform 1 0 19688 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_200
timestamp 1606821651
transform 1 0 19504 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1606821651
transform 1 0 20700 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606821651
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_211
timestamp 1606821651
transform 1 0 20516 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_217
timestamp 1606821651
transform 1 0 21068 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606821651
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1606821651
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1606821651
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606821651
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1606821651
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1606821651
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1606821651
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1606821651
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1606821651
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1606821651
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606821651
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1606821651
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 12052 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1606821651
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_117
timestamp 1606821651
transform 1 0 11868 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1606821651
transform 1 0 13708 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_135
timestamp 1606821651
transform 1 0 13524 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1606821651
transform 1 0 14076 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_145
timestamp 1606821651
transform 1 0 14444 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1606821651
transform 1 0 16284 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1606821651
transform 1 0 14536 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1606821651
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606821651
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_150
timestamp 1606821651
transform 1 0 14904 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_163
timestamp 1606821651
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1606821651
transform 1 0 16928 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1606821651
transform 1 0 17756 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_168
timestamp 1606821651
transform 1 0 16560 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_175
timestamp 1606821651
transform 1 0 17204 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1606821651
transform 1 0 19780 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1606821651
transform 1 0 18768 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_190
timestamp 1606821651
transform 1 0 18584 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_201
timestamp 1606821651
transform 1 0 19596 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606821651
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606821651
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1606821651
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1606821651
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1606821651
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606821651
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1606821651
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1606821651
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1606821651
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1606821651
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606821651
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1606821651
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1606821651
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1606821651
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1606821651
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10304 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1606821651
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_98
timestamp 1606821651
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1606821651
transform 1 0 11868 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1606821651
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606821651
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 11316 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_109
timestamp 1606821651
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_114
timestamp 1606821651
transform 1 0 11592 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1606821651
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13616 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_132
timestamp 1606821651
transform 1 0 13248 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1606821651
transform 1 0 15272 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 15824 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_152
timestamp 1606821651
transform 1 0 15088 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_157
timestamp 1606821651
transform 1 0 15548 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1606821651
transform 1 0 18032 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606821651
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_176
timestamp 1606821651
transform 1 0 17296 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_182
timestamp 1606821651
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_187
timestamp 1606821651
transform 1 0 18308 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 18492 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1606821651
transform 1 0 20148 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_205
timestamp 1606821651
transform 1 0 19964 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606821651
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_216
timestamp 1606821651
transform 1 0 20976 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606821651
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606821651
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1606821651
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1606821651
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1606821651
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1606821651
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606821651
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1606821651
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1606821651
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1606821651
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1606821651
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6808 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606821651
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1606821651
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1606821651
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1606821651
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1606821651
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 8464 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1606821651
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1606821651
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_78
timestamp 1606821651
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 9752 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1606821651
transform 1 0 10120 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606821651
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_93
timestamp 1606821651
transform 1 0 9660 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_103
timestamp 1606821651
transform 1 0 10580 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_96
timestamp 1606821651
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10856 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1606821651
transform 1 0 12512 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1606821651
transform 1 0 11132 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606821651
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_122
timestamp 1606821651
transform 1 0 12328 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_107
timestamp 1606821651
transform 1 0 10948 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1606821651
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1606821651
transform 1 0 14168 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1606821651
transform 1 0 13432 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1606821651
transform 1 0 14444 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_6_133
timestamp 1606821651
transform 1 0 13340 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_141
timestamp 1606821651
transform 1 0 14076 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_132
timestamp 1606821651
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_143
timestamp 1606821651
transform 1 0 14260 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15272 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1606821651
transform 1 0 15640 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606821651
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1606821651
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_154
timestamp 1606821651
transform 1 0 15272 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_167
timestamp 1606821651
transform 1 0 16468 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_174
timestamp 1606821651
transform 1 0 17112 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_170
timestamp 1606821651
transform 1 0 16744 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1606821651
transform 1 0 16652 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_184
timestamp 1606821651
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_182
timestamp 1606821651
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_178
timestamp 1606821651
transform 1 0 17480 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606821651
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1606821651
transform 1 0 18216 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 17204 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 18860 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 19228 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_6_191
timestamp 1606821651
transform 1 0 18676 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_195
timestamp 1606821651
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1606821651
transform 1 0 20884 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606821651
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606821651
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606821651
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_209
timestamp 1606821651
transform 1 0 20332 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1606821651
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_218
timestamp 1606821651
transform 1 0 21160 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_213
timestamp 1606821651
transform 1 0 20700 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_219
timestamp 1606821651
transform 1 0 21252 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606821651
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1606821651
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1606821651
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606821651
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1606821651
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1606821651
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1606821651
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1606821651
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1606821651
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_80
timestamp 1606821651
transform 1 0 8464 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1606821651
transform 1 0 9108 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1606821651
transform 1 0 10672 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606821651
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_86
timestamp 1606821651
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1606821651
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_102
timestamp 1606821651
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 11776 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_8_113
timestamp 1606821651
transform 1 0 11500 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1606821651
transform 1 0 13432 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1606821651
transform 1 0 13892 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_132
timestamp 1606821651
transform 1 0 13248 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_137
timestamp 1606821651
transform 1 0 13708 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1606821651
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606821651
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 16284 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_148
timestamp 1606821651
transform 1 0 14720 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_152
timestamp 1606821651
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_163
timestamp 1606821651
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1606821651
transform 1 0 17848 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16836 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_8_168
timestamp 1606821651
transform 1 0 16560 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_180
timestamp 1606821651
transform 1 0 17664 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 19136 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_191
timestamp 1606821651
transform 1 0 18676 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1606821651
transform 1 0 19044 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606821651
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606821651
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1606821651
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1606821651
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1606821651
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606821651
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1606821651
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1606821651
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1606821651
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1606821651
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606821651
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1606821651
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1606821651
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1606821651
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 8372 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_74
timestamp 1606821651
transform 1 0 7912 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_78
timestamp 1606821651
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1606821651
transform 1 0 10304 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_95
timestamp 1606821651
transform 1 0 9844 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_99
timestamp 1606821651
transform 1 0 10212 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1606821651
transform 1 0 11316 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606821651
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_109
timestamp 1606821651
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1606821651
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_123
timestamp 1606821651
transform 1 0 12420 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 13800 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1606821651
transform 1 0 12788 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_136
timestamp 1606821651
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 15548 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_9_154
timestamp 1606821651
transform 1 0 15272 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1606821651
transform 1 0 17204 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1606821651
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606821651
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_173
timestamp 1606821651
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_178
timestamp 1606821651
transform 1 0 17480 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1606821651
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1606821651
transform 1 0 19872 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_193
timestamp 1606821651
transform 1 0 18860 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_201
timestamp 1606821651
transform 1 0 19596 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606821651
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_213
timestamp 1606821651
transform 1 0 20700 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_219
timestamp 1606821651
transform 1 0 21252 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606821651
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1606821651
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1606821651
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606821651
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1606821651
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1606821651
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1606821651
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1606821651
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1606821651
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1606821651
transform 1 0 8464 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 8832 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10028 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606821651
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1606821651
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_93
timestamp 1606821651
transform 1 0 9660 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 11040 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_106
timestamp 1606821651
transform 1 0 10856 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_124
timestamp 1606821651
transform 1 0 12512 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1606821651
transform 1 0 13892 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12880 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_137
timestamp 1606821651
transform 1 0 13708 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1606821651
transform 1 0 15732 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606821651
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_148
timestamp 1606821651
transform 1 0 14720 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1606821651
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_154
timestamp 1606821651
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_158
timestamp 1606821651
transform 1 0 15640 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 16744 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_168
timestamp 1606821651
transform 1 0 16560 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_186
timestamp 1606821651
transform 1 0 18216 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 18952 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1606821651
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606821651
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606821651
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_210
timestamp 1606821651
transform 1 0 20424 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_218
timestamp 1606821651
transform 1 0 21160 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606821651
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1606821651
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1606821651
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1606821651
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1606821651
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606821651
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1606821651
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1606821651
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1606821651
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1606821651
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 9200 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_86
timestamp 1606821651
transform 1 0 9016 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_104
timestamp 1606821651
transform 1 0 10672 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1606821651
transform 1 0 10856 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606821651
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 11868 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_115
timestamp 1606821651
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1606821651
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13800 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_11_132
timestamp 1606821651
transform 1 0 13248 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1606821651
transform 1 0 15732 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 15180 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_147
timestamp 1606821651
transform 1 0 14628 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_11_156
timestamp 1606821651
transform 1 0 15456 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1606821651
transform 1 0 16744 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606821651
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_168
timestamp 1606821651
transform 1 0 16560 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_179
timestamp 1606821651
transform 1 0 17572 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_184
timestamp 1606821651
transform 1 0 18032 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1606821651
transform 1 0 19688 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1606821651
transform 1 0 18676 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_190
timestamp 1606821651
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_200
timestamp 1606821651
transform 1 0 19504 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606821651
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_211
timestamp 1606821651
transform 1 0 20516 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_219
timestamp 1606821651
transform 1 0 21252 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606821651
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1606821651
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1606821651
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606821651
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1606821651
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1606821651
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1606821651
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1606821651
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8556 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1606821651
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_80
timestamp 1606821651
transform 1 0 8464 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9660 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606821651
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1606821651
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1606821651
transform 1 0 11316 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_109
timestamp 1606821651
transform 1 0 11132 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_120
timestamp 1606821651
transform 1 0 12144 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 12972 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_12_128
timestamp 1606821651
transform 1 0 12880 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_145
timestamp 1606821651
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 15732 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606821651
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_154
timestamp 1606821651
transform 1 0 15272 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_158
timestamp 1606821651
transform 1 0 15640 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1606821651
transform 1 0 17572 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_175
timestamp 1606821651
transform 1 0 17204 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 18584 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_188
timestamp 1606821651
transform 1 0 18400 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_206
timestamp 1606821651
transform 1 0 20056 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606821651
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606821651
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1606821651
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1606821651
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606821651
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606821651
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1606821651
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1606821651
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1606821651
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1606821651
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606821651
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1606821651
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1606821651
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1606821651
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1606821651
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606821651
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1606821651
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1606821651
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1606821651
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1606821651
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1606821651
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 8188 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_13_74
timestamp 1606821651
transform 1 0 7912 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1606821651
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_80
timestamp 1606821651
transform 1 0 8464 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1606821651
transform 1 0 9108 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 10028 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10672 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606821651
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_93
timestamp 1606821651
transform 1 0 9660 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_86
timestamp 1606821651
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1606821651
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_102
timestamp 1606821651
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1606821651
transform 1 0 11684 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 12420 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 12328 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606821651
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1606821651
transform 1 0 11500 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_118
timestamp 1606821651
transform 1 0 11960 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_120
timestamp 1606821651
transform 1 0 12144 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 14444 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1606821651
transform 1 0 14168 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1606821651
transform 1 0 13156 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 14076 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_139
timestamp 1606821651
transform 1 0 13892 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_144
timestamp 1606821651
transform 1 0 14352 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_128
timestamp 1606821651
transform 1 0 12880 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_140
timestamp 1606821651
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1606821651
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1606821651
transform 1 0 16100 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 16100 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606821651
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_161
timestamp 1606821651
transform 1 0 15916 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1606821651
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_169
timestamp 1606821651
transform 1 0 16652 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_175
timestamp 1606821651
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 17388 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1606821651
transform 1 0 16744 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1606821651
transform 1 0 16928 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_183
timestamp 1606821651
transform 1 0 17940 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_179
timestamp 1606821651
transform 1 0 17572 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_180
timestamp 1606821651
transform 1 0 17664 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606821651
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1606821651
transform 1 0 18032 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 18032 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 19044 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1606821651
transform 1 0 20056 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_13_200
timestamp 1606821651
transform 1 0 19504 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_193
timestamp 1606821651
transform 1 0 18860 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1606821651
transform 1 0 20884 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606821651
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606821651
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606821651
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_215
timestamp 1606821651
transform 1 0 20884 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_219
timestamp 1606821651
transform 1 0 21252 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_211
timestamp 1606821651
transform 1 0 20516 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_218
timestamp 1606821651
transform 1 0 21160 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606821651
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1606821651
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1606821651
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1606821651
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1606821651
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606821651
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1606821651
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1606821651
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1606821651
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 8004 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_74
timestamp 1606821651
transform 1 0 7912 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 9660 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 10396 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_91
timestamp 1606821651
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_99
timestamp 1606821651
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_104
timestamp 1606821651
transform 1 0 10672 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1606821651
transform 1 0 11316 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1606821651
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606821651
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_110
timestamp 1606821651
transform 1 0 11224 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1606821651
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1606821651
transform 1 0 13432 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_132
timestamp 1606821651
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_143
timestamp 1606821651
transform 1 0 14260 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 16284 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1606821651
transform 1 0 14536 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1606821651
transform 1 0 15364 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_164
timestamp 1606821651
transform 1 0 16192 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1606821651
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606821651
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1606821651
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_187
timestamp 1606821651
transform 1 0 18308 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 19596 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1606821651
transform 1 0 18584 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_199
timestamp 1606821651
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606821651
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_217
timestamp 1606821651
transform 1 0 21068 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606821651
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1606821651
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1606821651
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606821651
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1606821651
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1606821651
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1606821651
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1606821651
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8556 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1606821651
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_80
timestamp 1606821651
transform 1 0 8464 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606821651
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1606821651
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_102
timestamp 1606821651
transform 1 0 10488 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10948 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_16_106
timestamp 1606821651
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_123
timestamp 1606821651
transform 1 0 12420 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 12880 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_16_127
timestamp 1606821651
transform 1 0 12788 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1606821651
transform 1 0 15548 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606821651
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_148
timestamp 1606821651
transform 1 0 14720 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1606821651
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_154
timestamp 1606821651
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_166
timestamp 1606821651
transform 1 0 16376 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 16560 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1606821651
transform 1 0 18216 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_184
timestamp 1606821651
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1606821651
transform 1 0 19504 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_195
timestamp 1606821651
transform 1 0 19044 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_199
timestamp 1606821651
transform 1 0 19412 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606821651
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606821651
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_209
timestamp 1606821651
transform 1 0 20332 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1606821651
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1606821651
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1606821651
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606821651
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1606821651
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1606821651
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1606821651
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1606821651
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606821651
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1606821651
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1606821651
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1606821651
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 8188 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_17_74
timestamp 1606821651
transform 1 0 7912 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1606821651
transform 1 0 9844 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_93
timestamp 1606821651
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_98
timestamp 1606821651
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1606821651
transform 1 0 11224 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12604 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1606821651
transform 1 0 11500 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606821651
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_123
timestamp 1606821651
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13524 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1606821651
transform 1 0 14352 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_134
timestamp 1606821651
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1606821651
transform 1 0 15548 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_153
timestamp 1606821651
transform 1 0 15180 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_166
timestamp 1606821651
transform 1 0 16376 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1606821651
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16928 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1606821651
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1606821651
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1606821651
transform 1 0 19136 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 19688 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_17_193
timestamp 1606821651
transform 1 0 18860 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_200
timestamp 1606821651
transform 1 0 19504 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606821651
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_218
timestamp 1606821651
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606821651
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1606821651
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1606821651
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1606821651
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1606821651
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1606821651
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1606821651
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1606821651
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7728 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_68
timestamp 1606821651
transform 1 0 7360 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 9660 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1606821651
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_88
timestamp 1606821651
transform 1 0 9200 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_99
timestamp 1606821651
transform 1 0 10212 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 11316 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 12972 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_127
timestamp 1606821651
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_145
timestamp 1606821651
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1606821651
transform 1 0 14628 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1606821651
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 15824 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1606821651
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_150
timestamp 1606821651
transform 1 0 14904 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_157
timestamp 1606821651
transform 1 0 15548 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1606821651
transform 1 0 17572 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_18_176
timestamp 1606821651
transform 1 0 17296 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1606821651
transform 1 0 20240 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 18584 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_188
timestamp 1606821651
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_206
timestamp 1606821651
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1606821651
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606821651
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1606821651
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1606821651
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_218
timestamp 1606821651
transform 1 0 21160 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606821651
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606821651
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1606821651
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1606821651
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1606821651
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1606821651
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1606821651
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1606821651
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1606821651
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1606821651
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1606821651
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1606821651
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1606821651
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1606821651
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1606821651
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1606821651
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1606821651
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 8740 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_19_74
timestamp 1606821651
transform 1 0 7912 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_82
timestamp 1606821651
transform 1 0 8648 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1606821651
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_80
timestamp 1606821651
transform 1 0 8464 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1606821651
transform 1 0 10396 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1606821651
transform 1 0 9844 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1606821651
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_99
timestamp 1606821651
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_88
timestamp 1606821651
transform 1 0 9200 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_93
timestamp 1606821651
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_104
timestamp 1606821651
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1606821651
transform 1 0 11224 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10856 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1606821651
transform 1 0 11408 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_115
timestamp 1606821651
transform 1 0 11684 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 1606821651
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_115
timestamp 1606821651
transform 1 0 11684 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1606821651
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 12052 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_125
timestamp 1606821651
transform 1 0 12604 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 13432 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 13156 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1606821651
transform 1 0 14168 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 12788 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_132
timestamp 1606821651
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_130
timestamp 1606821651
transform 1 0 13064 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_137
timestamp 1606821651
transform 1 0 13708 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_141
timestamp 1606821651
transform 1 0 14076 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1606821651
transform 1 0 16284 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 15088 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1606821651
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1606821651
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_150
timestamp 1606821651
transform 1 0 14904 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1606821651
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_163
timestamp 1606821651
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 17848 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1606821651
transform 1 0 16744 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1606821651
transform 1 0 16652 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 18032 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1606821651
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1606821651
transform 1 0 17664 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_168
timestamp 1606821651
transform 1 0 16560 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_179
timestamp 1606821651
transform 1 0 17572 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_178
timestamp 1606821651
transform 1 0 17480 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1606821651
transform 1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 18768 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1606821651
transform 1 0 19320 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_190
timestamp 1606821651
transform 1 0 18584 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_208
timestamp 1606821651
transform 1 0 20240 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_191
timestamp 1606821651
transform 1 0 18676 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_196
timestamp 1606821651
transform 1 0 19136 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_207
timestamp 1606821651
transform 1 0 20148 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 20424 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606821651
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606821651
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1606821651
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_216
timestamp 1606821651
transform 1 0 20976 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1606821651
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1606821651
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1606821651
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606821651
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1606821651
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1606821651
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1606821651
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1606821651
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1606821651
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1606821651
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1606821651
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1606821651
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1606821651
transform 1 0 8740 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_74
timestamp 1606821651
transform 1 0 7912 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_82
timestamp 1606821651
transform 1 0 8648 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9476 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_21_86
timestamp 1606821651
transform 1 0 9016 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_90
timestamp 1606821651
transform 1 0 9384 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1606821651
transform 1 0 11132 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1606821651
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1606821651
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_107
timestamp 1606821651
transform 1 0 10948 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_118
timestamp 1606821651
transform 1 0 11960 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1606821651
transform 1 0 14444 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1606821651
transform 1 0 13432 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_132
timestamp 1606821651
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_143
timestamp 1606821651
transform 1 0 14260 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1606821651
transform 1 0 15732 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 16284 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 15456 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_154
timestamp 1606821651
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_163
timestamp 1606821651
transform 1 0 16100 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1606821651
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1606821651
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1606821651
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19044 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_1_
timestamp 1606821651
transform 1 0 19780 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_193
timestamp 1606821651
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_201
timestamp 1606821651
transform 1 0 19596 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1606821651
transform 1 0 20792 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606821651
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_212
timestamp 1606821651
transform 1 0 20608 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_218
timestamp 1606821651
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606821651
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1606821651
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1606821651
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1606821651
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1606821651
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1606821651
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6716 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1606821651
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_56
timestamp 1606821651
transform 1 0 6256 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_60
timestamp 1606821651
transform 1 0 6624 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1606821651
transform 1 0 8372 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_77
timestamp 1606821651
transform 1 0 8188 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 9660 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1606821651
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_88
timestamp 1606821651
transform 1 0 9200 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 11684 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 11316 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_109
timestamp 1606821651
transform 1 0 11132 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_114
timestamp 1606821651
transform 1 0 11592 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1606821651
transform 1 0 13340 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 14352 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_131
timestamp 1606821651
transform 1 0 13156 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_142
timestamp 1606821651
transform 1 0 14168 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 16100 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 15272 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1606821651
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_150
timestamp 1606821651
transform 1 0 14904 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_160
timestamp 1606821651
transform 1 0 15824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 17756 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_179
timestamp 1606821651
transform 1 0 17572 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1606821651
transform 1 0 19044 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1606821651
transform 1 0 19596 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_190
timestamp 1606821651
transform 1 0 18584 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_194
timestamp 1606821651
transform 1 0 18952 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_199
timestamp 1606821651
transform 1 0 19412 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1606821651
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606821651
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1606821651
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_210
timestamp 1606821651
transform 1 0 20424 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_218
timestamp 1606821651
transform 1 0 21160 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606821651
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1606821651
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1606821651
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1606821651
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_39
timestamp 1606821651
transform 1 0 4692 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5704 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1606821651
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_47
timestamp 1606821651
transform 1 0 5428 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1606821651
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_62
timestamp 1606821651
transform 1 0 6808 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 7452 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_23_68
timestamp 1606821651
transform 1 0 7360 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10304 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1606821651
transform 1 0 9108 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_85
timestamp 1606821651
transform 1 0 8924 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_96
timestamp 1606821651
transform 1 0 9936 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 12420 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1606821651
transform 1 0 11316 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1606821651
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_109
timestamp 1606821651
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1606821651
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 14352 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 14076 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_139
timestamp 1606821651
transform 1 0 13892 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1606821651
transform 1 0 16192 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_160
timestamp 1606821651
transform 1 0 15824 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1606821651
transform 1 0 16744 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1606821651
transform 1 0 18124 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1606821651
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_168
timestamp 1606821651
transform 1 0 16560 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_179
timestamp 1606821651
transform 1 0 17572 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_184
timestamp 1606821651
transform 1 0 18032 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 19136 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_194
timestamp 1606821651
transform 1 0 18952 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1606821651
transform 1 0 20792 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606821651
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_212
timestamp 1606821651
transform 1 0 20608 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_218
timestamp 1606821651
transform 1 0 21160 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606821651
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1606821651
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1606821651
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1606821651
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1606821651
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1606821651
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6072 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_24_44
timestamp 1606821651
transform 1 0 5152 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_52
timestamp 1606821651
transform 1 0 5888 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1606821651
transform 1 0 7912 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8372 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_70
timestamp 1606821651
transform 1 0 7544 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_77
timestamp 1606821651
transform 1 0 8188 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1606821651
transform 1 0 10488 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 9660 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1606821651
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_88
timestamp 1606821651
transform 1 0 9200 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_99
timestamp 1606821651
transform 1 0 10212 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1606821651
transform 1 0 11868 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_24_111
timestamp 1606821651
transform 1 0 11316 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1606821651
transform 1 0 14168 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_2_
timestamp 1606821651
transform 1 0 12972 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_24_126
timestamp 1606821651
transform 1 0 12696 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_138
timestamp 1606821651
transform 1 0 13800 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 16376 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1606821651
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1606821651
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1606821651
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_163
timestamp 1606821651
transform 1 0 16100 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1606821651
transform 1 0 18032 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_182
timestamp 1606821651
transform 1 0 17848 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_187
timestamp 1606821651
transform 1 0 18308 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1606821651
transform 1 0 20240 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 18492 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_24_205
timestamp 1606821651
transform 1 0 19964 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606821651
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1606821651
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1606821651
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1606821651
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1606821651
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606821651
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1606821651
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1606821651
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1606821651
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1606821651
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6808 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1606821651
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1606821651
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1606821651
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 8740 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_78
timestamp 1606821651
transform 1 0 8280 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_82
timestamp 1606821651
transform 1 0 8648 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 9476 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_89
timestamp 1606821651
transform 1 0 9292 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 12420 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1606821651
transform 1 0 11132 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1606821651
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_107
timestamp 1606821651
transform 1 0 10948 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_118
timestamp 1606821651
transform 1 0 11960 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 14076 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_139
timestamp 1606821651
transform 1 0 13892 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1606821651
transform 1 0 15732 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_157
timestamp 1606821651
transform 1 0 15548 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 18032 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1606821651
transform 1 0 16744 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1606821651
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_168
timestamp 1606821651
transform 1 0 16560 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_179
timestamp 1606821651
transform 1 0 17572 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1606821651
transform 1 0 19780 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_25_200
timestamp 1606821651
transform 1 0 19504 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1606821651
transform 1 0 20792 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606821651
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_212
timestamp 1606821651
transform 1 0 20608 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_218
timestamp 1606821651
transform 1 0 21160 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606821651
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606821651
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1606821651
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1606821651
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1606821651
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1606821651
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1606821651
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1606821651
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1606821651
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1606821651
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1606821651
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1606821651
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1606821651
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_56
timestamp 1606821651
transform 1 0 6256 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1606821651
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1606821651
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_62
timestamp 1606821651
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6992 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1606821651
transform 1 0 6992 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8188 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_1_
timestamp 1606821651
transform 1 0 8648 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_26_73
timestamp 1606821651
transform 1 0 7820 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_80
timestamp 1606821651
transform 1 0 8464 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10396 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l3_in_0_
timestamp 1606821651
transform 1 0 9660 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 9660 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1606821651
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 9292 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_86
timestamp 1606821651
transform 1 0 9016 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_99
timestamp 1606821651
transform 1 0 10212 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_91
timestamp 1606821651
transform 1 0 9476 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_102
timestamp 1606821651
transform 1 0 10488 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1606821651
transform 1 0 11776 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12512 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1606821651
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_3_
timestamp 1606821651
transform 1 0 12052 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1606821651
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_117
timestamp 1606821651
transform 1 0 11868 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_114
timestamp 1606821651
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1606821651
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_123
timestamp 1606821651
transform 1 0 12420 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1606821651
transform 1 0 13064 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 13524 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13708 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_128
timestamp 1606821651
transform 1 0 12880 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_133
timestamp 1606821651
transform 1 0 13340 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_133
timestamp 1606821651
transform 1 0 13340 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1606821651
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1606821651
transform 1 0 15732 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1606821651
transform 1 0 14720 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1606821651
transform 1 0 15732 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1606821651
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_151
timestamp 1606821651
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_157
timestamp 1606821651
transform 1 0 15548 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_146
timestamp 1606821651
transform 1 0 14536 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_157
timestamp 1606821651
transform 1 0 15548 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_175
timestamp 1606821651
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_168
timestamp 1606821651
transform 1 0 16560 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_176
timestamp 1606821651
transform 1 0 17296 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_168
timestamp 1606821651
transform 1 0 16560 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1606821651
transform 1 0 16928 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1606821651
transform 1 0 16836 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1606821651
transform 1 0 17388 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 1606821651
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_187
timestamp 1606821651
transform 1 0 18308 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1606821651
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1606821651
transform 1 0 17480 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 18032 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19688 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1606821651
transform 1 0 18492 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_1_
timestamp 1606821651
transform 1 0 19504 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_198
timestamp 1606821651
transform 1 0 19320 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_200
timestamp 1606821651
transform 1 0 19504 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_208
timestamp 1606821651
transform 1 0 20240 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 20424 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606821651
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606821651
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1606821651
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_209
timestamp 1606821651
transform 1 0 20332 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_213
timestamp 1606821651
transform 1 0 20700 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1606821651
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1606821651
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_216
timestamp 1606821651
transform 1 0 20976 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606821651
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1606821651
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1606821651
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1606821651
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1606821651
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1606821651
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1606821651
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1606821651
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 7544 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_68
timestamp 1606821651
transform 1 0 7360 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1606821651
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_86
timestamp 1606821651
transform 1 0 9016 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_28_102
timestamp 1606821651
transform 1 0 10488 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1606821651
transform 1 0 12512 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 10764 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1606821651
transform 1 0 11500 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_111
timestamp 1606821651
transform 1 0 11316 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_122
timestamp 1606821651
transform 1 0 12328 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_1_
timestamp 1606821651
transform 1 0 12972 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1606821651
transform 1 0 14168 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_127
timestamp 1606821651
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_138
timestamp 1606821651
transform 1 0 13800 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1606821651
transform 1 0 15272 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1606821651
transform 1 0 15732 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1606821651
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1606821651
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_157
timestamp 1606821651
transform 1 0 15548 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 17112 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 16744 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_168
timestamp 1606821651
transform 1 0 16560 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_173
timestamp 1606821651
transform 1 0 17020 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1606821651
transform 1 0 19780 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1606821651
transform 1 0 18768 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_190
timestamp 1606821651
transform 1 0 18584 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_201
timestamp 1606821651
transform 1 0 19596 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1606821651
transform 1 0 20884 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606821651
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1606821651
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_212
timestamp 1606821651
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_218
timestamp 1606821651
transform 1 0 21160 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606821651
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1606821651
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1606821651
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1606821651
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1606821651
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1606821651
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1606821651
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1606821651
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1606821651
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_74
timestamp 1606821651
transform 1 0 7912 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_82
timestamp 1606821651
transform 1 0 8648 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8832 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l3_in_0_
timestamp 1606821651
transform 1 0 9936 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_29_93
timestamp 1606821651
transform 1 0 9660 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1606821651
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1606821651
transform 1 0 11776 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 10948 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1606821651
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_105
timestamp 1606821651
transform 1 0 10764 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_113
timestamp 1606821651
transform 1 0 11500 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1606821651
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13892 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l3_in_0_
timestamp 1606821651
transform 1 0 12880 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_126
timestamp 1606821651
transform 1 0 12696 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_137
timestamp 1606821651
transform 1 0 13708 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1606821651
transform 1 0 15548 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 16284 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_155
timestamp 1606821651
transform 1 0 15364 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_161
timestamp 1606821651
transform 1 0 15916 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_1_
timestamp 1606821651
transform 1 0 18124 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1606821651
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1606821651
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_184
timestamp 1606821651
transform 1 0 18032 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1606821651
transform 1 0 19228 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19780 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_29_194
timestamp 1606821651
transform 1 0 18952 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_201
timestamp 1606821651
transform 1 0 19596 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 20516 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606821651
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_209
timestamp 1606821651
transform 1 0 20332 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_217
timestamp 1606821651
transform 1 0 21068 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606821651
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1606821651
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1606821651
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1606821651
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1606821651
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1606821651
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1606821651
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1606821651
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7728 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_30_68
timestamp 1606821651
transform 1 0 7360 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1606821651
transform 1 0 9936 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10488 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1606821651
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_88
timestamp 1606821651
transform 1 0 9200 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_93
timestamp 1606821651
transform 1 0 9660 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_100
timestamp 1606821651
transform 1 0 10304 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1606821651
transform 1 0 12144 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_118
timestamp 1606821651
transform 1 0 11960 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_124
timestamp 1606821651
transform 1 0 12512 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 12696 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 14352 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_142
timestamp 1606821651
transform 1 0 14168 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15272 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1606821651
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_150
timestamp 1606821651
transform 1 0 14904 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1606821651
transform 1 0 17756 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1606821651
transform 1 0 16928 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_170
timestamp 1606821651
transform 1 0 16744 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_176
timestamp 1606821651
transform 1 0 17296 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_180
timestamp 1606821651
transform 1 0 17664 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_185
timestamp 1606821651
transform 1 0 18124 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1606821651
transform 1 0 19136 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1606821651
transform 1 0 18584 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19688 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_189
timestamp 1606821651
transform 1 0 18492 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1606821651
transform 1 0 18952 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_200
timestamp 1606821651
transform 1 0 19504 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_208
timestamp 1606821651
transform 1 0 20240 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606821651
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1606821651
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1606821651
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1606821651
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606821651
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1606821651
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1606821651
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1606821651
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1606821651
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1606821651
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1606821651
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1606821651
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1606821651
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 8464 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_31_74
timestamp 1606821651
transform 1 0 7912 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 10120 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_96
timestamp 1606821651
transform 1 0 9936 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1606821651
transform 1 0 11776 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 12420 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1606821651
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_114
timestamp 1606821651
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_120
timestamp 1606821651
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1606821651
transform 1 0 14076 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_139
timestamp 1606821651
transform 1 0 13892 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_145
timestamp 1606821651
transform 1 0 14444 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1606821651
transform 1 0 15732 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 14720 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_154
timestamp 1606821651
transform 1 0 15272 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_158
timestamp 1606821651
transform 1 0 15640 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 17020 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 18216 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1606821651
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_168
timestamp 1606821651
transform 1 0 16560 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_172
timestamp 1606821651
transform 1 0 16928 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_179
timestamp 1606821651
transform 1 0 17572 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_184
timestamp 1606821651
transform 1 0 18032 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1606821651
transform 1 0 19044 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 19688 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_192
timestamp 1606821651
transform 1 0 18768 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_199
timestamp 1606821651
transform 1 0 19412 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606821651
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_214
timestamp 1606821651
transform 1 0 20792 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606821651
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1606821651
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1606821651
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1606821651
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1606821651
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1606821651
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1606821651
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1606821651
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_56
timestamp 1606821651
transform 1 0 6256 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1606821651
transform 1 0 6900 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_75
timestamp 1606821651
transform 1 0 8004 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_1_
timestamp 1606821651
transform 1 0 9936 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1606821651
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_87
timestamp 1606821651
transform 1 0 9108 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_94
timestamp 1606821651
transform 1 0 9752 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1606821651
transform 1 0 12604 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1606821651
transform 1 0 10948 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1606821651
transform 1 0 11500 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1606821651
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_105
timestamp 1606821651
transform 1 0 10764 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_111
timestamp 1606821651
transform 1 0 11316 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_122
timestamp 1606821651
transform 1 0 12328 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1606821651
transform 1 0 13524 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1606821651
transform 1 0 14076 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_129
timestamp 1606821651
transform 1 0 12972 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_139
timestamp 1606821651
transform 1 0 13892 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_145
timestamp 1606821651
transform 1 0 14444 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1606821651
transform 1 0 15548 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1606821651
transform 1 0 16100 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1606821651
transform 1 0 14628 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1606821651
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_151
timestamp 1606821651
transform 1 0 14996 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_156
timestamp 1606821651
transform 1 0 15456 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_161
timestamp 1606821651
transform 1 0 15916 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1606821651
transform 1 0 18308 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1606821651
transform 1 0 17204 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1606821651
transform 1 0 16652 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1606821651
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_167
timestamp 1606821651
transform 1 0 16468 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_173
timestamp 1606821651
transform 1 0 17020 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_179
timestamp 1606821651
transform 1 0 17572 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_185
timestamp 1606821651
transform 1 0 18124 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1606821651
transform 1 0 19964 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1606821651
transform 1 0 19412 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1606821651
transform 1 0 18860 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_191
timestamp 1606821651
transform 1 0 18676 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1606821651
transform 1 0 19228 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_203
timestamp 1606821651
transform 1 0 19780 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1606821651
transform 1 0 20516 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606821651
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1606821651
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_209
timestamp 1606821651
transform 1 0 20332 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1606821651
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1606821651
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
<< labels >>
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_1_
port 0 nsew default input
rlabel metal3 s 0 5720 480 5840 6 ccff_head
port 1 nsew default input
rlabel metal3 s 0 17144 480 17264 6 ccff_tail
port 2 nsew default tristate
rlabel metal3 s 22320 3816 22800 3936 6 chanx_right_in[0]
port 3 nsew default input
rlabel metal3 s 22320 8440 22800 8560 6 chanx_right_in[10]
port 4 nsew default input
rlabel metal3 s 22320 8984 22800 9104 6 chanx_right_in[11]
port 5 nsew default input
rlabel metal3 s 22320 9392 22800 9512 6 chanx_right_in[12]
port 6 nsew default input
rlabel metal3 s 22320 9936 22800 10056 6 chanx_right_in[13]
port 7 nsew default input
rlabel metal3 s 22320 10344 22800 10464 6 chanx_right_in[14]
port 8 nsew default input
rlabel metal3 s 22320 10752 22800 10872 6 chanx_right_in[15]
port 9 nsew default input
rlabel metal3 s 22320 11296 22800 11416 6 chanx_right_in[16]
port 10 nsew default input
rlabel metal3 s 22320 11704 22800 11824 6 chanx_right_in[17]
port 11 nsew default input
rlabel metal3 s 22320 12248 22800 12368 6 chanx_right_in[18]
port 12 nsew default input
rlabel metal3 s 22320 12656 22800 12776 6 chanx_right_in[19]
port 13 nsew default input
rlabel metal3 s 22320 4224 22800 4344 6 chanx_right_in[1]
port 14 nsew default input
rlabel metal3 s 22320 4768 22800 4888 6 chanx_right_in[2]
port 15 nsew default input
rlabel metal3 s 22320 5176 22800 5296 6 chanx_right_in[3]
port 16 nsew default input
rlabel metal3 s 22320 5720 22800 5840 6 chanx_right_in[4]
port 17 nsew default input
rlabel metal3 s 22320 6128 22800 6248 6 chanx_right_in[5]
port 18 nsew default input
rlabel metal3 s 22320 6672 22800 6792 6 chanx_right_in[6]
port 19 nsew default input
rlabel metal3 s 22320 7080 22800 7200 6 chanx_right_in[7]
port 20 nsew default input
rlabel metal3 s 22320 7488 22800 7608 6 chanx_right_in[8]
port 21 nsew default input
rlabel metal3 s 22320 8032 22800 8152 6 chanx_right_in[9]
port 22 nsew default input
rlabel metal3 s 22320 13200 22800 13320 6 chanx_right_out[0]
port 23 nsew default tristate
rlabel metal3 s 22320 17824 22800 17944 6 chanx_right_out[10]
port 24 nsew default tristate
rlabel metal3 s 22320 18232 22800 18352 6 chanx_right_out[11]
port 25 nsew default tristate
rlabel metal3 s 22320 18776 22800 18896 6 chanx_right_out[12]
port 26 nsew default tristate
rlabel metal3 s 22320 19184 22800 19304 6 chanx_right_out[13]
port 27 nsew default tristate
rlabel metal3 s 22320 19728 22800 19848 6 chanx_right_out[14]
port 28 nsew default tristate
rlabel metal3 s 22320 20136 22800 20256 6 chanx_right_out[15]
port 29 nsew default tristate
rlabel metal3 s 22320 20544 22800 20664 6 chanx_right_out[16]
port 30 nsew default tristate
rlabel metal3 s 22320 21088 22800 21208 6 chanx_right_out[17]
port 31 nsew default tristate
rlabel metal3 s 22320 21496 22800 21616 6 chanx_right_out[18]
port 32 nsew default tristate
rlabel metal3 s 22320 22040 22800 22160 6 chanx_right_out[19]
port 33 nsew default tristate
rlabel metal3 s 22320 13608 22800 13728 6 chanx_right_out[1]
port 34 nsew default tristate
rlabel metal3 s 22320 14016 22800 14136 6 chanx_right_out[2]
port 35 nsew default tristate
rlabel metal3 s 22320 14560 22800 14680 6 chanx_right_out[3]
port 36 nsew default tristate
rlabel metal3 s 22320 14968 22800 15088 6 chanx_right_out[4]
port 37 nsew default tristate
rlabel metal3 s 22320 15512 22800 15632 6 chanx_right_out[5]
port 38 nsew default tristate
rlabel metal3 s 22320 15920 22800 16040 6 chanx_right_out[6]
port 39 nsew default tristate
rlabel metal3 s 22320 16464 22800 16584 6 chanx_right_out[7]
port 40 nsew default tristate
rlabel metal3 s 22320 16872 22800 16992 6 chanx_right_out[8]
port 41 nsew default tristate
rlabel metal3 s 22320 17280 22800 17400 6 chanx_right_out[9]
port 42 nsew default tristate
rlabel metal2 s 846 0 902 480 6 chany_bottom_in[0]
port 43 nsew default input
rlabel metal2 s 6366 0 6422 480 6 chany_bottom_in[10]
port 44 nsew default input
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_in[11]
port 45 nsew default input
rlabel metal2 s 7470 0 7526 480 6 chany_bottom_in[12]
port 46 nsew default input
rlabel metal2 s 8022 0 8078 480 6 chany_bottom_in[13]
port 47 nsew default input
rlabel metal2 s 8574 0 8630 480 6 chany_bottom_in[14]
port 48 nsew default input
rlabel metal2 s 9126 0 9182 480 6 chany_bottom_in[15]
port 49 nsew default input
rlabel metal2 s 9678 0 9734 480 6 chany_bottom_in[16]
port 50 nsew default input
rlabel metal2 s 10230 0 10286 480 6 chany_bottom_in[17]
port 51 nsew default input
rlabel metal2 s 10782 0 10838 480 6 chany_bottom_in[18]
port 52 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[19]
port 53 nsew default input
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_in[1]
port 54 nsew default input
rlabel metal2 s 1950 0 2006 480 6 chany_bottom_in[2]
port 55 nsew default input
rlabel metal2 s 2502 0 2558 480 6 chany_bottom_in[3]
port 56 nsew default input
rlabel metal2 s 3054 0 3110 480 6 chany_bottom_in[4]
port 57 nsew default input
rlabel metal2 s 3606 0 3662 480 6 chany_bottom_in[5]
port 58 nsew default input
rlabel metal2 s 4158 0 4214 480 6 chany_bottom_in[6]
port 59 nsew default input
rlabel metal2 s 4710 0 4766 480 6 chany_bottom_in[7]
port 60 nsew default input
rlabel metal2 s 5262 0 5318 480 6 chany_bottom_in[8]
port 61 nsew default input
rlabel metal2 s 5814 0 5870 480 6 chany_bottom_in[9]
port 62 nsew default input
rlabel metal2 s 11978 0 12034 480 6 chany_bottom_out[0]
port 63 nsew default tristate
rlabel metal2 s 17498 0 17554 480 6 chany_bottom_out[10]
port 64 nsew default tristate
rlabel metal2 s 18050 0 18106 480 6 chany_bottom_out[11]
port 65 nsew default tristate
rlabel metal2 s 18602 0 18658 480 6 chany_bottom_out[12]
port 66 nsew default tristate
rlabel metal2 s 19154 0 19210 480 6 chany_bottom_out[13]
port 67 nsew default tristate
rlabel metal2 s 19706 0 19762 480 6 chany_bottom_out[14]
port 68 nsew default tristate
rlabel metal2 s 20258 0 20314 480 6 chany_bottom_out[15]
port 69 nsew default tristate
rlabel metal2 s 20810 0 20866 480 6 chany_bottom_out[16]
port 70 nsew default tristate
rlabel metal2 s 21362 0 21418 480 6 chany_bottom_out[17]
port 71 nsew default tristate
rlabel metal2 s 21914 0 21970 480 6 chany_bottom_out[18]
port 72 nsew default tristate
rlabel metal2 s 22466 0 22522 480 6 chany_bottom_out[19]
port 73 nsew default tristate
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_out[1]
port 74 nsew default tristate
rlabel metal2 s 13082 0 13138 480 6 chany_bottom_out[2]
port 75 nsew default tristate
rlabel metal2 s 13634 0 13690 480 6 chany_bottom_out[3]
port 76 nsew default tristate
rlabel metal2 s 14186 0 14242 480 6 chany_bottom_out[4]
port 77 nsew default tristate
rlabel metal2 s 14738 0 14794 480 6 chany_bottom_out[5]
port 78 nsew default tristate
rlabel metal2 s 15290 0 15346 480 6 chany_bottom_out[6]
port 79 nsew default tristate
rlabel metal2 s 15842 0 15898 480 6 chany_bottom_out[7]
port 80 nsew default tristate
rlabel metal2 s 16394 0 16450 480 6 chany_bottom_out[8]
port 81 nsew default tristate
rlabel metal2 s 16946 0 17002 480 6 chany_bottom_out[9]
port 82 nsew default tristate
rlabel metal2 s 846 22320 902 22800 6 chany_top_in[0]
port 83 nsew default input
rlabel metal2 s 6366 22320 6422 22800 6 chany_top_in[10]
port 84 nsew default input
rlabel metal2 s 6918 22320 6974 22800 6 chany_top_in[11]
port 85 nsew default input
rlabel metal2 s 7470 22320 7526 22800 6 chany_top_in[12]
port 86 nsew default input
rlabel metal2 s 8022 22320 8078 22800 6 chany_top_in[13]
port 87 nsew default input
rlabel metal2 s 8574 22320 8630 22800 6 chany_top_in[14]
port 88 nsew default input
rlabel metal2 s 9126 22320 9182 22800 6 chany_top_in[15]
port 89 nsew default input
rlabel metal2 s 9678 22320 9734 22800 6 chany_top_in[16]
port 90 nsew default input
rlabel metal2 s 10230 22320 10286 22800 6 chany_top_in[17]
port 91 nsew default input
rlabel metal2 s 10782 22320 10838 22800 6 chany_top_in[18]
port 92 nsew default input
rlabel metal2 s 11334 22320 11390 22800 6 chany_top_in[19]
port 93 nsew default input
rlabel metal2 s 1398 22320 1454 22800 6 chany_top_in[1]
port 94 nsew default input
rlabel metal2 s 1950 22320 2006 22800 6 chany_top_in[2]
port 95 nsew default input
rlabel metal2 s 2502 22320 2558 22800 6 chany_top_in[3]
port 96 nsew default input
rlabel metal2 s 3054 22320 3110 22800 6 chany_top_in[4]
port 97 nsew default input
rlabel metal2 s 3606 22320 3662 22800 6 chany_top_in[5]
port 98 nsew default input
rlabel metal2 s 4158 22320 4214 22800 6 chany_top_in[6]
port 99 nsew default input
rlabel metal2 s 4710 22320 4766 22800 6 chany_top_in[7]
port 100 nsew default input
rlabel metal2 s 5262 22320 5318 22800 6 chany_top_in[8]
port 101 nsew default input
rlabel metal2 s 5814 22320 5870 22800 6 chany_top_in[9]
port 102 nsew default input
rlabel metal2 s 11978 22320 12034 22800 6 chany_top_out[0]
port 103 nsew default tristate
rlabel metal2 s 17498 22320 17554 22800 6 chany_top_out[10]
port 104 nsew default tristate
rlabel metal2 s 18050 22320 18106 22800 6 chany_top_out[11]
port 105 nsew default tristate
rlabel metal2 s 18602 22320 18658 22800 6 chany_top_out[12]
port 106 nsew default tristate
rlabel metal2 s 19154 22320 19210 22800 6 chany_top_out[13]
port 107 nsew default tristate
rlabel metal2 s 19706 22320 19762 22800 6 chany_top_out[14]
port 108 nsew default tristate
rlabel metal2 s 20258 22320 20314 22800 6 chany_top_out[15]
port 109 nsew default tristate
rlabel metal2 s 20810 22320 20866 22800 6 chany_top_out[16]
port 110 nsew default tristate
rlabel metal2 s 21362 22320 21418 22800 6 chany_top_out[17]
port 111 nsew default tristate
rlabel metal2 s 21914 22320 21970 22800 6 chany_top_out[18]
port 112 nsew default tristate
rlabel metal2 s 22466 22320 22522 22800 6 chany_top_out[19]
port 113 nsew default tristate
rlabel metal2 s 12530 22320 12586 22800 6 chany_top_out[1]
port 114 nsew default tristate
rlabel metal2 s 13082 22320 13138 22800 6 chany_top_out[2]
port 115 nsew default tristate
rlabel metal2 s 13634 22320 13690 22800 6 chany_top_out[3]
port 116 nsew default tristate
rlabel metal2 s 14186 22320 14242 22800 6 chany_top_out[4]
port 117 nsew default tristate
rlabel metal2 s 14738 22320 14794 22800 6 chany_top_out[5]
port 118 nsew default tristate
rlabel metal2 s 15290 22320 15346 22800 6 chany_top_out[6]
port 119 nsew default tristate
rlabel metal2 s 15842 22320 15898 22800 6 chany_top_out[7]
port 120 nsew default tristate
rlabel metal2 s 16394 22320 16450 22800 6 chany_top_out[8]
port 121 nsew default tristate
rlabel metal2 s 16946 22320 17002 22800 6 chany_top_out[9]
port 122 nsew default tristate
rlabel metal3 s 22320 22448 22800 22568 6 prog_clk_0_E_in
port 123 nsew default input
rlabel metal3 s 22320 144 22800 264 6 right_bottom_grid_pin_34_
port 124 nsew default input
rlabel metal3 s 22320 552 22800 672 6 right_bottom_grid_pin_35_
port 125 nsew default input
rlabel metal3 s 22320 960 22800 1080 6 right_bottom_grid_pin_36_
port 126 nsew default input
rlabel metal3 s 22320 1504 22800 1624 6 right_bottom_grid_pin_37_
port 127 nsew default input
rlabel metal3 s 22320 1912 22800 2032 6 right_bottom_grid_pin_38_
port 128 nsew default input
rlabel metal3 s 22320 2456 22800 2576 6 right_bottom_grid_pin_39_
port 129 nsew default input
rlabel metal3 s 22320 2864 22800 2984 6 right_bottom_grid_pin_40_
port 130 nsew default input
rlabel metal3 s 22320 3408 22800 3528 6 right_bottom_grid_pin_41_
port 131 nsew default input
rlabel metal2 s 294 22320 350 22800 6 top_left_grid_pin_1_
port 132 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 133 nsew default input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 134 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22800
<< end >>
