magic
tech EFS8A
magscale 1 2
timestamp 1604337009
<< locali >>
rect 5273 22559 5307 22661
rect 19901 21879 19935 22117
rect 23765 21335 23799 21641
rect 6469 20247 6503 20349
rect 19533 20247 19567 20349
rect 16129 18139 16163 18377
rect 13185 13923 13219 14025
rect 12081 10455 12115 10761
<< viali >>
rect 13001 25449 13035 25483
rect 14105 25449 14139 25483
rect 18521 25449 18555 25483
rect 21373 25449 21407 25483
rect 24225 25449 24259 25483
rect 25329 25449 25363 25483
rect 5089 25381 5123 25415
rect 8493 25381 8527 25415
rect 15761 25381 15795 25415
rect 4813 25313 4847 25347
rect 8585 25313 8619 25347
rect 11069 25313 11103 25347
rect 11345 25313 11379 25347
rect 12817 25313 12851 25347
rect 13921 25313 13955 25347
rect 15485 25313 15519 25347
rect 16957 25313 16991 25347
rect 18337 25313 18371 25347
rect 19441 25313 19475 25347
rect 21189 25313 21223 25347
rect 22293 25313 22327 25347
rect 24041 25313 24075 25347
rect 25145 25313 25179 25347
rect 1685 25245 1719 25279
rect 8493 25245 8527 25279
rect 13461 25245 13495 25279
rect 17141 25245 17175 25279
rect 19625 25177 19659 25211
rect 22477 25177 22511 25211
rect 4353 25109 4387 25143
rect 7757 25109 7791 25143
rect 8033 25109 8067 25143
rect 10885 25109 10919 25143
rect 14473 25109 14507 25143
rect 8677 24905 8711 24939
rect 22661 24905 22695 24939
rect 10885 24837 10919 24871
rect 12541 24837 12575 24871
rect 21557 24837 21591 24871
rect 1593 24769 1627 24803
rect 2881 24769 2915 24803
rect 3893 24769 3927 24803
rect 4537 24769 4571 24803
rect 4721 24769 4755 24803
rect 7573 24769 7607 24803
rect 10609 24769 10643 24803
rect 11437 24769 11471 24803
rect 15577 24769 15611 24803
rect 16037 24769 16071 24803
rect 18337 24769 18371 24803
rect 23489 24769 23523 24803
rect 2145 24701 2179 24735
rect 12265 24701 12299 24735
rect 13093 24701 13127 24735
rect 14841 24701 14875 24735
rect 15761 24701 15795 24735
rect 16497 24701 16531 24735
rect 18061 24701 18095 24735
rect 18797 24701 18831 24735
rect 19349 24701 19383 24735
rect 20085 24701 20119 24735
rect 20637 24701 20671 24735
rect 21189 24701 21223 24735
rect 21741 24701 21775 24735
rect 22293 24701 22327 24735
rect 23673 24701 23707 24735
rect 24777 24701 24811 24735
rect 25329 24701 25363 24735
rect 2421 24633 2455 24667
rect 3617 24633 3651 24667
rect 4629 24633 4663 24667
rect 8033 24633 8067 24667
rect 8309 24633 8343 24667
rect 10333 24633 10367 24667
rect 11161 24633 11195 24667
rect 11345 24633 11379 24667
rect 11897 24633 11931 24667
rect 12817 24633 12851 24667
rect 14013 24633 14047 24667
rect 14565 24633 14599 24667
rect 19165 24633 19199 24667
rect 19625 24633 19659 24667
rect 1961 24565 1995 24599
rect 4159 24565 4193 24599
rect 5089 24565 5123 24599
rect 5641 24565 5675 24599
rect 7113 24565 7147 24599
rect 7747 24565 7781 24599
rect 8217 24565 8251 24599
rect 9137 24565 9171 24599
rect 13001 24565 13035 24599
rect 13645 24565 13679 24599
rect 14279 24565 14313 24599
rect 14749 24565 14783 24599
rect 15301 24565 15335 24599
rect 16957 24565 16991 24599
rect 17877 24565 17911 24599
rect 20821 24565 20855 24599
rect 21925 24565 21959 24599
rect 23857 24565 23891 24599
rect 24225 24565 24259 24599
rect 24961 24565 24995 24599
rect 25697 24565 25731 24599
rect 2513 24361 2547 24395
rect 8401 24361 8435 24395
rect 10057 24361 10091 24395
rect 10885 24361 10919 24395
rect 12449 24361 12483 24395
rect 19441 24361 19475 24395
rect 24869 24361 24903 24395
rect 1869 24293 1903 24327
rect 2053 24293 2087 24327
rect 2881 24293 2915 24327
rect 7297 24293 7331 24327
rect 7941 24293 7975 24327
rect 8033 24293 8067 24327
rect 11336 24293 11370 24327
rect 14197 24293 14231 24327
rect 17509 24293 17543 24327
rect 18797 24293 18831 24327
rect 23673 24293 23707 24327
rect 5172 24225 5206 24259
rect 7757 24225 7791 24259
rect 14289 24225 14323 24259
rect 15577 24225 15611 24259
rect 16865 24225 16899 24259
rect 18521 24225 18555 24259
rect 21833 24225 21867 24259
rect 22569 24225 22603 24259
rect 24685 24225 24719 24259
rect 2145 24157 2179 24191
rect 4905 24157 4939 24191
rect 11069 24157 11103 24191
rect 13553 24157 13587 24191
rect 14105 24157 14139 24191
rect 15853 24157 15887 24191
rect 17509 24157 17543 24191
rect 17601 24157 17635 24191
rect 19809 24157 19843 24191
rect 22109 24157 22143 24191
rect 23581 24157 23615 24191
rect 23765 24157 23799 24191
rect 1593 24089 1627 24123
rect 13093 24089 13127 24123
rect 16497 24089 16531 24123
rect 24133 24089 24167 24123
rect 4353 24021 4387 24055
rect 6285 24021 6319 24055
rect 7481 24021 7515 24055
rect 13737 24021 13771 24055
rect 14749 24021 14783 24055
rect 17049 24021 17083 24055
rect 18153 24021 18187 24055
rect 20361 24021 20395 24055
rect 22937 24021 22971 24055
rect 23213 24021 23247 24055
rect 4169 23817 4203 23851
rect 7389 23817 7423 23851
rect 8861 23817 8895 23851
rect 9413 23817 9447 23851
rect 10057 23817 10091 23851
rect 12725 23817 12759 23851
rect 16497 23817 16531 23851
rect 21465 23817 21499 23851
rect 23121 23817 23155 23851
rect 24041 23817 24075 23851
rect 9781 23749 9815 23783
rect 16313 23749 16347 23783
rect 18153 23749 18187 23783
rect 19165 23749 19199 23783
rect 20085 23749 20119 23783
rect 22109 23749 22143 23783
rect 1409 23681 1443 23715
rect 4261 23681 4295 23715
rect 10609 23681 10643 23715
rect 19533 23681 19567 23715
rect 20545 23681 20579 23715
rect 22477 23681 22511 23715
rect 24133 23681 24167 23715
rect 4528 23613 4562 23647
rect 7481 23613 7515 23647
rect 11161 23613 11195 23647
rect 12173 23613 12207 23647
rect 12541 23613 12575 23647
rect 13645 23613 13679 23647
rect 15945 23613 15979 23647
rect 21833 23613 21867 23647
rect 1654 23545 1688 23579
rect 3801 23545 3835 23579
rect 6653 23545 6687 23579
rect 7748 23545 7782 23579
rect 10333 23545 10367 23579
rect 10517 23545 10551 23579
rect 13912 23545 13946 23579
rect 16773 23545 16807 23579
rect 16957 23545 16991 23579
rect 17049 23545 17083 23579
rect 17877 23545 17911 23579
rect 18429 23545 18463 23579
rect 18705 23545 18739 23579
rect 20637 23545 20671 23579
rect 21189 23545 21223 23579
rect 22661 23545 22695 23579
rect 24378 23545 24412 23579
rect 2789 23477 2823 23511
rect 3433 23477 3467 23511
rect 5641 23477 5675 23511
rect 6193 23477 6227 23511
rect 11529 23477 11563 23511
rect 13093 23477 13127 23511
rect 13553 23477 13587 23511
rect 15025 23477 15059 23511
rect 17509 23477 17543 23511
rect 18613 23477 18647 23511
rect 19901 23477 19935 23511
rect 20545 23477 20579 23511
rect 22569 23477 22603 23511
rect 25513 23477 25547 23511
rect 2881 23273 2915 23307
rect 4261 23273 4295 23307
rect 5825 23273 5859 23307
rect 6929 23273 6963 23307
rect 16221 23273 16255 23307
rect 16681 23273 16715 23307
rect 23213 23273 23247 23307
rect 24869 23273 24903 23307
rect 1768 23205 1802 23239
rect 4712 23205 4746 23239
rect 7021 23205 7055 23239
rect 7481 23205 7515 23239
rect 8401 23205 8435 23239
rect 8585 23205 8619 23239
rect 9505 23205 9539 23239
rect 11152 23205 11186 23239
rect 14013 23205 14047 23239
rect 14197 23205 14231 23239
rect 14657 23205 14691 23239
rect 15761 23205 15795 23239
rect 17325 23205 17359 23239
rect 19809 23205 19843 23239
rect 21158 23205 21192 23239
rect 23765 23205 23799 23239
rect 23949 23205 23983 23239
rect 25237 23205 25271 23239
rect 1501 23137 1535 23171
rect 3525 23137 3559 23171
rect 4445 23137 4479 23171
rect 7941 23137 7975 23171
rect 10885 23137 10919 23171
rect 14289 23137 14323 23171
rect 15485 23137 15519 23171
rect 17141 23137 17175 23171
rect 20913 23137 20947 23171
rect 24961 23137 24995 23171
rect 8677 23069 8711 23103
rect 9689 23069 9723 23103
rect 13553 23069 13587 23103
rect 17417 23069 17451 23103
rect 19809 23069 19843 23103
rect 19901 23069 19935 23103
rect 24041 23069 24075 23103
rect 8125 23001 8159 23035
rect 10149 23001 10183 23035
rect 13737 23001 13771 23035
rect 16865 23001 16899 23035
rect 3801 22933 3835 22967
rect 10609 22933 10643 22967
rect 12265 22933 12299 22967
rect 13185 22933 13219 22967
rect 15025 22933 15059 22967
rect 18153 22933 18187 22967
rect 18797 22933 18831 22967
rect 19165 22933 19199 22967
rect 19349 22933 19383 22967
rect 20361 22933 20395 22967
rect 22293 22933 22327 22967
rect 23489 22933 23523 22967
rect 24409 22933 24443 22967
rect 1501 22729 1535 22763
rect 4169 22729 4203 22763
rect 4445 22729 4479 22763
rect 5457 22729 5491 22763
rect 5733 22729 5767 22763
rect 7757 22729 7791 22763
rect 9597 22729 9631 22763
rect 10241 22729 10275 22763
rect 10609 22729 10643 22763
rect 10885 22729 10919 22763
rect 14105 22729 14139 22763
rect 16313 22729 16347 22763
rect 17693 22729 17727 22763
rect 18613 22729 18647 22763
rect 21649 22729 21683 22763
rect 23029 22729 23063 22763
rect 25421 22729 25455 22763
rect 5273 22661 5307 22695
rect 8125 22661 8159 22695
rect 12541 22661 12575 22695
rect 18797 22661 18831 22695
rect 24133 22661 24167 22695
rect 2881 22593 2915 22627
rect 3249 22593 3283 22627
rect 4905 22593 4939 22627
rect 8217 22593 8251 22627
rect 14657 22593 14691 22627
rect 15025 22593 15059 22627
rect 16129 22593 16163 22627
rect 16773 22593 16807 22627
rect 16865 22593 16899 22627
rect 19349 22593 19383 22627
rect 24593 22593 24627 22627
rect 25053 22593 25087 22627
rect 25605 22593 25639 22627
rect 1777 22525 1811 22559
rect 2421 22525 2455 22559
rect 2973 22525 3007 22559
rect 4997 22525 5031 22559
rect 5273 22525 5307 22559
rect 6469 22525 6503 22559
rect 6837 22525 6871 22559
rect 11161 22525 11195 22559
rect 13461 22525 13495 22559
rect 15761 22525 15795 22559
rect 19073 22525 19107 22559
rect 20269 22525 20303 22559
rect 20536 22525 20570 22559
rect 23489 22525 23523 22559
rect 23949 22525 23983 22559
rect 2053 22457 2087 22491
rect 4905 22457 4939 22491
rect 7113 22457 7147 22491
rect 8462 22457 8496 22491
rect 11437 22457 11471 22491
rect 12265 22457 12299 22491
rect 12817 22457 12851 22491
rect 13093 22457 13127 22491
rect 13921 22457 13955 22491
rect 14381 22457 14415 22491
rect 14565 22457 14599 22491
rect 16773 22457 16807 22491
rect 19257 22457 19291 22491
rect 20177 22457 20211 22491
rect 24593 22457 24627 22491
rect 24685 22457 24719 22491
rect 1961 22389 1995 22423
rect 3801 22389 3835 22423
rect 6193 22389 6227 22423
rect 11345 22389 11379 22423
rect 11805 22389 11839 22423
rect 13001 22389 13035 22423
rect 17233 22389 17267 22423
rect 19809 22389 19843 22423
rect 22293 22389 22327 22423
rect 3801 22185 3835 22219
rect 5181 22185 5215 22219
rect 5457 22185 5491 22219
rect 8953 22185 8987 22219
rect 10241 22185 10275 22219
rect 11161 22185 11195 22219
rect 11253 22185 11287 22219
rect 13645 22185 13679 22219
rect 14933 22185 14967 22219
rect 16773 22185 16807 22219
rect 20085 22185 20119 22219
rect 22845 22185 22879 22219
rect 23489 22185 23523 22219
rect 6561 22117 6595 22151
rect 8125 22117 8159 22151
rect 12081 22117 12115 22151
rect 14289 22117 14323 22151
rect 15853 22117 15887 22151
rect 17110 22117 17144 22151
rect 19901 22117 19935 22151
rect 21557 22117 21591 22151
rect 24102 22117 24136 22151
rect 1501 22049 1535 22083
rect 1768 22049 1802 22083
rect 4353 22049 4387 22083
rect 6653 22049 6687 22083
rect 7389 22049 7423 22083
rect 8585 22049 8619 22083
rect 9505 22049 9539 22083
rect 12521 22049 12555 22083
rect 15945 22049 15979 22083
rect 16865 22049 16899 22083
rect 19349 22049 19383 22083
rect 19625 22049 19659 22083
rect 4629 21981 4663 22015
rect 6561 21981 6595 22015
rect 8125 21981 8159 22015
rect 8217 21981 8251 22015
rect 10241 21981 10275 22015
rect 10333 21981 10367 22015
rect 12265 21981 12299 22015
rect 15853 21981 15887 22015
rect 3433 21913 3467 21947
rect 7665 21913 7699 21947
rect 9781 21913 9815 21947
rect 16405 21913 16439 21947
rect 20913 22049 20947 22083
rect 22661 22049 22695 22083
rect 22937 21981 22971 22015
rect 23857 21981 23891 22015
rect 22385 21913 22419 21947
rect 2881 21845 2915 21879
rect 5825 21845 5859 21879
rect 6101 21845 6135 21879
rect 7021 21845 7055 21879
rect 10793 21845 10827 21879
rect 11713 21845 11747 21879
rect 14657 21845 14691 21879
rect 15393 21845 15427 21879
rect 18245 21845 18279 21879
rect 18981 21845 19015 21879
rect 19901 21845 19935 21879
rect 20545 21845 20579 21879
rect 21097 21845 21131 21879
rect 22109 21845 22143 21879
rect 25237 21845 25271 21879
rect 2881 21641 2915 21675
rect 3985 21641 4019 21675
rect 8861 21641 8895 21675
rect 10425 21641 10459 21675
rect 10609 21641 10643 21675
rect 11897 21641 11931 21675
rect 12541 21641 12575 21675
rect 14197 21641 14231 21675
rect 16497 21641 16531 21675
rect 17785 21641 17819 21675
rect 18981 21641 19015 21675
rect 19901 21641 19935 21675
rect 21925 21641 21959 21675
rect 23121 21641 23155 21675
rect 23765 21641 23799 21675
rect 23857 21641 23891 21675
rect 24685 21641 24719 21675
rect 1501 21573 1535 21607
rect 3065 21573 3099 21607
rect 5273 21573 5307 21607
rect 8217 21573 8251 21607
rect 20545 21573 20579 21607
rect 22109 21573 22143 21607
rect 3525 21505 3559 21539
rect 5733 21505 5767 21539
rect 11161 21505 11195 21539
rect 13461 21505 13495 21539
rect 14657 21505 14691 21539
rect 16865 21505 16899 21539
rect 18797 21505 18831 21539
rect 19441 21505 19475 21539
rect 21097 21505 21131 21539
rect 22569 21505 22603 21539
rect 2421 21437 2455 21471
rect 3617 21437 3651 21471
rect 5089 21437 5123 21471
rect 5825 21437 5859 21471
rect 6193 21437 6227 21471
rect 6837 21437 6871 21471
rect 12265 21437 12299 21471
rect 12817 21437 12851 21471
rect 15301 21437 15335 21471
rect 19533 21437 19567 21471
rect 22661 21437 22695 21471
rect 1777 21369 1811 21403
rect 2053 21369 2087 21403
rect 3525 21369 3559 21403
rect 4721 21369 4755 21403
rect 5733 21369 5767 21403
rect 7082 21369 7116 21403
rect 10885 21369 10919 21403
rect 13093 21369 13127 21403
rect 14657 21369 14691 21403
rect 14749 21369 14783 21403
rect 15761 21369 15795 21403
rect 16957 21369 16991 21403
rect 17049 21369 17083 21403
rect 18429 21369 18463 21403
rect 19441 21369 19475 21403
rect 20821 21369 20855 21403
rect 21557 21369 21591 21403
rect 23489 21369 23523 21403
rect 24961 21437 24995 21471
rect 25237 21369 25271 21403
rect 1961 21301 1995 21335
rect 6653 21301 6687 21335
rect 9137 21301 9171 21335
rect 9505 21301 9539 21335
rect 10057 21301 10091 21335
rect 11069 21301 11103 21335
rect 13001 21301 13035 21335
rect 14013 21301 14047 21335
rect 16313 21301 16347 21335
rect 17417 21301 17451 21335
rect 20269 21301 20303 21335
rect 21005 21301 21039 21335
rect 22569 21301 22603 21335
rect 23765 21301 23799 21335
rect 24409 21301 24443 21335
rect 25145 21301 25179 21335
rect 2605 21097 2639 21131
rect 2973 21097 3007 21131
rect 3433 21097 3467 21131
rect 6469 21097 6503 21131
rect 7665 21097 7699 21131
rect 9965 21097 9999 21131
rect 11989 21097 12023 21131
rect 13645 21097 13679 21131
rect 14105 21097 14139 21131
rect 14565 21097 14599 21131
rect 16405 21097 16439 21131
rect 16865 21097 16899 21131
rect 18521 21097 18555 21131
rect 19809 21097 19843 21131
rect 20453 21097 20487 21131
rect 22293 21097 22327 21131
rect 22937 21097 22971 21131
rect 25421 21097 25455 21131
rect 2145 21029 2179 21063
rect 8401 21029 8435 21063
rect 8493 21029 8527 21063
rect 10854 21029 10888 21063
rect 15853 21029 15887 21063
rect 19441 21029 19475 21063
rect 24225 21029 24259 21063
rect 24777 21029 24811 21063
rect 1961 20961 1995 20995
rect 4077 20961 4111 20995
rect 5345 20961 5379 20995
rect 7297 20961 7331 20995
rect 10609 20961 10643 20995
rect 13737 20961 13771 20995
rect 15669 20961 15703 20995
rect 17397 20961 17431 20995
rect 19625 20961 19659 20995
rect 21169 20961 21203 20995
rect 24317 20961 24351 20995
rect 25237 20961 25271 20995
rect 2237 20893 2271 20927
rect 5089 20893 5123 20927
rect 8401 20893 8435 20927
rect 13553 20893 13587 20927
rect 15945 20893 15979 20927
rect 17141 20893 17175 20927
rect 20913 20893 20947 20927
rect 24133 20893 24167 20927
rect 1685 20825 1719 20859
rect 4629 20825 4663 20859
rect 7941 20825 7975 20859
rect 13185 20825 13219 20859
rect 15393 20825 15427 20859
rect 23765 20825 23799 20859
rect 3709 20757 3743 20791
rect 4905 20757 4939 20791
rect 10333 20757 10367 20791
rect 12633 20757 12667 20791
rect 13001 20757 13035 20791
rect 15025 20757 15059 20791
rect 19073 20757 19107 20791
rect 23489 20757 23523 20791
rect 25145 20757 25179 20791
rect 3065 20553 3099 20587
rect 3617 20553 3651 20587
rect 5273 20553 5307 20587
rect 7297 20553 7331 20587
rect 9321 20553 9355 20587
rect 11897 20553 11931 20587
rect 13277 20553 13311 20587
rect 15117 20553 15151 20587
rect 18337 20553 18371 20587
rect 21189 20553 21223 20587
rect 22201 20553 22235 20587
rect 22661 20553 22695 20587
rect 25881 20553 25915 20587
rect 3985 20485 4019 20519
rect 16313 20485 16347 20519
rect 1685 20417 1719 20451
rect 5733 20417 5767 20451
rect 6285 20417 6319 20451
rect 23029 20417 23063 20451
rect 1952 20349 1986 20383
rect 6469 20349 6503 20383
rect 7389 20349 7423 20383
rect 7656 20349 7690 20383
rect 9781 20349 9815 20383
rect 9873 20349 9907 20383
rect 12173 20349 12207 20383
rect 13645 20349 13679 20383
rect 13737 20349 13771 20383
rect 13993 20349 14027 20383
rect 16589 20349 16623 20383
rect 17233 20349 17267 20383
rect 17877 20349 17911 20383
rect 19533 20349 19567 20383
rect 19809 20349 19843 20383
rect 22477 20349 22511 20383
rect 23489 20349 23523 20383
rect 23949 20349 23983 20383
rect 24205 20349 24239 20383
rect 4169 20281 4203 20315
rect 4721 20281 4755 20315
rect 5825 20281 5859 20315
rect 10140 20281 10174 20315
rect 12725 20281 12759 20315
rect 16865 20281 16899 20315
rect 18613 20281 18647 20315
rect 18889 20281 18923 20315
rect 19349 20281 19383 20315
rect 20076 20281 20110 20315
rect 4997 20213 5031 20247
rect 5733 20213 5767 20247
rect 6469 20213 6503 20247
rect 6561 20213 6595 20247
rect 8769 20213 8803 20247
rect 11253 20213 11287 20247
rect 15761 20213 15795 20247
rect 16129 20213 16163 20247
rect 16773 20213 16807 20247
rect 18797 20213 18831 20247
rect 19533 20213 19567 20247
rect 19717 20213 19751 20247
rect 21833 20213 21867 20247
rect 25329 20213 25363 20247
rect 1685 20009 1719 20043
rect 2053 20009 2087 20043
rect 3525 20009 3559 20043
rect 3801 20009 3835 20043
rect 6101 20009 6135 20043
rect 10885 20009 10919 20043
rect 13737 20009 13771 20043
rect 14749 20009 14783 20043
rect 15117 20009 15151 20043
rect 16681 20009 16715 20043
rect 17049 20009 17083 20043
rect 18521 20009 18555 20043
rect 19625 20009 19659 20043
rect 21097 20009 21131 20043
rect 22201 20009 22235 20043
rect 24685 20009 24719 20043
rect 25421 20009 25455 20043
rect 2973 19941 3007 19975
rect 6377 19941 6411 19975
rect 8401 19941 8435 19975
rect 8493 19941 8527 19975
rect 10701 19941 10735 19975
rect 12624 19941 12658 19975
rect 16129 19941 16163 19975
rect 16221 19941 16255 19975
rect 17408 19941 17442 19975
rect 20453 19941 20487 19975
rect 21465 19941 21499 19975
rect 24317 19941 24351 19975
rect 25237 19941 25271 19975
rect 4077 19873 4111 19907
rect 4344 19873 4378 19907
rect 6561 19873 6595 19907
rect 9965 19873 9999 19907
rect 12357 19873 12391 19907
rect 20913 19873 20947 19907
rect 22385 19873 22419 19907
rect 22652 19873 22686 19907
rect 2973 19805 3007 19839
rect 3065 19805 3099 19839
rect 6745 19805 6779 19839
rect 8401 19805 8435 19839
rect 10977 19805 11011 19839
rect 16129 19805 16163 19839
rect 17141 19805 17175 19839
rect 25513 19805 25547 19839
rect 2513 19737 2547 19771
rect 7941 19737 7975 19771
rect 10425 19737 10459 19771
rect 5457 19669 5491 19703
rect 7573 19669 7607 19703
rect 9137 19669 9171 19703
rect 11345 19669 11379 19703
rect 12173 19669 12207 19703
rect 15669 19669 15703 19703
rect 19073 19669 19107 19703
rect 20177 19669 20211 19703
rect 23765 19669 23799 19703
rect 24961 19669 24995 19703
rect 1961 19465 1995 19499
rect 6193 19465 6227 19499
rect 8861 19465 8895 19499
rect 10241 19465 10275 19499
rect 10517 19465 10551 19499
rect 12173 19465 12207 19499
rect 13921 19465 13955 19499
rect 19993 19465 20027 19499
rect 22385 19465 22419 19499
rect 23029 19465 23063 19499
rect 24317 19465 24351 19499
rect 25973 19465 26007 19499
rect 4169 19397 4203 19431
rect 25237 19397 25271 19431
rect 2145 19329 2179 19363
rect 6653 19329 6687 19363
rect 8125 19329 8159 19363
rect 11069 19329 11103 19363
rect 12523 19329 12557 19363
rect 19165 19329 19199 19363
rect 20085 19329 20119 19363
rect 25605 19329 25639 19363
rect 2412 19261 2446 19295
rect 7555 19261 7589 19295
rect 9137 19261 9171 19295
rect 9413 19261 9447 19295
rect 9965 19261 9999 19295
rect 10793 19261 10827 19295
rect 11805 19261 11839 19295
rect 13093 19261 13127 19295
rect 14381 19261 14415 19295
rect 14637 19261 14671 19295
rect 16865 19261 16899 19295
rect 17877 19261 17911 19295
rect 19625 19261 19659 19295
rect 20341 19261 20375 19295
rect 24869 19261 24903 19295
rect 1685 19193 1719 19227
rect 4997 19193 5031 19227
rect 5181 19193 5215 19227
rect 5273 19193 5307 19227
rect 5641 19193 5675 19227
rect 7389 19193 7423 19227
rect 7849 19193 7883 19227
rect 8033 19193 8067 19227
rect 12817 19193 12851 19227
rect 14289 19193 14323 19227
rect 17325 19193 17359 19227
rect 18337 19193 18371 19227
rect 18889 19193 18923 19227
rect 19073 19193 19107 19227
rect 23489 19193 23523 19227
rect 24593 19193 24627 19227
rect 3525 19125 3559 19159
rect 4445 19125 4479 19159
rect 4703 19125 4737 19159
rect 8493 19125 8527 19159
rect 10977 19125 11011 19159
rect 11437 19125 11471 19159
rect 13001 19125 13035 19159
rect 13553 19125 13587 19159
rect 15761 19125 15795 19159
rect 16313 19125 16347 19159
rect 16773 19125 16807 19159
rect 18603 19125 18637 19159
rect 21465 19125 21499 19159
rect 22569 19125 22603 19159
rect 24041 19125 24075 19159
rect 24777 19125 24811 19159
rect 3341 18921 3375 18955
rect 3709 18921 3743 18955
rect 4353 18921 4387 18955
rect 7665 18921 7699 18955
rect 8309 18921 8343 18955
rect 9505 18921 9539 18955
rect 10149 18921 10183 18955
rect 10885 18921 10919 18955
rect 11345 18921 11379 18955
rect 12909 18921 12943 18955
rect 13277 18921 13311 18955
rect 14565 18921 14599 18955
rect 15577 18921 15611 18955
rect 17141 18921 17175 18955
rect 18613 18921 18647 18955
rect 21097 18921 21131 18955
rect 21465 18921 21499 18955
rect 2881 18853 2915 18887
rect 2973 18853 3007 18887
rect 5273 18853 5307 18887
rect 11713 18853 11747 18887
rect 12449 18853 12483 18887
rect 14013 18853 14047 18887
rect 16221 18853 16255 18887
rect 17500 18853 17534 18887
rect 22652 18853 22686 18887
rect 25421 18853 25455 18887
rect 5365 18785 5399 18819
rect 6552 18785 6586 18819
rect 10701 18785 10735 18819
rect 14105 18785 14139 18819
rect 16037 18785 16071 18819
rect 21281 18785 21315 18819
rect 22385 18785 22419 18819
rect 25237 18785 25271 18819
rect 2789 18717 2823 18751
rect 5273 18717 5307 18751
rect 6285 18717 6319 18751
rect 10977 18717 11011 18751
rect 12357 18717 12391 18751
rect 12541 18717 12575 18751
rect 14013 18717 14047 18751
rect 16313 18717 16347 18751
rect 17233 18717 17267 18751
rect 19809 18717 19843 18751
rect 25513 18717 25547 18751
rect 2421 18649 2455 18683
rect 4813 18649 4847 18683
rect 10425 18649 10459 18683
rect 15761 18649 15795 18683
rect 24409 18649 24443 18683
rect 24961 18649 24995 18683
rect 1593 18581 1627 18615
rect 1961 18581 1995 18615
rect 5733 18581 5767 18615
rect 6101 18581 6135 18615
rect 8677 18581 8711 18615
rect 9045 18581 9079 18615
rect 11989 18581 12023 18615
rect 13553 18581 13587 18615
rect 14841 18581 14875 18615
rect 16773 18581 16807 18615
rect 19533 18581 19567 18615
rect 22109 18581 22143 18615
rect 23765 18581 23799 18615
rect 2973 18377 3007 18411
rect 7021 18377 7055 18411
rect 10241 18377 10275 18411
rect 11161 18377 11195 18411
rect 11621 18377 11655 18411
rect 12817 18377 12851 18411
rect 13185 18377 13219 18411
rect 14381 18377 14415 18411
rect 14933 18377 14967 18411
rect 16129 18377 16163 18411
rect 16221 18377 16255 18411
rect 16497 18377 16531 18411
rect 17877 18377 17911 18411
rect 19441 18377 19475 18411
rect 20913 18377 20947 18411
rect 21465 18377 21499 18411
rect 22109 18377 22143 18411
rect 25053 18377 25087 18411
rect 25513 18377 25547 18411
rect 9965 18309 9999 18343
rect 13369 18309 13403 18343
rect 10701 18241 10735 18275
rect 13921 18241 13955 18275
rect 15393 18241 15427 18275
rect 1593 18173 1627 18207
rect 1860 18173 1894 18207
rect 4169 18173 4203 18207
rect 4261 18173 4295 18207
rect 7665 18173 7699 18207
rect 9689 18173 9723 18207
rect 13645 18173 13679 18207
rect 14749 18173 14783 18207
rect 15485 18173 15519 18207
rect 18245 18309 18279 18343
rect 23029 18309 23063 18343
rect 24133 18309 24167 18343
rect 16957 18241 16991 18275
rect 19533 18241 19567 18275
rect 21925 18241 21959 18275
rect 22569 18241 22603 18275
rect 23489 18241 23523 18275
rect 23857 18241 23891 18275
rect 17049 18173 17083 18207
rect 4506 18105 4540 18139
rect 7910 18105 7944 18139
rect 10701 18105 10735 18139
rect 10793 18105 10827 18139
rect 13829 18105 13863 18139
rect 15393 18105 15427 18139
rect 16129 18105 16163 18139
rect 16957 18105 16991 18139
rect 19778 18105 19812 18139
rect 22569 18105 22603 18139
rect 22661 18105 22695 18139
rect 24409 18105 24443 18139
rect 24685 18105 24719 18139
rect 3617 18037 3651 18071
rect 5641 18037 5675 18071
rect 6285 18037 6319 18071
rect 7481 18037 7515 18071
rect 9045 18037 9079 18071
rect 11989 18037 12023 18071
rect 15945 18037 15979 18071
rect 17417 18037 17451 18071
rect 18613 18037 18647 18071
rect 24593 18037 24627 18071
rect 25789 18037 25823 18071
rect 2789 17833 2823 17867
rect 3433 17833 3467 17867
rect 3893 17833 3927 17867
rect 4353 17833 4387 17867
rect 4445 17833 4479 17867
rect 5273 17833 5307 17867
rect 6837 17833 6871 17867
rect 8585 17833 8619 17867
rect 9321 17833 9355 17867
rect 10149 17833 10183 17867
rect 13369 17833 13403 17867
rect 14197 17833 14231 17867
rect 16129 17833 16163 17867
rect 16497 17833 16531 17867
rect 21281 17833 21315 17867
rect 22109 17833 22143 17867
rect 2237 17765 2271 17799
rect 4905 17765 4939 17799
rect 7757 17765 7791 17799
rect 15577 17765 15611 17799
rect 19809 17765 19843 17799
rect 19901 17765 19935 17799
rect 24133 17765 24167 17799
rect 25237 17765 25271 17799
rect 5713 17697 5747 17731
rect 11060 17697 11094 17731
rect 14289 17697 14323 17731
rect 15301 17697 15335 17731
rect 16948 17697 16982 17731
rect 22457 17697 22491 17731
rect 2237 17629 2271 17663
rect 2329 17629 2363 17663
rect 3065 17629 3099 17663
rect 5457 17629 5491 17663
rect 8493 17629 8527 17663
rect 8677 17629 8711 17663
rect 9689 17629 9723 17663
rect 10793 17629 10827 17663
rect 14197 17629 14231 17663
rect 16681 17629 16715 17663
rect 19809 17629 19843 17663
rect 22201 17629 22235 17663
rect 25145 17629 25179 17663
rect 25329 17629 25363 17663
rect 1777 17561 1811 17595
rect 8125 17561 8159 17595
rect 13737 17561 13771 17595
rect 24501 17561 24535 17595
rect 24777 17561 24811 17595
rect 10609 17493 10643 17527
rect 12173 17493 12207 17527
rect 12725 17493 12759 17527
rect 14841 17493 14875 17527
rect 18061 17493 18095 17527
rect 19349 17493 19383 17527
rect 23581 17493 23615 17527
rect 4997 17289 5031 17323
rect 8769 17289 8803 17323
rect 10701 17289 10735 17323
rect 11621 17289 11655 17323
rect 16497 17289 16531 17323
rect 17417 17289 17451 17323
rect 21465 17289 21499 17323
rect 23029 17289 23063 17323
rect 4445 17221 4479 17255
rect 19993 17221 20027 17255
rect 22109 17221 22143 17255
rect 23765 17221 23799 17255
rect 22569 17153 22603 17187
rect 25237 17153 25271 17187
rect 2421 17085 2455 17119
rect 2688 17085 2722 17119
rect 6837 17085 6871 17119
rect 7093 17085 7127 17119
rect 9321 17085 9355 17119
rect 9577 17085 9611 17119
rect 12633 17085 12667 17119
rect 15117 17085 15151 17119
rect 18061 17085 18095 17119
rect 18317 17085 18351 17119
rect 1777 17017 1811 17051
rect 5273 17017 5307 17051
rect 5549 17017 5583 17051
rect 6009 17017 6043 17051
rect 6653 17017 6687 17051
rect 12900 17017 12934 17051
rect 15362 17017 15396 17051
rect 21097 17017 21131 17051
rect 22569 17017 22603 17051
rect 22661 17017 22695 17051
rect 24041 17017 24075 17051
rect 24225 17017 24259 17051
rect 24317 17017 24351 17051
rect 24777 17017 24811 17051
rect 2237 16949 2271 16983
rect 3801 16949 3835 16983
rect 4721 16949 4755 16983
rect 5457 16949 5491 16983
rect 8217 16949 8251 16983
rect 9137 16949 9171 16983
rect 11253 16949 11287 16983
rect 12173 16949 12207 16983
rect 14013 16949 14047 16983
rect 14565 16949 14599 16983
rect 15025 16949 15059 16983
rect 17049 16949 17083 16983
rect 17785 16949 17819 16983
rect 19441 16949 19475 16983
rect 21833 16949 21867 16983
rect 23397 16949 23431 16983
rect 25053 16949 25087 16983
rect 25697 16949 25731 16983
rect 1685 16745 1719 16779
rect 3525 16745 3559 16779
rect 5457 16745 5491 16779
rect 6009 16745 6043 16779
rect 6929 16745 6963 16779
rect 8585 16745 8619 16779
rect 9137 16745 9171 16779
rect 11989 16745 12023 16779
rect 12623 16745 12657 16779
rect 14657 16745 14691 16779
rect 18889 16745 18923 16779
rect 19625 16745 19659 16779
rect 21649 16745 21683 16779
rect 23121 16745 23155 16779
rect 24685 16745 24719 16779
rect 2329 16677 2363 16711
rect 2421 16677 2455 16711
rect 4322 16677 4356 16711
rect 7941 16677 7975 16711
rect 10241 16677 10275 16711
rect 10701 16677 10735 16711
rect 12265 16677 12299 16711
rect 13093 16677 13127 16711
rect 13921 16677 13955 16711
rect 15025 16677 15059 16711
rect 15568 16677 15602 16711
rect 18153 16677 18187 16711
rect 18337 16677 18371 16711
rect 19349 16677 19383 16711
rect 22293 16677 22327 16711
rect 22845 16677 22879 16711
rect 23550 16677 23584 16711
rect 1851 16609 1885 16643
rect 2145 16609 2179 16643
rect 2881 16609 2915 16643
rect 3249 16609 3283 16643
rect 4077 16609 4111 16643
rect 8401 16609 8435 16643
rect 8677 16609 8711 16643
rect 10057 16609 10091 16643
rect 14381 16609 14415 16643
rect 17233 16609 17267 16643
rect 18429 16609 18463 16643
rect 22385 16609 22419 16643
rect 25237 16609 25271 16643
rect 10333 16541 10367 16575
rect 13001 16541 13035 16575
rect 13185 16541 13219 16575
rect 13645 16541 13679 16575
rect 15301 16541 15335 16575
rect 22293 16541 22327 16575
rect 23305 16541 23339 16575
rect 9781 16473 9815 16507
rect 6469 16405 6503 16439
rect 7297 16405 7331 16439
rect 8125 16405 8159 16439
rect 11161 16405 11195 16439
rect 16681 16405 16715 16439
rect 17877 16405 17911 16439
rect 21833 16405 21867 16439
rect 2513 16201 2547 16235
rect 3433 16201 3467 16235
rect 4445 16201 4479 16235
rect 8953 16201 8987 16235
rect 9229 16201 9263 16235
rect 10149 16201 10183 16235
rect 12265 16201 12299 16235
rect 14289 16201 14323 16235
rect 14657 16201 14691 16235
rect 14933 16201 14967 16235
rect 16497 16201 16531 16235
rect 17509 16201 17543 16235
rect 17877 16201 17911 16235
rect 18337 16201 18371 16235
rect 23305 16201 23339 16235
rect 23857 16201 23891 16235
rect 2329 16133 2363 16167
rect 5273 16133 5307 16167
rect 6653 16133 6687 16167
rect 7389 16133 7423 16167
rect 10885 16133 10919 16167
rect 13369 16133 13403 16167
rect 18889 16133 18923 16167
rect 2973 16065 3007 16099
rect 3065 16065 3099 16099
rect 5733 16065 5767 16099
rect 7205 16065 7239 16099
rect 7849 16065 7883 16099
rect 9597 16065 9631 16099
rect 9781 16065 9815 16099
rect 10701 16065 10735 16099
rect 11437 16065 11471 16099
rect 15301 16065 15335 16099
rect 16313 16065 16347 16099
rect 16957 16065 16991 16099
rect 24409 16065 24443 16099
rect 24777 16065 24811 16099
rect 1961 15997 1995 16031
rect 5089 15997 5123 16031
rect 5825 15997 5859 16031
rect 13185 15997 13219 16031
rect 13921 15997 13955 16031
rect 19165 15997 19199 16031
rect 20821 15997 20855 16031
rect 24133 15997 24167 16031
rect 25329 15997 25363 16031
rect 25881 15997 25915 16031
rect 7941 15929 7975 15963
rect 9689 15929 9723 15963
rect 11161 15929 11195 15963
rect 12817 15929 12851 15963
rect 13645 15929 13679 15963
rect 13829 15929 13863 15963
rect 15485 15929 15519 15963
rect 17049 15929 17083 15963
rect 19441 15929 19475 15963
rect 19809 15929 19843 15963
rect 20361 15929 20395 15963
rect 21088 15929 21122 15963
rect 22937 15929 22971 15963
rect 1409 15861 1443 15895
rect 2973 15861 3007 15895
rect 4169 15861 4203 15895
rect 5733 15861 5767 15895
rect 6285 15861 6319 15895
rect 7849 15861 7883 15895
rect 8401 15861 8435 15895
rect 11345 15861 11379 15895
rect 11897 15861 11931 15895
rect 15393 15861 15427 15895
rect 15853 15861 15887 15895
rect 16957 15861 16991 15895
rect 18613 15861 18647 15895
rect 19349 15861 19383 15895
rect 20729 15861 20763 15895
rect 22201 15861 22235 15895
rect 24317 15861 24351 15895
rect 25513 15861 25547 15895
rect 2881 15657 2915 15691
rect 6653 15657 6687 15691
rect 7297 15657 7331 15691
rect 8309 15657 8343 15691
rect 8769 15657 8803 15691
rect 9229 15657 9263 15691
rect 11069 15657 11103 15691
rect 11989 15657 12023 15691
rect 13829 15657 13863 15691
rect 14565 15657 14599 15691
rect 15761 15657 15795 15691
rect 17325 15657 17359 15691
rect 19533 15657 19567 15691
rect 21465 15657 21499 15691
rect 22017 15657 22051 15691
rect 22385 15657 22419 15691
rect 23765 15657 23799 15691
rect 4721 15589 4755 15623
rect 10241 15589 10275 15623
rect 14841 15589 14875 15623
rect 15669 15589 15703 15623
rect 18889 15589 18923 15623
rect 19073 15589 19107 15623
rect 22845 15589 22879 15623
rect 23029 15589 23063 15623
rect 24409 15589 24443 15623
rect 24593 15589 24627 15623
rect 1501 15521 1535 15555
rect 1768 15521 1802 15555
rect 4077 15521 4111 15555
rect 5273 15521 5307 15555
rect 5540 15521 5574 15555
rect 8401 15521 8435 15555
rect 10057 15521 10091 15555
rect 12357 15521 12391 15555
rect 12716 15521 12750 15555
rect 16405 15521 16439 15555
rect 17141 15521 17175 15555
rect 21281 15521 21315 15555
rect 23121 15521 23155 15555
rect 24685 15521 24719 15555
rect 25053 15521 25087 15555
rect 8217 15453 8251 15487
rect 10333 15453 10367 15487
rect 12449 15453 12483 15487
rect 17417 15453 17451 15487
rect 18061 15453 18095 15487
rect 19165 15453 19199 15487
rect 21557 15453 21591 15487
rect 3893 15385 3927 15419
rect 9781 15385 9815 15419
rect 16865 15385 16899 15419
rect 20269 15385 20303 15419
rect 21005 15385 21039 15419
rect 3433 15317 3467 15351
rect 4261 15317 4295 15351
rect 5089 15317 5123 15351
rect 7849 15317 7883 15351
rect 10701 15317 10735 15351
rect 18613 15317 18647 15351
rect 20637 15317 20671 15351
rect 22569 15317 22603 15351
rect 24133 15317 24167 15351
rect 1501 15113 1535 15147
rect 2881 15113 2915 15147
rect 3617 15113 3651 15147
rect 4169 15113 4203 15147
rect 5641 15113 5675 15147
rect 6193 15113 6227 15147
rect 6929 15113 6963 15147
rect 7941 15113 7975 15147
rect 12173 15113 12207 15147
rect 13461 15113 13495 15147
rect 16497 15113 16531 15147
rect 16773 15113 16807 15147
rect 17417 15113 17451 15147
rect 19993 15113 20027 15147
rect 20453 15113 20487 15147
rect 21557 15113 21591 15147
rect 21925 15113 21959 15147
rect 22661 15113 22695 15147
rect 23489 15113 23523 15147
rect 24685 15113 24719 15147
rect 11805 15045 11839 15079
rect 12541 15045 12575 15079
rect 15117 15045 15151 15079
rect 20637 15045 20671 15079
rect 23765 15045 23799 15079
rect 1961 14977 1995 15011
rect 2053 14977 2087 15011
rect 12909 14977 12943 15011
rect 13093 14977 13127 15011
rect 13921 14977 13955 15011
rect 15577 14977 15611 15011
rect 16037 14977 16071 15011
rect 21005 14977 21039 15011
rect 22109 14977 22143 15011
rect 2973 14909 3007 14943
rect 4261 14909 4295 14943
rect 7205 14909 7239 14943
rect 9045 14909 9079 14943
rect 9873 14909 9907 14943
rect 14013 14909 14047 14943
rect 14933 14909 14967 14943
rect 15669 14909 15703 14943
rect 18061 14909 18095 14943
rect 18317 14909 18351 14943
rect 24041 14909 24075 14943
rect 25237 14909 25271 14943
rect 25789 14909 25823 14943
rect 1961 14841 1995 14875
rect 4506 14841 4540 14875
rect 6561 14841 6595 14875
rect 7389 14841 7423 14875
rect 7481 14841 7515 14875
rect 8309 14841 8343 14875
rect 10118 14841 10152 14875
rect 13001 14841 13035 14875
rect 15577 14841 15611 14875
rect 17785 14841 17819 14875
rect 21097 14841 21131 14875
rect 21189 14841 21223 14875
rect 24225 14841 24259 14875
rect 24317 14841 24351 14875
rect 25053 14841 25087 14875
rect 2421 14773 2455 14807
rect 3157 14773 3191 14807
rect 8493 14773 8527 14807
rect 9413 14773 9447 14807
rect 9781 14773 9815 14807
rect 11253 14773 11287 14807
rect 14473 14773 14507 14807
rect 16957 14773 16991 14807
rect 19441 14773 19475 14807
rect 22937 14773 22971 14807
rect 25421 14773 25455 14807
rect 2789 14569 2823 14603
rect 3065 14569 3099 14603
rect 5457 14569 5491 14603
rect 6009 14569 6043 14603
rect 6469 14569 6503 14603
rect 6837 14569 6871 14603
rect 8401 14569 8435 14603
rect 9413 14569 9447 14603
rect 10425 14569 10459 14603
rect 12817 14569 12851 14603
rect 15853 14569 15887 14603
rect 18061 14569 18095 14603
rect 18889 14569 18923 14603
rect 19809 14569 19843 14603
rect 20637 14569 20671 14603
rect 22845 14569 22879 14603
rect 25329 14569 25363 14603
rect 2053 14501 2087 14535
rect 2237 14501 2271 14535
rect 2329 14501 2363 14535
rect 7757 14501 7791 14535
rect 11253 14501 11287 14535
rect 17417 14501 17451 14535
rect 18613 14501 18647 14535
rect 23642 14501 23676 14535
rect 4333 14433 4367 14467
rect 7849 14433 7883 14467
rect 10241 14433 10275 14467
rect 11693 14433 11727 14467
rect 13461 14433 13495 14467
rect 15669 14433 15703 14467
rect 17509 14433 17543 14467
rect 19625 14433 19659 14467
rect 21169 14433 21203 14467
rect 4077 14365 4111 14399
rect 7757 14365 7791 14399
rect 10517 14365 10551 14399
rect 11437 14365 11471 14399
rect 15117 14365 15151 14399
rect 15945 14365 15979 14399
rect 16773 14365 16807 14399
rect 17417 14365 17451 14399
rect 19901 14365 19935 14399
rect 20913 14365 20947 14399
rect 23397 14365 23431 14399
rect 1777 14297 1811 14331
rect 9965 14297 9999 14331
rect 15393 14297 15427 14331
rect 3525 14229 3559 14263
rect 3893 14229 3927 14263
rect 7297 14229 7331 14263
rect 8861 14229 8895 14263
rect 10885 14229 10919 14263
rect 16957 14229 16991 14263
rect 19349 14229 19383 14263
rect 22293 14229 22327 14263
rect 23305 14229 23339 14263
rect 24777 14229 24811 14263
rect 1501 14025 1535 14059
rect 2789 14025 2823 14059
rect 3341 14025 3375 14059
rect 4445 14025 4479 14059
rect 6653 14025 6687 14059
rect 6929 14025 6963 14059
rect 9965 14025 9999 14059
rect 12173 14025 12207 14059
rect 13185 14025 13219 14059
rect 13277 14025 13311 14059
rect 13553 14025 13587 14059
rect 16405 14025 16439 14059
rect 16957 14025 16991 14059
rect 17325 14025 17359 14059
rect 18153 14025 18187 14059
rect 19165 14025 19199 14059
rect 21005 14025 21039 14059
rect 25053 14025 25087 14059
rect 2513 13957 2547 13991
rect 3525 13957 3559 13991
rect 5181 13957 5215 13991
rect 8493 13957 8527 13991
rect 10241 13957 10275 13991
rect 10885 13957 10919 13991
rect 13001 13957 13035 13991
rect 14841 13957 14875 13991
rect 17785 13957 17819 13991
rect 19533 13957 19567 13991
rect 2053 13889 2087 13923
rect 3893 13889 3927 13923
rect 4997 13889 5031 13923
rect 5641 13889 5675 13923
rect 7389 13889 7423 13923
rect 9413 13889 9447 13923
rect 11437 13889 11471 13923
rect 13185 13889 13219 13923
rect 13921 13889 13955 13923
rect 14105 13889 14139 13923
rect 14565 13889 14599 13923
rect 18705 13889 18739 13923
rect 1777 13821 1811 13855
rect 5733 13821 5767 13855
rect 7481 13821 7515 13855
rect 7941 13821 7975 13855
rect 8309 13821 8343 13855
rect 8769 13821 8803 13855
rect 9045 13821 9079 13855
rect 10701 13821 10735 13855
rect 15025 13821 15059 13855
rect 15292 13821 15326 13855
rect 18429 13821 18463 13855
rect 19625 13821 19659 13855
rect 21557 13821 21591 13855
rect 23029 13821 23063 13855
rect 23397 13821 23431 13855
rect 23673 13821 23707 13855
rect 23940 13821 23974 13855
rect 4077 13753 4111 13787
rect 6193 13753 6227 13787
rect 8953 13753 8987 13787
rect 11161 13753 11195 13787
rect 14013 13753 14047 13787
rect 18613 13753 18647 13787
rect 19892 13753 19926 13787
rect 1961 13685 1995 13719
rect 3985 13685 4019 13719
rect 5641 13685 5675 13719
rect 7389 13685 7423 13719
rect 11345 13685 11379 13719
rect 11805 13685 11839 13719
rect 1685 13481 1719 13515
rect 3525 13481 3559 13515
rect 5089 13481 5123 13515
rect 5457 13481 5491 13515
rect 6929 13481 6963 13515
rect 7481 13481 7515 13515
rect 7849 13481 7883 13515
rect 8585 13481 8619 13515
rect 10517 13481 10551 13515
rect 12081 13481 12115 13515
rect 18245 13481 18279 13515
rect 19165 13481 19199 13515
rect 20269 13481 20303 13515
rect 21097 13481 21131 13515
rect 23397 13481 23431 13515
rect 2789 13413 2823 13447
rect 2973 13413 3007 13447
rect 3801 13413 3835 13447
rect 5816 13413 5850 13447
rect 8401 13413 8435 13447
rect 10946 13413 10980 13447
rect 13737 13413 13771 13447
rect 15577 13413 15611 13447
rect 16466 13413 16500 13447
rect 18797 13413 18831 13447
rect 19809 13413 19843 13447
rect 22569 13413 22603 13447
rect 22661 13413 22695 13447
rect 24133 13413 24167 13447
rect 24225 13413 24259 13447
rect 4077 13345 4111 13379
rect 13093 13345 13127 13379
rect 19901 13345 19935 13379
rect 22385 13345 22419 13379
rect 25145 13345 25179 13379
rect 3065 13277 3099 13311
rect 5549 13277 5583 13311
rect 8677 13277 8711 13311
rect 9689 13277 9723 13311
rect 10701 13277 10735 13311
rect 13737 13277 13771 13311
rect 13829 13277 13863 13311
rect 15025 13277 15059 13311
rect 16221 13277 16255 13311
rect 19717 13277 19751 13311
rect 24041 13277 24075 13311
rect 2513 13209 2547 13243
rect 4721 13209 4755 13243
rect 8125 13209 8159 13243
rect 13277 13209 13311 13243
rect 22109 13209 22143 13243
rect 23121 13209 23155 13243
rect 23673 13209 23707 13243
rect 1961 13141 1995 13175
rect 4261 13141 4295 13175
rect 9229 13141 9263 13175
rect 10149 13141 10183 13175
rect 17601 13141 17635 13175
rect 19349 13141 19383 13175
rect 21465 13141 21499 13175
rect 1685 12937 1719 12971
rect 3525 12937 3559 12971
rect 4721 12937 4755 12971
rect 6009 12937 6043 12971
rect 13093 12937 13127 12971
rect 13369 12937 13403 12971
rect 14381 12937 14415 12971
rect 15393 12937 15427 12971
rect 17233 12937 17267 12971
rect 18981 12937 19015 12971
rect 19349 12937 19383 12971
rect 22109 12937 22143 12971
rect 22845 12937 22879 12971
rect 24685 12937 24719 12971
rect 25053 12937 25087 12971
rect 2053 12869 2087 12903
rect 7021 12869 7055 12903
rect 8033 12869 8067 12903
rect 16037 12869 16071 12903
rect 16313 12869 16347 12903
rect 19533 12869 19567 12903
rect 21097 12869 21131 12903
rect 22477 12869 22511 12903
rect 23765 12869 23799 12903
rect 4169 12801 4203 12835
rect 4537 12801 4571 12835
rect 5181 12801 5215 12835
rect 5273 12801 5307 12835
rect 7481 12801 7515 12835
rect 8493 12801 8527 12835
rect 13737 12801 13771 12835
rect 13921 12801 13955 12835
rect 14657 12801 14691 12835
rect 16773 12801 16807 12835
rect 21649 12801 21683 12835
rect 2145 12733 2179 12767
rect 9413 12733 9447 12767
rect 9597 12733 9631 12767
rect 15761 12733 15795 12767
rect 16865 12733 16899 12767
rect 19809 12733 19843 12767
rect 24041 12733 24075 12767
rect 25237 12733 25271 12767
rect 25789 12733 25823 12767
rect 2412 12665 2446 12699
rect 5181 12665 5215 12699
rect 6653 12665 6687 12699
rect 7573 12665 7607 12699
rect 9137 12665 9171 12699
rect 9864 12665 9898 12699
rect 12817 12665 12851 12699
rect 13829 12665 13863 12699
rect 16773 12665 16807 12699
rect 18613 12665 18647 12699
rect 19993 12665 20027 12699
rect 20085 12665 20119 12699
rect 20545 12665 20579 12699
rect 21373 12665 21407 12699
rect 21557 12665 21591 12699
rect 23489 12665 23523 12699
rect 24317 12665 24351 12699
rect 5733 12597 5767 12631
rect 7481 12597 7515 12631
rect 10977 12597 11011 12631
rect 11621 12597 11655 12631
rect 20913 12597 20947 12631
rect 24225 12597 24259 12631
rect 25421 12597 25455 12631
rect 2973 12393 3007 12427
rect 3433 12393 3467 12427
rect 8493 12393 8527 12427
rect 8769 12393 8803 12427
rect 11161 12393 11195 12427
rect 13829 12393 13863 12427
rect 16773 12393 16807 12427
rect 19993 12393 20027 12427
rect 22293 12393 22327 12427
rect 23305 12393 23339 12427
rect 3065 12325 3099 12359
rect 7941 12325 7975 12359
rect 10241 12325 10275 12359
rect 16221 12325 16255 12359
rect 17500 12325 17534 12359
rect 23673 12325 23707 12359
rect 24124 12325 24158 12359
rect 2237 12257 2271 12291
rect 4077 12257 4111 12291
rect 4344 12257 4378 12291
rect 7757 12257 7791 12291
rect 10057 12257 10091 12291
rect 12164 12257 12198 12291
rect 19349 12257 19383 12291
rect 21180 12257 21214 12291
rect 1409 12189 1443 12223
rect 2973 12189 3007 12223
rect 6009 12189 6043 12223
rect 8033 12189 8067 12223
rect 10333 12189 10367 12223
rect 11897 12189 11931 12223
rect 16129 12189 16163 12223
rect 16313 12189 16347 12223
rect 17233 12189 17267 12223
rect 20913 12189 20947 12223
rect 23857 12189 23891 12223
rect 6653 12121 6687 12155
rect 13277 12121 13311 12155
rect 2513 12053 2547 12087
rect 3893 12053 3927 12087
rect 5457 12053 5491 12087
rect 7021 12053 7055 12087
rect 7481 12053 7515 12087
rect 9137 12053 9171 12087
rect 9781 12053 9815 12087
rect 10701 12053 10735 12087
rect 11713 12053 11747 12087
rect 15761 12053 15795 12087
rect 18613 12053 18647 12087
rect 19717 12053 19751 12087
rect 25237 12053 25271 12087
rect 2789 11849 2823 11883
rect 3341 11849 3375 11883
rect 5917 11849 5951 11883
rect 6285 11849 6319 11883
rect 7389 11849 7423 11883
rect 7665 11849 7699 11883
rect 11805 11849 11839 11883
rect 15669 11849 15703 11883
rect 16221 11849 16255 11883
rect 17601 11849 17635 11883
rect 18889 11849 18923 11883
rect 20637 11849 20671 11883
rect 23121 11849 23155 11883
rect 25513 11849 25547 11883
rect 1777 11781 1811 11815
rect 9229 11781 9263 11815
rect 10885 11781 10919 11815
rect 12817 11781 12851 11815
rect 20821 11781 20855 11815
rect 23489 11781 23523 11815
rect 23949 11781 23983 11815
rect 3801 11713 3835 11747
rect 5457 11713 5491 11747
rect 8125 11713 8159 11747
rect 8585 11713 8619 11747
rect 11437 11713 11471 11747
rect 13185 11713 13219 11747
rect 18337 11713 18371 11747
rect 19441 11713 19475 11747
rect 19901 11713 19935 11747
rect 21189 11713 21223 11747
rect 24133 11713 24167 11747
rect 3157 11645 3191 11679
rect 3893 11645 3927 11679
rect 4353 11645 4387 11679
rect 5181 11645 5215 11679
rect 9505 11645 9539 11679
rect 14105 11645 14139 11679
rect 14289 11645 14323 11679
rect 24400 11645 24434 11679
rect 2053 11577 2087 11611
rect 2329 11577 2363 11611
rect 4887 11577 4921 11611
rect 7113 11577 7147 11611
rect 8217 11577 8251 11611
rect 9781 11577 9815 11611
rect 10149 11577 10183 11611
rect 11161 11577 11195 11611
rect 11345 11577 11379 11611
rect 12173 11577 12207 11611
rect 13369 11577 13403 11611
rect 13737 11577 13771 11611
rect 14534 11577 14568 11611
rect 19165 11577 19199 11611
rect 20269 11577 20303 11611
rect 21373 11577 21407 11611
rect 2237 11509 2271 11543
rect 3801 11509 3835 11543
rect 4721 11509 4755 11543
rect 5365 11509 5399 11543
rect 6653 11509 6687 11543
rect 8125 11509 8159 11543
rect 9045 11509 9079 11543
rect 9689 11509 9723 11543
rect 10609 11509 10643 11543
rect 13277 11509 13311 11543
rect 17233 11509 17267 11543
rect 18613 11509 18647 11543
rect 19349 11509 19383 11543
rect 21281 11509 21315 11543
rect 21833 11509 21867 11543
rect 2237 11305 2271 11339
rect 2881 11305 2915 11339
rect 3893 11305 3927 11339
rect 5457 11305 5491 11339
rect 6469 11305 6503 11339
rect 8309 11305 8343 11339
rect 8953 11305 8987 11339
rect 11161 11305 11195 11339
rect 11621 11305 11655 11339
rect 14381 11305 14415 11339
rect 15761 11305 15795 11339
rect 18797 11305 18831 11339
rect 21097 11305 21131 11339
rect 23213 11305 23247 11339
rect 23765 11305 23799 11339
rect 24225 11305 24259 11339
rect 4445 11237 4479 11271
rect 4629 11237 4663 11271
rect 4721 11237 4755 11271
rect 8125 11237 8159 11271
rect 10057 11237 10091 11271
rect 10241 11237 10275 11271
rect 11980 11237 12014 11271
rect 19717 11237 19751 11271
rect 24685 11237 24719 11271
rect 24869 11237 24903 11271
rect 24961 11237 24995 11271
rect 1409 11169 1443 11203
rect 2697 11169 2731 11203
rect 6285 11169 6319 11203
rect 7021 11169 7055 11203
rect 8401 11169 8435 11203
rect 9321 11169 9355 11203
rect 16129 11169 16163 11203
rect 16948 11169 16982 11203
rect 19809 11169 19843 11203
rect 22100 11169 22134 11203
rect 1685 11101 1719 11135
rect 3525 11101 3559 11135
rect 6561 11101 6595 11135
rect 7665 11101 7699 11135
rect 10333 11101 10367 11135
rect 11713 11101 11747 11135
rect 16681 11101 16715 11135
rect 19625 11101 19659 11135
rect 21833 11101 21867 11135
rect 2513 11033 2547 11067
rect 6009 11033 6043 11067
rect 7849 11033 7883 11067
rect 9781 11033 9815 11067
rect 10885 11033 10919 11067
rect 19257 11033 19291 11067
rect 24409 11033 24443 11067
rect 4169 10965 4203 10999
rect 5181 10965 5215 10999
rect 13093 10965 13127 10999
rect 18061 10965 18095 10999
rect 21465 10965 21499 10999
rect 3801 10761 3835 10795
rect 4537 10761 4571 10795
rect 6009 10761 6043 10795
rect 7021 10761 7055 10795
rect 8033 10761 8067 10795
rect 9321 10761 9355 10795
rect 10333 10761 10367 10795
rect 12081 10761 12115 10795
rect 12173 10761 12207 10795
rect 14381 10761 14415 10795
rect 16681 10761 16715 10795
rect 19625 10761 19659 10795
rect 20821 10761 20855 10795
rect 22385 10761 22419 10795
rect 23397 10761 23431 10795
rect 25053 10761 25087 10795
rect 2697 10693 2731 10727
rect 3525 10693 3559 10727
rect 4813 10693 4847 10727
rect 8309 10693 8343 10727
rect 10885 10693 10919 10727
rect 5365 10625 5399 10659
rect 7481 10625 7515 10659
rect 9137 10625 9171 10659
rect 9781 10625 9815 10659
rect 11345 10625 11379 10659
rect 1409 10557 1443 10591
rect 2513 10557 2547 10591
rect 3617 10557 3651 10591
rect 5089 10557 5123 10591
rect 11897 10557 11931 10591
rect 3157 10489 3191 10523
rect 6653 10489 6687 10523
rect 7481 10489 7515 10523
rect 7573 10489 7607 10523
rect 8769 10489 8803 10523
rect 9873 10489 9907 10523
rect 11345 10489 11379 10523
rect 11437 10489 11471 10523
rect 12541 10693 12575 10727
rect 18153 10693 18187 10727
rect 19901 10693 19935 10727
rect 21465 10693 21499 10727
rect 25605 10693 25639 10727
rect 13829 10625 13863 10659
rect 14565 10625 14599 10659
rect 21281 10625 21315 10659
rect 22017 10625 22051 10659
rect 23673 10625 23707 10659
rect 12817 10557 12851 10591
rect 17509 10557 17543 10591
rect 19349 10557 19383 10591
rect 23929 10557 23963 10591
rect 13093 10489 13127 10523
rect 14810 10489 14844 10523
rect 17141 10489 17175 10523
rect 18429 10489 18463 10523
rect 18705 10489 18739 10523
rect 20177 10489 20211 10523
rect 20453 10489 20487 10523
rect 21741 10489 21775 10523
rect 1593 10421 1627 10455
rect 2053 10421 2087 10455
rect 2329 10421 2363 10455
rect 4169 10421 4203 10455
rect 5273 10421 5307 10455
rect 9781 10421 9815 10455
rect 10701 10421 10735 10455
rect 12081 10421 12115 10455
rect 13001 10421 13035 10455
rect 13461 10421 13495 10455
rect 15945 10421 15979 10455
rect 17785 10421 17819 10455
rect 18613 10421 18647 10455
rect 20361 10421 20395 10455
rect 21925 10421 21959 10455
rect 22753 10421 22787 10455
rect 1961 10217 1995 10251
rect 2421 10217 2455 10251
rect 3341 10217 3375 10251
rect 3617 10217 3651 10251
rect 4353 10217 4387 10251
rect 6193 10217 6227 10251
rect 7021 10217 7055 10251
rect 7665 10217 7699 10251
rect 8861 10217 8895 10251
rect 9965 10217 9999 10251
rect 12449 10217 12483 10251
rect 13093 10217 13127 10251
rect 14657 10217 14691 10251
rect 15853 10217 15887 10251
rect 17417 10217 17451 10251
rect 18889 10217 18923 10251
rect 19533 10217 19567 10251
rect 23305 10217 23339 10251
rect 23949 10217 23983 10251
rect 24501 10217 24535 10251
rect 25145 10217 25179 10251
rect 5080 10149 5114 10183
rect 8309 10149 8343 10183
rect 8401 10149 8435 10183
rect 11529 10149 11563 10183
rect 14933 10149 14967 10183
rect 15669 10149 15703 10183
rect 15945 10149 15979 10183
rect 17754 10149 17788 10183
rect 23765 10149 23799 10183
rect 1409 10081 1443 10115
rect 2513 10081 2547 10115
rect 8125 10081 8159 10115
rect 9321 10081 9355 10115
rect 11345 10081 11379 10115
rect 12909 10081 12943 10115
rect 14105 10081 14139 10115
rect 21180 10081 21214 10115
rect 24041 10081 24075 10115
rect 24961 10081 24995 10115
rect 4813 10013 4847 10047
rect 11621 10013 11655 10047
rect 13185 10013 13219 10047
rect 17509 10013 17543 10047
rect 20913 10013 20947 10047
rect 2697 9945 2731 9979
rect 11989 9945 12023 9979
rect 23489 9945 23523 9979
rect 1593 9877 1627 9911
rect 4721 9877 4755 9911
rect 7849 9877 7883 9911
rect 10241 9877 10275 9911
rect 10793 9877 10827 9911
rect 11069 9877 11103 9911
rect 12633 9877 12667 9911
rect 15393 9877 15427 9911
rect 19901 9877 19935 9911
rect 22293 9877 22327 9911
rect 22937 9877 22971 9911
rect 24869 9877 24903 9911
rect 7665 9673 7699 9707
rect 11897 9673 11931 9707
rect 15945 9673 15979 9707
rect 17509 9673 17543 9707
rect 20729 9673 20763 9707
rect 20913 9673 20947 9707
rect 23489 9673 23523 9707
rect 24961 9673 24995 9707
rect 2697 9605 2731 9639
rect 3525 9605 3559 9639
rect 5641 9605 5675 9639
rect 10425 9605 10459 9639
rect 13829 9605 13863 9639
rect 15025 9605 15059 9639
rect 18153 9605 18187 9639
rect 19165 9605 19199 9639
rect 19533 9605 19567 9639
rect 20361 9605 20395 9639
rect 23029 9605 23063 9639
rect 23765 9605 23799 9639
rect 25421 9605 25455 9639
rect 2421 9537 2455 9571
rect 9873 9537 9907 9571
rect 11529 9537 11563 9571
rect 14473 9537 14507 9571
rect 15393 9537 15427 9571
rect 15577 9537 15611 9571
rect 16957 9537 16991 9571
rect 18705 9537 18739 9571
rect 19993 9537 20027 9571
rect 21465 9537 21499 9571
rect 22385 9537 22419 9571
rect 24317 9537 24351 9571
rect 1409 9469 1443 9503
rect 2519 9469 2553 9503
rect 4169 9469 4203 9503
rect 4261 9469 4295 9503
rect 4528 9469 4562 9503
rect 7849 9469 7883 9503
rect 8116 9469 8150 9503
rect 12173 9469 12207 9503
rect 12449 9469 12483 9503
rect 14841 9469 14875 9503
rect 16865 9469 16899 9503
rect 21189 9469 21223 9503
rect 22201 9469 22235 9503
rect 25237 9469 25271 9503
rect 25789 9469 25823 9503
rect 2053 9401 2087 9435
rect 7389 9401 7423 9435
rect 10701 9401 10735 9435
rect 10885 9401 10919 9435
rect 10977 9401 11011 9435
rect 12716 9401 12750 9435
rect 15485 9401 15519 9435
rect 18429 9401 18463 9435
rect 24041 9401 24075 9435
rect 24225 9401 24259 9435
rect 1593 9333 1627 9367
rect 3157 9333 3191 9367
rect 6285 9333 6319 9367
rect 6837 9333 6871 9367
rect 9229 9333 9263 9367
rect 10149 9333 10183 9367
rect 18613 9333 18647 9367
rect 21373 9333 21407 9367
rect 21833 9333 21867 9367
rect 1961 9129 1995 9163
rect 4353 9129 4387 9163
rect 5181 9129 5215 9163
rect 7665 9129 7699 9163
rect 8217 9129 8251 9163
rect 9505 9129 9539 9163
rect 10149 9129 10183 9163
rect 11989 9129 12023 9163
rect 13645 9129 13679 9163
rect 14197 9129 14231 9163
rect 15025 9129 15059 9163
rect 15577 9129 15611 9163
rect 17233 9129 17267 9163
rect 17601 9129 17635 9163
rect 18153 9129 18187 9163
rect 23121 9129 23155 9163
rect 24225 9129 24259 9163
rect 24961 9129 24995 9163
rect 4813 9061 4847 9095
rect 8677 9061 8711 9095
rect 10517 9061 10551 9095
rect 13461 9061 13495 9095
rect 18797 9061 18831 9095
rect 21557 9061 21591 9095
rect 23581 9061 23615 9095
rect 23765 9061 23799 9095
rect 1409 8993 1443 9027
rect 6541 8993 6575 9027
rect 10876 8993 10910 9027
rect 12541 8993 12575 9027
rect 21373 8993 21407 9027
rect 24777 8993 24811 9027
rect 6285 8925 6319 8959
rect 10609 8925 10643 8959
rect 13737 8925 13771 8959
rect 18705 8925 18739 8959
rect 18889 8925 18923 8959
rect 21649 8925 21683 8959
rect 23857 8925 23891 8959
rect 13185 8857 13219 8891
rect 18337 8857 18371 8891
rect 21097 8857 21131 8891
rect 23305 8857 23339 8891
rect 1593 8789 1627 8823
rect 13001 8789 13035 8823
rect 1593 8585 1627 8619
rect 2053 8585 2087 8619
rect 5641 8585 5675 8619
rect 5917 8585 5951 8619
rect 6929 8585 6963 8619
rect 9229 8585 9263 8619
rect 10793 8585 10827 8619
rect 11805 8585 11839 8619
rect 13553 8585 13587 8619
rect 17877 8585 17911 8619
rect 21373 8585 21407 8619
rect 21741 8585 21775 8619
rect 23213 8585 23247 8619
rect 24869 8585 24903 8619
rect 25145 8585 25179 8619
rect 11437 8517 11471 8551
rect 12541 8517 12575 8551
rect 14105 8517 14139 8551
rect 22937 8517 22971 8551
rect 7481 8449 7515 8483
rect 13093 8449 13127 8483
rect 14657 8449 14691 8483
rect 21097 8449 21131 8483
rect 1409 8381 1443 8415
rect 2329 8381 2363 8415
rect 6285 8381 6319 8415
rect 7205 8381 7239 8415
rect 9413 8381 9447 8415
rect 12265 8381 12299 8415
rect 12817 8381 12851 8415
rect 14381 8381 14415 8415
rect 17509 8381 17543 8415
rect 18245 8381 18279 8415
rect 23673 8381 23707 8415
rect 24409 8381 24443 8415
rect 24961 8381 24995 8415
rect 25513 8381 25547 8415
rect 9658 8313 9692 8347
rect 13001 8313 13035 8347
rect 13921 8313 13955 8347
rect 14565 8313 14599 8347
rect 18521 8313 18555 8347
rect 19073 8313 19107 8347
rect 23949 8313 23983 8347
rect 7389 8245 7423 8279
rect 1593 8041 1627 8075
rect 6469 8041 6503 8075
rect 7021 8041 7055 8075
rect 7389 8041 7423 8075
rect 8115 8041 8149 8075
rect 10241 8041 10275 8075
rect 10793 8041 10827 8075
rect 14013 8041 14047 8075
rect 14473 8041 14507 8075
rect 18337 8041 18371 8075
rect 23305 8041 23339 8075
rect 24777 8041 24811 8075
rect 6561 7973 6595 8007
rect 8585 7973 8619 8007
rect 9505 7973 9539 8007
rect 12449 7973 12483 8007
rect 13535 7973 13569 8007
rect 1409 7905 1443 7939
rect 8401 7905 8435 7939
rect 10057 7905 10091 7939
rect 12265 7905 12299 7939
rect 16957 7905 16991 7939
rect 23489 7905 23523 7939
rect 24593 7905 24627 7939
rect 6469 7837 6503 7871
rect 8677 7837 8711 7871
rect 10333 7837 10367 7871
rect 12541 7837 12575 7871
rect 13185 7837 13219 7871
rect 14013 7837 14047 7871
rect 14105 7837 14139 7871
rect 17233 7837 17267 7871
rect 6009 7769 6043 7803
rect 9781 7769 9815 7803
rect 11989 7701 12023 7735
rect 23673 7701 23707 7735
rect 2053 7497 2087 7531
rect 6009 7497 6043 7531
rect 7941 7497 7975 7531
rect 8309 7497 8343 7531
rect 8493 7497 8527 7531
rect 9781 7497 9815 7531
rect 11621 7497 11655 7531
rect 11989 7497 12023 7531
rect 12725 7497 12759 7531
rect 13093 7497 13127 7531
rect 13461 7497 13495 7531
rect 13921 7497 13955 7531
rect 14197 7497 14231 7531
rect 16957 7497 16991 7531
rect 23949 7497 23983 7531
rect 24409 7497 24443 7531
rect 24777 7497 24811 7531
rect 1593 7429 1627 7463
rect 5641 7429 5675 7463
rect 10701 7429 10735 7463
rect 6377 7361 6411 7395
rect 8953 7361 8987 7395
rect 10149 7361 10183 7395
rect 1409 7293 1443 7327
rect 7573 7293 7607 7327
rect 9045 7293 9079 7327
rect 9965 7293 9999 7327
rect 18061 7293 18095 7327
rect 18613 7293 18647 7327
rect 24593 7293 24627 7327
rect 25145 7293 25179 7327
rect 8953 7225 8987 7259
rect 18245 7157 18279 7191
rect 1593 6953 1627 6987
rect 8493 6953 8527 6987
rect 8769 6953 8803 6987
rect 9873 6953 9907 6987
rect 10241 6953 10275 6987
rect 11989 6953 12023 6987
rect 24777 6953 24811 6987
rect 4629 6817 4663 6851
rect 8125 6817 8159 6851
rect 24593 6817 24627 6851
rect 4813 6749 4847 6783
rect 4721 6409 4755 6443
rect 4997 6409 5031 6443
rect 9321 6409 9355 6443
rect 24777 6409 24811 6443
rect 24501 6341 24535 6375
rect 4077 6205 4111 6239
rect 8677 6205 8711 6239
rect 24593 6205 24627 6239
rect 25145 6205 25179 6239
rect 4261 6069 4295 6103
rect 8861 6069 8895 6103
rect 24777 5865 24811 5899
rect 20913 5729 20947 5763
rect 24593 5729 24627 5763
rect 21097 5661 21131 5695
rect 20913 5321 20947 5355
rect 24777 5321 24811 5355
rect 24501 5253 24535 5287
rect 24593 5117 24627 5151
rect 25145 5117 25179 5151
rect 21281 4777 21315 4811
rect 21097 4641 21131 4675
rect 21097 4233 21131 4267
rect 2421 4097 2455 4131
rect 1685 4029 1719 4063
rect 1961 3961 1995 3995
rect 1409 3553 1443 3587
rect 23581 3553 23615 3587
rect 24869 3553 24903 3587
rect 23857 3485 23891 3519
rect 1593 3417 1627 3451
rect 25053 3349 25087 3383
rect 1593 3145 1627 3179
rect 4537 3145 4571 3179
rect 23121 3145 23155 3179
rect 24869 3145 24903 3179
rect 3709 2941 3743 2975
rect 8125 2941 8159 2975
rect 8861 2941 8895 2975
rect 23489 2941 23523 2975
rect 23857 2941 23891 2975
rect 24133 2941 24167 2975
rect 25145 2941 25179 2975
rect 25697 2941 25731 2975
rect 3985 2873 4019 2907
rect 8401 2873 8435 2907
rect 25329 2805 25363 2839
rect 2053 2601 2087 2635
rect 8033 2601 8067 2635
rect 1409 2465 1443 2499
rect 7389 2465 7423 2499
rect 22845 2465 22879 2499
rect 24041 2465 24075 2499
rect 24777 2465 24811 2499
rect 25329 2465 25363 2499
rect 25881 2465 25915 2499
rect 23489 2397 23523 2431
rect 24225 2397 24259 2431
rect 1593 2261 1627 2295
rect 7573 2261 7607 2295
rect 23029 2261 23063 2295
rect 25513 2261 25547 2295
<< metal1 >>
rect 9766 26392 9772 26444
rect 9824 26432 9830 26444
rect 24762 26432 24768 26444
rect 9824 26404 24768 26432
rect 9824 26392 9830 26404
rect 24762 26392 24768 26404
rect 24820 26392 24826 26444
rect 8202 26324 8208 26376
rect 8260 26364 8266 26376
rect 23566 26364 23572 26376
rect 8260 26336 23572 26364
rect 8260 26324 8266 26336
rect 23566 26324 23572 26336
rect 23624 26324 23630 26376
rect 7374 26256 7380 26308
rect 7432 26296 7438 26308
rect 24302 26296 24308 26308
rect 7432 26268 24308 26296
rect 7432 26256 7438 26268
rect 24302 26256 24308 26268
rect 24360 26256 24366 26308
rect 4062 25780 4068 25832
rect 4120 25820 4126 25832
rect 13722 25820 13728 25832
rect 4120 25792 13728 25820
rect 4120 25780 4126 25792
rect 13722 25780 13728 25792
rect 13780 25780 13786 25832
rect 12894 25712 12900 25764
rect 12952 25752 12958 25764
rect 21726 25752 21732 25764
rect 12952 25724 21732 25752
rect 12952 25712 12958 25724
rect 21726 25712 21732 25724
rect 21784 25712 21790 25764
rect 8570 25644 8576 25696
rect 8628 25684 8634 25696
rect 25958 25684 25964 25696
rect 8628 25656 25964 25684
rect 8628 25644 8634 25656
rect 25958 25644 25964 25656
rect 26016 25644 26022 25696
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 12894 25480 12900 25492
rect 5092 25452 12900 25480
rect 5092 25421 5120 25452
rect 12894 25440 12900 25452
rect 12952 25440 12958 25492
rect 12989 25483 13047 25489
rect 12989 25449 13001 25483
rect 13035 25449 13047 25483
rect 12989 25443 13047 25449
rect 14093 25483 14151 25489
rect 14093 25449 14105 25483
rect 14139 25480 14151 25483
rect 15654 25480 15660 25492
rect 14139 25452 15660 25480
rect 14139 25449 14151 25452
rect 14093 25443 14151 25449
rect 5077 25415 5135 25421
rect 5077 25381 5089 25415
rect 5123 25381 5135 25415
rect 5077 25375 5135 25381
rect 8386 25372 8392 25424
rect 8444 25412 8450 25424
rect 8481 25415 8539 25421
rect 8481 25412 8493 25415
rect 8444 25384 8493 25412
rect 8444 25372 8450 25384
rect 8481 25381 8493 25384
rect 8527 25381 8539 25415
rect 13004 25412 13032 25443
rect 15654 25440 15660 25452
rect 15712 25440 15718 25492
rect 16850 25440 16856 25492
rect 16908 25480 16914 25492
rect 18509 25483 18567 25489
rect 18509 25480 18521 25483
rect 16908 25452 18521 25480
rect 16908 25440 16914 25452
rect 18509 25449 18521 25452
rect 18555 25449 18567 25483
rect 18509 25443 18567 25449
rect 20070 25440 20076 25492
rect 20128 25480 20134 25492
rect 21361 25483 21419 25489
rect 21361 25480 21373 25483
rect 20128 25452 21373 25480
rect 20128 25440 20134 25452
rect 21361 25449 21373 25452
rect 21407 25449 21419 25483
rect 21361 25443 21419 25449
rect 22186 25440 22192 25492
rect 22244 25480 22250 25492
rect 24213 25483 24271 25489
rect 24213 25480 24225 25483
rect 22244 25452 24225 25480
rect 22244 25440 22250 25452
rect 24213 25449 24225 25452
rect 24259 25449 24271 25483
rect 24213 25443 24271 25449
rect 25317 25483 25375 25489
rect 25317 25449 25329 25483
rect 25363 25480 25375 25483
rect 25406 25480 25412 25492
rect 25363 25452 25412 25480
rect 25363 25449 25375 25452
rect 25317 25443 25375 25449
rect 25406 25440 25412 25452
rect 25464 25440 25470 25492
rect 15749 25415 15807 25421
rect 13004 25384 15608 25412
rect 8481 25375 8539 25381
rect 4801 25347 4859 25353
rect 4801 25313 4813 25347
rect 4847 25344 4859 25347
rect 4847 25316 5120 25344
rect 4847 25313 4859 25316
rect 4801 25307 4859 25313
rect 5092 25288 5120 25316
rect 7098 25304 7104 25356
rect 7156 25344 7162 25356
rect 8573 25347 8631 25353
rect 8573 25344 8585 25347
rect 7156 25316 8585 25344
rect 7156 25304 7162 25316
rect 8573 25313 8585 25316
rect 8619 25313 8631 25347
rect 8573 25307 8631 25313
rect 10686 25304 10692 25356
rect 10744 25344 10750 25356
rect 11057 25347 11115 25353
rect 11057 25344 11069 25347
rect 10744 25316 11069 25344
rect 10744 25304 10750 25316
rect 11057 25313 11069 25316
rect 11103 25313 11115 25347
rect 11330 25344 11336 25356
rect 11291 25316 11336 25344
rect 11057 25307 11115 25313
rect 11330 25304 11336 25316
rect 11388 25304 11394 25356
rect 12805 25347 12863 25353
rect 12805 25313 12817 25347
rect 12851 25313 12863 25347
rect 12805 25307 12863 25313
rect 13909 25347 13967 25353
rect 13909 25313 13921 25347
rect 13955 25344 13967 25347
rect 14734 25344 14740 25356
rect 13955 25316 14740 25344
rect 13955 25313 13967 25316
rect 13909 25307 13967 25313
rect 1670 25276 1676 25288
rect 1631 25248 1676 25276
rect 1670 25236 1676 25248
rect 1728 25236 1734 25288
rect 5074 25236 5080 25288
rect 5132 25236 5138 25288
rect 8478 25276 8484 25288
rect 8439 25248 8484 25276
rect 8478 25236 8484 25248
rect 8536 25276 8542 25288
rect 8754 25276 8760 25288
rect 8536 25248 8760 25276
rect 8536 25236 8542 25248
rect 8754 25236 8760 25248
rect 8812 25236 8818 25288
rect 12820 25276 12848 25307
rect 14734 25304 14740 25316
rect 14792 25304 14798 25356
rect 15286 25304 15292 25356
rect 15344 25344 15350 25356
rect 15473 25347 15531 25353
rect 15473 25344 15485 25347
rect 15344 25316 15485 25344
rect 15344 25304 15350 25316
rect 15473 25313 15485 25316
rect 15519 25313 15531 25347
rect 15580 25344 15608 25384
rect 15749 25381 15761 25415
rect 15795 25412 15807 25415
rect 23474 25412 23480 25424
rect 15795 25384 23480 25412
rect 15795 25381 15807 25384
rect 15749 25375 15807 25381
rect 23474 25372 23480 25384
rect 23532 25372 23538 25424
rect 16298 25344 16304 25356
rect 15580 25316 16304 25344
rect 15473 25307 15531 25313
rect 16298 25304 16304 25316
rect 16356 25304 16362 25356
rect 16942 25344 16948 25356
rect 16903 25316 16948 25344
rect 16942 25304 16948 25316
rect 17000 25304 17006 25356
rect 18230 25304 18236 25356
rect 18288 25344 18294 25356
rect 18325 25347 18383 25353
rect 18325 25344 18337 25347
rect 18288 25316 18337 25344
rect 18288 25304 18294 25316
rect 18325 25313 18337 25316
rect 18371 25313 18383 25347
rect 19426 25344 19432 25356
rect 19387 25316 19432 25344
rect 18325 25307 18383 25313
rect 19426 25304 19432 25316
rect 19484 25304 19490 25356
rect 21082 25304 21088 25356
rect 21140 25344 21146 25356
rect 21177 25347 21235 25353
rect 21177 25344 21189 25347
rect 21140 25316 21189 25344
rect 21140 25304 21146 25316
rect 21177 25313 21189 25316
rect 21223 25313 21235 25347
rect 21177 25307 21235 25313
rect 22281 25347 22339 25353
rect 22281 25313 22293 25347
rect 22327 25344 22339 25347
rect 22646 25344 22652 25356
rect 22327 25316 22652 25344
rect 22327 25313 22339 25316
rect 22281 25307 22339 25313
rect 13449 25279 13507 25285
rect 13449 25276 13461 25279
rect 12820 25248 13461 25276
rect 13449 25245 13461 25248
rect 13495 25276 13507 25279
rect 15654 25276 15660 25288
rect 13495 25248 15660 25276
rect 13495 25245 13507 25248
rect 13449 25239 13507 25245
rect 15654 25236 15660 25248
rect 15712 25236 15718 25288
rect 17129 25279 17187 25285
rect 17129 25245 17141 25279
rect 17175 25245 17187 25279
rect 17129 25239 17187 25245
rect 3970 25168 3976 25220
rect 4028 25208 4034 25220
rect 10594 25208 10600 25220
rect 4028 25180 10600 25208
rect 4028 25168 4034 25180
rect 10594 25168 10600 25180
rect 10652 25168 10658 25220
rect 4341 25143 4399 25149
rect 4341 25109 4353 25143
rect 4387 25140 4399 25143
rect 4706 25140 4712 25152
rect 4387 25112 4712 25140
rect 4387 25109 4399 25112
rect 4341 25103 4399 25109
rect 4706 25100 4712 25112
rect 4764 25100 4770 25152
rect 7745 25143 7803 25149
rect 7745 25109 7757 25143
rect 7791 25140 7803 25143
rect 7834 25140 7840 25152
rect 7791 25112 7840 25140
rect 7791 25109 7803 25112
rect 7745 25103 7803 25109
rect 7834 25100 7840 25112
rect 7892 25100 7898 25152
rect 8021 25143 8079 25149
rect 8021 25109 8033 25143
rect 8067 25140 8079 25143
rect 9398 25140 9404 25152
rect 8067 25112 9404 25140
rect 8067 25109 8079 25112
rect 8021 25103 8079 25109
rect 9398 25100 9404 25112
rect 9456 25100 9462 25152
rect 10873 25143 10931 25149
rect 10873 25109 10885 25143
rect 10919 25140 10931 25143
rect 11330 25140 11336 25152
rect 10919 25112 11336 25140
rect 10919 25109 10931 25112
rect 10873 25103 10931 25109
rect 11330 25100 11336 25112
rect 11388 25100 11394 25152
rect 14090 25100 14096 25152
rect 14148 25140 14154 25152
rect 14461 25143 14519 25149
rect 14461 25140 14473 25143
rect 14148 25112 14473 25140
rect 14148 25100 14154 25112
rect 14461 25109 14473 25112
rect 14507 25109 14519 25143
rect 17144 25140 17172 25239
rect 17218 25236 17224 25288
rect 17276 25276 17282 25288
rect 22296 25276 22324 25307
rect 22646 25304 22652 25316
rect 22704 25304 22710 25356
rect 24026 25344 24032 25356
rect 23987 25316 24032 25344
rect 24026 25304 24032 25316
rect 24084 25304 24090 25356
rect 25133 25347 25191 25353
rect 25133 25313 25145 25347
rect 25179 25344 25191 25347
rect 25682 25344 25688 25356
rect 25179 25316 25688 25344
rect 25179 25313 25191 25316
rect 25133 25307 25191 25313
rect 25682 25304 25688 25316
rect 25740 25304 25746 25356
rect 17276 25248 22324 25276
rect 17276 25236 17282 25248
rect 17402 25168 17408 25220
rect 17460 25208 17466 25220
rect 19613 25211 19671 25217
rect 19613 25208 19625 25211
rect 17460 25180 19625 25208
rect 17460 25168 17466 25180
rect 19613 25177 19625 25180
rect 19659 25177 19671 25211
rect 19613 25171 19671 25177
rect 20622 25168 20628 25220
rect 20680 25208 20686 25220
rect 22465 25211 22523 25217
rect 22465 25208 22477 25211
rect 20680 25180 22477 25208
rect 20680 25168 20686 25180
rect 22465 25177 22477 25180
rect 22511 25177 22523 25211
rect 22465 25171 22523 25177
rect 20162 25140 20168 25152
rect 17144 25112 20168 25140
rect 14461 25103 14519 25109
rect 20162 25100 20168 25112
rect 20220 25100 20226 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 8386 24896 8392 24948
rect 8444 24936 8450 24948
rect 8665 24939 8723 24945
rect 8665 24936 8677 24939
rect 8444 24908 8677 24936
rect 8444 24896 8450 24908
rect 8665 24905 8677 24908
rect 8711 24905 8723 24939
rect 8665 24899 8723 24905
rect 13078 24896 13084 24948
rect 13136 24936 13142 24948
rect 22646 24936 22652 24948
rect 13136 24908 22508 24936
rect 22607 24908 22652 24936
rect 13136 24896 13142 24908
rect 8478 24868 8484 24880
rect 8312 24840 8484 24868
rect 1578 24800 1584 24812
rect 1539 24772 1584 24800
rect 1578 24760 1584 24772
rect 1636 24760 1642 24812
rect 2869 24803 2927 24809
rect 2869 24800 2881 24803
rect 2148 24772 2881 24800
rect 1762 24692 1768 24744
rect 1820 24732 1826 24744
rect 2148 24741 2176 24772
rect 2869 24769 2881 24772
rect 2915 24769 2927 24803
rect 2869 24763 2927 24769
rect 3786 24760 3792 24812
rect 3844 24800 3850 24812
rect 3881 24803 3939 24809
rect 3881 24800 3893 24803
rect 3844 24772 3893 24800
rect 3844 24760 3850 24772
rect 3881 24769 3893 24772
rect 3927 24800 3939 24803
rect 4525 24803 4583 24809
rect 4525 24800 4537 24803
rect 3927 24772 4537 24800
rect 3927 24769 3939 24772
rect 3881 24763 3939 24769
rect 4525 24769 4537 24772
rect 4571 24769 4583 24803
rect 4706 24800 4712 24812
rect 4667 24772 4712 24800
rect 4525 24763 4583 24769
rect 4706 24760 4712 24772
rect 4764 24760 4770 24812
rect 7561 24803 7619 24809
rect 7561 24769 7573 24803
rect 7607 24800 7619 24803
rect 8312 24800 8340 24840
rect 8478 24828 8484 24840
rect 8536 24828 8542 24880
rect 10873 24871 10931 24877
rect 10873 24837 10885 24871
rect 10919 24837 10931 24871
rect 10873 24831 10931 24837
rect 12529 24871 12587 24877
rect 12529 24837 12541 24871
rect 12575 24837 12587 24871
rect 21082 24868 21088 24880
rect 12529 24831 12587 24837
rect 16040 24840 21088 24868
rect 10594 24800 10600 24812
rect 7607 24772 8340 24800
rect 10555 24772 10600 24800
rect 7607 24769 7619 24772
rect 7561 24763 7619 24769
rect 10594 24760 10600 24772
rect 10652 24760 10658 24812
rect 10888 24800 10916 24831
rect 10962 24800 10968 24812
rect 10888 24772 10968 24800
rect 10962 24760 10968 24772
rect 11020 24760 11026 24812
rect 11330 24760 11336 24812
rect 11388 24800 11394 24812
rect 11425 24803 11483 24809
rect 11425 24800 11437 24803
rect 11388 24772 11437 24800
rect 11388 24760 11394 24772
rect 11425 24769 11437 24772
rect 11471 24800 11483 24803
rect 11606 24800 11612 24812
rect 11471 24772 11612 24800
rect 11471 24769 11483 24772
rect 11425 24763 11483 24769
rect 11606 24760 11612 24772
rect 11664 24760 11670 24812
rect 12544 24800 12572 24831
rect 15562 24800 15568 24812
rect 12544 24772 15568 24800
rect 15562 24760 15568 24772
rect 15620 24760 15626 24812
rect 16040 24809 16068 24840
rect 21082 24828 21088 24840
rect 21140 24868 21146 24880
rect 21545 24871 21603 24877
rect 21545 24868 21557 24871
rect 21140 24840 21557 24868
rect 21140 24828 21146 24840
rect 21545 24837 21557 24840
rect 21591 24837 21603 24871
rect 22480 24868 22508 24908
rect 22646 24896 22652 24908
rect 22704 24896 22710 24948
rect 24762 24868 24768 24880
rect 22480 24840 24768 24868
rect 21545 24831 21603 24837
rect 24762 24828 24768 24840
rect 24820 24828 24826 24880
rect 16025 24803 16083 24809
rect 16025 24769 16037 24803
rect 16071 24769 16083 24803
rect 16025 24763 16083 24769
rect 18325 24803 18383 24809
rect 18325 24769 18337 24803
rect 18371 24800 18383 24803
rect 23474 24800 23480 24812
rect 18371 24772 21772 24800
rect 23435 24772 23480 24800
rect 18371 24769 18383 24772
rect 18325 24763 18383 24769
rect 2133 24735 2191 24741
rect 2133 24732 2145 24735
rect 1820 24704 2145 24732
rect 1820 24692 1826 24704
rect 2133 24701 2145 24704
rect 2179 24701 2191 24735
rect 10612 24732 10640 24760
rect 12253 24735 12311 24741
rect 10612 24704 11376 24732
rect 2133 24695 2191 24701
rect 2406 24664 2412 24676
rect 2367 24636 2412 24664
rect 2406 24624 2412 24636
rect 2464 24624 2470 24676
rect 3605 24667 3663 24673
rect 3605 24633 3617 24667
rect 3651 24664 3663 24667
rect 3694 24664 3700 24676
rect 3651 24636 3700 24664
rect 3651 24633 3663 24636
rect 3605 24627 3663 24633
rect 3694 24624 3700 24636
rect 3752 24664 3758 24676
rect 4617 24667 4675 24673
rect 4617 24664 4629 24667
rect 3752 24636 4629 24664
rect 3752 24624 3758 24636
rect 4617 24633 4629 24636
rect 4663 24633 4675 24667
rect 4617 24627 4675 24633
rect 7006 24624 7012 24676
rect 7064 24664 7070 24676
rect 7834 24664 7840 24676
rect 7064 24636 7840 24664
rect 7064 24624 7070 24636
rect 7834 24624 7840 24636
rect 7892 24664 7898 24676
rect 8021 24667 8079 24673
rect 8021 24664 8033 24667
rect 7892 24636 8033 24664
rect 7892 24624 7898 24636
rect 8021 24633 8033 24636
rect 8067 24633 8079 24667
rect 8294 24664 8300 24676
rect 8255 24636 8300 24664
rect 8021 24627 8079 24633
rect 8294 24624 8300 24636
rect 8352 24624 8358 24676
rect 10321 24667 10379 24673
rect 8588 24636 9168 24664
rect 1394 24556 1400 24608
rect 1452 24596 1458 24608
rect 1949 24599 2007 24605
rect 1949 24596 1961 24599
rect 1452 24568 1961 24596
rect 1452 24556 1458 24568
rect 1949 24565 1961 24568
rect 1995 24565 2007 24599
rect 1949 24559 2007 24565
rect 4147 24599 4205 24605
rect 4147 24565 4159 24599
rect 4193 24596 4205 24599
rect 4338 24596 4344 24608
rect 4193 24568 4344 24596
rect 4193 24565 4205 24568
rect 4147 24559 4205 24565
rect 4338 24556 4344 24568
rect 4396 24556 4402 24608
rect 5074 24596 5080 24608
rect 5035 24568 5080 24596
rect 5074 24556 5080 24568
rect 5132 24556 5138 24608
rect 5534 24556 5540 24608
rect 5592 24596 5598 24608
rect 5629 24599 5687 24605
rect 5629 24596 5641 24599
rect 5592 24568 5641 24596
rect 5592 24556 5598 24568
rect 5629 24565 5641 24568
rect 5675 24565 5687 24599
rect 7098 24596 7104 24608
rect 7059 24568 7104 24596
rect 5629 24559 5687 24565
rect 7098 24556 7104 24568
rect 7156 24556 7162 24608
rect 7742 24605 7748 24608
rect 7735 24599 7748 24605
rect 7735 24596 7747 24599
rect 7703 24568 7747 24596
rect 7735 24565 7747 24568
rect 7735 24559 7748 24565
rect 7742 24556 7748 24559
rect 7800 24556 7806 24608
rect 8205 24599 8263 24605
rect 8205 24565 8217 24599
rect 8251 24596 8263 24599
rect 8588 24596 8616 24636
rect 9140 24605 9168 24636
rect 10321 24633 10333 24667
rect 10367 24664 10379 24667
rect 10686 24664 10692 24676
rect 10367 24636 10692 24664
rect 10367 24633 10379 24636
rect 10321 24627 10379 24633
rect 10686 24624 10692 24636
rect 10744 24624 10750 24676
rect 10870 24624 10876 24676
rect 10928 24664 10934 24676
rect 11348 24673 11376 24704
rect 12253 24701 12265 24735
rect 12299 24732 12311 24735
rect 13081 24735 13139 24741
rect 13081 24732 13093 24735
rect 12299 24704 13093 24732
rect 12299 24701 12311 24704
rect 12253 24695 12311 24701
rect 13081 24701 13093 24704
rect 13127 24732 13139 24735
rect 13446 24732 13452 24744
rect 13127 24704 13452 24732
rect 13127 24701 13139 24704
rect 13081 24695 13139 24701
rect 13446 24692 13452 24704
rect 13504 24692 13510 24744
rect 14090 24692 14096 24744
rect 14148 24732 14154 24744
rect 14829 24735 14887 24741
rect 14829 24732 14841 24735
rect 14148 24704 14841 24732
rect 14148 24692 14154 24704
rect 14829 24701 14841 24704
rect 14875 24701 14887 24735
rect 14829 24695 14887 24701
rect 15378 24692 15384 24744
rect 15436 24732 15442 24744
rect 15749 24735 15807 24741
rect 15749 24732 15761 24735
rect 15436 24704 15761 24732
rect 15436 24692 15442 24704
rect 15749 24701 15761 24704
rect 15795 24732 15807 24735
rect 16485 24735 16543 24741
rect 16485 24732 16497 24735
rect 15795 24704 16497 24732
rect 15795 24701 15807 24704
rect 15749 24695 15807 24701
rect 16485 24701 16497 24704
rect 16531 24701 16543 24735
rect 18046 24732 18052 24744
rect 18007 24704 18052 24732
rect 16485 24695 16543 24701
rect 18046 24692 18052 24704
rect 18104 24732 18110 24744
rect 18785 24735 18843 24741
rect 18785 24732 18797 24735
rect 18104 24704 18797 24732
rect 18104 24692 18110 24704
rect 18785 24701 18797 24704
rect 18831 24701 18843 24735
rect 18785 24695 18843 24701
rect 19334 24692 19340 24744
rect 19392 24732 19398 24744
rect 20073 24735 20131 24741
rect 20073 24732 20085 24735
rect 19392 24704 20085 24732
rect 19392 24692 19398 24704
rect 20073 24701 20085 24704
rect 20119 24701 20131 24735
rect 20622 24732 20628 24744
rect 20583 24704 20628 24732
rect 20073 24695 20131 24701
rect 20622 24692 20628 24704
rect 20680 24732 20686 24744
rect 21744 24741 21772 24772
rect 23474 24760 23480 24772
rect 23532 24760 23538 24812
rect 21177 24735 21235 24741
rect 21177 24732 21189 24735
rect 20680 24704 21189 24732
rect 20680 24692 20686 24704
rect 21177 24701 21189 24704
rect 21223 24701 21235 24735
rect 21177 24695 21235 24701
rect 21729 24735 21787 24741
rect 21729 24701 21741 24735
rect 21775 24732 21787 24735
rect 22281 24735 22339 24741
rect 22281 24732 22293 24735
rect 21775 24704 22293 24732
rect 21775 24701 21787 24704
rect 21729 24695 21787 24701
rect 22281 24701 22293 24704
rect 22327 24701 22339 24735
rect 23492 24732 23520 24760
rect 23661 24735 23719 24741
rect 23661 24732 23673 24735
rect 23492 24704 23673 24732
rect 22281 24695 22339 24701
rect 23661 24701 23673 24704
rect 23707 24701 23719 24735
rect 24762 24732 24768 24744
rect 24723 24704 24768 24732
rect 23661 24695 23719 24701
rect 24762 24692 24768 24704
rect 24820 24732 24826 24744
rect 25317 24735 25375 24741
rect 25317 24732 25329 24735
rect 24820 24704 25329 24732
rect 24820 24692 24826 24704
rect 25317 24701 25329 24704
rect 25363 24701 25375 24735
rect 25317 24695 25375 24701
rect 11149 24667 11207 24673
rect 11149 24664 11161 24667
rect 10928 24636 11161 24664
rect 10928 24624 10934 24636
rect 11149 24633 11161 24636
rect 11195 24633 11207 24667
rect 11149 24627 11207 24633
rect 11333 24667 11391 24673
rect 11333 24633 11345 24667
rect 11379 24664 11391 24667
rect 11698 24664 11704 24676
rect 11379 24636 11704 24664
rect 11379 24633 11391 24636
rect 11333 24627 11391 24633
rect 11698 24624 11704 24636
rect 11756 24624 11762 24676
rect 11885 24667 11943 24673
rect 11885 24633 11897 24667
rect 11931 24664 11943 24667
rect 12526 24664 12532 24676
rect 11931 24636 12532 24664
rect 11931 24633 11943 24636
rect 11885 24627 11943 24633
rect 12526 24624 12532 24636
rect 12584 24624 12590 24676
rect 12802 24664 12808 24676
rect 12763 24636 12808 24664
rect 12802 24624 12808 24636
rect 12860 24624 12866 24676
rect 14001 24667 14059 24673
rect 14001 24633 14013 24667
rect 14047 24664 14059 24667
rect 14553 24667 14611 24673
rect 14553 24664 14565 24667
rect 14047 24636 14565 24664
rect 14047 24633 14059 24636
rect 14001 24627 14059 24633
rect 14553 24633 14565 24636
rect 14599 24664 14611 24667
rect 15470 24664 15476 24676
rect 14599 24636 15476 24664
rect 14599 24633 14611 24636
rect 14553 24627 14611 24633
rect 15470 24624 15476 24636
rect 15528 24624 15534 24676
rect 18230 24624 18236 24676
rect 18288 24664 18294 24676
rect 19153 24667 19211 24673
rect 19153 24664 19165 24667
rect 18288 24636 19165 24664
rect 18288 24624 18294 24636
rect 19153 24633 19165 24636
rect 19199 24633 19211 24667
rect 19153 24627 19211 24633
rect 19613 24667 19671 24673
rect 19613 24633 19625 24667
rect 19659 24664 19671 24667
rect 20530 24664 20536 24676
rect 19659 24636 20536 24664
rect 19659 24633 19671 24636
rect 19613 24627 19671 24633
rect 20530 24624 20536 24636
rect 20588 24624 20594 24676
rect 8251 24568 8616 24596
rect 9125 24599 9183 24605
rect 8251 24565 8263 24568
rect 8205 24559 8263 24565
rect 9125 24565 9137 24599
rect 9171 24596 9183 24599
rect 9582 24596 9588 24608
rect 9171 24568 9588 24596
rect 9171 24565 9183 24568
rect 9125 24559 9183 24565
rect 9582 24556 9588 24568
rect 9640 24556 9646 24608
rect 12544 24596 12572 24624
rect 12989 24599 13047 24605
rect 12989 24596 13001 24599
rect 12544 24568 13001 24596
rect 12989 24565 13001 24568
rect 13035 24565 13047 24599
rect 12989 24559 13047 24565
rect 13354 24556 13360 24608
rect 13412 24596 13418 24608
rect 13633 24599 13691 24605
rect 13633 24596 13645 24599
rect 13412 24568 13645 24596
rect 13412 24556 13418 24568
rect 13633 24565 13645 24568
rect 13679 24565 13691 24599
rect 13633 24559 13691 24565
rect 14267 24599 14325 24605
rect 14267 24565 14279 24599
rect 14313 24596 14325 24599
rect 14458 24596 14464 24608
rect 14313 24568 14464 24596
rect 14313 24565 14325 24568
rect 14267 24559 14325 24565
rect 14458 24556 14464 24568
rect 14516 24556 14522 24608
rect 14737 24599 14795 24605
rect 14737 24565 14749 24599
rect 14783 24596 14795 24599
rect 14826 24596 14832 24608
rect 14783 24568 14832 24596
rect 14783 24565 14795 24568
rect 14737 24559 14795 24565
rect 14826 24556 14832 24568
rect 14884 24556 14890 24608
rect 15286 24596 15292 24608
rect 15247 24568 15292 24596
rect 15286 24556 15292 24568
rect 15344 24556 15350 24608
rect 16390 24556 16396 24608
rect 16448 24596 16454 24608
rect 16942 24596 16948 24608
rect 16448 24568 16948 24596
rect 16448 24556 16454 24568
rect 16942 24556 16948 24568
rect 17000 24556 17006 24608
rect 17865 24599 17923 24605
rect 17865 24565 17877 24599
rect 17911 24596 17923 24599
rect 18322 24596 18328 24608
rect 17911 24568 18328 24596
rect 17911 24565 17923 24568
rect 17865 24559 17923 24565
rect 18322 24556 18328 24568
rect 18380 24556 18386 24608
rect 20806 24596 20812 24608
rect 20767 24568 20812 24596
rect 20806 24556 20812 24568
rect 20864 24556 20870 24608
rect 21910 24596 21916 24608
rect 21871 24568 21916 24596
rect 21910 24556 21916 24568
rect 21968 24556 21974 24608
rect 23842 24596 23848 24608
rect 23803 24568 23848 24596
rect 23842 24556 23848 24568
rect 23900 24556 23906 24608
rect 24026 24556 24032 24608
rect 24084 24596 24090 24608
rect 24213 24599 24271 24605
rect 24213 24596 24225 24599
rect 24084 24568 24225 24596
rect 24084 24556 24090 24568
rect 24213 24565 24225 24568
rect 24259 24565 24271 24599
rect 24946 24596 24952 24608
rect 24907 24568 24952 24596
rect 24213 24559 24271 24565
rect 24946 24556 24952 24568
rect 25004 24556 25010 24608
rect 25682 24596 25688 24608
rect 25643 24568 25688 24596
rect 25682 24556 25688 24568
rect 25740 24556 25746 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 2501 24395 2559 24401
rect 2501 24392 2513 24395
rect 1872 24364 2513 24392
rect 1670 24284 1676 24336
rect 1728 24324 1734 24336
rect 1872 24333 1900 24364
rect 2501 24361 2513 24364
rect 2547 24361 2559 24395
rect 2501 24355 2559 24361
rect 8294 24352 8300 24404
rect 8352 24392 8358 24404
rect 8389 24395 8447 24401
rect 8389 24392 8401 24395
rect 8352 24364 8401 24392
rect 8352 24352 8358 24364
rect 8389 24361 8401 24364
rect 8435 24361 8447 24395
rect 8389 24355 8447 24361
rect 10045 24395 10103 24401
rect 10045 24361 10057 24395
rect 10091 24392 10103 24395
rect 10870 24392 10876 24404
rect 10091 24364 10876 24392
rect 10091 24361 10103 24364
rect 10045 24355 10103 24361
rect 10870 24352 10876 24364
rect 10928 24352 10934 24404
rect 11606 24352 11612 24404
rect 11664 24392 11670 24404
rect 12437 24395 12495 24401
rect 12437 24392 12449 24395
rect 11664 24364 12449 24392
rect 11664 24352 11670 24364
rect 12437 24361 12449 24364
rect 12483 24361 12495 24395
rect 12437 24355 12495 24361
rect 13354 24352 13360 24404
rect 13412 24392 13418 24404
rect 14826 24392 14832 24404
rect 13412 24364 14832 24392
rect 13412 24352 13418 24364
rect 14826 24352 14832 24364
rect 14884 24352 14890 24404
rect 19426 24392 19432 24404
rect 18800 24364 19432 24392
rect 1857 24327 1915 24333
rect 1857 24324 1869 24327
rect 1728 24296 1869 24324
rect 1728 24284 1734 24296
rect 1857 24293 1869 24296
rect 1903 24293 1915 24327
rect 2038 24324 2044 24336
rect 1999 24296 2044 24324
rect 1857 24287 1915 24293
rect 2038 24284 2044 24296
rect 2096 24324 2102 24336
rect 2869 24327 2927 24333
rect 2869 24324 2881 24327
rect 2096 24296 2881 24324
rect 2096 24284 2102 24296
rect 2869 24293 2881 24296
rect 2915 24293 2927 24327
rect 2869 24287 2927 24293
rect 7285 24327 7343 24333
rect 7285 24293 7297 24327
rect 7331 24324 7343 24327
rect 7926 24324 7932 24336
rect 7331 24296 7932 24324
rect 7331 24293 7343 24296
rect 7285 24287 7343 24293
rect 7926 24284 7932 24296
rect 7984 24284 7990 24336
rect 8021 24327 8079 24333
rect 8021 24293 8033 24327
rect 8067 24324 8079 24327
rect 8110 24324 8116 24336
rect 8067 24296 8116 24324
rect 8067 24293 8079 24296
rect 8021 24287 8079 24293
rect 8110 24284 8116 24296
rect 8168 24324 8174 24336
rect 8570 24324 8576 24336
rect 8168 24296 8576 24324
rect 8168 24284 8174 24296
rect 8570 24284 8576 24296
rect 8628 24284 8634 24336
rect 11324 24327 11382 24333
rect 11324 24293 11336 24327
rect 11370 24324 11382 24327
rect 11514 24324 11520 24336
rect 11370 24296 11520 24324
rect 11370 24293 11382 24296
rect 11324 24287 11382 24293
rect 11514 24284 11520 24296
rect 11572 24284 11578 24336
rect 13814 24284 13820 24336
rect 13872 24324 13878 24336
rect 14185 24327 14243 24333
rect 14185 24324 14197 24327
rect 13872 24296 14197 24324
rect 13872 24284 13878 24296
rect 14185 24293 14197 24296
rect 14231 24293 14243 24327
rect 14185 24287 14243 24293
rect 17497 24327 17555 24333
rect 17497 24293 17509 24327
rect 17543 24324 17555 24327
rect 17586 24324 17592 24336
rect 17543 24296 17592 24324
rect 17543 24293 17555 24296
rect 17497 24287 17555 24293
rect 17586 24284 17592 24296
rect 17644 24284 17650 24336
rect 18800 24333 18828 24364
rect 19426 24352 19432 24364
rect 19484 24352 19490 24404
rect 24854 24392 24860 24404
rect 24815 24364 24860 24392
rect 24854 24352 24860 24364
rect 24912 24352 24918 24404
rect 18785 24327 18843 24333
rect 18785 24293 18797 24327
rect 18831 24293 18843 24327
rect 18785 24287 18843 24293
rect 19334 24284 19340 24336
rect 19392 24284 19398 24336
rect 23106 24284 23112 24336
rect 23164 24324 23170 24336
rect 23661 24327 23719 24333
rect 23661 24324 23673 24327
rect 23164 24296 23673 24324
rect 23164 24284 23170 24296
rect 23661 24293 23673 24296
rect 23707 24293 23719 24327
rect 23661 24287 23719 24293
rect 658 24216 664 24268
rect 716 24256 722 24268
rect 4982 24256 4988 24268
rect 716 24228 4988 24256
rect 716 24216 722 24228
rect 4982 24216 4988 24228
rect 5040 24216 5046 24268
rect 5166 24265 5172 24268
rect 5160 24256 5172 24265
rect 5127 24228 5172 24256
rect 5160 24219 5172 24228
rect 5166 24216 5172 24219
rect 5224 24216 5230 24268
rect 7742 24256 7748 24268
rect 7703 24228 7748 24256
rect 7742 24216 7748 24228
rect 7800 24216 7806 24268
rect 13170 24216 13176 24268
rect 13228 24256 13234 24268
rect 13630 24256 13636 24268
rect 13228 24228 13636 24256
rect 13228 24216 13234 24228
rect 13630 24216 13636 24228
rect 13688 24216 13694 24268
rect 14277 24259 14335 24265
rect 14277 24256 14289 24259
rect 13924 24228 14289 24256
rect 13924 24200 13952 24228
rect 14277 24225 14289 24228
rect 14323 24225 14335 24259
rect 15562 24256 15568 24268
rect 15523 24228 15568 24256
rect 14277 24219 14335 24225
rect 15562 24216 15568 24228
rect 15620 24216 15626 24268
rect 16853 24259 16911 24265
rect 16853 24225 16865 24259
rect 16899 24256 16911 24259
rect 16899 24228 17632 24256
rect 16899 24225 16911 24228
rect 16853 24219 16911 24225
rect 2133 24191 2191 24197
rect 2133 24157 2145 24191
rect 2179 24188 2191 24191
rect 3418 24188 3424 24200
rect 2179 24160 3424 24188
rect 2179 24157 2191 24160
rect 2133 24151 2191 24157
rect 3418 24148 3424 24160
rect 3476 24148 3482 24200
rect 4154 24148 4160 24200
rect 4212 24188 4218 24200
rect 4893 24191 4951 24197
rect 4893 24188 4905 24191
rect 4212 24160 4905 24188
rect 4212 24148 4218 24160
rect 4893 24157 4905 24160
rect 4939 24157 4951 24191
rect 11054 24188 11060 24200
rect 11015 24160 11060 24188
rect 4893 24151 4951 24157
rect 11054 24148 11060 24160
rect 11112 24148 11118 24200
rect 13541 24191 13599 24197
rect 13541 24157 13553 24191
rect 13587 24188 13599 24191
rect 13906 24188 13912 24200
rect 13587 24160 13912 24188
rect 13587 24157 13599 24160
rect 13541 24151 13599 24157
rect 13906 24148 13912 24160
rect 13964 24148 13970 24200
rect 13998 24148 14004 24200
rect 14056 24188 14062 24200
rect 14093 24191 14151 24197
rect 14093 24188 14105 24191
rect 14056 24160 14105 24188
rect 14056 24148 14062 24160
rect 14093 24157 14105 24160
rect 14139 24157 14151 24191
rect 14093 24151 14151 24157
rect 15841 24191 15899 24197
rect 15841 24157 15853 24191
rect 15887 24188 15899 24191
rect 16022 24188 16028 24200
rect 15887 24160 16028 24188
rect 15887 24157 15899 24160
rect 15841 24151 15899 24157
rect 16022 24148 16028 24160
rect 16080 24148 16086 24200
rect 17494 24188 17500 24200
rect 17455 24160 17500 24188
rect 17494 24148 17500 24160
rect 17552 24148 17558 24200
rect 17604 24197 17632 24228
rect 18322 24216 18328 24268
rect 18380 24256 18386 24268
rect 18509 24259 18567 24265
rect 18509 24256 18521 24259
rect 18380 24228 18521 24256
rect 18380 24216 18386 24228
rect 18509 24225 18521 24228
rect 18555 24225 18567 24259
rect 18509 24219 18567 24225
rect 17589 24191 17647 24197
rect 17589 24157 17601 24191
rect 17635 24157 17647 24191
rect 17589 24151 17647 24157
rect 1581 24123 1639 24129
rect 1581 24089 1593 24123
rect 1627 24120 1639 24123
rect 1762 24120 1768 24132
rect 1627 24092 1768 24120
rect 1627 24089 1639 24092
rect 1581 24083 1639 24089
rect 1762 24080 1768 24092
rect 1820 24080 1826 24132
rect 12802 24080 12808 24132
rect 12860 24120 12866 24132
rect 13081 24123 13139 24129
rect 13081 24120 13093 24123
rect 12860 24092 13093 24120
rect 12860 24080 12866 24092
rect 13081 24089 13093 24092
rect 13127 24120 13139 24123
rect 13630 24120 13636 24132
rect 13127 24092 13636 24120
rect 13127 24089 13139 24092
rect 13081 24083 13139 24089
rect 13630 24080 13636 24092
rect 13688 24080 13694 24132
rect 14182 24080 14188 24132
rect 14240 24120 14246 24132
rect 14550 24120 14556 24132
rect 14240 24092 14556 24120
rect 14240 24080 14246 24092
rect 14550 24080 14556 24092
rect 14608 24080 14614 24132
rect 16485 24123 16543 24129
rect 16485 24089 16497 24123
rect 16531 24120 16543 24123
rect 17126 24120 17132 24132
rect 16531 24092 17132 24120
rect 16531 24089 16543 24092
rect 16485 24083 16543 24089
rect 17126 24080 17132 24092
rect 17184 24080 17190 24132
rect 4341 24055 4399 24061
rect 4341 24021 4353 24055
rect 4387 24052 4399 24055
rect 4522 24052 4528 24064
rect 4387 24024 4528 24052
rect 4387 24021 4399 24024
rect 4341 24015 4399 24021
rect 4522 24012 4528 24024
rect 4580 24012 4586 24064
rect 6270 24052 6276 24064
rect 6231 24024 6276 24052
rect 6270 24012 6276 24024
rect 6328 24012 6334 24064
rect 7190 24012 7196 24064
rect 7248 24052 7254 24064
rect 7469 24055 7527 24061
rect 7469 24052 7481 24055
rect 7248 24024 7481 24052
rect 7248 24012 7254 24024
rect 7469 24021 7481 24024
rect 7515 24021 7527 24055
rect 13722 24052 13728 24064
rect 13683 24024 13728 24052
rect 7469 24015 7527 24021
rect 13722 24012 13728 24024
rect 13780 24012 13786 24064
rect 14734 24052 14740 24064
rect 14695 24024 14740 24052
rect 14734 24012 14740 24024
rect 14792 24012 14798 24064
rect 16942 24012 16948 24064
rect 17000 24052 17006 24064
rect 17037 24055 17095 24061
rect 17037 24052 17049 24055
rect 17000 24024 17049 24052
rect 17000 24012 17006 24024
rect 17037 24021 17049 24024
rect 17083 24021 17095 24055
rect 17604 24052 17632 24151
rect 19352 24064 19380 24284
rect 21821 24259 21879 24265
rect 21821 24225 21833 24259
rect 21867 24256 21879 24259
rect 21910 24256 21916 24268
rect 21867 24228 21916 24256
rect 21867 24225 21879 24228
rect 21821 24219 21879 24225
rect 21910 24216 21916 24228
rect 21968 24256 21974 24268
rect 22557 24259 22615 24265
rect 22557 24256 22569 24259
rect 21968 24228 22569 24256
rect 21968 24216 21974 24228
rect 22557 24225 22569 24228
rect 22603 24225 22615 24259
rect 22557 24219 22615 24225
rect 24210 24216 24216 24268
rect 24268 24256 24274 24268
rect 24673 24259 24731 24265
rect 24673 24256 24685 24259
rect 24268 24228 24685 24256
rect 24268 24216 24274 24228
rect 24673 24225 24685 24228
rect 24719 24256 24731 24259
rect 24946 24256 24952 24268
rect 24719 24228 24952 24256
rect 24719 24225 24731 24228
rect 24673 24219 24731 24225
rect 24946 24216 24952 24228
rect 25004 24216 25010 24268
rect 19426 24148 19432 24200
rect 19484 24148 19490 24200
rect 19794 24188 19800 24200
rect 19755 24160 19800 24188
rect 19794 24148 19800 24160
rect 19852 24148 19858 24200
rect 22094 24148 22100 24200
rect 22152 24188 22158 24200
rect 23566 24188 23572 24200
rect 22152 24160 22197 24188
rect 23527 24160 23572 24188
rect 22152 24148 22158 24160
rect 23566 24148 23572 24160
rect 23624 24148 23630 24200
rect 23753 24191 23811 24197
rect 23753 24157 23765 24191
rect 23799 24157 23811 24191
rect 23753 24151 23811 24157
rect 19444 24120 19472 24148
rect 20438 24120 20444 24132
rect 19444 24092 20444 24120
rect 20438 24080 20444 24092
rect 20496 24080 20502 24132
rect 23768 24120 23796 24151
rect 24121 24123 24179 24129
rect 24121 24120 24133 24123
rect 22940 24092 24133 24120
rect 22940 24064 22968 24092
rect 24121 24089 24133 24092
rect 24167 24089 24179 24123
rect 24121 24083 24179 24089
rect 18141 24055 18199 24061
rect 18141 24052 18153 24055
rect 17604 24024 18153 24052
rect 17037 24015 17095 24021
rect 18141 24021 18153 24024
rect 18187 24052 18199 24055
rect 18506 24052 18512 24064
rect 18187 24024 18512 24052
rect 18187 24021 18199 24024
rect 18141 24015 18199 24021
rect 18506 24012 18512 24024
rect 18564 24012 18570 24064
rect 19334 24012 19340 24064
rect 19392 24012 19398 24064
rect 20346 24052 20352 24064
rect 20307 24024 20352 24052
rect 20346 24012 20352 24024
rect 20404 24012 20410 24064
rect 22922 24052 22928 24064
rect 22883 24024 22928 24052
rect 22922 24012 22928 24024
rect 22980 24012 22986 24064
rect 23201 24055 23259 24061
rect 23201 24021 23213 24055
rect 23247 24052 23259 24055
rect 23382 24052 23388 24064
rect 23247 24024 23388 24052
rect 23247 24021 23259 24024
rect 23201 24015 23259 24021
rect 23382 24012 23388 24024
rect 23440 24012 23446 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 4154 23848 4160 23860
rect 4115 23820 4160 23848
rect 4154 23808 4160 23820
rect 4212 23808 4218 23860
rect 7377 23851 7435 23857
rect 7377 23817 7389 23851
rect 7423 23848 7435 23851
rect 8110 23848 8116 23860
rect 7423 23820 8116 23848
rect 7423 23817 7435 23820
rect 7377 23811 7435 23817
rect 8110 23808 8116 23820
rect 8168 23808 8174 23860
rect 8386 23808 8392 23860
rect 8444 23848 8450 23860
rect 8849 23851 8907 23857
rect 8849 23848 8861 23851
rect 8444 23820 8861 23848
rect 8444 23808 8450 23820
rect 8849 23817 8861 23820
rect 8895 23817 8907 23851
rect 9398 23848 9404 23860
rect 9359 23820 9404 23848
rect 8849 23811 8907 23817
rect 1394 23712 1400 23724
rect 1355 23684 1400 23712
rect 1394 23672 1400 23684
rect 1452 23672 1458 23724
rect 4172 23712 4200 23808
rect 8864 23780 8892 23811
rect 9398 23808 9404 23820
rect 9456 23808 9462 23860
rect 10042 23848 10048 23860
rect 10003 23820 10048 23848
rect 10042 23808 10048 23820
rect 10100 23808 10106 23860
rect 12710 23848 12716 23860
rect 12671 23820 12716 23848
rect 12710 23808 12716 23820
rect 12768 23808 12774 23860
rect 16482 23848 16488 23860
rect 16443 23820 16488 23848
rect 16482 23808 16488 23820
rect 16540 23808 16546 23860
rect 21450 23848 21456 23860
rect 21411 23820 21456 23848
rect 21450 23808 21456 23820
rect 21508 23808 21514 23860
rect 23106 23848 23112 23860
rect 23067 23820 23112 23848
rect 23106 23808 23112 23820
rect 23164 23808 23170 23860
rect 24029 23851 24087 23857
rect 24029 23817 24041 23851
rect 24075 23848 24087 23851
rect 25406 23848 25412 23860
rect 24075 23820 25412 23848
rect 24075 23817 24087 23820
rect 24029 23811 24087 23817
rect 9769 23783 9827 23789
rect 9769 23780 9781 23783
rect 8864 23752 9781 23780
rect 9769 23749 9781 23752
rect 9815 23780 9827 23783
rect 16301 23783 16359 23789
rect 9815 23752 10640 23780
rect 9815 23749 9827 23752
rect 9769 23743 9827 23749
rect 10612 23721 10640 23752
rect 16301 23749 16313 23783
rect 16347 23780 16359 23783
rect 17494 23780 17500 23792
rect 16347 23752 17500 23780
rect 16347 23749 16359 23752
rect 16301 23743 16359 23749
rect 17494 23740 17500 23752
rect 17552 23740 17558 23792
rect 18141 23783 18199 23789
rect 18141 23749 18153 23783
rect 18187 23749 18199 23783
rect 18141 23743 18199 23749
rect 4249 23715 4307 23721
rect 4249 23712 4261 23715
rect 4172 23684 4261 23712
rect 4249 23681 4261 23684
rect 4295 23681 4307 23715
rect 4249 23675 4307 23681
rect 10597 23715 10655 23721
rect 10597 23681 10609 23715
rect 10643 23681 10655 23715
rect 10597 23675 10655 23681
rect 4522 23653 4528 23656
rect 4516 23644 4528 23653
rect 4483 23616 4528 23644
rect 4516 23607 4528 23616
rect 4522 23604 4528 23607
rect 4580 23604 4586 23656
rect 7466 23644 7472 23656
rect 7427 23616 7472 23644
rect 7466 23604 7472 23616
rect 7524 23604 7530 23656
rect 9398 23604 9404 23656
rect 9456 23644 9462 23656
rect 9456 23616 10548 23644
rect 9456 23604 9462 23616
rect 1578 23536 1584 23588
rect 1636 23585 1642 23588
rect 1636 23579 1700 23585
rect 1636 23545 1654 23579
rect 1688 23545 1700 23579
rect 1636 23539 1700 23545
rect 3789 23579 3847 23585
rect 3789 23545 3801 23579
rect 3835 23576 3847 23579
rect 4338 23576 4344 23588
rect 3835 23548 4344 23576
rect 3835 23545 3847 23548
rect 3789 23539 3847 23545
rect 1636 23536 1642 23539
rect 4338 23536 4344 23548
rect 4396 23536 4402 23588
rect 5166 23536 5172 23588
rect 5224 23576 5230 23588
rect 6641 23579 6699 23585
rect 5224 23548 5856 23576
rect 5224 23536 5230 23548
rect 5828 23520 5856 23548
rect 6641 23545 6653 23579
rect 6687 23576 6699 23579
rect 7098 23576 7104 23588
rect 6687 23548 7104 23576
rect 6687 23545 6699 23548
rect 6641 23539 6699 23545
rect 7098 23536 7104 23548
rect 7156 23576 7162 23588
rect 7736 23579 7794 23585
rect 7736 23576 7748 23579
rect 7156 23548 7748 23576
rect 7156 23536 7162 23548
rect 7736 23545 7748 23548
rect 7782 23576 7794 23579
rect 7926 23576 7932 23588
rect 7782 23548 7932 23576
rect 7782 23545 7794 23548
rect 7736 23539 7794 23545
rect 7926 23536 7932 23548
rect 7984 23536 7990 23588
rect 10042 23536 10048 23588
rect 10100 23576 10106 23588
rect 10520 23585 10548 23616
rect 10870 23604 10876 23656
rect 10928 23644 10934 23656
rect 11054 23644 11060 23656
rect 10928 23616 11060 23644
rect 10928 23604 10934 23616
rect 11054 23604 11060 23616
rect 11112 23644 11118 23656
rect 11149 23647 11207 23653
rect 11149 23644 11161 23647
rect 11112 23616 11161 23644
rect 11112 23604 11118 23616
rect 11149 23613 11161 23616
rect 11195 23644 11207 23647
rect 11882 23644 11888 23656
rect 11195 23616 11888 23644
rect 11195 23613 11207 23616
rect 11149 23607 11207 23613
rect 11882 23604 11888 23616
rect 11940 23604 11946 23656
rect 12158 23644 12164 23656
rect 12119 23616 12164 23644
rect 12158 23604 12164 23616
rect 12216 23644 12222 23656
rect 12529 23647 12587 23653
rect 12529 23644 12541 23647
rect 12216 23616 12541 23644
rect 12216 23604 12222 23616
rect 12529 23613 12541 23616
rect 12575 23613 12587 23647
rect 13633 23647 13691 23653
rect 13633 23644 13645 23647
rect 12529 23607 12587 23613
rect 13096 23616 13645 23644
rect 10321 23579 10379 23585
rect 10321 23576 10333 23579
rect 10100 23548 10333 23576
rect 10100 23536 10106 23548
rect 10321 23545 10333 23548
rect 10367 23545 10379 23579
rect 10321 23539 10379 23545
rect 10505 23579 10563 23585
rect 10505 23545 10517 23579
rect 10551 23545 10563 23579
rect 10505 23539 10563 23545
rect 2774 23468 2780 23520
rect 2832 23508 2838 23520
rect 3418 23508 3424 23520
rect 2832 23480 2877 23508
rect 3379 23480 3424 23508
rect 2832 23468 2838 23480
rect 3418 23468 3424 23480
rect 3476 23468 3482 23520
rect 4706 23468 4712 23520
rect 4764 23508 4770 23520
rect 5626 23508 5632 23520
rect 4764 23480 5632 23508
rect 4764 23468 4770 23480
rect 5626 23468 5632 23480
rect 5684 23468 5690 23520
rect 5810 23468 5816 23520
rect 5868 23508 5874 23520
rect 6181 23511 6239 23517
rect 6181 23508 6193 23511
rect 5868 23480 6193 23508
rect 5868 23468 5874 23480
rect 6181 23477 6193 23480
rect 6227 23477 6239 23511
rect 11514 23508 11520 23520
rect 11475 23480 11520 23508
rect 6181 23471 6239 23477
rect 11514 23468 11520 23480
rect 11572 23468 11578 23520
rect 11882 23468 11888 23520
rect 11940 23508 11946 23520
rect 13096 23517 13124 23616
rect 13633 23613 13645 23616
rect 13679 23613 13691 23647
rect 13633 23607 13691 23613
rect 15933 23647 15991 23653
rect 15933 23613 15945 23647
rect 15979 23644 15991 23647
rect 16298 23644 16304 23656
rect 15979 23616 16304 23644
rect 15979 23613 15991 23616
rect 15933 23607 15991 23613
rect 16298 23604 16304 23616
rect 16356 23644 16362 23656
rect 16356 23616 16988 23644
rect 16356 23604 16362 23616
rect 13906 23585 13912 23588
rect 13900 23576 13912 23585
rect 13867 23548 13912 23576
rect 13900 23539 13912 23548
rect 13906 23536 13912 23539
rect 13964 23536 13970 23588
rect 15470 23576 15476 23588
rect 14200 23548 15476 23576
rect 13081 23511 13139 23517
rect 13081 23508 13093 23511
rect 11940 23480 13093 23508
rect 11940 23468 11946 23480
rect 13081 23477 13093 23480
rect 13127 23477 13139 23511
rect 13081 23471 13139 23477
rect 13541 23511 13599 23517
rect 13541 23477 13553 23511
rect 13587 23508 13599 23511
rect 13814 23508 13820 23520
rect 13587 23480 13820 23508
rect 13587 23477 13599 23480
rect 13541 23471 13599 23477
rect 13814 23468 13820 23480
rect 13872 23508 13878 23520
rect 14200 23508 14228 23548
rect 15470 23536 15476 23548
rect 15528 23536 15534 23588
rect 16666 23536 16672 23588
rect 16724 23576 16730 23588
rect 16960 23585 16988 23616
rect 17494 23604 17500 23656
rect 17552 23644 17558 23656
rect 18156 23644 18184 23743
rect 18874 23740 18880 23792
rect 18932 23780 18938 23792
rect 19153 23783 19211 23789
rect 19153 23780 19165 23783
rect 18932 23752 19165 23780
rect 18932 23740 18938 23752
rect 19153 23749 19165 23752
rect 19199 23780 19211 23783
rect 20073 23783 20131 23789
rect 20073 23780 20085 23783
rect 19199 23752 20085 23780
rect 19199 23749 19211 23752
rect 19153 23743 19211 23749
rect 20073 23749 20085 23752
rect 20119 23749 20131 23783
rect 20073 23743 20131 23749
rect 19521 23715 19579 23721
rect 19521 23681 19533 23715
rect 19567 23712 19579 23715
rect 20530 23712 20536 23724
rect 19567 23684 20536 23712
rect 19567 23681 19579 23684
rect 19521 23675 19579 23681
rect 20530 23672 20536 23684
rect 20588 23672 20594 23724
rect 21468 23712 21496 23808
rect 22097 23783 22155 23789
rect 22097 23749 22109 23783
rect 22143 23780 22155 23783
rect 23014 23780 23020 23792
rect 22143 23752 23020 23780
rect 22143 23749 22155 23752
rect 22097 23743 22155 23749
rect 23014 23740 23020 23752
rect 23072 23740 23078 23792
rect 24136 23721 24164 23820
rect 25406 23808 25412 23820
rect 25464 23848 25470 23860
rect 27614 23848 27620 23860
rect 25464 23820 27620 23848
rect 25464 23808 25470 23820
rect 27614 23808 27620 23820
rect 27672 23808 27678 23860
rect 22465 23715 22523 23721
rect 22465 23712 22477 23715
rect 21468 23684 22477 23712
rect 22465 23681 22477 23684
rect 22511 23681 22523 23715
rect 22465 23675 22523 23681
rect 24121 23715 24179 23721
rect 24121 23681 24133 23715
rect 24167 23681 24179 23715
rect 24121 23675 24179 23681
rect 21818 23644 21824 23656
rect 17552 23616 18184 23644
rect 21779 23616 21824 23644
rect 17552 23604 17558 23616
rect 21818 23604 21824 23616
rect 21876 23604 21882 23656
rect 16761 23579 16819 23585
rect 16761 23576 16773 23579
rect 16724 23548 16773 23576
rect 16724 23536 16730 23548
rect 16761 23545 16773 23548
rect 16807 23545 16819 23579
rect 16761 23539 16819 23545
rect 16945 23579 17003 23585
rect 16945 23545 16957 23579
rect 16991 23545 17003 23579
rect 16945 23539 17003 23545
rect 17037 23579 17095 23585
rect 17037 23545 17049 23579
rect 17083 23576 17095 23579
rect 17126 23576 17132 23588
rect 17083 23548 17132 23576
rect 17083 23545 17095 23548
rect 17037 23539 17095 23545
rect 17126 23536 17132 23548
rect 17184 23576 17190 23588
rect 17770 23576 17776 23588
rect 17184 23548 17776 23576
rect 17184 23536 17190 23548
rect 17770 23536 17776 23548
rect 17828 23536 17834 23588
rect 17865 23579 17923 23585
rect 17865 23545 17877 23579
rect 17911 23576 17923 23579
rect 18414 23576 18420 23588
rect 17911 23548 18420 23576
rect 17911 23545 17923 23548
rect 17865 23539 17923 23545
rect 18414 23536 18420 23548
rect 18472 23536 18478 23588
rect 18506 23536 18512 23588
rect 18564 23576 18570 23588
rect 18693 23579 18751 23585
rect 18693 23576 18705 23579
rect 18564 23548 18705 23576
rect 18564 23536 18570 23548
rect 18693 23545 18705 23548
rect 18739 23545 18751 23579
rect 18693 23539 18751 23545
rect 20346 23536 20352 23588
rect 20404 23576 20410 23588
rect 20625 23579 20683 23585
rect 20625 23576 20637 23579
rect 20404 23548 20637 23576
rect 20404 23536 20410 23548
rect 20625 23545 20637 23548
rect 20671 23545 20683 23579
rect 20625 23539 20683 23545
rect 21177 23579 21235 23585
rect 21177 23545 21189 23579
rect 21223 23576 21235 23579
rect 22002 23576 22008 23588
rect 21223 23548 22008 23576
rect 21223 23545 21235 23548
rect 21177 23539 21235 23545
rect 22002 23536 22008 23548
rect 22060 23576 22066 23588
rect 22649 23579 22707 23585
rect 22649 23576 22661 23579
rect 22060 23548 22661 23576
rect 22060 23536 22066 23548
rect 22649 23545 22661 23548
rect 22695 23576 22707 23579
rect 22922 23576 22928 23588
rect 22695 23548 22928 23576
rect 22695 23545 22707 23548
rect 22649 23539 22707 23545
rect 22922 23536 22928 23548
rect 22980 23576 22986 23588
rect 24366 23579 24424 23585
rect 24366 23576 24378 23579
rect 22980 23548 24378 23576
rect 22980 23536 22986 23548
rect 24366 23545 24378 23548
rect 24412 23545 24424 23579
rect 24366 23539 24424 23545
rect 13872 23480 14228 23508
rect 13872 23468 13878 23480
rect 14274 23468 14280 23520
rect 14332 23508 14338 23520
rect 15013 23511 15071 23517
rect 15013 23508 15025 23511
rect 14332 23480 15025 23508
rect 14332 23468 14338 23480
rect 15013 23477 15025 23480
rect 15059 23477 15071 23511
rect 15013 23471 15071 23477
rect 17497 23511 17555 23517
rect 17497 23477 17509 23511
rect 17543 23508 17555 23511
rect 17586 23508 17592 23520
rect 17543 23480 17592 23508
rect 17543 23477 17555 23480
rect 17497 23471 17555 23477
rect 17586 23468 17592 23480
rect 17644 23468 17650 23520
rect 18138 23468 18144 23520
rect 18196 23508 18202 23520
rect 18601 23511 18659 23517
rect 18601 23508 18613 23511
rect 18196 23480 18613 23508
rect 18196 23468 18202 23480
rect 18601 23477 18613 23480
rect 18647 23477 18659 23511
rect 18601 23471 18659 23477
rect 19889 23511 19947 23517
rect 19889 23477 19901 23511
rect 19935 23508 19947 23511
rect 19978 23508 19984 23520
rect 19935 23480 19984 23508
rect 19935 23477 19947 23480
rect 19889 23471 19947 23477
rect 19978 23468 19984 23480
rect 20036 23508 20042 23520
rect 20533 23511 20591 23517
rect 20533 23508 20545 23511
rect 20036 23480 20545 23508
rect 20036 23468 20042 23480
rect 20533 23477 20545 23480
rect 20579 23477 20591 23511
rect 20533 23471 20591 23477
rect 21818 23468 21824 23520
rect 21876 23508 21882 23520
rect 22557 23511 22615 23517
rect 22557 23508 22569 23511
rect 21876 23480 22569 23508
rect 21876 23468 21882 23480
rect 22557 23477 22569 23480
rect 22603 23477 22615 23511
rect 22557 23471 22615 23477
rect 25038 23468 25044 23520
rect 25096 23508 25102 23520
rect 25501 23511 25559 23517
rect 25501 23508 25513 23511
rect 25096 23480 25513 23508
rect 25096 23468 25102 23480
rect 25501 23477 25513 23480
rect 25547 23477 25559 23511
rect 25501 23471 25559 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 2869 23307 2927 23313
rect 2869 23273 2881 23307
rect 2915 23304 2927 23307
rect 3418 23304 3424 23316
rect 2915 23276 3424 23304
rect 2915 23273 2927 23276
rect 2869 23267 2927 23273
rect 3418 23264 3424 23276
rect 3476 23264 3482 23316
rect 4154 23264 4160 23316
rect 4212 23304 4218 23316
rect 4249 23307 4307 23313
rect 4249 23304 4261 23307
rect 4212 23276 4261 23304
rect 4212 23264 4218 23276
rect 4249 23273 4261 23276
rect 4295 23273 4307 23307
rect 5810 23304 5816 23316
rect 5771 23276 5816 23304
rect 4249 23267 4307 23273
rect 1756 23239 1814 23245
rect 1756 23205 1768 23239
rect 1802 23236 1814 23239
rect 1854 23236 1860 23248
rect 1802 23208 1860 23236
rect 1802 23205 1814 23208
rect 1756 23199 1814 23205
rect 1854 23196 1860 23208
rect 1912 23196 1918 23248
rect 1394 23128 1400 23180
rect 1452 23168 1458 23180
rect 1489 23171 1547 23177
rect 1489 23168 1501 23171
rect 1452 23140 1501 23168
rect 1452 23128 1458 23140
rect 1489 23137 1501 23140
rect 1535 23137 1547 23171
rect 3510 23168 3516 23180
rect 3471 23140 3516 23168
rect 1489 23131 1547 23137
rect 3510 23128 3516 23140
rect 3568 23128 3574 23180
rect 4264 23168 4292 23267
rect 5810 23264 5816 23276
rect 5868 23264 5874 23316
rect 6917 23307 6975 23313
rect 6917 23273 6929 23307
rect 6963 23304 6975 23307
rect 7742 23304 7748 23316
rect 6963 23276 7748 23304
rect 6963 23273 6975 23276
rect 6917 23267 6975 23273
rect 7742 23264 7748 23276
rect 7800 23264 7806 23316
rect 12802 23264 12808 23316
rect 12860 23304 12866 23316
rect 16206 23304 16212 23316
rect 12860 23276 16212 23304
rect 12860 23264 12866 23276
rect 16206 23264 16212 23276
rect 16264 23264 16270 23316
rect 16666 23304 16672 23316
rect 16627 23276 16672 23304
rect 16666 23264 16672 23276
rect 16724 23264 16730 23316
rect 23201 23307 23259 23313
rect 23201 23273 23213 23307
rect 23247 23304 23259 23307
rect 23566 23304 23572 23316
rect 23247 23276 23572 23304
rect 23247 23273 23259 23276
rect 23201 23267 23259 23273
rect 23400 23248 23428 23276
rect 23566 23264 23572 23276
rect 23624 23264 23630 23316
rect 24857 23307 24915 23313
rect 24857 23273 24869 23307
rect 24903 23304 24915 23307
rect 24946 23304 24952 23316
rect 24903 23276 24952 23304
rect 24903 23273 24915 23276
rect 24857 23267 24915 23273
rect 24946 23264 24952 23276
rect 25004 23264 25010 23316
rect 4706 23245 4712 23248
rect 4700 23236 4712 23245
rect 4667 23208 4712 23236
rect 4700 23199 4712 23208
rect 4706 23196 4712 23199
rect 4764 23196 4770 23248
rect 7006 23236 7012 23248
rect 6967 23208 7012 23236
rect 7006 23196 7012 23208
rect 7064 23196 7070 23248
rect 7466 23236 7472 23248
rect 7427 23208 7472 23236
rect 7466 23196 7472 23208
rect 7524 23196 7530 23248
rect 8110 23196 8116 23248
rect 8168 23236 8174 23248
rect 8389 23239 8447 23245
rect 8389 23236 8401 23239
rect 8168 23208 8401 23236
rect 8168 23196 8174 23208
rect 8389 23205 8401 23208
rect 8435 23205 8447 23239
rect 8570 23236 8576 23248
rect 8531 23208 8576 23236
rect 8389 23199 8447 23205
rect 8570 23196 8576 23208
rect 8628 23196 8634 23248
rect 9490 23236 9496 23248
rect 9451 23208 9496 23236
rect 9490 23196 9496 23208
rect 9548 23196 9554 23248
rect 11146 23245 11152 23248
rect 11140 23236 11152 23245
rect 11059 23208 11152 23236
rect 11140 23199 11152 23208
rect 11204 23236 11210 23248
rect 11606 23236 11612 23248
rect 11204 23208 11612 23236
rect 11146 23196 11152 23199
rect 11204 23196 11210 23208
rect 11606 23196 11612 23208
rect 11664 23196 11670 23248
rect 13814 23196 13820 23248
rect 13872 23236 13878 23248
rect 14001 23239 14059 23245
rect 14001 23236 14013 23239
rect 13872 23208 14013 23236
rect 13872 23196 13878 23208
rect 14001 23205 14013 23208
rect 14047 23205 14059 23239
rect 14182 23236 14188 23248
rect 14143 23208 14188 23236
rect 14001 23199 14059 23205
rect 14182 23196 14188 23208
rect 14240 23236 14246 23248
rect 14645 23239 14703 23245
rect 14645 23236 14657 23239
rect 14240 23208 14657 23236
rect 14240 23196 14246 23208
rect 14645 23205 14657 23208
rect 14691 23205 14703 23239
rect 15746 23236 15752 23248
rect 15707 23208 15752 23236
rect 14645 23199 14703 23205
rect 15746 23196 15752 23208
rect 15804 23196 15810 23248
rect 17218 23196 17224 23248
rect 17276 23236 17282 23248
rect 17313 23239 17371 23245
rect 17313 23236 17325 23239
rect 17276 23208 17325 23236
rect 17276 23196 17282 23208
rect 17313 23205 17325 23208
rect 17359 23205 17371 23239
rect 19794 23236 19800 23248
rect 19755 23208 19800 23236
rect 17313 23199 17371 23205
rect 19794 23196 19800 23208
rect 19852 23196 19858 23248
rect 20346 23196 20352 23248
rect 20404 23236 20410 23248
rect 21146 23239 21204 23245
rect 21146 23236 21158 23239
rect 20404 23208 21158 23236
rect 20404 23196 20410 23208
rect 21146 23205 21158 23208
rect 21192 23236 21204 23239
rect 22278 23236 22284 23248
rect 21192 23208 22284 23236
rect 21192 23205 21204 23208
rect 21146 23199 21204 23205
rect 22278 23196 22284 23208
rect 22336 23196 22342 23248
rect 23382 23196 23388 23248
rect 23440 23196 23446 23248
rect 23474 23196 23480 23248
rect 23532 23236 23538 23248
rect 23753 23239 23811 23245
rect 23753 23236 23765 23239
rect 23532 23208 23765 23236
rect 23532 23196 23538 23208
rect 23753 23205 23765 23208
rect 23799 23205 23811 23239
rect 23753 23199 23811 23205
rect 23937 23239 23995 23245
rect 23937 23205 23949 23239
rect 23983 23205 23995 23239
rect 23937 23199 23995 23205
rect 25225 23239 25283 23245
rect 25225 23205 25237 23239
rect 25271 23236 25283 23239
rect 25682 23236 25688 23248
rect 25271 23208 25688 23236
rect 25271 23205 25283 23208
rect 25225 23199 25283 23205
rect 4433 23171 4491 23177
rect 4433 23168 4445 23171
rect 4264 23140 4445 23168
rect 4433 23137 4445 23140
rect 4479 23137 4491 23171
rect 7926 23168 7932 23180
rect 7839 23140 7932 23168
rect 4433 23131 4491 23137
rect 7926 23128 7932 23140
rect 7984 23168 7990 23180
rect 7984 23140 8708 23168
rect 7984 23128 7990 23140
rect 8680 23112 8708 23140
rect 10594 23128 10600 23180
rect 10652 23168 10658 23180
rect 10870 23168 10876 23180
rect 10652 23140 10876 23168
rect 10652 23128 10658 23140
rect 10870 23128 10876 23140
rect 10928 23128 10934 23180
rect 14274 23168 14280 23180
rect 14235 23140 14280 23168
rect 14274 23128 14280 23140
rect 14332 23128 14338 23180
rect 15473 23171 15531 23177
rect 15473 23168 15485 23171
rect 15028 23140 15485 23168
rect 8662 23100 8668 23112
rect 8623 23072 8668 23100
rect 8662 23060 8668 23072
rect 8720 23060 8726 23112
rect 9582 23060 9588 23112
rect 9640 23100 9646 23112
rect 9677 23103 9735 23109
rect 9677 23100 9689 23103
rect 9640 23072 9689 23100
rect 9640 23060 9646 23072
rect 9677 23069 9689 23072
rect 9723 23069 9735 23103
rect 13538 23100 13544 23112
rect 13451 23072 13544 23100
rect 9677 23063 9735 23069
rect 13538 23060 13544 23072
rect 13596 23100 13602 23112
rect 13998 23100 14004 23112
rect 13596 23072 14004 23100
rect 13596 23060 13602 23072
rect 13998 23060 14004 23072
rect 14056 23060 14062 23112
rect 8113 23035 8171 23041
rect 8113 23001 8125 23035
rect 8159 23032 8171 23035
rect 10042 23032 10048 23044
rect 8159 23004 10048 23032
rect 8159 23001 8171 23004
rect 8113 22995 8171 23001
rect 10042 22992 10048 23004
rect 10100 23032 10106 23044
rect 10137 23035 10195 23041
rect 10137 23032 10149 23035
rect 10100 23004 10149 23032
rect 10100 22992 10106 23004
rect 10137 23001 10149 23004
rect 10183 23001 10195 23035
rect 13722 23032 13728 23044
rect 13683 23004 13728 23032
rect 10137 22995 10195 23001
rect 13722 22992 13728 23004
rect 13780 22992 13786 23044
rect 3786 22964 3792 22976
rect 3747 22936 3792 22964
rect 3786 22924 3792 22936
rect 3844 22924 3850 22976
rect 10597 22967 10655 22973
rect 10597 22933 10609 22967
rect 10643 22964 10655 22967
rect 10870 22964 10876 22976
rect 10643 22936 10876 22964
rect 10643 22933 10655 22936
rect 10597 22927 10655 22933
rect 10870 22924 10876 22936
rect 10928 22924 10934 22976
rect 12158 22924 12164 22976
rect 12216 22964 12222 22976
rect 12253 22967 12311 22973
rect 12253 22964 12265 22967
rect 12216 22936 12265 22964
rect 12216 22924 12222 22936
rect 12253 22933 12265 22936
rect 12299 22933 12311 22967
rect 12253 22927 12311 22933
rect 13173 22967 13231 22973
rect 13173 22933 13185 22967
rect 13219 22964 13231 22967
rect 13262 22964 13268 22976
rect 13219 22936 13268 22964
rect 13219 22933 13231 22936
rect 13173 22927 13231 22933
rect 13262 22924 13268 22936
rect 13320 22924 13326 22976
rect 14826 22924 14832 22976
rect 14884 22964 14890 22976
rect 15028 22973 15056 23140
rect 15473 23137 15485 23140
rect 15519 23137 15531 23171
rect 15473 23131 15531 23137
rect 17129 23171 17187 23177
rect 17129 23137 17141 23171
rect 17175 23168 17187 23171
rect 17678 23168 17684 23180
rect 17175 23140 17684 23168
rect 17175 23137 17187 23140
rect 17129 23131 17187 23137
rect 17678 23128 17684 23140
rect 17736 23128 17742 23180
rect 20901 23171 20959 23177
rect 20901 23137 20913 23171
rect 20947 23168 20959 23171
rect 21542 23168 21548 23180
rect 20947 23140 21548 23168
rect 20947 23137 20959 23140
rect 20901 23131 20959 23137
rect 21542 23128 21548 23140
rect 21600 23128 21606 23180
rect 23014 23128 23020 23180
rect 23072 23168 23078 23180
rect 23952 23168 23980 23199
rect 25682 23196 25688 23208
rect 25740 23196 25746 23248
rect 24946 23168 24952 23180
rect 23072 23140 23980 23168
rect 24907 23140 24952 23168
rect 23072 23128 23078 23140
rect 24946 23128 24952 23140
rect 25004 23128 25010 23180
rect 17402 23100 17408 23112
rect 17363 23072 17408 23100
rect 17402 23060 17408 23072
rect 17460 23060 17466 23112
rect 19797 23103 19855 23109
rect 19797 23069 19809 23103
rect 19843 23069 19855 23103
rect 19797 23063 19855 23069
rect 19889 23103 19947 23109
rect 19889 23069 19901 23103
rect 19935 23100 19947 23103
rect 20070 23100 20076 23112
rect 19935 23072 20076 23100
rect 19935 23069 19947 23072
rect 19889 23063 19947 23069
rect 16666 22992 16672 23044
rect 16724 23032 16730 23044
rect 16853 23035 16911 23041
rect 16853 23032 16865 23035
rect 16724 23004 16865 23032
rect 16724 22992 16730 23004
rect 16853 23001 16865 23004
rect 16899 23001 16911 23035
rect 19812 23032 19840 23063
rect 20070 23060 20076 23072
rect 20128 23060 20134 23112
rect 24026 23100 24032 23112
rect 23987 23072 24032 23100
rect 24026 23060 24032 23072
rect 24084 23060 24090 23112
rect 19978 23032 19984 23044
rect 19812 23004 19984 23032
rect 16853 22995 16911 23001
rect 19978 22992 19984 23004
rect 20036 22992 20042 23044
rect 15013 22967 15071 22973
rect 15013 22964 15025 22967
rect 14884 22936 15025 22964
rect 14884 22924 14890 22936
rect 15013 22933 15025 22936
rect 15059 22933 15071 22967
rect 18138 22964 18144 22976
rect 18099 22936 18144 22964
rect 15013 22927 15071 22933
rect 18138 22924 18144 22936
rect 18196 22924 18202 22976
rect 18785 22967 18843 22973
rect 18785 22933 18797 22967
rect 18831 22964 18843 22967
rect 18966 22964 18972 22976
rect 18831 22936 18972 22964
rect 18831 22933 18843 22936
rect 18785 22927 18843 22933
rect 18966 22924 18972 22936
rect 19024 22924 19030 22976
rect 19150 22964 19156 22976
rect 19111 22936 19156 22964
rect 19150 22924 19156 22936
rect 19208 22924 19214 22976
rect 19334 22964 19340 22976
rect 19295 22936 19340 22964
rect 19334 22924 19340 22936
rect 19392 22924 19398 22976
rect 20349 22967 20407 22973
rect 20349 22933 20361 22967
rect 20395 22964 20407 22967
rect 20530 22964 20536 22976
rect 20395 22936 20536 22964
rect 20395 22933 20407 22936
rect 20349 22927 20407 22933
rect 20530 22924 20536 22936
rect 20588 22964 20594 22976
rect 22281 22967 22339 22973
rect 22281 22964 22293 22967
rect 20588 22936 22293 22964
rect 20588 22924 20594 22936
rect 22281 22933 22293 22936
rect 22327 22933 22339 22967
rect 22281 22927 22339 22933
rect 23477 22967 23535 22973
rect 23477 22933 23489 22967
rect 23523 22964 23535 22967
rect 23566 22964 23572 22976
rect 23523 22936 23572 22964
rect 23523 22933 23535 22936
rect 23477 22927 23535 22933
rect 23566 22924 23572 22936
rect 23624 22924 23630 22976
rect 24210 22924 24216 22976
rect 24268 22964 24274 22976
rect 24397 22967 24455 22973
rect 24397 22964 24409 22967
rect 24268 22936 24409 22964
rect 24268 22924 24274 22936
rect 24397 22933 24409 22936
rect 24443 22933 24455 22967
rect 24397 22927 24455 22933
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1489 22763 1547 22769
rect 1489 22729 1501 22763
rect 1535 22760 1547 22763
rect 2038 22760 2044 22772
rect 1535 22732 2044 22760
rect 1535 22729 1547 22732
rect 1489 22723 1547 22729
rect 2038 22720 2044 22732
rect 2096 22720 2102 22772
rect 4154 22760 4160 22772
rect 4115 22732 4160 22760
rect 4154 22720 4160 22732
rect 4212 22720 4218 22772
rect 4433 22763 4491 22769
rect 4433 22729 4445 22763
rect 4479 22760 4491 22763
rect 5074 22760 5080 22772
rect 4479 22732 5080 22760
rect 4479 22729 4491 22732
rect 4433 22723 4491 22729
rect 5074 22720 5080 22732
rect 5132 22720 5138 22772
rect 5442 22760 5448 22772
rect 5403 22732 5448 22760
rect 5442 22720 5448 22732
rect 5500 22720 5506 22772
rect 5534 22720 5540 22772
rect 5592 22760 5598 22772
rect 5721 22763 5779 22769
rect 5721 22760 5733 22763
rect 5592 22732 5733 22760
rect 5592 22720 5598 22732
rect 5721 22729 5733 22732
rect 5767 22729 5779 22763
rect 5721 22723 5779 22729
rect 7745 22763 7803 22769
rect 7745 22729 7757 22763
rect 7791 22760 7803 22763
rect 8570 22760 8576 22772
rect 7791 22732 8576 22760
rect 7791 22729 7803 22732
rect 7745 22723 7803 22729
rect 8570 22720 8576 22732
rect 8628 22720 8634 22772
rect 8846 22720 8852 22772
rect 8904 22760 8910 22772
rect 9585 22763 9643 22769
rect 9585 22760 9597 22763
rect 8904 22732 9597 22760
rect 8904 22720 8910 22732
rect 9585 22729 9597 22732
rect 9631 22729 9643 22763
rect 9585 22723 9643 22729
rect 9950 22720 9956 22772
rect 10008 22760 10014 22772
rect 10229 22763 10287 22769
rect 10229 22760 10241 22763
rect 10008 22732 10241 22760
rect 10008 22720 10014 22732
rect 10229 22729 10241 22732
rect 10275 22729 10287 22763
rect 10594 22760 10600 22772
rect 10555 22732 10600 22760
rect 10229 22723 10287 22729
rect 566 22652 572 22704
rect 624 22692 630 22704
rect 5261 22695 5319 22701
rect 5261 22692 5273 22695
rect 624 22664 5273 22692
rect 624 22652 630 22664
rect 5261 22661 5273 22664
rect 5307 22661 5319 22695
rect 5261 22655 5319 22661
rect 1394 22584 1400 22636
rect 1452 22624 1458 22636
rect 2866 22624 2872 22636
rect 1452 22596 2872 22624
rect 1452 22584 1458 22596
rect 2866 22584 2872 22596
rect 2924 22584 2930 22636
rect 3234 22624 3240 22636
rect 3195 22596 3240 22624
rect 3234 22584 3240 22596
rect 3292 22584 3298 22636
rect 4893 22627 4951 22633
rect 4893 22593 4905 22627
rect 4939 22624 4951 22627
rect 5460 22624 5488 22720
rect 8110 22692 8116 22704
rect 8071 22664 8116 22692
rect 8110 22652 8116 22664
rect 8168 22652 8174 22704
rect 4939 22596 5488 22624
rect 4939 22593 4951 22596
rect 4893 22587 4951 22593
rect 7466 22584 7472 22636
rect 7524 22624 7530 22636
rect 8205 22627 8263 22633
rect 8205 22624 8217 22627
rect 7524 22596 8217 22624
rect 7524 22584 7530 22596
rect 8205 22593 8217 22596
rect 8251 22593 8263 22627
rect 8205 22587 8263 22593
rect 1762 22556 1768 22568
rect 1723 22528 1768 22556
rect 1762 22516 1768 22528
rect 1820 22556 1826 22568
rect 2409 22559 2467 22565
rect 2409 22556 2421 22559
rect 1820 22528 2421 22556
rect 1820 22516 1826 22528
rect 2409 22525 2421 22528
rect 2455 22525 2467 22559
rect 2958 22556 2964 22568
rect 2871 22528 2964 22556
rect 2409 22519 2467 22525
rect 2958 22516 2964 22528
rect 3016 22556 3022 22568
rect 3786 22556 3792 22568
rect 3016 22528 3792 22556
rect 3016 22516 3022 22528
rect 3786 22516 3792 22528
rect 3844 22516 3850 22568
rect 4985 22559 5043 22565
rect 4985 22525 4997 22559
rect 5031 22556 5043 22559
rect 5166 22556 5172 22568
rect 5031 22528 5172 22556
rect 5031 22525 5043 22528
rect 4985 22519 5043 22525
rect 5166 22516 5172 22528
rect 5224 22516 5230 22568
rect 5261 22559 5319 22565
rect 5261 22525 5273 22559
rect 5307 22556 5319 22559
rect 5442 22556 5448 22568
rect 5307 22528 5448 22556
rect 5307 22525 5319 22528
rect 5261 22519 5319 22525
rect 5442 22516 5448 22528
rect 5500 22516 5506 22568
rect 6178 22516 6184 22568
rect 6236 22556 6242 22568
rect 6457 22559 6515 22565
rect 6457 22556 6469 22559
rect 6236 22528 6469 22556
rect 6236 22516 6242 22528
rect 6457 22525 6469 22528
rect 6503 22525 6515 22559
rect 6822 22556 6828 22568
rect 6783 22528 6828 22556
rect 6457 22519 6515 22525
rect 6822 22516 6828 22528
rect 6880 22516 6886 22568
rect 1854 22448 1860 22500
rect 1912 22488 1918 22500
rect 2041 22491 2099 22497
rect 2041 22488 2053 22491
rect 1912 22460 2053 22488
rect 1912 22448 1918 22460
rect 2041 22457 2053 22460
rect 2087 22488 2099 22491
rect 2087 22460 3188 22488
rect 2087 22457 2099 22460
rect 2041 22451 2099 22457
rect 1949 22423 2007 22429
rect 1949 22389 1961 22423
rect 1995 22420 2007 22423
rect 2130 22420 2136 22432
rect 1995 22392 2136 22420
rect 1995 22389 2007 22392
rect 1949 22383 2007 22389
rect 2130 22380 2136 22392
rect 2188 22420 2194 22432
rect 3050 22420 3056 22432
rect 2188 22392 3056 22420
rect 2188 22380 2194 22392
rect 3050 22380 3056 22392
rect 3108 22380 3114 22432
rect 3160 22420 3188 22460
rect 4338 22448 4344 22500
rect 4396 22488 4402 22500
rect 4893 22491 4951 22497
rect 4893 22488 4905 22491
rect 4396 22460 4905 22488
rect 4396 22448 4402 22460
rect 4893 22457 4905 22460
rect 4939 22457 4951 22491
rect 7098 22488 7104 22500
rect 7059 22460 7104 22488
rect 4893 22451 4951 22457
rect 7098 22448 7104 22460
rect 7156 22448 7162 22500
rect 8386 22448 8392 22500
rect 8444 22497 8450 22500
rect 8444 22491 8508 22497
rect 8444 22457 8462 22491
rect 8496 22457 8508 22491
rect 10244 22488 10272 22723
rect 10594 22720 10600 22732
rect 10652 22720 10658 22772
rect 10873 22763 10931 22769
rect 10873 22729 10885 22763
rect 10919 22760 10931 22763
rect 10962 22760 10968 22772
rect 10919 22732 10968 22760
rect 10919 22729 10931 22732
rect 10873 22723 10931 22729
rect 10962 22720 10968 22732
rect 11020 22720 11026 22772
rect 14093 22763 14151 22769
rect 14093 22729 14105 22763
rect 14139 22760 14151 22763
rect 14182 22760 14188 22772
rect 14139 22732 14188 22760
rect 14139 22729 14151 22732
rect 14093 22723 14151 22729
rect 14182 22720 14188 22732
rect 14240 22720 14246 22772
rect 16298 22760 16304 22772
rect 16259 22732 16304 22760
rect 16298 22720 16304 22732
rect 16356 22720 16362 22772
rect 17678 22760 17684 22772
rect 17639 22732 17684 22760
rect 17678 22720 17684 22732
rect 17736 22720 17742 22772
rect 18046 22720 18052 22772
rect 18104 22760 18110 22772
rect 18601 22763 18659 22769
rect 18601 22760 18613 22763
rect 18104 22732 18613 22760
rect 18104 22720 18110 22732
rect 18601 22729 18613 22732
rect 18647 22760 18659 22763
rect 21634 22760 21640 22772
rect 18647 22732 19564 22760
rect 21595 22732 21640 22760
rect 18647 22729 18659 22732
rect 18601 22723 18659 22729
rect 10612 22624 10640 22720
rect 11330 22652 11336 22704
rect 11388 22692 11394 22704
rect 12529 22695 12587 22701
rect 12529 22692 12541 22695
rect 11388 22664 12541 22692
rect 11388 22652 11394 22664
rect 12529 22661 12541 22664
rect 12575 22661 12587 22695
rect 12529 22655 12587 22661
rect 14734 22652 14740 22704
rect 14792 22692 14798 22704
rect 14918 22692 14924 22704
rect 14792 22664 14924 22692
rect 14792 22652 14798 22664
rect 14918 22652 14924 22664
rect 14976 22652 14982 22704
rect 18782 22692 18788 22704
rect 18743 22664 18788 22692
rect 18782 22652 18788 22664
rect 18840 22652 18846 22704
rect 19536 22692 19564 22732
rect 21634 22720 21640 22732
rect 21692 22720 21698 22772
rect 23014 22760 23020 22772
rect 22975 22732 23020 22760
rect 23014 22720 23020 22732
rect 23072 22720 23078 22772
rect 24946 22720 24952 22772
rect 25004 22760 25010 22772
rect 25314 22760 25320 22772
rect 25004 22732 25320 22760
rect 25004 22720 25010 22732
rect 25314 22720 25320 22732
rect 25372 22760 25378 22772
rect 25409 22763 25467 22769
rect 25409 22760 25421 22763
rect 25372 22732 25421 22760
rect 25372 22720 25378 22732
rect 25409 22729 25421 22732
rect 25455 22729 25467 22763
rect 25409 22723 25467 22729
rect 19794 22692 19800 22704
rect 19536 22664 19800 22692
rect 19794 22652 19800 22664
rect 19852 22652 19858 22704
rect 23750 22652 23756 22704
rect 23808 22692 23814 22704
rect 24121 22695 24179 22701
rect 24121 22692 24133 22695
rect 23808 22664 24133 22692
rect 23808 22652 23814 22664
rect 24121 22661 24133 22664
rect 24167 22661 24179 22695
rect 24121 22655 24179 22661
rect 10962 22624 10968 22636
rect 10612 22596 10968 22624
rect 10962 22584 10968 22596
rect 11020 22584 11026 22636
rect 12250 22584 12256 22636
rect 12308 22624 12314 22636
rect 12618 22624 12624 22636
rect 12308 22596 12624 22624
rect 12308 22584 12314 22596
rect 12618 22584 12624 22596
rect 12676 22584 12682 22636
rect 13262 22584 13268 22636
rect 13320 22624 13326 22636
rect 13722 22624 13728 22636
rect 13320 22596 13728 22624
rect 13320 22584 13326 22596
rect 13722 22584 13728 22596
rect 13780 22624 13786 22636
rect 13906 22624 13912 22636
rect 13780 22596 13912 22624
rect 13780 22584 13786 22596
rect 13906 22584 13912 22596
rect 13964 22624 13970 22636
rect 14645 22627 14703 22633
rect 14645 22624 14657 22627
rect 13964 22596 14657 22624
rect 13964 22584 13970 22596
rect 14645 22593 14657 22596
rect 14691 22624 14703 22627
rect 15013 22627 15071 22633
rect 15013 22624 15025 22627
rect 14691 22596 15025 22624
rect 14691 22593 14703 22596
rect 14645 22587 14703 22593
rect 15013 22593 15025 22596
rect 15059 22593 15071 22627
rect 15013 22587 15071 22593
rect 16117 22627 16175 22633
rect 16117 22593 16129 22627
rect 16163 22624 16175 22627
rect 16758 22624 16764 22636
rect 16163 22596 16764 22624
rect 16163 22593 16175 22596
rect 16117 22587 16175 22593
rect 16758 22584 16764 22596
rect 16816 22584 16822 22636
rect 16850 22584 16856 22636
rect 16908 22624 16914 22636
rect 17402 22624 17408 22636
rect 16908 22596 17408 22624
rect 16908 22584 16914 22596
rect 17402 22584 17408 22596
rect 17460 22584 17466 22636
rect 18966 22584 18972 22636
rect 19024 22624 19030 22636
rect 19337 22627 19395 22633
rect 19337 22624 19349 22627
rect 19024 22596 19349 22624
rect 19024 22584 19030 22596
rect 19337 22593 19349 22596
rect 19383 22624 19395 22627
rect 24581 22627 24639 22633
rect 19383 22596 20392 22624
rect 19383 22593 19395 22596
rect 19337 22587 19395 22593
rect 11054 22516 11060 22568
rect 11112 22556 11118 22568
rect 11149 22559 11207 22565
rect 11149 22556 11161 22559
rect 11112 22528 11161 22556
rect 11112 22516 11118 22528
rect 11149 22525 11161 22528
rect 11195 22525 11207 22559
rect 11149 22519 11207 22525
rect 12986 22516 12992 22568
rect 13044 22556 13050 22568
rect 13449 22559 13507 22565
rect 13449 22556 13461 22559
rect 13044 22528 13461 22556
rect 13044 22516 13050 22528
rect 13449 22525 13461 22528
rect 13495 22556 13507 22559
rect 13495 22528 14596 22556
rect 13495 22525 13507 22528
rect 13449 22519 13507 22525
rect 11425 22491 11483 22497
rect 11425 22488 11437 22491
rect 10244 22460 11437 22488
rect 8444 22451 8508 22457
rect 11425 22457 11437 22460
rect 11471 22488 11483 22491
rect 12158 22488 12164 22500
rect 11471 22460 12164 22488
rect 11471 22457 11483 22460
rect 11425 22451 11483 22457
rect 8444 22448 8450 22451
rect 12158 22448 12164 22460
rect 12216 22448 12222 22500
rect 12253 22491 12311 22497
rect 12253 22457 12265 22491
rect 12299 22488 12311 22491
rect 12434 22488 12440 22500
rect 12299 22460 12440 22488
rect 12299 22457 12311 22460
rect 12253 22451 12311 22457
rect 12434 22448 12440 22460
rect 12492 22488 12498 22500
rect 12805 22491 12863 22497
rect 12805 22488 12817 22491
rect 12492 22460 12817 22488
rect 12492 22448 12498 22460
rect 12805 22457 12817 22460
rect 12851 22457 12863 22491
rect 12805 22451 12863 22457
rect 12894 22448 12900 22500
rect 12952 22488 12958 22500
rect 13081 22491 13139 22497
rect 13081 22488 13093 22491
rect 12952 22460 13093 22488
rect 12952 22448 12958 22460
rect 13081 22457 13093 22460
rect 13127 22457 13139 22491
rect 13081 22451 13139 22457
rect 13909 22491 13967 22497
rect 13909 22457 13921 22491
rect 13955 22488 13967 22491
rect 14182 22488 14188 22500
rect 13955 22460 14188 22488
rect 13955 22457 13967 22460
rect 13909 22451 13967 22457
rect 14182 22448 14188 22460
rect 14240 22488 14246 22500
rect 14568 22497 14596 22528
rect 14734 22516 14740 22568
rect 14792 22556 14798 22568
rect 15378 22556 15384 22568
rect 14792 22528 15384 22556
rect 14792 22516 14798 22528
rect 15378 22516 15384 22528
rect 15436 22516 15442 22568
rect 15749 22559 15807 22565
rect 15749 22525 15761 22559
rect 15795 22556 15807 22559
rect 16868 22556 16896 22584
rect 15795 22528 16896 22556
rect 15795 22525 15807 22528
rect 15749 22519 15807 22525
rect 18874 22516 18880 22568
rect 18932 22556 18938 22568
rect 19061 22559 19119 22565
rect 19061 22556 19073 22559
rect 18932 22528 19073 22556
rect 18932 22516 18938 22528
rect 19061 22525 19073 22528
rect 19107 22525 19119 22559
rect 19061 22519 19119 22525
rect 20257 22559 20315 22565
rect 20257 22525 20269 22559
rect 20303 22525 20315 22559
rect 20364 22556 20392 22596
rect 24581 22593 24593 22627
rect 24627 22624 24639 22627
rect 24670 22624 24676 22636
rect 24627 22596 24676 22624
rect 24627 22593 24639 22596
rect 24581 22587 24639 22593
rect 24670 22584 24676 22596
rect 24728 22624 24734 22636
rect 25041 22627 25099 22633
rect 25041 22624 25053 22627
rect 24728 22596 25053 22624
rect 24728 22584 24734 22596
rect 25041 22593 25053 22596
rect 25087 22593 25099 22627
rect 25590 22624 25596 22636
rect 25551 22596 25596 22624
rect 25041 22587 25099 22593
rect 25590 22584 25596 22596
rect 25648 22584 25654 22636
rect 20530 22565 20536 22568
rect 20524 22556 20536 22565
rect 20364 22528 20536 22556
rect 20257 22519 20315 22525
rect 20524 22519 20536 22528
rect 14369 22491 14427 22497
rect 14369 22488 14381 22491
rect 14240 22460 14381 22488
rect 14240 22448 14246 22460
rect 14369 22457 14381 22460
rect 14415 22457 14427 22491
rect 14369 22451 14427 22457
rect 14553 22491 14611 22497
rect 14553 22457 14565 22491
rect 14599 22457 14611 22491
rect 14553 22451 14611 22457
rect 16206 22448 16212 22500
rect 16264 22488 16270 22500
rect 16761 22491 16819 22497
rect 16761 22488 16773 22491
rect 16264 22460 16773 22488
rect 16264 22448 16270 22460
rect 16761 22457 16773 22460
rect 16807 22457 16819 22491
rect 16761 22451 16819 22457
rect 18966 22448 18972 22500
rect 19024 22488 19030 22500
rect 19150 22488 19156 22500
rect 19024 22460 19156 22488
rect 19024 22448 19030 22460
rect 19150 22448 19156 22460
rect 19208 22488 19214 22500
rect 19245 22491 19303 22497
rect 19245 22488 19257 22491
rect 19208 22460 19257 22488
rect 19208 22448 19214 22460
rect 19245 22457 19257 22460
rect 19291 22457 19303 22491
rect 19245 22451 19303 22457
rect 20165 22491 20223 22497
rect 20165 22457 20177 22491
rect 20211 22488 20223 22491
rect 20272 22488 20300 22519
rect 20530 22516 20536 22519
rect 20588 22516 20594 22568
rect 23477 22559 23535 22565
rect 23477 22525 23489 22559
rect 23523 22556 23535 22559
rect 23937 22559 23995 22565
rect 23937 22556 23949 22559
rect 23523 22528 23949 22556
rect 23523 22525 23535 22528
rect 23477 22519 23535 22525
rect 23937 22525 23949 22528
rect 23983 22556 23995 22559
rect 24026 22556 24032 22568
rect 23983 22528 24032 22556
rect 23983 22525 23995 22528
rect 23937 22519 23995 22525
rect 24026 22516 24032 22528
rect 24084 22556 24090 22568
rect 24084 22528 24716 22556
rect 24084 22516 24090 22528
rect 21542 22488 21548 22500
rect 20211 22460 21548 22488
rect 20211 22457 20223 22460
rect 20165 22451 20223 22457
rect 21542 22448 21548 22460
rect 21600 22448 21606 22500
rect 23658 22448 23664 22500
rect 23716 22488 23722 22500
rect 24210 22488 24216 22500
rect 23716 22460 24216 22488
rect 23716 22448 23722 22460
rect 24210 22448 24216 22460
rect 24268 22488 24274 22500
rect 24688 22497 24716 22528
rect 24581 22491 24639 22497
rect 24581 22488 24593 22491
rect 24268 22460 24593 22488
rect 24268 22448 24274 22460
rect 24581 22457 24593 22460
rect 24627 22457 24639 22491
rect 24581 22451 24639 22457
rect 24673 22491 24731 22497
rect 24673 22457 24685 22491
rect 24719 22488 24731 22491
rect 25038 22488 25044 22500
rect 24719 22460 25044 22488
rect 24719 22457 24731 22460
rect 24673 22451 24731 22457
rect 25038 22448 25044 22460
rect 25096 22448 25102 22500
rect 3510 22420 3516 22432
rect 3160 22392 3516 22420
rect 3510 22380 3516 22392
rect 3568 22380 3574 22432
rect 3786 22420 3792 22432
rect 3747 22392 3792 22420
rect 3786 22380 3792 22392
rect 3844 22380 3850 22432
rect 6181 22423 6239 22429
rect 6181 22389 6193 22423
rect 6227 22420 6239 22423
rect 6362 22420 6368 22432
rect 6227 22392 6368 22420
rect 6227 22389 6239 22392
rect 6181 22383 6239 22389
rect 6362 22380 6368 22392
rect 6420 22380 6426 22432
rect 11330 22420 11336 22432
rect 11291 22392 11336 22420
rect 11330 22380 11336 22392
rect 11388 22380 11394 22432
rect 11606 22380 11612 22432
rect 11664 22420 11670 22432
rect 11793 22423 11851 22429
rect 11793 22420 11805 22423
rect 11664 22392 11805 22420
rect 11664 22380 11670 22392
rect 11793 22389 11805 22392
rect 11839 22420 11851 22423
rect 12989 22423 13047 22429
rect 12989 22420 13001 22423
rect 11839 22392 13001 22420
rect 11839 22389 11851 22392
rect 11793 22383 11851 22389
rect 12989 22389 13001 22392
rect 13035 22389 13047 22423
rect 17218 22420 17224 22432
rect 17179 22392 17224 22420
rect 12989 22383 13047 22389
rect 17218 22380 17224 22392
rect 17276 22380 17282 22432
rect 19797 22423 19855 22429
rect 19797 22389 19809 22423
rect 19843 22420 19855 22423
rect 19978 22420 19984 22432
rect 19843 22392 19984 22420
rect 19843 22389 19855 22392
rect 19797 22383 19855 22389
rect 19978 22380 19984 22392
rect 20036 22380 20042 22432
rect 22278 22420 22284 22432
rect 22239 22392 22284 22420
rect 22278 22380 22284 22392
rect 22336 22380 22342 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 3510 22176 3516 22228
rect 3568 22216 3574 22228
rect 3789 22219 3847 22225
rect 3789 22216 3801 22219
rect 3568 22188 3801 22216
rect 3568 22176 3574 22188
rect 3789 22185 3801 22188
rect 3835 22185 3847 22219
rect 5166 22216 5172 22228
rect 5127 22188 5172 22216
rect 3789 22179 3847 22185
rect 5166 22176 5172 22188
rect 5224 22176 5230 22228
rect 5442 22216 5448 22228
rect 5403 22188 5448 22216
rect 5442 22176 5448 22188
rect 5500 22176 5506 22228
rect 5552 22188 6960 22216
rect 2866 22108 2872 22160
rect 2924 22148 2930 22160
rect 4246 22148 4252 22160
rect 2924 22120 4252 22148
rect 2924 22108 2930 22120
rect 4246 22108 4252 22120
rect 4304 22108 4310 22160
rect 5552 22148 5580 22188
rect 5460 22120 5580 22148
rect 1394 22040 1400 22092
rect 1452 22080 1458 22092
rect 1489 22083 1547 22089
rect 1489 22080 1501 22083
rect 1452 22052 1501 22080
rect 1452 22040 1458 22052
rect 1489 22049 1501 22052
rect 1535 22049 1547 22083
rect 1489 22043 1547 22049
rect 1756 22083 1814 22089
rect 1756 22049 1768 22083
rect 1802 22080 1814 22083
rect 3418 22080 3424 22092
rect 1802 22052 3424 22080
rect 1802 22049 1814 22052
rect 1756 22043 1814 22049
rect 3418 22040 3424 22052
rect 3476 22040 3482 22092
rect 4338 22080 4344 22092
rect 4299 22052 4344 22080
rect 4338 22040 4344 22052
rect 4396 22080 4402 22092
rect 5460 22080 5488 22120
rect 5626 22108 5632 22160
rect 5684 22148 5690 22160
rect 6549 22151 6607 22157
rect 6549 22148 6561 22151
rect 5684 22120 6561 22148
rect 5684 22108 5690 22120
rect 6549 22117 6561 22120
rect 6595 22148 6607 22151
rect 6822 22148 6828 22160
rect 6595 22120 6828 22148
rect 6595 22117 6607 22120
rect 6549 22111 6607 22117
rect 6822 22108 6828 22120
rect 6880 22108 6886 22160
rect 6641 22083 6699 22089
rect 6641 22080 6653 22083
rect 4396 22052 5488 22080
rect 5828 22052 6653 22080
rect 4396 22040 4402 22052
rect 4614 22012 4620 22024
rect 4575 21984 4620 22012
rect 4614 21972 4620 21984
rect 4672 21972 4678 22024
rect 2774 21904 2780 21956
rect 2832 21944 2838 21956
rect 3421 21947 3479 21953
rect 3421 21944 3433 21947
rect 2832 21916 3433 21944
rect 2832 21904 2838 21916
rect 3421 21913 3433 21916
rect 3467 21913 3479 21947
rect 3421 21907 3479 21913
rect 2222 21836 2228 21888
rect 2280 21876 2286 21888
rect 2869 21879 2927 21885
rect 2869 21876 2881 21879
rect 2280 21848 2881 21876
rect 2280 21836 2286 21848
rect 2869 21845 2881 21848
rect 2915 21845 2927 21879
rect 2869 21839 2927 21845
rect 4890 21836 4896 21888
rect 4948 21876 4954 21888
rect 5828 21885 5856 22052
rect 6641 22049 6653 22052
rect 6687 22049 6699 22083
rect 6932 22080 6960 22188
rect 7466 22176 7472 22228
rect 7524 22216 7530 22228
rect 7524 22188 8248 22216
rect 7524 22176 7530 22188
rect 7926 22108 7932 22160
rect 7984 22148 7990 22160
rect 8110 22148 8116 22160
rect 7984 22120 8116 22148
rect 7984 22108 7990 22120
rect 8110 22108 8116 22120
rect 8168 22108 8174 22160
rect 7377 22083 7435 22089
rect 7377 22080 7389 22083
rect 6932 22052 7389 22080
rect 6641 22043 6699 22049
rect 7377 22049 7389 22052
rect 7423 22049 7435 22083
rect 7377 22043 7435 22049
rect 7742 22040 7748 22092
rect 7800 22080 7806 22092
rect 8018 22080 8024 22092
rect 7800 22052 8024 22080
rect 7800 22040 7806 22052
rect 8018 22040 8024 22052
rect 8076 22040 8082 22092
rect 8220 22080 8248 22188
rect 8386 22176 8392 22228
rect 8444 22216 8450 22228
rect 8941 22219 8999 22225
rect 8941 22216 8953 22219
rect 8444 22188 8953 22216
rect 8444 22176 8450 22188
rect 8941 22185 8953 22188
rect 8987 22185 8999 22219
rect 8941 22179 8999 22185
rect 9766 22176 9772 22228
rect 9824 22216 9830 22228
rect 10229 22219 10287 22225
rect 10229 22216 10241 22219
rect 9824 22188 10241 22216
rect 9824 22176 9830 22188
rect 10229 22185 10241 22188
rect 10275 22185 10287 22219
rect 11146 22216 11152 22228
rect 11107 22188 11152 22216
rect 10229 22179 10287 22185
rect 11146 22176 11152 22188
rect 11204 22176 11210 22228
rect 11241 22219 11299 22225
rect 11241 22185 11253 22219
rect 11287 22216 11299 22219
rect 13538 22216 13544 22228
rect 11287 22188 13544 22216
rect 11287 22185 11299 22188
rect 11241 22179 11299 22185
rect 13538 22176 13544 22188
rect 13596 22176 13602 22228
rect 13633 22219 13691 22225
rect 13633 22185 13645 22219
rect 13679 22216 13691 22219
rect 13722 22216 13728 22228
rect 13679 22188 13728 22216
rect 13679 22185 13691 22188
rect 13633 22179 13691 22185
rect 13722 22176 13728 22188
rect 13780 22176 13786 22228
rect 13814 22176 13820 22228
rect 13872 22216 13878 22228
rect 14921 22219 14979 22225
rect 14921 22216 14933 22219
rect 13872 22188 14933 22216
rect 13872 22176 13878 22188
rect 14921 22185 14933 22188
rect 14967 22185 14979 22219
rect 14921 22179 14979 22185
rect 16666 22176 16672 22228
rect 16724 22216 16730 22228
rect 16761 22219 16819 22225
rect 16761 22216 16773 22219
rect 16724 22188 16773 22216
rect 16724 22176 16730 22188
rect 16761 22185 16773 22188
rect 16807 22216 16819 22219
rect 16850 22216 16856 22228
rect 16807 22188 16856 22216
rect 16807 22185 16819 22188
rect 16761 22179 16819 22185
rect 16850 22176 16856 22188
rect 16908 22176 16914 22228
rect 20070 22216 20076 22228
rect 20031 22188 20076 22216
rect 20070 22176 20076 22188
rect 20128 22176 20134 22228
rect 22833 22219 22891 22225
rect 22833 22185 22845 22219
rect 22879 22216 22891 22219
rect 23106 22216 23112 22228
rect 22879 22188 23112 22216
rect 22879 22185 22891 22188
rect 22833 22179 22891 22185
rect 23106 22176 23112 22188
rect 23164 22176 23170 22228
rect 23474 22216 23480 22228
rect 23435 22188 23480 22216
rect 23474 22176 23480 22188
rect 23532 22176 23538 22228
rect 10042 22108 10048 22160
rect 10100 22148 10106 22160
rect 11164 22148 11192 22176
rect 12069 22151 12127 22157
rect 12069 22148 12081 22151
rect 10100 22120 11100 22148
rect 11164 22120 12081 22148
rect 10100 22108 10106 22120
rect 8573 22083 8631 22089
rect 8573 22080 8585 22083
rect 8220 22052 8585 22080
rect 8573 22049 8585 22052
rect 8619 22049 8631 22083
rect 9490 22080 9496 22092
rect 9451 22052 9496 22080
rect 8573 22043 8631 22049
rect 9490 22040 9496 22052
rect 9548 22040 9554 22092
rect 10778 22080 10784 22092
rect 10060 22052 10784 22080
rect 10060 22024 10088 22052
rect 10778 22040 10784 22052
rect 10836 22040 10842 22092
rect 11072 22080 11100 22120
rect 12069 22117 12081 22120
rect 12115 22148 12127 22151
rect 12894 22148 12900 22160
rect 12115 22120 12900 22148
rect 12115 22117 12127 22120
rect 12069 22111 12127 22117
rect 12894 22108 12900 22120
rect 12952 22108 12958 22160
rect 13446 22108 13452 22160
rect 13504 22108 13510 22160
rect 14274 22148 14280 22160
rect 14235 22120 14280 22148
rect 14274 22108 14280 22120
rect 14332 22108 14338 22160
rect 15286 22108 15292 22160
rect 15344 22148 15350 22160
rect 15841 22151 15899 22157
rect 15841 22148 15853 22151
rect 15344 22120 15853 22148
rect 15344 22108 15350 22120
rect 15841 22117 15853 22120
rect 15887 22117 15899 22151
rect 16868 22148 16896 22176
rect 17098 22151 17156 22157
rect 17098 22148 17110 22151
rect 16868 22120 17110 22148
rect 15841 22111 15899 22117
rect 17098 22117 17110 22120
rect 17144 22117 17156 22151
rect 17098 22111 17156 22117
rect 18782 22108 18788 22160
rect 18840 22148 18846 22160
rect 18840 22120 19288 22148
rect 18840 22108 18846 22120
rect 11698 22080 11704 22092
rect 11072 22052 11704 22080
rect 11698 22040 11704 22052
rect 11756 22040 11762 22092
rect 11974 22040 11980 22092
rect 12032 22080 12038 22092
rect 12509 22083 12567 22089
rect 12509 22080 12521 22083
rect 12032 22052 12521 22080
rect 12032 22040 12038 22052
rect 12509 22049 12521 22052
rect 12555 22049 12567 22083
rect 13464 22080 13492 22108
rect 13722 22080 13728 22092
rect 13464 22052 13728 22080
rect 12509 22043 12567 22049
rect 13722 22040 13728 22052
rect 13780 22040 13786 22092
rect 15562 22040 15568 22092
rect 15620 22080 15626 22092
rect 15933 22083 15991 22089
rect 15933 22080 15945 22083
rect 15620 22052 15945 22080
rect 15620 22040 15626 22052
rect 15933 22049 15945 22052
rect 15979 22049 15991 22083
rect 15933 22043 15991 22049
rect 16853 22083 16911 22089
rect 16853 22049 16865 22083
rect 16899 22080 16911 22083
rect 17402 22080 17408 22092
rect 16899 22052 17408 22080
rect 16899 22049 16911 22052
rect 16853 22043 16911 22049
rect 17402 22040 17408 22052
rect 17460 22040 17466 22092
rect 19260 22080 19288 22120
rect 19518 22108 19524 22160
rect 19576 22108 19582 22160
rect 19889 22151 19947 22157
rect 19889 22117 19901 22151
rect 19935 22148 19947 22151
rect 19978 22148 19984 22160
rect 19935 22120 19984 22148
rect 19935 22117 19947 22120
rect 19889 22111 19947 22117
rect 19978 22108 19984 22120
rect 20036 22108 20042 22160
rect 21542 22148 21548 22160
rect 21455 22120 21548 22148
rect 21542 22108 21548 22120
rect 21600 22148 21606 22160
rect 21600 22120 23428 22148
rect 21600 22108 21606 22120
rect 19337 22083 19395 22089
rect 19337 22080 19349 22083
rect 19260 22052 19349 22080
rect 19337 22049 19349 22052
rect 19383 22049 19395 22083
rect 19337 22043 19395 22049
rect 6362 21972 6368 22024
rect 6420 22012 6426 22024
rect 6549 22015 6607 22021
rect 6549 22012 6561 22015
rect 6420 21984 6561 22012
rect 6420 21972 6426 21984
rect 6549 21981 6561 21984
rect 6595 21981 6607 22015
rect 8110 22012 8116 22024
rect 8071 21984 8116 22012
rect 6549 21975 6607 21981
rect 6564 21944 6592 21975
rect 8110 21972 8116 21984
rect 8168 21972 8174 22024
rect 8205 22015 8263 22021
rect 8205 21981 8217 22015
rect 8251 22012 8263 22015
rect 8478 22012 8484 22024
rect 8251 21984 8484 22012
rect 8251 21981 8263 21984
rect 8205 21975 8263 21981
rect 8478 21972 8484 21984
rect 8536 21972 8542 22024
rect 10042 21972 10048 22024
rect 10100 21972 10106 22024
rect 10226 22012 10232 22024
rect 10187 21984 10232 22012
rect 10226 21972 10232 21984
rect 10284 21972 10290 22024
rect 10321 22015 10379 22021
rect 10321 21981 10333 22015
rect 10367 21981 10379 22015
rect 10321 21975 10379 21981
rect 7653 21947 7711 21953
rect 7653 21944 7665 21947
rect 6564 21916 7665 21944
rect 7653 21913 7665 21916
rect 7699 21913 7711 21947
rect 7653 21907 7711 21913
rect 9674 21904 9680 21956
rect 9732 21944 9738 21956
rect 9769 21947 9827 21953
rect 9769 21944 9781 21947
rect 9732 21916 9781 21944
rect 9732 21904 9738 21916
rect 9769 21913 9781 21916
rect 9815 21913 9827 21947
rect 9769 21907 9827 21913
rect 9950 21904 9956 21956
rect 10008 21944 10014 21956
rect 10336 21944 10364 21975
rect 10962 21972 10968 22024
rect 11020 22012 11026 22024
rect 11146 22012 11152 22024
rect 11020 21984 11152 22012
rect 11020 21972 11026 21984
rect 11146 21972 11152 21984
rect 11204 22012 11210 22024
rect 11882 22012 11888 22024
rect 11204 21984 11888 22012
rect 11204 21972 11210 21984
rect 11882 21972 11888 21984
rect 11940 22012 11946 22024
rect 12253 22015 12311 22021
rect 12253 22012 12265 22015
rect 11940 21984 12265 22012
rect 11940 21972 11946 21984
rect 12253 21981 12265 21984
rect 12299 21981 12311 22015
rect 15838 22012 15844 22024
rect 15799 21984 15844 22012
rect 12253 21975 12311 21981
rect 15838 21972 15844 21984
rect 15896 21972 15902 22024
rect 19352 22012 19380 22043
rect 19426 22040 19432 22092
rect 19484 22080 19490 22092
rect 19536 22080 19564 22108
rect 19484 22052 19564 22080
rect 19613 22083 19671 22089
rect 19484 22040 19490 22052
rect 19613 22049 19625 22083
rect 19659 22080 19671 22083
rect 20622 22080 20628 22092
rect 19659 22052 20628 22080
rect 19659 22049 19671 22052
rect 19613 22043 19671 22049
rect 20622 22040 20628 22052
rect 20680 22040 20686 22092
rect 20898 22080 20904 22092
rect 20859 22052 20904 22080
rect 20898 22040 20904 22052
rect 20956 22040 20962 22092
rect 21910 22040 21916 22092
rect 21968 22080 21974 22092
rect 22649 22083 22707 22089
rect 22649 22080 22661 22083
rect 21968 22052 22661 22080
rect 21968 22040 21974 22052
rect 22649 22049 22661 22052
rect 22695 22080 22707 22083
rect 23290 22080 23296 22092
rect 22695 22052 23296 22080
rect 22695 22049 22707 22052
rect 22649 22043 22707 22049
rect 23290 22040 23296 22052
rect 23348 22040 23354 22092
rect 23400 22080 23428 22120
rect 23842 22108 23848 22160
rect 23900 22148 23906 22160
rect 24026 22148 24032 22160
rect 23900 22120 24032 22148
rect 23900 22108 23906 22120
rect 24026 22108 24032 22120
rect 24084 22157 24090 22160
rect 24084 22151 24148 22157
rect 24084 22117 24102 22151
rect 24136 22117 24148 22151
rect 24084 22111 24148 22117
rect 24084 22108 24090 22111
rect 24210 22108 24216 22160
rect 24268 22108 24274 22160
rect 24578 22108 24584 22160
rect 24636 22148 24642 22160
rect 24762 22148 24768 22160
rect 24636 22120 24768 22148
rect 24636 22108 24642 22120
rect 24762 22108 24768 22120
rect 24820 22108 24826 22160
rect 24228 22080 24256 22108
rect 25406 22080 25412 22092
rect 23400 22052 25412 22080
rect 19886 22012 19892 22024
rect 19352 21984 19892 22012
rect 19886 21972 19892 21984
rect 19944 21972 19950 22024
rect 20254 21972 20260 22024
rect 20312 22012 20318 22024
rect 20916 22012 20944 22040
rect 20312 21984 20944 22012
rect 22925 22015 22983 22021
rect 20312 21972 20318 21984
rect 22925 21981 22937 22015
rect 22971 22012 22983 22015
rect 23014 22012 23020 22024
rect 22971 21984 23020 22012
rect 22971 21981 22983 21984
rect 22925 21975 22983 21981
rect 23014 21972 23020 21984
rect 23072 21972 23078 22024
rect 23860 22021 23888 22052
rect 25406 22040 25412 22052
rect 25464 22040 25470 22092
rect 23845 22015 23903 22021
rect 23845 21981 23857 22015
rect 23891 21981 23903 22015
rect 23845 21975 23903 21981
rect 10008 21916 10364 21944
rect 10008 21904 10014 21916
rect 14274 21904 14280 21956
rect 14332 21944 14338 21956
rect 14918 21944 14924 21956
rect 14332 21916 14924 21944
rect 14332 21904 14338 21916
rect 14918 21904 14924 21916
rect 14976 21904 14982 21956
rect 16393 21947 16451 21953
rect 16393 21913 16405 21947
rect 16439 21944 16451 21947
rect 16850 21944 16856 21956
rect 16439 21916 16856 21944
rect 16439 21913 16451 21916
rect 16393 21907 16451 21913
rect 16850 21904 16856 21916
rect 16908 21904 16914 21956
rect 22373 21947 22431 21953
rect 22373 21913 22385 21947
rect 22419 21944 22431 21947
rect 23658 21944 23664 21956
rect 22419 21916 23664 21944
rect 22419 21913 22431 21916
rect 22373 21907 22431 21913
rect 23658 21904 23664 21916
rect 23716 21904 23722 21956
rect 5813 21879 5871 21885
rect 5813 21876 5825 21879
rect 4948 21848 5825 21876
rect 4948 21836 4954 21848
rect 5813 21845 5825 21848
rect 5859 21845 5871 21879
rect 6086 21876 6092 21888
rect 6047 21848 6092 21876
rect 5813 21839 5871 21845
rect 6086 21836 6092 21848
rect 6144 21836 6150 21888
rect 7006 21876 7012 21888
rect 6967 21848 7012 21876
rect 7006 21836 7012 21848
rect 7064 21836 7070 21888
rect 10778 21876 10784 21888
rect 10739 21848 10784 21876
rect 10778 21836 10784 21848
rect 10836 21836 10842 21888
rect 11054 21836 11060 21888
rect 11112 21876 11118 21888
rect 11701 21879 11759 21885
rect 11701 21876 11713 21879
rect 11112 21848 11713 21876
rect 11112 21836 11118 21848
rect 11701 21845 11713 21848
rect 11747 21845 11759 21879
rect 11701 21839 11759 21845
rect 12894 21836 12900 21888
rect 12952 21876 12958 21888
rect 13170 21876 13176 21888
rect 12952 21848 13176 21876
rect 12952 21836 12958 21848
rect 13170 21836 13176 21848
rect 13228 21836 13234 21888
rect 13906 21836 13912 21888
rect 13964 21876 13970 21888
rect 14182 21876 14188 21888
rect 13964 21848 14188 21876
rect 13964 21836 13970 21848
rect 14182 21836 14188 21848
rect 14240 21836 14246 21888
rect 14642 21876 14648 21888
rect 14603 21848 14648 21876
rect 14642 21836 14648 21848
rect 14700 21836 14706 21888
rect 15378 21876 15384 21888
rect 15339 21848 15384 21876
rect 15378 21836 15384 21848
rect 15436 21836 15442 21888
rect 17770 21836 17776 21888
rect 17828 21876 17834 21888
rect 18233 21879 18291 21885
rect 18233 21876 18245 21879
rect 17828 21848 18245 21876
rect 17828 21836 17834 21848
rect 18233 21845 18245 21848
rect 18279 21845 18291 21879
rect 18233 21839 18291 21845
rect 18969 21879 19027 21885
rect 18969 21845 18981 21879
rect 19015 21876 19027 21879
rect 19058 21876 19064 21888
rect 19015 21848 19064 21876
rect 19015 21845 19027 21848
rect 18969 21839 19027 21845
rect 19058 21836 19064 21848
rect 19116 21836 19122 21888
rect 19426 21836 19432 21888
rect 19484 21876 19490 21888
rect 19889 21879 19947 21885
rect 19889 21876 19901 21879
rect 19484 21848 19901 21876
rect 19484 21836 19490 21848
rect 19889 21845 19901 21848
rect 19935 21845 19947 21879
rect 19889 21839 19947 21845
rect 20533 21879 20591 21885
rect 20533 21845 20545 21879
rect 20579 21876 20591 21879
rect 20714 21876 20720 21888
rect 20579 21848 20720 21876
rect 20579 21845 20591 21848
rect 20533 21839 20591 21845
rect 20714 21836 20720 21848
rect 20772 21836 20778 21888
rect 21082 21876 21088 21888
rect 21043 21848 21088 21876
rect 21082 21836 21088 21848
rect 21140 21836 21146 21888
rect 22097 21879 22155 21885
rect 22097 21845 22109 21879
rect 22143 21876 22155 21879
rect 22646 21876 22652 21888
rect 22143 21848 22652 21876
rect 22143 21845 22155 21848
rect 22097 21839 22155 21845
rect 22646 21836 22652 21848
rect 22704 21836 22710 21888
rect 22922 21836 22928 21888
rect 22980 21876 22986 21888
rect 23290 21876 23296 21888
rect 22980 21848 23296 21876
rect 22980 21836 22986 21848
rect 23290 21836 23296 21848
rect 23348 21836 23354 21888
rect 24026 21836 24032 21888
rect 24084 21876 24090 21888
rect 25225 21879 25283 21885
rect 25225 21876 25237 21879
rect 24084 21848 25237 21876
rect 24084 21836 24090 21848
rect 25225 21845 25237 21848
rect 25271 21845 25283 21879
rect 25225 21839 25283 21845
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 2866 21672 2872 21684
rect 2827 21644 2872 21672
rect 2866 21632 2872 21644
rect 2924 21632 2930 21684
rect 3418 21632 3424 21684
rect 3476 21672 3482 21684
rect 3973 21675 4031 21681
rect 3973 21672 3985 21675
rect 3476 21644 3985 21672
rect 3476 21632 3482 21644
rect 3973 21641 3985 21644
rect 4019 21641 4031 21675
rect 3973 21635 4031 21641
rect 8110 21632 8116 21684
rect 8168 21672 8174 21684
rect 8849 21675 8907 21681
rect 8849 21672 8861 21675
rect 8168 21644 8861 21672
rect 8168 21632 8174 21644
rect 8849 21641 8861 21644
rect 8895 21672 8907 21675
rect 9582 21672 9588 21684
rect 8895 21644 9588 21672
rect 8895 21641 8907 21644
rect 8849 21635 8907 21641
rect 9582 21632 9588 21644
rect 9640 21632 9646 21684
rect 10410 21672 10416 21684
rect 10371 21644 10416 21672
rect 10410 21632 10416 21644
rect 10468 21632 10474 21684
rect 10597 21675 10655 21681
rect 10597 21641 10609 21675
rect 10643 21672 10655 21675
rect 10686 21672 10692 21684
rect 10643 21644 10692 21672
rect 10643 21641 10655 21644
rect 10597 21635 10655 21641
rect 10686 21632 10692 21644
rect 10744 21632 10750 21684
rect 11882 21672 11888 21684
rect 11843 21644 11888 21672
rect 11882 21632 11888 21644
rect 11940 21632 11946 21684
rect 12526 21672 12532 21684
rect 12487 21644 12532 21672
rect 12526 21632 12532 21644
rect 12584 21632 12590 21684
rect 14185 21675 14243 21681
rect 14185 21641 14197 21675
rect 14231 21672 14243 21675
rect 14734 21672 14740 21684
rect 14231 21644 14740 21672
rect 14231 21641 14243 21644
rect 14185 21635 14243 21641
rect 14734 21632 14740 21644
rect 14792 21632 14798 21684
rect 16390 21632 16396 21684
rect 16448 21672 16454 21684
rect 16485 21675 16543 21681
rect 16485 21672 16497 21675
rect 16448 21644 16497 21672
rect 16448 21632 16454 21644
rect 16485 21641 16497 21644
rect 16531 21641 16543 21675
rect 16485 21635 16543 21641
rect 17494 21632 17500 21684
rect 17552 21672 17558 21684
rect 17773 21675 17831 21681
rect 17773 21672 17785 21675
rect 17552 21644 17785 21672
rect 17552 21632 17558 21644
rect 17773 21641 17785 21644
rect 17819 21641 17831 21675
rect 18966 21672 18972 21684
rect 18927 21644 18972 21672
rect 17773 21635 17831 21641
rect 18966 21632 18972 21644
rect 19024 21632 19030 21684
rect 19886 21672 19892 21684
rect 19847 21644 19892 21672
rect 19886 21632 19892 21644
rect 19944 21632 19950 21684
rect 21910 21672 21916 21684
rect 21871 21644 21916 21672
rect 21910 21632 21916 21644
rect 21968 21632 21974 21684
rect 23106 21672 23112 21684
rect 23067 21644 23112 21672
rect 23106 21632 23112 21644
rect 23164 21632 23170 21684
rect 23753 21675 23811 21681
rect 23753 21641 23765 21675
rect 23799 21672 23811 21675
rect 23845 21675 23903 21681
rect 23845 21672 23857 21675
rect 23799 21644 23857 21672
rect 23799 21641 23811 21644
rect 23753 21635 23811 21641
rect 23845 21641 23857 21644
rect 23891 21672 23903 21675
rect 24210 21672 24216 21684
rect 23891 21644 24216 21672
rect 23891 21641 23903 21644
rect 23845 21635 23903 21641
rect 24210 21632 24216 21644
rect 24268 21632 24274 21684
rect 24670 21672 24676 21684
rect 24631 21644 24676 21672
rect 24670 21632 24676 21644
rect 24728 21632 24734 21684
rect 1486 21604 1492 21616
rect 1447 21576 1492 21604
rect 1486 21564 1492 21576
rect 1544 21564 1550 21616
rect 3053 21607 3111 21613
rect 3053 21573 3065 21607
rect 3099 21604 3111 21607
rect 3786 21604 3792 21616
rect 3099 21576 3792 21604
rect 3099 21573 3111 21576
rect 3053 21567 3111 21573
rect 3786 21564 3792 21576
rect 3844 21564 3850 21616
rect 5261 21607 5319 21613
rect 5261 21573 5273 21607
rect 5307 21604 5319 21607
rect 5534 21604 5540 21616
rect 5307 21576 5540 21604
rect 5307 21573 5319 21576
rect 5261 21567 5319 21573
rect 5534 21564 5540 21576
rect 5592 21564 5598 21616
rect 8202 21604 8208 21616
rect 8163 21576 8208 21604
rect 8202 21564 8208 21576
rect 8260 21564 8266 21616
rect 12342 21564 12348 21616
rect 12400 21604 12406 21616
rect 14550 21604 14556 21616
rect 12400 21576 14136 21604
rect 12400 21564 12406 21576
rect 3513 21539 3571 21545
rect 3513 21505 3525 21539
rect 3559 21536 3571 21539
rect 3694 21536 3700 21548
rect 3559 21508 3700 21536
rect 3559 21505 3571 21508
rect 3513 21499 3571 21505
rect 3694 21496 3700 21508
rect 3752 21496 3758 21548
rect 5721 21539 5779 21545
rect 5721 21505 5733 21539
rect 5767 21536 5779 21539
rect 6086 21536 6092 21548
rect 5767 21508 6092 21536
rect 5767 21505 5779 21508
rect 5721 21499 5779 21505
rect 6086 21496 6092 21508
rect 6144 21496 6150 21548
rect 10778 21496 10784 21548
rect 10836 21536 10842 21548
rect 11149 21539 11207 21545
rect 11149 21536 11161 21539
rect 10836 21508 11161 21536
rect 10836 21496 10842 21508
rect 11149 21505 11161 21508
rect 11195 21536 11207 21539
rect 11974 21536 11980 21548
rect 11195 21508 11980 21536
rect 11195 21505 11207 21508
rect 11149 21499 11207 21505
rect 11974 21496 11980 21508
rect 12032 21536 12038 21548
rect 13449 21539 13507 21545
rect 13449 21536 13461 21539
rect 12032 21508 13461 21536
rect 12032 21496 12038 21508
rect 13449 21505 13461 21508
rect 13495 21505 13507 21539
rect 13449 21499 13507 21505
rect 2409 21471 2467 21477
rect 2409 21468 2421 21471
rect 1780 21440 2421 21468
rect 1780 21412 1808 21440
rect 2409 21437 2421 21440
rect 2455 21437 2467 21471
rect 2409 21431 2467 21437
rect 2498 21428 2504 21480
rect 2556 21468 2562 21480
rect 2774 21468 2780 21480
rect 2556 21440 2780 21468
rect 2556 21428 2562 21440
rect 2774 21428 2780 21440
rect 2832 21468 2838 21480
rect 3605 21471 3663 21477
rect 3605 21468 3617 21471
rect 2832 21440 3617 21468
rect 2832 21428 2838 21440
rect 3605 21437 3617 21440
rect 3651 21437 3663 21471
rect 3605 21431 3663 21437
rect 5077 21471 5135 21477
rect 5077 21437 5089 21471
rect 5123 21468 5135 21471
rect 5813 21471 5871 21477
rect 5813 21468 5825 21471
rect 5123 21440 5825 21468
rect 5123 21437 5135 21440
rect 5077 21431 5135 21437
rect 5813 21437 5825 21440
rect 5859 21468 5871 21471
rect 6181 21471 6239 21477
rect 6181 21468 6193 21471
rect 5859 21440 6193 21468
rect 5859 21437 5871 21440
rect 5813 21431 5871 21437
rect 6181 21437 6193 21440
rect 6227 21468 6239 21471
rect 6454 21468 6460 21480
rect 6227 21440 6460 21468
rect 6227 21437 6239 21440
rect 6181 21431 6239 21437
rect 6454 21428 6460 21440
rect 6512 21428 6518 21480
rect 6638 21428 6644 21480
rect 6696 21468 6702 21480
rect 6825 21471 6883 21477
rect 6825 21468 6837 21471
rect 6696 21440 6837 21468
rect 6696 21428 6702 21440
rect 6825 21437 6837 21440
rect 6871 21468 6883 21471
rect 7466 21468 7472 21480
rect 6871 21440 7472 21468
rect 6871 21437 6883 21440
rect 6825 21431 6883 21437
rect 7466 21428 7472 21440
rect 7524 21428 7530 21480
rect 12253 21471 12311 21477
rect 12253 21437 12265 21471
rect 12299 21468 12311 21471
rect 12805 21471 12863 21477
rect 12805 21468 12817 21471
rect 12299 21440 12817 21468
rect 12299 21437 12311 21440
rect 12253 21431 12311 21437
rect 12805 21437 12817 21440
rect 12851 21468 12863 21471
rect 14108 21468 14136 21576
rect 14200 21576 14556 21604
rect 14200 21548 14228 21576
rect 14550 21564 14556 21576
rect 14608 21564 14614 21616
rect 19978 21564 19984 21616
rect 20036 21604 20042 21616
rect 20533 21607 20591 21613
rect 20533 21604 20545 21607
rect 20036 21576 20545 21604
rect 20036 21564 20042 21576
rect 20533 21573 20545 21576
rect 20579 21573 20591 21607
rect 20533 21567 20591 21573
rect 22097 21607 22155 21613
rect 22097 21573 22109 21607
rect 22143 21604 22155 21607
rect 23290 21604 23296 21616
rect 22143 21576 23296 21604
rect 22143 21573 22155 21576
rect 22097 21567 22155 21573
rect 23290 21564 23296 21576
rect 23348 21564 23354 21616
rect 23658 21564 23664 21616
rect 23716 21604 23722 21616
rect 23934 21604 23940 21616
rect 23716 21576 23940 21604
rect 23716 21564 23722 21576
rect 23934 21564 23940 21576
rect 23992 21564 23998 21616
rect 14182 21496 14188 21548
rect 14240 21496 14246 21548
rect 14642 21536 14648 21548
rect 14603 21508 14648 21536
rect 14642 21496 14648 21508
rect 14700 21496 14706 21548
rect 16850 21536 16856 21548
rect 16811 21508 16856 21536
rect 16850 21496 16856 21508
rect 16908 21496 16914 21548
rect 18785 21539 18843 21545
rect 18785 21505 18797 21539
rect 18831 21536 18843 21539
rect 19429 21539 19487 21545
rect 19429 21536 19441 21539
rect 18831 21508 19441 21536
rect 18831 21505 18843 21508
rect 18785 21499 18843 21505
rect 19429 21505 19441 21508
rect 19475 21536 19487 21539
rect 20070 21536 20076 21548
rect 19475 21508 20076 21536
rect 19475 21505 19487 21508
rect 19429 21499 19487 21505
rect 20070 21496 20076 21508
rect 20128 21496 20134 21548
rect 20714 21496 20720 21548
rect 20772 21536 20778 21548
rect 21085 21539 21143 21545
rect 21085 21536 21097 21539
rect 20772 21508 21097 21536
rect 20772 21496 20778 21508
rect 21085 21505 21097 21508
rect 21131 21536 21143 21539
rect 21358 21536 21364 21548
rect 21131 21508 21364 21536
rect 21131 21505 21143 21508
rect 21085 21499 21143 21505
rect 21358 21496 21364 21508
rect 21416 21496 21422 21548
rect 22186 21496 22192 21548
rect 22244 21536 22250 21548
rect 22557 21539 22615 21545
rect 22557 21536 22569 21539
rect 22244 21508 22569 21536
rect 22244 21496 22250 21508
rect 22557 21505 22569 21508
rect 22603 21536 22615 21539
rect 23750 21536 23756 21548
rect 22603 21508 23756 21536
rect 22603 21505 22615 21508
rect 22557 21499 22615 21505
rect 23750 21496 23756 21508
rect 23808 21496 23814 21548
rect 15286 21468 15292 21480
rect 12851 21440 13492 21468
rect 14108 21440 15292 21468
rect 12851 21437 12863 21440
rect 12805 21431 12863 21437
rect 1762 21400 1768 21412
rect 1723 21372 1768 21400
rect 1762 21360 1768 21372
rect 1820 21360 1826 21412
rect 2041 21403 2099 21409
rect 2041 21369 2053 21403
rect 2087 21400 2099 21403
rect 2222 21400 2228 21412
rect 2087 21372 2228 21400
rect 2087 21369 2099 21372
rect 2041 21363 2099 21369
rect 2222 21360 2228 21372
rect 2280 21360 2286 21412
rect 2958 21360 2964 21412
rect 3016 21400 3022 21412
rect 3513 21403 3571 21409
rect 3513 21400 3525 21403
rect 3016 21372 3525 21400
rect 3016 21360 3022 21372
rect 3513 21369 3525 21372
rect 3559 21369 3571 21403
rect 3513 21363 3571 21369
rect 4709 21403 4767 21409
rect 4709 21369 4721 21403
rect 4755 21400 4767 21403
rect 5258 21400 5264 21412
rect 4755 21372 5264 21400
rect 4755 21369 4767 21372
rect 4709 21363 4767 21369
rect 5258 21360 5264 21372
rect 5316 21400 5322 21412
rect 5721 21403 5779 21409
rect 5721 21400 5733 21403
rect 5316 21372 5733 21400
rect 5316 21360 5322 21372
rect 5721 21369 5733 21372
rect 5767 21369 5779 21403
rect 6472 21400 6500 21428
rect 13464 21412 13492 21440
rect 15286 21428 15292 21440
rect 15344 21468 15350 21480
rect 15930 21468 15936 21480
rect 15344 21440 15936 21468
rect 15344 21428 15350 21440
rect 15930 21428 15936 21440
rect 15988 21428 15994 21480
rect 17494 21468 17500 21480
rect 16960 21440 17500 21468
rect 7070 21403 7128 21409
rect 7070 21400 7082 21403
rect 6472 21372 7082 21400
rect 5721 21363 5779 21369
rect 7070 21369 7082 21372
rect 7116 21369 7128 21403
rect 7070 21363 7128 21369
rect 7558 21360 7564 21412
rect 7616 21400 7622 21412
rect 7742 21400 7748 21412
rect 7616 21372 7748 21400
rect 7616 21360 7622 21372
rect 7742 21360 7748 21372
rect 7800 21360 7806 21412
rect 10870 21400 10876 21412
rect 10831 21372 10876 21400
rect 10870 21360 10876 21372
rect 10928 21360 10934 21412
rect 13078 21400 13084 21412
rect 13039 21372 13084 21400
rect 13078 21360 13084 21372
rect 13136 21360 13142 21412
rect 13446 21360 13452 21412
rect 13504 21360 13510 21412
rect 14550 21360 14556 21412
rect 14608 21400 14614 21412
rect 14645 21403 14703 21409
rect 14645 21400 14657 21403
rect 14608 21372 14657 21400
rect 14608 21360 14614 21372
rect 14645 21369 14657 21372
rect 14691 21369 14703 21403
rect 14645 21363 14703 21369
rect 14737 21403 14795 21409
rect 14737 21369 14749 21403
rect 14783 21400 14795 21403
rect 15102 21400 15108 21412
rect 14783 21372 15108 21400
rect 14783 21369 14795 21372
rect 14737 21363 14795 21369
rect 1949 21335 2007 21341
rect 1949 21301 1961 21335
rect 1995 21332 2007 21335
rect 2314 21332 2320 21344
rect 1995 21304 2320 21332
rect 1995 21301 2007 21304
rect 1949 21295 2007 21301
rect 2314 21292 2320 21304
rect 2372 21292 2378 21344
rect 6638 21332 6644 21344
rect 6599 21304 6644 21332
rect 6638 21292 6644 21304
rect 6696 21292 6702 21344
rect 8478 21292 8484 21344
rect 8536 21332 8542 21344
rect 9125 21335 9183 21341
rect 9125 21332 9137 21335
rect 8536 21304 9137 21332
rect 8536 21292 8542 21304
rect 9125 21301 9137 21304
rect 9171 21301 9183 21335
rect 9125 21295 9183 21301
rect 9493 21335 9551 21341
rect 9493 21301 9505 21335
rect 9539 21332 9551 21335
rect 9674 21332 9680 21344
rect 9539 21304 9680 21332
rect 9539 21301 9551 21304
rect 9493 21295 9551 21301
rect 9674 21292 9680 21304
rect 9732 21292 9738 21344
rect 9766 21292 9772 21344
rect 9824 21332 9830 21344
rect 10045 21335 10103 21341
rect 10045 21332 10057 21335
rect 9824 21304 10057 21332
rect 9824 21292 9830 21304
rect 10045 21301 10057 21304
rect 10091 21332 10103 21335
rect 10686 21332 10692 21344
rect 10091 21304 10692 21332
rect 10091 21301 10103 21304
rect 10045 21295 10103 21301
rect 10686 21292 10692 21304
rect 10744 21292 10750 21344
rect 11054 21332 11060 21344
rect 11015 21304 11060 21332
rect 11054 21292 11060 21304
rect 11112 21292 11118 21344
rect 12618 21292 12624 21344
rect 12676 21332 12682 21344
rect 12989 21335 13047 21341
rect 12989 21332 13001 21335
rect 12676 21304 13001 21332
rect 12676 21292 12682 21304
rect 12989 21301 13001 21304
rect 13035 21301 13047 21335
rect 13998 21332 14004 21344
rect 13911 21304 14004 21332
rect 12989 21295 13047 21301
rect 13998 21292 14004 21304
rect 14056 21332 14062 21344
rect 14752 21332 14780 21363
rect 15102 21360 15108 21372
rect 15160 21360 15166 21412
rect 15749 21403 15807 21409
rect 15749 21369 15761 21403
rect 15795 21400 15807 21403
rect 15838 21400 15844 21412
rect 15795 21372 15844 21400
rect 15795 21369 15807 21372
rect 15749 21363 15807 21369
rect 15838 21360 15844 21372
rect 15896 21400 15902 21412
rect 16482 21400 16488 21412
rect 15896 21372 16488 21400
rect 15896 21360 15902 21372
rect 16482 21360 16488 21372
rect 16540 21360 16546 21412
rect 16960 21409 16988 21440
rect 17494 21428 17500 21440
rect 17552 21428 17558 21480
rect 19058 21428 19064 21480
rect 19116 21468 19122 21480
rect 19521 21471 19579 21477
rect 19521 21468 19533 21471
rect 19116 21440 19533 21468
rect 19116 21428 19122 21440
rect 19521 21437 19533 21440
rect 19567 21468 19579 21471
rect 20346 21468 20352 21480
rect 19567 21440 20352 21468
rect 19567 21437 19579 21440
rect 19521 21431 19579 21437
rect 20346 21428 20352 21440
rect 20404 21428 20410 21480
rect 22646 21468 22652 21480
rect 22607 21440 22652 21468
rect 22646 21428 22652 21440
rect 22704 21428 22710 21480
rect 24118 21428 24124 21480
rect 24176 21468 24182 21480
rect 24670 21468 24676 21480
rect 24176 21440 24676 21468
rect 24176 21428 24182 21440
rect 24670 21428 24676 21440
rect 24728 21428 24734 21480
rect 24854 21428 24860 21480
rect 24912 21468 24918 21480
rect 24949 21471 25007 21477
rect 24949 21468 24961 21471
rect 24912 21440 24961 21468
rect 24912 21428 24918 21440
rect 24949 21437 24961 21440
rect 24995 21437 25007 21471
rect 24949 21431 25007 21437
rect 16945 21403 17003 21409
rect 16945 21369 16957 21403
rect 16991 21369 17003 21403
rect 16945 21363 17003 21369
rect 17037 21403 17095 21409
rect 17037 21369 17049 21403
rect 17083 21400 17095 21403
rect 17954 21400 17960 21412
rect 17083 21372 17960 21400
rect 17083 21369 17095 21372
rect 17037 21363 17095 21369
rect 14056 21304 14780 21332
rect 16301 21335 16359 21341
rect 14056 21292 14062 21304
rect 16301 21301 16313 21335
rect 16347 21332 16359 21335
rect 17052 21332 17080 21363
rect 17954 21360 17960 21372
rect 18012 21360 18018 21412
rect 18417 21403 18475 21409
rect 18417 21369 18429 21403
rect 18463 21400 18475 21403
rect 19334 21400 19340 21412
rect 18463 21372 19340 21400
rect 18463 21369 18475 21372
rect 18417 21363 18475 21369
rect 19334 21360 19340 21372
rect 19392 21400 19398 21412
rect 19429 21403 19487 21409
rect 19429 21400 19441 21403
rect 19392 21372 19441 21400
rect 19392 21360 19398 21372
rect 19429 21369 19441 21372
rect 19475 21369 19487 21403
rect 19429 21363 19487 21369
rect 20438 21360 20444 21412
rect 20496 21400 20502 21412
rect 20809 21403 20867 21409
rect 20809 21400 20821 21403
rect 20496 21372 20821 21400
rect 20496 21360 20502 21372
rect 20809 21369 20821 21372
rect 20855 21369 20867 21403
rect 20809 21363 20867 21369
rect 21545 21403 21603 21409
rect 21545 21369 21557 21403
rect 21591 21400 21603 21403
rect 22002 21400 22008 21412
rect 21591 21372 22008 21400
rect 21591 21369 21603 21372
rect 21545 21363 21603 21369
rect 22002 21360 22008 21372
rect 22060 21400 22066 21412
rect 23014 21400 23020 21412
rect 22060 21372 23020 21400
rect 22060 21360 22066 21372
rect 23014 21360 23020 21372
rect 23072 21360 23078 21412
rect 23477 21403 23535 21409
rect 23477 21369 23489 21403
rect 23523 21400 23535 21403
rect 23934 21400 23940 21412
rect 23523 21372 23940 21400
rect 23523 21369 23535 21372
rect 23477 21363 23535 21369
rect 23934 21360 23940 21372
rect 23992 21360 23998 21412
rect 25038 21360 25044 21412
rect 25096 21400 25102 21412
rect 25225 21403 25283 21409
rect 25225 21400 25237 21403
rect 25096 21372 25237 21400
rect 25096 21360 25102 21372
rect 25225 21369 25237 21372
rect 25271 21369 25283 21403
rect 25225 21363 25283 21369
rect 16347 21304 17080 21332
rect 16347 21301 16359 21304
rect 16301 21295 16359 21301
rect 17126 21292 17132 21344
rect 17184 21332 17190 21344
rect 17402 21332 17408 21344
rect 17184 21304 17408 21332
rect 17184 21292 17190 21304
rect 17402 21292 17408 21304
rect 17460 21292 17466 21344
rect 20254 21332 20260 21344
rect 20215 21304 20260 21332
rect 20254 21292 20260 21304
rect 20312 21332 20318 21344
rect 20993 21335 21051 21341
rect 20993 21332 21005 21335
rect 20312 21304 21005 21332
rect 20312 21292 20318 21304
rect 20993 21301 21005 21304
rect 21039 21301 21051 21335
rect 22554 21332 22560 21344
rect 22515 21304 22560 21332
rect 20993 21295 21051 21301
rect 22554 21292 22560 21304
rect 22612 21292 22618 21344
rect 23750 21332 23756 21344
rect 23711 21304 23756 21332
rect 23750 21292 23756 21304
rect 23808 21292 23814 21344
rect 24118 21292 24124 21344
rect 24176 21332 24182 21344
rect 24397 21335 24455 21341
rect 24397 21332 24409 21335
rect 24176 21304 24409 21332
rect 24176 21292 24182 21304
rect 24397 21301 24409 21304
rect 24443 21332 24455 21335
rect 25130 21332 25136 21344
rect 24443 21304 25136 21332
rect 24443 21301 24455 21304
rect 24397 21295 24455 21301
rect 25130 21292 25136 21304
rect 25188 21292 25194 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 2314 21088 2320 21140
rect 2372 21128 2378 21140
rect 2593 21131 2651 21137
rect 2593 21128 2605 21131
rect 2372 21100 2605 21128
rect 2372 21088 2378 21100
rect 2593 21097 2605 21100
rect 2639 21097 2651 21131
rect 2958 21128 2964 21140
rect 2919 21100 2964 21128
rect 2593 21091 2651 21097
rect 2958 21088 2964 21100
rect 3016 21088 3022 21140
rect 3421 21131 3479 21137
rect 3421 21097 3433 21131
rect 3467 21128 3479 21131
rect 3694 21128 3700 21140
rect 3467 21100 3700 21128
rect 3467 21097 3479 21100
rect 3421 21091 3479 21097
rect 3694 21088 3700 21100
rect 3752 21088 3758 21140
rect 6454 21128 6460 21140
rect 6415 21100 6460 21128
rect 6454 21088 6460 21100
rect 6512 21088 6518 21140
rect 7653 21131 7711 21137
rect 7653 21097 7665 21131
rect 7699 21128 7711 21131
rect 7926 21128 7932 21140
rect 7699 21100 7932 21128
rect 7699 21097 7711 21100
rect 7653 21091 7711 21097
rect 7926 21088 7932 21100
rect 7984 21088 7990 21140
rect 9950 21128 9956 21140
rect 9911 21100 9956 21128
rect 9950 21088 9956 21100
rect 10008 21088 10014 21140
rect 11974 21128 11980 21140
rect 11935 21100 11980 21128
rect 11974 21088 11980 21100
rect 12032 21088 12038 21140
rect 13354 21088 13360 21140
rect 13412 21128 13418 21140
rect 13633 21131 13691 21137
rect 13633 21128 13645 21131
rect 13412 21100 13645 21128
rect 13412 21088 13418 21100
rect 13633 21097 13645 21100
rect 13679 21097 13691 21131
rect 13633 21091 13691 21097
rect 13722 21088 13728 21140
rect 13780 21128 13786 21140
rect 14093 21131 14151 21137
rect 14093 21128 14105 21131
rect 13780 21100 14105 21128
rect 13780 21088 13786 21100
rect 14093 21097 14105 21100
rect 14139 21097 14151 21131
rect 14550 21128 14556 21140
rect 14511 21100 14556 21128
rect 14093 21091 14151 21097
rect 14550 21088 14556 21100
rect 14608 21088 14614 21140
rect 16390 21128 16396 21140
rect 16351 21100 16396 21128
rect 16390 21088 16396 21100
rect 16448 21128 16454 21140
rect 16574 21128 16580 21140
rect 16448 21100 16580 21128
rect 16448 21088 16454 21100
rect 16574 21088 16580 21100
rect 16632 21088 16638 21140
rect 16666 21088 16672 21140
rect 16724 21128 16730 21140
rect 16853 21131 16911 21137
rect 16853 21128 16865 21131
rect 16724 21100 16865 21128
rect 16724 21088 16730 21100
rect 16853 21097 16865 21100
rect 16899 21097 16911 21131
rect 16853 21091 16911 21097
rect 17862 21088 17868 21140
rect 17920 21128 17926 21140
rect 18506 21128 18512 21140
rect 17920 21100 18512 21128
rect 17920 21088 17926 21100
rect 18506 21088 18512 21100
rect 18564 21088 18570 21140
rect 19518 21088 19524 21140
rect 19576 21128 19582 21140
rect 19797 21131 19855 21137
rect 19797 21128 19809 21131
rect 19576 21100 19809 21128
rect 19576 21088 19582 21100
rect 19797 21097 19809 21100
rect 19843 21097 19855 21131
rect 20438 21128 20444 21140
rect 20399 21100 20444 21128
rect 19797 21091 19855 21097
rect 20438 21088 20444 21100
rect 20496 21088 20502 21140
rect 22278 21128 22284 21140
rect 22239 21100 22284 21128
rect 22278 21088 22284 21100
rect 22336 21088 22342 21140
rect 22554 21088 22560 21140
rect 22612 21128 22618 21140
rect 22925 21131 22983 21137
rect 22925 21128 22937 21131
rect 22612 21100 22937 21128
rect 22612 21088 22618 21100
rect 22925 21097 22937 21100
rect 22971 21128 22983 21131
rect 23382 21128 23388 21140
rect 22971 21100 23388 21128
rect 22971 21097 22983 21100
rect 22925 21091 22983 21097
rect 23382 21088 23388 21100
rect 23440 21088 23446 21140
rect 24854 21088 24860 21140
rect 24912 21128 24918 21140
rect 25409 21131 25467 21137
rect 25409 21128 25421 21131
rect 24912 21100 25421 21128
rect 24912 21088 24918 21100
rect 25409 21097 25421 21100
rect 25455 21097 25467 21131
rect 25409 21091 25467 21097
rect 1486 21020 1492 21072
rect 1544 21060 1550 21072
rect 2133 21063 2191 21069
rect 2133 21060 2145 21063
rect 1544 21032 2145 21060
rect 1544 21020 1550 21032
rect 2133 21029 2145 21032
rect 2179 21060 2191 21063
rect 2682 21060 2688 21072
rect 2179 21032 2688 21060
rect 2179 21029 2191 21032
rect 2133 21023 2191 21029
rect 2682 21020 2688 21032
rect 2740 21020 2746 21072
rect 8110 21020 8116 21072
rect 8168 21060 8174 21072
rect 8386 21060 8392 21072
rect 8168 21032 8392 21060
rect 8168 21020 8174 21032
rect 8386 21020 8392 21032
rect 8444 21020 8450 21072
rect 8478 21020 8484 21072
rect 8536 21060 8542 21072
rect 8536 21032 8581 21060
rect 8536 21020 8542 21032
rect 10778 21020 10784 21072
rect 10836 21069 10842 21072
rect 10836 21063 10900 21069
rect 10836 21029 10854 21063
rect 10888 21029 10900 21063
rect 10836 21023 10900 21029
rect 10836 21020 10842 21023
rect 11698 21020 11704 21072
rect 11756 21060 11762 21072
rect 12802 21060 12808 21072
rect 11756 21032 12808 21060
rect 11756 21020 11762 21032
rect 12802 21020 12808 21032
rect 12860 21020 12866 21072
rect 15746 21020 15752 21072
rect 15804 21060 15810 21072
rect 15841 21063 15899 21069
rect 15841 21060 15853 21063
rect 15804 21032 15853 21060
rect 15804 21020 15810 21032
rect 15841 21029 15853 21032
rect 15887 21029 15899 21063
rect 15841 21023 15899 21029
rect 19429 21063 19487 21069
rect 19429 21029 19441 21063
rect 19475 21060 19487 21063
rect 20898 21060 20904 21072
rect 19475 21032 20904 21060
rect 19475 21029 19487 21032
rect 19429 21023 19487 21029
rect 20898 21020 20904 21032
rect 20956 21020 20962 21072
rect 24210 21060 24216 21072
rect 24171 21032 24216 21060
rect 24210 21020 24216 21032
rect 24268 21020 24274 21072
rect 24765 21063 24823 21069
rect 24765 21029 24777 21063
rect 24811 21060 24823 21063
rect 24946 21060 24952 21072
rect 24811 21032 24952 21060
rect 24811 21029 24823 21032
rect 24765 21023 24823 21029
rect 1949 20995 2007 21001
rect 1949 20961 1961 20995
rect 1995 20992 2007 20995
rect 2038 20992 2044 21004
rect 1995 20964 2044 20992
rect 1995 20961 2007 20964
rect 1949 20955 2007 20961
rect 2038 20952 2044 20964
rect 2096 20992 2102 21004
rect 4065 20995 4123 21001
rect 4065 20992 4077 20995
rect 2096 20964 4077 20992
rect 2096 20952 2102 20964
rect 4065 20961 4077 20964
rect 4111 20961 4123 20995
rect 4065 20955 4123 20961
rect 4890 20952 4896 21004
rect 4948 20992 4954 21004
rect 5333 20995 5391 21001
rect 5333 20992 5345 20995
rect 4948 20964 5345 20992
rect 4948 20952 4954 20964
rect 5333 20961 5345 20964
rect 5379 20961 5391 20995
rect 5333 20955 5391 20961
rect 7285 20995 7343 21001
rect 7285 20961 7297 20995
rect 7331 20992 7343 20995
rect 7650 20992 7656 21004
rect 7331 20964 7656 20992
rect 7331 20961 7343 20964
rect 7285 20955 7343 20961
rect 7650 20952 7656 20964
rect 7708 20992 7714 21004
rect 8496 20992 8524 21020
rect 7708 20964 8524 20992
rect 10597 20995 10655 21001
rect 7708 20952 7714 20964
rect 10597 20961 10609 20995
rect 10643 20992 10655 20995
rect 11146 20992 11152 21004
rect 10643 20964 11152 20992
rect 10643 20961 10655 20964
rect 10597 20955 10655 20961
rect 11146 20952 11152 20964
rect 11204 20952 11210 21004
rect 12434 20952 12440 21004
rect 12492 20992 12498 21004
rect 13722 20992 13728 21004
rect 12492 20964 13728 20992
rect 12492 20952 12498 20964
rect 13722 20952 13728 20964
rect 13780 20952 13786 21004
rect 15286 20952 15292 21004
rect 15344 20992 15350 21004
rect 15657 20995 15715 21001
rect 15657 20992 15669 20995
rect 15344 20964 15669 20992
rect 15344 20952 15350 20964
rect 15657 20961 15669 20964
rect 15703 20961 15715 20995
rect 15657 20955 15715 20961
rect 17034 20952 17040 21004
rect 17092 20992 17098 21004
rect 17385 20995 17443 21001
rect 17385 20992 17397 20995
rect 17092 20964 17397 20992
rect 17092 20952 17098 20964
rect 17385 20961 17397 20964
rect 17431 20992 17443 20995
rect 17770 20992 17776 21004
rect 17431 20964 17776 20992
rect 17431 20961 17443 20964
rect 17385 20955 17443 20961
rect 17770 20952 17776 20964
rect 17828 20952 17834 21004
rect 19334 20952 19340 21004
rect 19392 20992 19398 21004
rect 19613 20995 19671 21001
rect 19613 20992 19625 20995
rect 19392 20964 19625 20992
rect 19392 20952 19398 20964
rect 19613 20961 19625 20964
rect 19659 20961 19671 20995
rect 19613 20955 19671 20961
rect 20162 20952 20168 21004
rect 20220 20992 20226 21004
rect 20990 20992 20996 21004
rect 20220 20964 20996 20992
rect 20220 20952 20226 20964
rect 20990 20952 20996 20964
rect 21048 20992 21054 21004
rect 21157 20995 21215 21001
rect 21157 20992 21169 20995
rect 21048 20964 21169 20992
rect 21048 20952 21054 20964
rect 21157 20961 21169 20964
rect 21203 20961 21215 20995
rect 21157 20955 21215 20961
rect 24026 20952 24032 21004
rect 24084 20992 24090 21004
rect 24305 20995 24363 21001
rect 24305 20992 24317 20995
rect 24084 20964 24317 20992
rect 24084 20952 24090 20964
rect 24305 20961 24317 20964
rect 24351 20961 24363 20995
rect 24305 20955 24363 20961
rect 2225 20927 2283 20933
rect 2225 20893 2237 20927
rect 2271 20924 2283 20927
rect 2682 20924 2688 20936
rect 2271 20896 2688 20924
rect 2271 20893 2283 20896
rect 2225 20887 2283 20893
rect 2682 20884 2688 20896
rect 2740 20884 2746 20936
rect 5074 20924 5080 20936
rect 5035 20896 5080 20924
rect 5074 20884 5080 20896
rect 5132 20884 5138 20936
rect 8389 20927 8447 20933
rect 8389 20893 8401 20927
rect 8435 20924 8447 20927
rect 9306 20924 9312 20936
rect 8435 20896 9312 20924
rect 8435 20893 8447 20896
rect 8389 20887 8447 20893
rect 9306 20884 9312 20896
rect 9364 20884 9370 20936
rect 12158 20884 12164 20936
rect 12216 20924 12222 20936
rect 12986 20924 12992 20936
rect 12216 20896 12992 20924
rect 12216 20884 12222 20896
rect 12986 20884 12992 20896
rect 13044 20924 13050 20936
rect 13541 20927 13599 20933
rect 13541 20924 13553 20927
rect 13044 20896 13553 20924
rect 13044 20884 13050 20896
rect 13541 20893 13553 20896
rect 13587 20893 13599 20927
rect 13541 20887 13599 20893
rect 14734 20884 14740 20936
rect 14792 20924 14798 20936
rect 15933 20927 15991 20933
rect 15933 20924 15945 20927
rect 14792 20896 15945 20924
rect 14792 20884 14798 20896
rect 15933 20893 15945 20896
rect 15979 20893 15991 20927
rect 15933 20887 15991 20893
rect 16942 20884 16948 20936
rect 17000 20924 17006 20936
rect 17126 20924 17132 20936
rect 17000 20896 17132 20924
rect 17000 20884 17006 20896
rect 17126 20884 17132 20896
rect 17184 20884 17190 20936
rect 20898 20924 20904 20936
rect 20859 20896 20904 20924
rect 20898 20884 20904 20896
rect 20956 20884 20962 20936
rect 24121 20927 24179 20933
rect 24121 20924 24133 20927
rect 23492 20896 24133 20924
rect 1670 20856 1676 20868
rect 1631 20828 1676 20856
rect 1670 20816 1676 20828
rect 1728 20816 1734 20868
rect 4617 20859 4675 20865
rect 4617 20825 4629 20859
rect 4663 20856 4675 20859
rect 4663 20828 5120 20856
rect 4663 20825 4675 20828
rect 4617 20819 4675 20825
rect 3694 20788 3700 20800
rect 3655 20760 3700 20788
rect 3694 20748 3700 20760
rect 3752 20748 3758 20800
rect 4890 20788 4896 20800
rect 4851 20760 4896 20788
rect 4890 20748 4896 20760
rect 4948 20748 4954 20800
rect 5092 20788 5120 20828
rect 6822 20816 6828 20868
rect 6880 20856 6886 20868
rect 7929 20859 7987 20865
rect 7929 20856 7941 20859
rect 6880 20828 7941 20856
rect 6880 20816 6886 20828
rect 7929 20825 7941 20828
rect 7975 20825 7987 20859
rect 7929 20819 7987 20825
rect 12434 20816 12440 20868
rect 12492 20856 12498 20868
rect 13173 20859 13231 20865
rect 13173 20856 13185 20859
rect 12492 20828 13185 20856
rect 12492 20816 12498 20828
rect 13173 20825 13185 20828
rect 13219 20825 13231 20859
rect 13173 20819 13231 20825
rect 14642 20816 14648 20868
rect 14700 20856 14706 20868
rect 15381 20859 15439 20865
rect 15381 20856 15393 20859
rect 14700 20828 15393 20856
rect 14700 20816 14706 20828
rect 15381 20825 15393 20828
rect 15427 20825 15439 20859
rect 15381 20819 15439 20825
rect 23492 20800 23520 20896
rect 24121 20893 24133 20896
rect 24167 20893 24179 20927
rect 24121 20887 24179 20893
rect 24670 20884 24676 20936
rect 24728 20924 24734 20936
rect 24780 20924 24808 21023
rect 24946 21020 24952 21032
rect 25004 21020 25010 21072
rect 25222 20992 25228 21004
rect 25183 20964 25228 20992
rect 25222 20952 25228 20964
rect 25280 20952 25286 21004
rect 24728 20896 24808 20924
rect 24728 20884 24734 20896
rect 23753 20859 23811 20865
rect 23753 20825 23765 20859
rect 23799 20856 23811 20859
rect 24854 20856 24860 20868
rect 23799 20828 24860 20856
rect 23799 20825 23811 20828
rect 23753 20819 23811 20825
rect 24854 20816 24860 20828
rect 24912 20816 24918 20868
rect 5442 20788 5448 20800
rect 5092 20760 5448 20788
rect 5442 20748 5448 20760
rect 5500 20748 5506 20800
rect 10318 20788 10324 20800
rect 10279 20760 10324 20788
rect 10318 20748 10324 20760
rect 10376 20748 10382 20800
rect 12618 20788 12624 20800
rect 12579 20760 12624 20788
rect 12618 20748 12624 20760
rect 12676 20748 12682 20800
rect 12989 20791 13047 20797
rect 12989 20757 13001 20791
rect 13035 20788 13047 20791
rect 13078 20788 13084 20800
rect 13035 20760 13084 20788
rect 13035 20757 13047 20760
rect 12989 20751 13047 20757
rect 13078 20748 13084 20760
rect 13136 20788 13142 20800
rect 13538 20788 13544 20800
rect 13136 20760 13544 20788
rect 13136 20748 13142 20760
rect 13538 20748 13544 20760
rect 13596 20788 13602 20800
rect 15013 20791 15071 20797
rect 15013 20788 15025 20791
rect 13596 20760 15025 20788
rect 13596 20748 13602 20760
rect 15013 20757 15025 20760
rect 15059 20788 15071 20791
rect 15562 20788 15568 20800
rect 15059 20760 15568 20788
rect 15059 20757 15071 20760
rect 15013 20751 15071 20757
rect 15562 20748 15568 20760
rect 15620 20748 15626 20800
rect 18598 20748 18604 20800
rect 18656 20788 18662 20800
rect 19061 20791 19119 20797
rect 19061 20788 19073 20791
rect 18656 20760 19073 20788
rect 18656 20748 18662 20760
rect 19061 20757 19073 20760
rect 19107 20757 19119 20791
rect 23474 20788 23480 20800
rect 23435 20760 23480 20788
rect 19061 20751 19119 20757
rect 23474 20748 23480 20760
rect 23532 20748 23538 20800
rect 25130 20788 25136 20800
rect 25091 20760 25136 20788
rect 25130 20748 25136 20760
rect 25188 20748 25194 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 2774 20544 2780 20596
rect 2832 20584 2838 20596
rect 3053 20587 3111 20593
rect 3053 20584 3065 20587
rect 2832 20556 3065 20584
rect 2832 20544 2838 20556
rect 3053 20553 3065 20556
rect 3099 20584 3111 20587
rect 3605 20587 3663 20593
rect 3605 20584 3617 20587
rect 3099 20556 3617 20584
rect 3099 20553 3111 20556
rect 3053 20547 3111 20553
rect 3605 20553 3617 20556
rect 3651 20553 3663 20587
rect 5258 20584 5264 20596
rect 5219 20556 5264 20584
rect 3605 20547 3663 20553
rect 5258 20544 5264 20556
rect 5316 20544 5322 20596
rect 7282 20584 7288 20596
rect 7195 20556 7288 20584
rect 7282 20544 7288 20556
rect 7340 20584 7346 20596
rect 8110 20584 8116 20596
rect 7340 20556 8116 20584
rect 7340 20544 7346 20556
rect 8110 20544 8116 20556
rect 8168 20544 8174 20596
rect 9306 20584 9312 20596
rect 9267 20556 9312 20584
rect 9306 20544 9312 20556
rect 9364 20544 9370 20596
rect 11885 20587 11943 20593
rect 11885 20553 11897 20587
rect 11931 20584 11943 20587
rect 12342 20584 12348 20596
rect 11931 20556 12348 20584
rect 11931 20553 11943 20556
rect 11885 20547 11943 20553
rect 12342 20544 12348 20556
rect 12400 20544 12406 20596
rect 13265 20587 13323 20593
rect 13265 20553 13277 20587
rect 13311 20584 13323 20587
rect 13354 20584 13360 20596
rect 13311 20556 13360 20584
rect 13311 20553 13323 20556
rect 13265 20547 13323 20553
rect 13354 20544 13360 20556
rect 13412 20544 13418 20596
rect 14090 20544 14096 20596
rect 14148 20584 14154 20596
rect 14734 20584 14740 20596
rect 14148 20556 14740 20584
rect 14148 20544 14154 20556
rect 14734 20544 14740 20556
rect 14792 20584 14798 20596
rect 15105 20587 15163 20593
rect 15105 20584 15117 20587
rect 14792 20556 15117 20584
rect 14792 20544 14798 20556
rect 15105 20553 15117 20556
rect 15151 20553 15163 20587
rect 18322 20584 18328 20596
rect 18283 20556 18328 20584
rect 15105 20547 15163 20553
rect 18322 20544 18328 20556
rect 18380 20544 18386 20596
rect 20990 20544 20996 20596
rect 21048 20584 21054 20596
rect 21177 20587 21235 20593
rect 21177 20584 21189 20587
rect 21048 20556 21189 20584
rect 21048 20544 21054 20556
rect 21177 20553 21189 20556
rect 21223 20553 21235 20587
rect 22186 20584 22192 20596
rect 22147 20556 22192 20584
rect 21177 20547 21235 20553
rect 22186 20544 22192 20556
rect 22244 20544 22250 20596
rect 22649 20587 22707 20593
rect 22649 20553 22661 20587
rect 22695 20584 22707 20587
rect 22830 20584 22836 20596
rect 22695 20556 22836 20584
rect 22695 20553 22707 20556
rect 22649 20547 22707 20553
rect 22830 20544 22836 20556
rect 22888 20544 22894 20596
rect 25222 20544 25228 20596
rect 25280 20584 25286 20596
rect 25869 20587 25927 20593
rect 25869 20584 25881 20587
rect 25280 20556 25881 20584
rect 25280 20544 25286 20556
rect 25869 20553 25881 20556
rect 25915 20553 25927 20587
rect 25869 20547 25927 20553
rect 2866 20476 2872 20528
rect 2924 20516 2930 20528
rect 3973 20519 4031 20525
rect 3973 20516 3985 20519
rect 2924 20488 3985 20516
rect 2924 20476 2930 20488
rect 3973 20485 3985 20488
rect 4019 20485 4031 20519
rect 3973 20479 4031 20485
rect 16301 20519 16359 20525
rect 16301 20485 16313 20519
rect 16347 20485 16359 20519
rect 16301 20479 16359 20485
rect 1394 20408 1400 20460
rect 1452 20448 1458 20460
rect 1673 20451 1731 20457
rect 1673 20448 1685 20451
rect 1452 20420 1685 20448
rect 1452 20408 1458 20420
rect 1673 20417 1685 20420
rect 1719 20417 1731 20451
rect 1673 20411 1731 20417
rect 5442 20408 5448 20460
rect 5500 20448 5506 20460
rect 5721 20451 5779 20457
rect 5721 20448 5733 20451
rect 5500 20420 5733 20448
rect 5500 20408 5506 20420
rect 5721 20417 5733 20420
rect 5767 20448 5779 20451
rect 5810 20448 5816 20460
rect 5767 20420 5816 20448
rect 5767 20417 5779 20420
rect 5721 20411 5779 20417
rect 5810 20408 5816 20420
rect 5868 20408 5874 20460
rect 6273 20451 6331 20457
rect 6273 20417 6285 20451
rect 6319 20448 6331 20451
rect 6319 20420 7512 20448
rect 6319 20417 6331 20420
rect 6273 20411 6331 20417
rect 1940 20383 1998 20389
rect 1940 20349 1952 20383
rect 1986 20380 1998 20383
rect 2222 20380 2228 20392
rect 1986 20352 2228 20380
rect 1986 20349 1998 20352
rect 1940 20343 1998 20349
rect 2222 20340 2228 20352
rect 2280 20380 2286 20392
rect 3694 20380 3700 20392
rect 2280 20352 3700 20380
rect 2280 20340 2286 20352
rect 3694 20340 3700 20352
rect 3752 20340 3758 20392
rect 6457 20383 6515 20389
rect 6457 20349 6469 20383
rect 6503 20380 6515 20383
rect 6638 20380 6644 20392
rect 6503 20352 6644 20380
rect 6503 20349 6515 20352
rect 6457 20343 6515 20349
rect 6638 20340 6644 20352
rect 6696 20380 6702 20392
rect 7377 20383 7435 20389
rect 7377 20380 7389 20383
rect 6696 20352 7389 20380
rect 6696 20340 6702 20352
rect 7377 20349 7389 20352
rect 7423 20349 7435 20383
rect 7484 20380 7512 20420
rect 7650 20389 7656 20392
rect 7644 20380 7656 20389
rect 7484 20352 7656 20380
rect 7377 20343 7435 20349
rect 7644 20343 7656 20352
rect 7650 20340 7656 20343
rect 7708 20340 7714 20392
rect 9769 20383 9827 20389
rect 9769 20349 9781 20383
rect 9815 20380 9827 20383
rect 9858 20380 9864 20392
rect 9815 20352 9864 20380
rect 9815 20349 9827 20352
rect 9769 20343 9827 20349
rect 9858 20340 9864 20352
rect 9916 20340 9922 20392
rect 12158 20380 12164 20392
rect 10060 20352 12164 20380
rect 2958 20272 2964 20324
rect 3016 20312 3022 20324
rect 4157 20315 4215 20321
rect 4157 20312 4169 20315
rect 3016 20284 4169 20312
rect 3016 20272 3022 20284
rect 4157 20281 4169 20284
rect 4203 20281 4215 20315
rect 4157 20275 4215 20281
rect 4709 20315 4767 20321
rect 4709 20281 4721 20315
rect 4755 20312 4767 20315
rect 4890 20312 4896 20324
rect 4755 20284 4896 20312
rect 4755 20281 4767 20284
rect 4709 20275 4767 20281
rect 4890 20272 4896 20284
rect 4948 20312 4954 20324
rect 5813 20315 5871 20321
rect 5813 20312 5825 20315
rect 4948 20284 5825 20312
rect 4948 20272 4954 20284
rect 5813 20281 5825 20284
rect 5859 20312 5871 20315
rect 5859 20284 7512 20312
rect 5859 20281 5871 20284
rect 5813 20275 5871 20281
rect 4246 20204 4252 20256
rect 4304 20244 4310 20256
rect 4985 20247 5043 20253
rect 4985 20244 4997 20247
rect 4304 20216 4997 20244
rect 4304 20204 4310 20216
rect 4985 20213 4997 20216
rect 5031 20244 5043 20247
rect 5074 20244 5080 20256
rect 5031 20216 5080 20244
rect 5031 20213 5043 20216
rect 4985 20207 5043 20213
rect 5074 20204 5080 20216
rect 5132 20204 5138 20256
rect 5718 20244 5724 20256
rect 5679 20216 5724 20244
rect 5718 20204 5724 20216
rect 5776 20204 5782 20256
rect 6270 20204 6276 20256
rect 6328 20244 6334 20256
rect 6457 20247 6515 20253
rect 6457 20244 6469 20247
rect 6328 20216 6469 20244
rect 6328 20204 6334 20216
rect 6457 20213 6469 20216
rect 6503 20244 6515 20247
rect 6549 20247 6607 20253
rect 6549 20244 6561 20247
rect 6503 20216 6561 20244
rect 6503 20213 6515 20216
rect 6457 20207 6515 20213
rect 6549 20213 6561 20216
rect 6595 20213 6607 20247
rect 7484 20244 7512 20284
rect 8757 20247 8815 20253
rect 8757 20244 8769 20247
rect 7484 20216 8769 20244
rect 6549 20207 6607 20213
rect 8757 20213 8769 20216
rect 8803 20213 8815 20247
rect 8757 20207 8815 20213
rect 9582 20204 9588 20256
rect 9640 20244 9646 20256
rect 10060 20244 10088 20352
rect 12158 20340 12164 20352
rect 12216 20340 12222 20392
rect 13630 20380 13636 20392
rect 13591 20352 13636 20380
rect 13630 20340 13636 20352
rect 13688 20380 13694 20392
rect 13725 20383 13783 20389
rect 13725 20380 13737 20383
rect 13688 20352 13737 20380
rect 13688 20340 13694 20352
rect 13725 20349 13737 20352
rect 13771 20349 13783 20383
rect 13725 20343 13783 20349
rect 13814 20340 13820 20392
rect 13872 20380 13878 20392
rect 13981 20383 14039 20389
rect 13981 20380 13993 20383
rect 13872 20352 13993 20380
rect 13872 20340 13878 20352
rect 13981 20349 13993 20352
rect 14027 20349 14039 20383
rect 13981 20343 14039 20349
rect 14550 20340 14556 20392
rect 14608 20380 14614 20392
rect 16316 20380 16344 20479
rect 22646 20408 22652 20460
rect 22704 20448 22710 20460
rect 23017 20451 23075 20457
rect 23017 20448 23029 20451
rect 22704 20420 23029 20448
rect 22704 20408 22710 20420
rect 23017 20417 23029 20420
rect 23063 20448 23075 20451
rect 23063 20420 24072 20448
rect 23063 20417 23075 20420
rect 23017 20411 23075 20417
rect 24044 20392 24072 20420
rect 16574 20380 16580 20392
rect 14608 20352 16344 20380
rect 16535 20352 16580 20380
rect 14608 20340 14614 20352
rect 16574 20340 16580 20352
rect 16632 20340 16638 20392
rect 16942 20340 16948 20392
rect 17000 20380 17006 20392
rect 17221 20383 17279 20389
rect 17221 20380 17233 20383
rect 17000 20352 17233 20380
rect 17000 20340 17006 20352
rect 17221 20349 17233 20352
rect 17267 20349 17279 20383
rect 17221 20343 17279 20349
rect 17865 20383 17923 20389
rect 17865 20349 17877 20383
rect 17911 20380 17923 20383
rect 19521 20383 19579 20389
rect 17911 20352 18920 20380
rect 17911 20349 17923 20352
rect 17865 20343 17923 20349
rect 10128 20315 10186 20321
rect 10128 20281 10140 20315
rect 10174 20312 10186 20315
rect 10318 20312 10324 20324
rect 10174 20284 10324 20312
rect 10174 20281 10186 20284
rect 10128 20275 10186 20281
rect 10318 20272 10324 20284
rect 10376 20272 10382 20324
rect 12713 20315 12771 20321
rect 12713 20281 12725 20315
rect 12759 20312 12771 20315
rect 15010 20312 15016 20324
rect 12759 20284 15016 20312
rect 12759 20281 12771 20284
rect 12713 20275 12771 20281
rect 15010 20272 15016 20284
rect 15068 20272 15074 20324
rect 16850 20312 16856 20324
rect 15212 20284 16160 20312
rect 16811 20284 16856 20312
rect 9640 20216 10088 20244
rect 9640 20204 9646 20216
rect 10778 20204 10784 20256
rect 10836 20244 10842 20256
rect 11241 20247 11299 20253
rect 11241 20244 11253 20247
rect 10836 20216 11253 20244
rect 10836 20204 10842 20216
rect 11241 20213 11253 20216
rect 11287 20244 11299 20247
rect 11330 20244 11336 20256
rect 11287 20216 11336 20244
rect 11287 20213 11299 20216
rect 11241 20207 11299 20213
rect 11330 20204 11336 20216
rect 11388 20204 11394 20256
rect 14642 20204 14648 20256
rect 14700 20244 14706 20256
rect 15212 20244 15240 20284
rect 15746 20244 15752 20256
rect 14700 20216 15240 20244
rect 15707 20216 15752 20244
rect 14700 20204 14706 20216
rect 15746 20204 15752 20216
rect 15804 20204 15810 20256
rect 16132 20253 16160 20284
rect 16850 20272 16856 20284
rect 16908 20272 16914 20324
rect 18046 20312 18052 20324
rect 16960 20284 18052 20312
rect 16117 20247 16175 20253
rect 16117 20213 16129 20247
rect 16163 20244 16175 20247
rect 16761 20247 16819 20253
rect 16761 20244 16773 20247
rect 16163 20216 16773 20244
rect 16163 20213 16175 20216
rect 16117 20207 16175 20213
rect 16761 20213 16773 20216
rect 16807 20244 16819 20247
rect 16960 20244 16988 20284
rect 18046 20272 18052 20284
rect 18104 20272 18110 20324
rect 18598 20312 18604 20324
rect 18559 20284 18604 20312
rect 18598 20272 18604 20284
rect 18656 20272 18662 20324
rect 18892 20321 18920 20352
rect 19521 20349 19533 20383
rect 19567 20380 19579 20383
rect 19797 20383 19855 20389
rect 19797 20380 19809 20383
rect 19567 20352 19809 20380
rect 19567 20349 19579 20352
rect 19521 20343 19579 20349
rect 19797 20349 19809 20352
rect 19843 20349 19855 20383
rect 19797 20343 19855 20349
rect 22094 20340 22100 20392
rect 22152 20380 22158 20392
rect 22465 20383 22523 20389
rect 22465 20380 22477 20383
rect 22152 20352 22477 20380
rect 22152 20340 22158 20352
rect 22465 20349 22477 20352
rect 22511 20349 22523 20383
rect 22465 20343 22523 20349
rect 23477 20383 23535 20389
rect 23477 20349 23489 20383
rect 23523 20380 23535 20383
rect 23750 20380 23756 20392
rect 23523 20352 23756 20380
rect 23523 20349 23535 20352
rect 23477 20343 23535 20349
rect 23750 20340 23756 20352
rect 23808 20380 23814 20392
rect 23937 20383 23995 20389
rect 23937 20380 23949 20383
rect 23808 20352 23949 20380
rect 23808 20340 23814 20352
rect 23937 20349 23949 20352
rect 23983 20349 23995 20383
rect 23937 20343 23995 20349
rect 24026 20340 24032 20392
rect 24084 20380 24090 20392
rect 24193 20383 24251 20389
rect 24193 20380 24205 20383
rect 24084 20352 24205 20380
rect 24084 20340 24090 20352
rect 24193 20349 24205 20352
rect 24239 20349 24251 20383
rect 24193 20343 24251 20349
rect 18877 20315 18935 20321
rect 18877 20281 18889 20315
rect 18923 20312 18935 20315
rect 19337 20315 19395 20321
rect 19337 20312 19349 20315
rect 18923 20284 19349 20312
rect 18923 20281 18935 20284
rect 18877 20275 18935 20281
rect 19337 20281 19349 20284
rect 19383 20312 19395 20315
rect 20064 20315 20122 20321
rect 20064 20312 20076 20315
rect 19383 20284 20076 20312
rect 19383 20281 19395 20284
rect 19337 20275 19395 20281
rect 20064 20281 20076 20284
rect 20110 20312 20122 20315
rect 20622 20312 20628 20324
rect 20110 20284 20628 20312
rect 20110 20281 20122 20284
rect 20064 20275 20122 20281
rect 20622 20272 20628 20284
rect 20680 20272 20686 20324
rect 16807 20216 16988 20244
rect 18785 20247 18843 20253
rect 16807 20213 16819 20216
rect 16761 20207 16819 20213
rect 18785 20213 18797 20247
rect 18831 20244 18843 20247
rect 19058 20244 19064 20256
rect 18831 20216 19064 20244
rect 18831 20213 18843 20216
rect 18785 20207 18843 20213
rect 19058 20204 19064 20216
rect 19116 20204 19122 20256
rect 19521 20247 19579 20253
rect 19521 20213 19533 20247
rect 19567 20244 19579 20247
rect 19705 20247 19763 20253
rect 19705 20244 19717 20247
rect 19567 20216 19717 20244
rect 19567 20213 19579 20216
rect 19521 20207 19579 20213
rect 19705 20213 19717 20216
rect 19751 20244 19763 20247
rect 20254 20244 20260 20256
rect 19751 20216 20260 20244
rect 19751 20213 19763 20216
rect 19705 20207 19763 20213
rect 20254 20204 20260 20216
rect 20312 20244 20318 20256
rect 20898 20244 20904 20256
rect 20312 20216 20904 20244
rect 20312 20204 20318 20216
rect 20898 20204 20904 20216
rect 20956 20244 20962 20256
rect 21821 20247 21879 20253
rect 21821 20244 21833 20247
rect 20956 20216 21833 20244
rect 20956 20204 20962 20216
rect 21821 20213 21833 20216
rect 21867 20244 21879 20247
rect 22370 20244 22376 20256
rect 21867 20216 22376 20244
rect 21867 20213 21879 20216
rect 21821 20207 21879 20213
rect 22370 20204 22376 20216
rect 22428 20204 22434 20256
rect 25317 20247 25375 20253
rect 25317 20213 25329 20247
rect 25363 20244 25375 20247
rect 25498 20244 25504 20256
rect 25363 20216 25504 20244
rect 25363 20213 25375 20216
rect 25317 20207 25375 20213
rect 25498 20204 25504 20216
rect 25556 20204 25562 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1394 20000 1400 20052
rect 1452 20040 1458 20052
rect 1673 20043 1731 20049
rect 1673 20040 1685 20043
rect 1452 20012 1685 20040
rect 1452 20000 1458 20012
rect 1673 20009 1685 20012
rect 1719 20009 1731 20043
rect 2038 20040 2044 20052
rect 1999 20012 2044 20040
rect 1673 20003 1731 20009
rect 2038 20000 2044 20012
rect 2096 20000 2102 20052
rect 3513 20043 3571 20049
rect 3513 20009 3525 20043
rect 3559 20040 3571 20043
rect 3694 20040 3700 20052
rect 3559 20012 3700 20040
rect 3559 20009 3571 20012
rect 3513 20003 3571 20009
rect 3694 20000 3700 20012
rect 3752 20000 3758 20052
rect 3786 20000 3792 20052
rect 3844 20040 3850 20052
rect 3844 20012 3889 20040
rect 3844 20000 3850 20012
rect 5718 20000 5724 20052
rect 5776 20040 5782 20052
rect 6089 20043 6147 20049
rect 6089 20040 6101 20043
rect 5776 20012 6101 20040
rect 5776 20000 5782 20012
rect 6089 20009 6101 20012
rect 6135 20040 6147 20043
rect 6822 20040 6828 20052
rect 6135 20012 6828 20040
rect 6135 20009 6147 20012
rect 6089 20003 6147 20009
rect 6822 20000 6828 20012
rect 6880 20000 6886 20052
rect 9766 20000 9772 20052
rect 9824 20040 9830 20052
rect 10873 20043 10931 20049
rect 10873 20040 10885 20043
rect 9824 20012 10885 20040
rect 9824 20000 9830 20012
rect 10873 20009 10885 20012
rect 10919 20009 10931 20043
rect 10873 20003 10931 20009
rect 13725 20043 13783 20049
rect 13725 20009 13737 20043
rect 13771 20040 13783 20043
rect 13814 20040 13820 20052
rect 13771 20012 13820 20040
rect 13771 20009 13783 20012
rect 13725 20003 13783 20009
rect 13814 20000 13820 20012
rect 13872 20000 13878 20052
rect 14734 20040 14740 20052
rect 14695 20012 14740 20040
rect 14734 20000 14740 20012
rect 14792 20000 14798 20052
rect 15102 20040 15108 20052
rect 15063 20012 15108 20040
rect 15102 20000 15108 20012
rect 15160 20000 15166 20052
rect 15838 20000 15844 20052
rect 15896 20040 15902 20052
rect 16669 20043 16727 20049
rect 16669 20040 16681 20043
rect 15896 20012 16681 20040
rect 15896 20000 15902 20012
rect 2774 19932 2780 19984
rect 2832 19972 2838 19984
rect 2961 19975 3019 19981
rect 2961 19972 2973 19975
rect 2832 19944 2973 19972
rect 2832 19932 2838 19944
rect 2961 19941 2973 19944
rect 3007 19972 3019 19975
rect 6365 19975 6423 19981
rect 6365 19972 6377 19975
rect 3007 19944 6377 19972
rect 3007 19941 3019 19944
rect 2961 19935 3019 19941
rect 6365 19941 6377 19944
rect 6411 19941 6423 19975
rect 8386 19972 8392 19984
rect 8347 19944 8392 19972
rect 6365 19935 6423 19941
rect 8386 19932 8392 19944
rect 8444 19932 8450 19984
rect 8478 19932 8484 19984
rect 8536 19972 8542 19984
rect 8536 19944 8581 19972
rect 8536 19932 8542 19944
rect 9674 19932 9680 19984
rect 9732 19972 9738 19984
rect 10689 19975 10747 19981
rect 10689 19972 10701 19975
rect 9732 19944 10701 19972
rect 9732 19932 9738 19944
rect 4065 19907 4123 19913
rect 4065 19873 4077 19907
rect 4111 19904 4123 19907
rect 4154 19904 4160 19916
rect 4111 19876 4160 19904
rect 4111 19873 4123 19876
rect 4065 19867 4123 19873
rect 4154 19864 4160 19876
rect 4212 19864 4218 19916
rect 4338 19913 4344 19916
rect 4332 19867 4344 19913
rect 4396 19904 4402 19916
rect 4396 19876 4432 19904
rect 4338 19864 4344 19867
rect 4396 19864 4402 19876
rect 5534 19864 5540 19916
rect 5592 19904 5598 19916
rect 6178 19904 6184 19916
rect 5592 19876 6184 19904
rect 5592 19864 5598 19876
rect 6178 19864 6184 19876
rect 6236 19904 6242 19916
rect 6549 19907 6607 19913
rect 6549 19904 6561 19907
rect 6236 19876 6561 19904
rect 6236 19864 6242 19876
rect 6549 19873 6561 19876
rect 6595 19873 6607 19907
rect 6549 19867 6607 19873
rect 2590 19796 2596 19848
rect 2648 19836 2654 19848
rect 2958 19836 2964 19848
rect 2648 19808 2964 19836
rect 2648 19796 2654 19808
rect 2958 19796 2964 19808
rect 3016 19796 3022 19848
rect 3053 19839 3111 19845
rect 3053 19805 3065 19839
rect 3099 19836 3111 19839
rect 3694 19836 3700 19848
rect 3099 19808 3700 19836
rect 3099 19805 3111 19808
rect 3053 19799 3111 19805
rect 3694 19796 3700 19808
rect 3752 19836 3758 19848
rect 6730 19836 6736 19848
rect 3752 19808 4016 19836
rect 6691 19808 6736 19836
rect 3752 19796 3758 19808
rect 2406 19728 2412 19780
rect 2464 19768 2470 19780
rect 2501 19771 2559 19777
rect 2501 19768 2513 19771
rect 2464 19740 2513 19768
rect 2464 19728 2470 19740
rect 2501 19737 2513 19740
rect 2547 19737 2559 19771
rect 2501 19731 2559 19737
rect 3988 19700 4016 19808
rect 6730 19796 6736 19808
rect 6788 19796 6794 19848
rect 8389 19839 8447 19845
rect 8389 19805 8401 19839
rect 8435 19836 8447 19839
rect 8570 19836 8576 19848
rect 8435 19808 8576 19836
rect 8435 19805 8447 19808
rect 8389 19799 8447 19805
rect 8570 19796 8576 19808
rect 8628 19796 8634 19848
rect 9784 19836 9812 19944
rect 10689 19941 10701 19944
rect 10735 19941 10747 19975
rect 10689 19935 10747 19941
rect 12612 19975 12670 19981
rect 12612 19941 12624 19975
rect 12658 19972 12670 19975
rect 13538 19972 13544 19984
rect 12658 19944 13544 19972
rect 12658 19941 12670 19944
rect 12612 19935 12670 19941
rect 13538 19932 13544 19944
rect 13596 19932 13602 19984
rect 16224 19981 16252 20012
rect 16669 20009 16681 20012
rect 16715 20040 16727 20043
rect 16850 20040 16856 20052
rect 16715 20012 16856 20040
rect 16715 20009 16727 20012
rect 16669 20003 16727 20009
rect 16850 20000 16856 20012
rect 16908 20000 16914 20052
rect 17034 20040 17040 20052
rect 16995 20012 17040 20040
rect 17034 20000 17040 20012
rect 17092 20000 17098 20052
rect 17954 20000 17960 20052
rect 18012 20040 18018 20052
rect 18509 20043 18567 20049
rect 18509 20040 18521 20043
rect 18012 20012 18521 20040
rect 18012 20000 18018 20012
rect 18509 20009 18521 20012
rect 18555 20009 18567 20043
rect 18509 20003 18567 20009
rect 19613 20043 19671 20049
rect 19613 20009 19625 20043
rect 19659 20040 19671 20043
rect 20530 20040 20536 20052
rect 19659 20012 20536 20040
rect 19659 20009 19671 20012
rect 19613 20003 19671 20009
rect 20530 20000 20536 20012
rect 20588 20000 20594 20052
rect 21085 20043 21143 20049
rect 21085 20009 21097 20043
rect 21131 20040 21143 20043
rect 21174 20040 21180 20052
rect 21131 20012 21180 20040
rect 21131 20009 21143 20012
rect 21085 20003 21143 20009
rect 21174 20000 21180 20012
rect 21232 20000 21238 20052
rect 22094 20000 22100 20052
rect 22152 20040 22158 20052
rect 22189 20043 22247 20049
rect 22189 20040 22201 20043
rect 22152 20012 22201 20040
rect 22152 20000 22158 20012
rect 22189 20009 22201 20012
rect 22235 20009 22247 20043
rect 22189 20003 22247 20009
rect 24210 20000 24216 20052
rect 24268 20040 24274 20052
rect 24673 20043 24731 20049
rect 24673 20040 24685 20043
rect 24268 20012 24685 20040
rect 24268 20000 24274 20012
rect 24673 20009 24685 20012
rect 24719 20009 24731 20043
rect 25406 20040 25412 20052
rect 25367 20012 25412 20040
rect 24673 20003 24731 20009
rect 25406 20000 25412 20012
rect 25464 20000 25470 20052
rect 16117 19975 16175 19981
rect 16117 19941 16129 19975
rect 16163 19941 16175 19975
rect 16117 19935 16175 19941
rect 16209 19975 16267 19981
rect 16209 19941 16221 19975
rect 16255 19941 16267 19975
rect 16209 19935 16267 19941
rect 9858 19864 9864 19916
rect 9916 19904 9922 19916
rect 9953 19907 10011 19913
rect 9953 19904 9965 19907
rect 9916 19876 9965 19904
rect 9916 19864 9922 19876
rect 9953 19873 9965 19876
rect 9999 19904 10011 19907
rect 11882 19904 11888 19916
rect 9999 19876 11888 19904
rect 9999 19873 10011 19876
rect 9953 19867 10011 19873
rect 11882 19864 11888 19876
rect 11940 19904 11946 19916
rect 12345 19907 12403 19913
rect 12345 19904 12357 19907
rect 11940 19876 12357 19904
rect 11940 19864 11946 19876
rect 12345 19873 12357 19876
rect 12391 19904 12403 19907
rect 13630 19904 13636 19916
rect 12391 19876 13636 19904
rect 12391 19873 12403 19876
rect 12345 19867 12403 19873
rect 13630 19864 13636 19876
rect 13688 19864 13694 19916
rect 16132 19904 16160 19935
rect 17126 19932 17132 19984
rect 17184 19972 17190 19984
rect 17396 19975 17454 19981
rect 17396 19972 17408 19975
rect 17184 19944 17408 19972
rect 17184 19932 17190 19944
rect 17396 19941 17408 19944
rect 17442 19972 17454 19975
rect 17862 19972 17868 19984
rect 17442 19944 17868 19972
rect 17442 19941 17454 19944
rect 17396 19935 17454 19941
rect 17862 19932 17868 19944
rect 17920 19932 17926 19984
rect 19334 19932 19340 19984
rect 19392 19972 19398 19984
rect 20441 19975 20499 19981
rect 20441 19972 20453 19975
rect 19392 19944 20453 19972
rect 19392 19932 19398 19944
rect 20441 19941 20453 19944
rect 20487 19941 20499 19975
rect 20441 19935 20499 19941
rect 20990 19932 20996 19984
rect 21048 19972 21054 19984
rect 21453 19975 21511 19981
rect 21453 19972 21465 19975
rect 21048 19944 21465 19972
rect 21048 19932 21054 19944
rect 21453 19941 21465 19944
rect 21499 19941 21511 19975
rect 23750 19972 23756 19984
rect 21453 19935 21511 19941
rect 22388 19944 23756 19972
rect 22388 19916 22416 19944
rect 23750 19932 23756 19944
rect 23808 19932 23814 19984
rect 24026 19932 24032 19984
rect 24084 19972 24090 19984
rect 24305 19975 24363 19981
rect 24305 19972 24317 19975
rect 24084 19944 24317 19972
rect 24084 19932 24090 19944
rect 24305 19941 24317 19944
rect 24351 19941 24363 19975
rect 24305 19935 24363 19941
rect 24854 19932 24860 19984
rect 24912 19972 24918 19984
rect 25225 19975 25283 19981
rect 25225 19972 25237 19975
rect 24912 19944 25237 19972
rect 24912 19932 24918 19944
rect 25225 19941 25237 19944
rect 25271 19941 25283 19975
rect 25225 19935 25283 19941
rect 16758 19904 16764 19916
rect 16132 19876 16764 19904
rect 16758 19864 16764 19876
rect 16816 19864 16822 19916
rect 20901 19907 20959 19913
rect 20901 19904 20913 19907
rect 20824 19876 20913 19904
rect 20824 19848 20852 19876
rect 20901 19873 20913 19876
rect 20947 19904 20959 19907
rect 21726 19904 21732 19916
rect 20947 19876 21732 19904
rect 20947 19873 20959 19876
rect 20901 19867 20959 19873
rect 21726 19864 21732 19876
rect 21784 19864 21790 19916
rect 22370 19904 22376 19916
rect 22283 19876 22376 19904
rect 22370 19864 22376 19876
rect 22428 19864 22434 19916
rect 22640 19907 22698 19913
rect 22640 19873 22652 19907
rect 22686 19904 22698 19907
rect 23014 19904 23020 19916
rect 22686 19876 23020 19904
rect 22686 19873 22698 19876
rect 22640 19867 22698 19873
rect 23014 19864 23020 19876
rect 23072 19864 23078 19916
rect 10134 19836 10140 19848
rect 9784 19808 10140 19836
rect 10134 19796 10140 19808
rect 10192 19796 10198 19848
rect 10965 19839 11023 19845
rect 10965 19805 10977 19839
rect 11011 19836 11023 19839
rect 16117 19839 16175 19845
rect 11011 19808 11376 19836
rect 11011 19805 11023 19808
rect 10965 19799 11023 19805
rect 5810 19728 5816 19780
rect 5868 19768 5874 19780
rect 7929 19771 7987 19777
rect 7929 19768 7941 19771
rect 5868 19740 7941 19768
rect 5868 19728 5874 19740
rect 7929 19737 7941 19740
rect 7975 19737 7987 19771
rect 7929 19731 7987 19737
rect 10413 19771 10471 19777
rect 10413 19737 10425 19771
rect 10459 19768 10471 19771
rect 10870 19768 10876 19780
rect 10459 19740 10876 19768
rect 10459 19737 10471 19740
rect 10413 19731 10471 19737
rect 10870 19728 10876 19740
rect 10928 19728 10934 19780
rect 11348 19712 11376 19808
rect 16117 19805 16129 19839
rect 16163 19836 16175 19839
rect 16298 19836 16304 19848
rect 16163 19808 16304 19836
rect 16163 19805 16175 19808
rect 16117 19799 16175 19805
rect 16298 19796 16304 19808
rect 16356 19796 16362 19848
rect 17034 19796 17040 19848
rect 17092 19836 17098 19848
rect 17129 19839 17187 19845
rect 17129 19836 17141 19839
rect 17092 19808 17141 19836
rect 17092 19796 17098 19808
rect 17129 19805 17141 19808
rect 17175 19805 17187 19839
rect 17129 19799 17187 19805
rect 20806 19796 20812 19848
rect 20864 19796 20870 19848
rect 25498 19836 25504 19848
rect 25459 19808 25504 19836
rect 25498 19796 25504 19808
rect 25556 19796 25562 19848
rect 5445 19703 5503 19709
rect 5445 19700 5457 19703
rect 3988 19672 5457 19700
rect 5445 19669 5457 19672
rect 5491 19669 5503 19703
rect 5445 19663 5503 19669
rect 7374 19660 7380 19712
rect 7432 19700 7438 19712
rect 7558 19700 7564 19712
rect 7432 19672 7564 19700
rect 7432 19660 7438 19672
rect 7558 19660 7564 19672
rect 7616 19660 7622 19712
rect 9122 19700 9128 19712
rect 9083 19672 9128 19700
rect 9122 19660 9128 19672
rect 9180 19660 9186 19712
rect 11330 19700 11336 19712
rect 11291 19672 11336 19700
rect 11330 19660 11336 19672
rect 11388 19660 11394 19712
rect 12066 19660 12072 19712
rect 12124 19700 12130 19712
rect 12161 19703 12219 19709
rect 12161 19700 12173 19703
rect 12124 19672 12173 19700
rect 12124 19660 12130 19672
rect 12161 19669 12173 19672
rect 12207 19669 12219 19703
rect 12161 19663 12219 19669
rect 15562 19660 15568 19712
rect 15620 19700 15626 19712
rect 15657 19703 15715 19709
rect 15657 19700 15669 19703
rect 15620 19672 15669 19700
rect 15620 19660 15626 19672
rect 15657 19669 15669 19672
rect 15703 19669 15715 19703
rect 19058 19700 19064 19712
rect 19019 19672 19064 19700
rect 15657 19663 15715 19669
rect 19058 19660 19064 19672
rect 19116 19660 19122 19712
rect 20162 19700 20168 19712
rect 20123 19672 20168 19700
rect 20162 19660 20168 19672
rect 20220 19660 20226 19712
rect 23382 19660 23388 19712
rect 23440 19700 23446 19712
rect 23753 19703 23811 19709
rect 23753 19700 23765 19703
rect 23440 19672 23765 19700
rect 23440 19660 23446 19672
rect 23753 19669 23765 19672
rect 23799 19669 23811 19703
rect 23753 19663 23811 19669
rect 24949 19703 25007 19709
rect 24949 19669 24961 19703
rect 24995 19700 25007 19703
rect 25866 19700 25872 19712
rect 24995 19672 25872 19700
rect 24995 19669 25007 19672
rect 24949 19663 25007 19669
rect 25866 19660 25872 19672
rect 25924 19660 25930 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 1394 19456 1400 19508
rect 1452 19496 1458 19508
rect 1949 19499 2007 19505
rect 1949 19496 1961 19499
rect 1452 19468 1961 19496
rect 1452 19456 1458 19468
rect 1949 19465 1961 19468
rect 1995 19465 2007 19499
rect 6178 19496 6184 19508
rect 6139 19468 6184 19496
rect 1949 19459 2007 19465
rect 1964 19360 1992 19459
rect 6178 19456 6184 19468
rect 6236 19456 6242 19508
rect 8478 19456 8484 19508
rect 8536 19496 8542 19508
rect 8849 19499 8907 19505
rect 8849 19496 8861 19499
rect 8536 19468 8861 19496
rect 8536 19456 8542 19468
rect 8849 19465 8861 19468
rect 8895 19465 8907 19499
rect 8849 19459 8907 19465
rect 9766 19456 9772 19508
rect 9824 19496 9830 19508
rect 10229 19499 10287 19505
rect 10229 19496 10241 19499
rect 9824 19468 10241 19496
rect 9824 19456 9830 19468
rect 10229 19465 10241 19468
rect 10275 19465 10287 19499
rect 10229 19459 10287 19465
rect 10505 19499 10563 19505
rect 10505 19465 10517 19499
rect 10551 19496 10563 19499
rect 10962 19496 10968 19508
rect 10551 19468 10968 19496
rect 10551 19465 10563 19468
rect 10505 19459 10563 19465
rect 10962 19456 10968 19468
rect 11020 19456 11026 19508
rect 11882 19456 11888 19508
rect 11940 19496 11946 19508
rect 12161 19499 12219 19505
rect 12161 19496 12173 19499
rect 11940 19468 12173 19496
rect 11940 19456 11946 19468
rect 12161 19465 12173 19468
rect 12207 19465 12219 19499
rect 12161 19459 12219 19465
rect 13909 19499 13967 19505
rect 13909 19465 13921 19499
rect 13955 19496 13967 19499
rect 14090 19496 14096 19508
rect 13955 19468 14096 19496
rect 13955 19465 13967 19468
rect 13909 19459 13967 19465
rect 14090 19456 14096 19468
rect 14148 19456 14154 19508
rect 19981 19499 20039 19505
rect 19981 19465 19993 19499
rect 20027 19496 20039 19499
rect 20254 19496 20260 19508
rect 20027 19468 20260 19496
rect 20027 19465 20039 19468
rect 19981 19459 20039 19465
rect 4157 19431 4215 19437
rect 4157 19397 4169 19431
rect 4203 19428 4215 19431
rect 4246 19428 4252 19440
rect 4203 19400 4252 19428
rect 4203 19397 4215 19400
rect 4157 19391 4215 19397
rect 4246 19388 4252 19400
rect 4304 19388 4310 19440
rect 2133 19363 2191 19369
rect 2133 19360 2145 19363
rect 1964 19332 2145 19360
rect 2133 19329 2145 19332
rect 2179 19329 2191 19363
rect 2133 19323 2191 19329
rect 3786 19320 3792 19372
rect 3844 19360 3850 19372
rect 6641 19363 6699 19369
rect 3844 19332 4200 19360
rect 3844 19320 3850 19332
rect 2400 19295 2458 19301
rect 2400 19261 2412 19295
rect 2446 19292 2458 19295
rect 2682 19292 2688 19304
rect 2446 19264 2688 19292
rect 2446 19261 2458 19264
rect 2400 19255 2458 19261
rect 2682 19252 2688 19264
rect 2740 19252 2746 19304
rect 4172 19292 4200 19332
rect 6641 19329 6653 19363
rect 6687 19360 6699 19363
rect 7650 19360 7656 19372
rect 6687 19332 7656 19360
rect 6687 19329 6699 19332
rect 6641 19323 6699 19329
rect 7650 19320 7656 19332
rect 7708 19360 7714 19372
rect 8113 19363 8171 19369
rect 8113 19360 8125 19363
rect 7708 19332 8125 19360
rect 7708 19320 7714 19332
rect 8113 19329 8125 19332
rect 8159 19360 8171 19363
rect 8496 19360 8524 19456
rect 11057 19363 11115 19369
rect 11057 19360 11069 19363
rect 8159 19332 8524 19360
rect 9600 19332 11069 19360
rect 8159 19329 8171 19332
rect 8113 19323 8171 19329
rect 4172 19264 5212 19292
rect 1673 19227 1731 19233
rect 1673 19193 1685 19227
rect 1719 19224 1731 19227
rect 2590 19224 2596 19236
rect 1719 19196 2596 19224
rect 1719 19193 1731 19196
rect 1673 19187 1731 19193
rect 2590 19184 2596 19196
rect 2648 19184 2654 19236
rect 4338 19224 4344 19236
rect 3528 19196 4344 19224
rect 2958 19116 2964 19168
rect 3016 19156 3022 19168
rect 3528 19165 3556 19196
rect 4338 19184 4344 19196
rect 4396 19184 4402 19236
rect 4982 19224 4988 19236
rect 4448 19196 4988 19224
rect 3513 19159 3571 19165
rect 3513 19156 3525 19159
rect 3016 19128 3525 19156
rect 3016 19116 3022 19128
rect 3513 19125 3525 19128
rect 3559 19125 3571 19159
rect 3513 19119 3571 19125
rect 4154 19116 4160 19168
rect 4212 19156 4218 19168
rect 4448 19165 4476 19196
rect 4982 19184 4988 19196
rect 5040 19184 5046 19236
rect 5184 19233 5212 19264
rect 6914 19252 6920 19304
rect 6972 19292 6978 19304
rect 7543 19295 7601 19301
rect 7543 19292 7555 19295
rect 6972 19264 7555 19292
rect 6972 19252 6978 19264
rect 7543 19261 7555 19264
rect 7589 19261 7601 19295
rect 7543 19255 7601 19261
rect 7668 19264 8064 19292
rect 5169 19227 5227 19233
rect 5169 19193 5181 19227
rect 5215 19193 5227 19227
rect 5169 19187 5227 19193
rect 5261 19227 5319 19233
rect 5261 19193 5273 19227
rect 5307 19224 5319 19227
rect 5350 19224 5356 19236
rect 5307 19196 5356 19224
rect 5307 19193 5319 19196
rect 5261 19187 5319 19193
rect 5350 19184 5356 19196
rect 5408 19224 5414 19236
rect 5629 19227 5687 19233
rect 5629 19224 5641 19227
rect 5408 19196 5641 19224
rect 5408 19184 5414 19196
rect 5629 19193 5641 19196
rect 5675 19193 5687 19227
rect 7374 19224 7380 19236
rect 7287 19196 7380 19224
rect 5629 19187 5687 19193
rect 7374 19184 7380 19196
rect 7432 19224 7438 19236
rect 7668 19224 7696 19264
rect 8036 19233 8064 19264
rect 8294 19252 8300 19304
rect 8352 19292 8358 19304
rect 9122 19292 9128 19304
rect 8352 19264 9128 19292
rect 8352 19252 8358 19264
rect 9122 19252 9128 19264
rect 9180 19252 9186 19304
rect 9398 19292 9404 19304
rect 9359 19264 9404 19292
rect 9398 19252 9404 19264
rect 9456 19252 9462 19304
rect 9490 19252 9496 19304
rect 9548 19292 9554 19304
rect 9600 19292 9628 19332
rect 11057 19329 11069 19332
rect 11103 19360 11115 19363
rect 11330 19360 11336 19372
rect 11103 19332 11336 19360
rect 11103 19329 11115 19332
rect 11057 19323 11115 19329
rect 11330 19320 11336 19332
rect 11388 19320 11394 19372
rect 12526 19369 12532 19372
rect 12511 19363 12532 19369
rect 12511 19329 12523 19363
rect 12511 19323 12532 19329
rect 12526 19320 12532 19323
rect 12584 19320 12590 19372
rect 14108 19360 14136 19456
rect 19153 19363 19211 19369
rect 19153 19360 19165 19363
rect 14108 19332 14504 19360
rect 9548 19264 9628 19292
rect 9548 19252 9554 19264
rect 9674 19252 9680 19304
rect 9732 19292 9738 19304
rect 9953 19295 10011 19301
rect 9953 19292 9965 19295
rect 9732 19264 9965 19292
rect 9732 19252 9738 19264
rect 9953 19261 9965 19264
rect 9999 19292 10011 19295
rect 10781 19295 10839 19301
rect 10781 19292 10793 19295
rect 9999 19264 10793 19292
rect 9999 19261 10011 19264
rect 9953 19255 10011 19261
rect 10781 19261 10793 19264
rect 10827 19292 10839 19295
rect 10962 19292 10968 19304
rect 10827 19264 10968 19292
rect 10827 19261 10839 19264
rect 10781 19255 10839 19261
rect 10962 19252 10968 19264
rect 11020 19252 11026 19304
rect 11606 19252 11612 19304
rect 11664 19292 11670 19304
rect 11793 19295 11851 19301
rect 11793 19292 11805 19295
rect 11664 19264 11805 19292
rect 11664 19252 11670 19264
rect 7432 19196 7696 19224
rect 7837 19227 7895 19233
rect 7432 19184 7438 19196
rect 7837 19193 7849 19227
rect 7883 19193 7895 19227
rect 7837 19187 7895 19193
rect 8021 19227 8079 19233
rect 8021 19193 8033 19227
rect 8067 19224 8079 19227
rect 8110 19224 8116 19236
rect 8067 19196 8116 19224
rect 8067 19193 8079 19196
rect 8021 19187 8079 19193
rect 4433 19159 4491 19165
rect 4433 19156 4445 19159
rect 4212 19128 4445 19156
rect 4212 19116 4218 19128
rect 4433 19125 4445 19128
rect 4479 19125 4491 19159
rect 4433 19119 4491 19125
rect 4522 19116 4528 19168
rect 4580 19156 4586 19168
rect 4691 19159 4749 19165
rect 4691 19156 4703 19159
rect 4580 19128 4703 19156
rect 4580 19116 4586 19128
rect 4691 19125 4703 19128
rect 4737 19125 4749 19159
rect 4691 19119 4749 19125
rect 7558 19116 7564 19168
rect 7616 19156 7622 19168
rect 7852 19156 7880 19187
rect 8110 19184 8116 19196
rect 8168 19184 8174 19236
rect 10226 19184 10232 19236
rect 10284 19224 10290 19236
rect 11146 19224 11152 19236
rect 10284 19196 11152 19224
rect 10284 19184 10290 19196
rect 11146 19184 11152 19196
rect 11204 19184 11210 19236
rect 8478 19156 8484 19168
rect 7616 19128 7880 19156
rect 8439 19128 8484 19156
rect 7616 19116 7622 19128
rect 8478 19116 8484 19128
rect 8536 19116 8542 19168
rect 9858 19116 9864 19168
rect 9916 19156 9922 19168
rect 10965 19159 11023 19165
rect 10965 19156 10977 19159
rect 9916 19128 10977 19156
rect 9916 19116 9922 19128
rect 10965 19125 10977 19128
rect 11011 19156 11023 19159
rect 11425 19159 11483 19165
rect 11425 19156 11437 19159
rect 11011 19128 11437 19156
rect 11011 19125 11023 19128
rect 10965 19119 11023 19125
rect 11425 19125 11437 19128
rect 11471 19125 11483 19159
rect 11716 19156 11744 19264
rect 11793 19261 11805 19264
rect 11839 19261 11851 19295
rect 13081 19295 13139 19301
rect 13081 19292 13093 19295
rect 11793 19255 11851 19261
rect 12452 19264 13093 19292
rect 12066 19184 12072 19236
rect 12124 19224 12130 19236
rect 12452 19224 12480 19264
rect 13081 19261 13093 19264
rect 13127 19261 13139 19295
rect 13081 19255 13139 19261
rect 14369 19295 14427 19301
rect 14369 19261 14381 19295
rect 14415 19261 14427 19295
rect 14476 19292 14504 19332
rect 18984 19332 19165 19360
rect 18984 19304 19012 19332
rect 19153 19329 19165 19332
rect 19199 19329 19211 19363
rect 19153 19323 19211 19329
rect 19426 19320 19432 19372
rect 19484 19360 19490 19372
rect 20088 19369 20116 19468
rect 20254 19456 20260 19468
rect 20312 19456 20318 19508
rect 22370 19496 22376 19508
rect 22331 19468 22376 19496
rect 22370 19456 22376 19468
rect 22428 19456 22434 19508
rect 23014 19496 23020 19508
rect 22975 19468 23020 19496
rect 23014 19456 23020 19468
rect 23072 19456 23078 19508
rect 24210 19456 24216 19508
rect 24268 19496 24274 19508
rect 24305 19499 24363 19505
rect 24305 19496 24317 19499
rect 24268 19468 24317 19496
rect 24268 19456 24274 19468
rect 24305 19465 24317 19468
rect 24351 19465 24363 19499
rect 24305 19459 24363 19465
rect 24854 19456 24860 19508
rect 24912 19496 24918 19508
rect 25961 19499 26019 19505
rect 25961 19496 25973 19499
rect 24912 19468 25973 19496
rect 24912 19456 24918 19468
rect 25961 19465 25973 19468
rect 26007 19465 26019 19499
rect 25961 19459 26019 19465
rect 23032 19428 23060 19456
rect 25225 19431 25283 19437
rect 25225 19428 25237 19431
rect 23032 19400 25237 19428
rect 25225 19397 25237 19400
rect 25271 19428 25283 19431
rect 25498 19428 25504 19440
rect 25271 19400 25504 19428
rect 25271 19397 25283 19400
rect 25225 19391 25283 19397
rect 25498 19388 25504 19400
rect 25556 19388 25562 19440
rect 20073 19363 20131 19369
rect 20073 19360 20085 19363
rect 19484 19332 20085 19360
rect 19484 19320 19490 19332
rect 20073 19329 20085 19332
rect 20119 19329 20131 19363
rect 20073 19323 20131 19329
rect 25406 19320 25412 19372
rect 25464 19360 25470 19372
rect 25593 19363 25651 19369
rect 25593 19360 25605 19363
rect 25464 19332 25605 19360
rect 25464 19320 25470 19332
rect 25593 19329 25605 19332
rect 25639 19329 25651 19363
rect 25593 19323 25651 19329
rect 14625 19295 14683 19301
rect 14625 19292 14637 19295
rect 14476 19264 14637 19292
rect 14369 19255 14427 19261
rect 14625 19261 14637 19264
rect 14671 19261 14683 19295
rect 14625 19255 14683 19261
rect 12124 19196 12480 19224
rect 12124 19184 12130 19196
rect 12802 19184 12808 19236
rect 12860 19224 12866 19236
rect 12860 19196 12905 19224
rect 12860 19184 12866 19196
rect 13630 19184 13636 19236
rect 13688 19224 13694 19236
rect 14277 19227 14335 19233
rect 14277 19224 14289 19227
rect 13688 19196 14289 19224
rect 13688 19184 13694 19196
rect 14277 19193 14289 19196
rect 14323 19224 14335 19227
rect 14384 19224 14412 19255
rect 16482 19252 16488 19304
rect 16540 19292 16546 19304
rect 16853 19295 16911 19301
rect 16853 19292 16865 19295
rect 16540 19264 16865 19292
rect 16540 19252 16546 19264
rect 16853 19261 16865 19264
rect 16899 19261 16911 19295
rect 16853 19255 16911 19261
rect 17865 19295 17923 19301
rect 17865 19261 17877 19295
rect 17911 19292 17923 19295
rect 18966 19292 18972 19304
rect 17911 19264 18972 19292
rect 17911 19261 17923 19264
rect 17865 19255 17923 19261
rect 18966 19252 18972 19264
rect 19024 19252 19030 19304
rect 19613 19295 19671 19301
rect 19613 19292 19625 19295
rect 19076 19264 19625 19292
rect 17034 19224 17040 19236
rect 14323 19196 17040 19224
rect 14323 19193 14335 19196
rect 14277 19187 14335 19193
rect 17034 19184 17040 19196
rect 17092 19224 17098 19236
rect 17313 19227 17371 19233
rect 17313 19224 17325 19227
rect 17092 19196 17325 19224
rect 17092 19184 17098 19196
rect 17313 19193 17325 19196
rect 17359 19193 17371 19227
rect 18322 19224 18328 19236
rect 18283 19196 18328 19224
rect 17313 19187 17371 19193
rect 18322 19184 18328 19196
rect 18380 19224 18386 19236
rect 19076 19233 19104 19264
rect 19613 19261 19625 19264
rect 19659 19292 19671 19295
rect 19978 19292 19984 19304
rect 19659 19264 19984 19292
rect 19659 19261 19671 19264
rect 19613 19255 19671 19261
rect 19978 19252 19984 19264
rect 20036 19252 20042 19304
rect 20162 19252 20168 19304
rect 20220 19292 20226 19304
rect 20329 19295 20387 19301
rect 20329 19292 20341 19295
rect 20220 19264 20341 19292
rect 20220 19252 20226 19264
rect 20329 19261 20341 19264
rect 20375 19261 20387 19295
rect 20329 19255 20387 19261
rect 24026 19252 24032 19304
rect 24084 19292 24090 19304
rect 24857 19295 24915 19301
rect 24857 19292 24869 19295
rect 24084 19264 24869 19292
rect 24084 19252 24090 19264
rect 24857 19261 24869 19264
rect 24903 19261 24915 19295
rect 24857 19255 24915 19261
rect 18877 19227 18935 19233
rect 18877 19224 18889 19227
rect 18380 19196 18889 19224
rect 18380 19184 18386 19196
rect 18877 19193 18889 19196
rect 18923 19193 18935 19227
rect 18877 19187 18935 19193
rect 19061 19227 19119 19233
rect 19061 19193 19073 19227
rect 19107 19193 19119 19227
rect 19061 19187 19119 19193
rect 19518 19184 19524 19236
rect 19576 19224 19582 19236
rect 20070 19224 20076 19236
rect 19576 19196 20076 19224
rect 19576 19184 19582 19196
rect 20070 19184 20076 19196
rect 20128 19184 20134 19236
rect 23477 19227 23535 19233
rect 23477 19193 23489 19227
rect 23523 19224 23535 19227
rect 24581 19227 24639 19233
rect 24581 19224 24593 19227
rect 23523 19196 24593 19224
rect 23523 19193 23535 19196
rect 23477 19187 23535 19193
rect 24581 19193 24593 19196
rect 24627 19224 24639 19227
rect 24670 19224 24676 19236
rect 24627 19196 24676 19224
rect 24627 19193 24639 19196
rect 24581 19187 24639 19193
rect 24670 19184 24676 19196
rect 24728 19184 24734 19236
rect 12989 19159 13047 19165
rect 12989 19156 13001 19159
rect 11716 19128 13001 19156
rect 11425 19119 11483 19125
rect 12989 19125 13001 19128
rect 13035 19156 13047 19159
rect 13262 19156 13268 19168
rect 13035 19128 13268 19156
rect 13035 19125 13047 19128
rect 12989 19119 13047 19125
rect 13262 19116 13268 19128
rect 13320 19116 13326 19168
rect 13538 19156 13544 19168
rect 13499 19128 13544 19156
rect 13538 19116 13544 19128
rect 13596 19116 13602 19168
rect 15378 19116 15384 19168
rect 15436 19156 15442 19168
rect 15749 19159 15807 19165
rect 15749 19156 15761 19159
rect 15436 19128 15761 19156
rect 15436 19116 15442 19128
rect 15749 19125 15761 19128
rect 15795 19125 15807 19159
rect 16298 19156 16304 19168
rect 16259 19128 16304 19156
rect 15749 19119 15807 19125
rect 16298 19116 16304 19128
rect 16356 19116 16362 19168
rect 16758 19156 16764 19168
rect 16719 19128 16764 19156
rect 16758 19116 16764 19128
rect 16816 19116 16822 19168
rect 18591 19159 18649 19165
rect 18591 19125 18603 19159
rect 18637 19156 18649 19159
rect 19242 19156 19248 19168
rect 18637 19128 19248 19156
rect 18637 19125 18649 19128
rect 18591 19119 18649 19125
rect 19242 19116 19248 19128
rect 19300 19116 19306 19168
rect 20714 19116 20720 19168
rect 20772 19156 20778 19168
rect 21453 19159 21511 19165
rect 21453 19156 21465 19159
rect 20772 19128 21465 19156
rect 20772 19116 20778 19128
rect 21453 19125 21465 19128
rect 21499 19125 21511 19159
rect 22554 19156 22560 19168
rect 22515 19128 22560 19156
rect 21453 19119 21511 19125
rect 22554 19116 22560 19128
rect 22612 19116 22618 19168
rect 24026 19156 24032 19168
rect 23987 19128 24032 19156
rect 24026 19116 24032 19128
rect 24084 19116 24090 19168
rect 24762 19156 24768 19168
rect 24723 19128 24768 19156
rect 24762 19116 24768 19128
rect 24820 19116 24826 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 2682 18912 2688 18964
rect 2740 18952 2746 18964
rect 3329 18955 3387 18961
rect 3329 18952 3341 18955
rect 2740 18924 3341 18952
rect 2740 18912 2746 18924
rect 3329 18921 3341 18924
rect 3375 18921 3387 18955
rect 3694 18952 3700 18964
rect 3655 18924 3700 18952
rect 3329 18915 3387 18921
rect 3694 18912 3700 18924
rect 3752 18912 3758 18964
rect 4338 18952 4344 18964
rect 4299 18924 4344 18952
rect 4338 18912 4344 18924
rect 4396 18912 4402 18964
rect 7650 18952 7656 18964
rect 7611 18924 7656 18952
rect 7650 18912 7656 18924
rect 7708 18912 7714 18964
rect 8297 18955 8355 18961
rect 8297 18921 8309 18955
rect 8343 18952 8355 18955
rect 8386 18952 8392 18964
rect 8343 18924 8392 18952
rect 8343 18921 8355 18924
rect 8297 18915 8355 18921
rect 8386 18912 8392 18924
rect 8444 18912 8450 18964
rect 9490 18952 9496 18964
rect 9451 18924 9496 18952
rect 9490 18912 9496 18924
rect 9548 18912 9554 18964
rect 10134 18952 10140 18964
rect 10095 18924 10140 18952
rect 10134 18912 10140 18924
rect 10192 18912 10198 18964
rect 10778 18912 10784 18964
rect 10836 18952 10842 18964
rect 10873 18955 10931 18961
rect 10873 18952 10885 18955
rect 10836 18924 10885 18952
rect 10836 18912 10842 18924
rect 10873 18921 10885 18924
rect 10919 18921 10931 18955
rect 11330 18952 11336 18964
rect 11291 18924 11336 18952
rect 10873 18915 10931 18921
rect 2869 18887 2927 18893
rect 2869 18853 2881 18887
rect 2915 18853 2927 18887
rect 2869 18847 2927 18853
rect 2884 18816 2912 18847
rect 2958 18844 2964 18896
rect 3016 18884 3022 18896
rect 5258 18884 5264 18896
rect 3016 18856 3061 18884
rect 5219 18856 5264 18884
rect 3016 18844 3022 18856
rect 5258 18844 5264 18856
rect 5316 18844 5322 18896
rect 10888 18884 10916 18915
rect 11330 18912 11336 18924
rect 11388 18912 11394 18964
rect 12618 18952 12624 18964
rect 11440 18924 12624 18952
rect 11440 18884 11468 18924
rect 12618 18912 12624 18924
rect 12676 18912 12682 18964
rect 12802 18912 12808 18964
rect 12860 18952 12866 18964
rect 12897 18955 12955 18961
rect 12897 18952 12909 18955
rect 12860 18924 12909 18952
rect 12860 18912 12866 18924
rect 12897 18921 12909 18924
rect 12943 18921 12955 18955
rect 12897 18915 12955 18921
rect 12986 18912 12992 18964
rect 13044 18952 13050 18964
rect 13265 18955 13323 18961
rect 13265 18952 13277 18955
rect 13044 18924 13277 18952
rect 13044 18912 13050 18924
rect 13265 18921 13277 18924
rect 13311 18921 13323 18955
rect 13265 18915 13323 18921
rect 13906 18912 13912 18964
rect 13964 18952 13970 18964
rect 14553 18955 14611 18961
rect 14553 18952 14565 18955
rect 13964 18924 14565 18952
rect 13964 18912 13970 18924
rect 14553 18921 14565 18924
rect 14599 18952 14611 18955
rect 15565 18955 15623 18961
rect 15565 18952 15577 18955
rect 14599 18924 15577 18952
rect 14599 18921 14611 18924
rect 14553 18915 14611 18921
rect 15565 18921 15577 18924
rect 15611 18952 15623 18955
rect 15838 18952 15844 18964
rect 15611 18924 15844 18952
rect 15611 18921 15623 18924
rect 15565 18915 15623 18921
rect 15838 18912 15844 18924
rect 15896 18912 15902 18964
rect 17126 18952 17132 18964
rect 17087 18924 17132 18952
rect 17126 18912 17132 18924
rect 17184 18912 17190 18964
rect 18598 18952 18604 18964
rect 18559 18924 18604 18952
rect 18598 18912 18604 18924
rect 18656 18912 18662 18964
rect 20806 18912 20812 18964
rect 20864 18952 20870 18964
rect 21085 18955 21143 18961
rect 21085 18952 21097 18955
rect 20864 18924 21097 18952
rect 20864 18912 20870 18924
rect 21085 18921 21097 18924
rect 21131 18921 21143 18955
rect 21450 18952 21456 18964
rect 21411 18924 21456 18952
rect 21085 18915 21143 18921
rect 21450 18912 21456 18924
rect 21508 18912 21514 18964
rect 11698 18884 11704 18896
rect 10888 18856 11468 18884
rect 11659 18856 11704 18884
rect 11698 18844 11704 18856
rect 11756 18844 11762 18896
rect 12342 18844 12348 18896
rect 12400 18884 12406 18896
rect 12437 18887 12495 18893
rect 12437 18884 12449 18887
rect 12400 18856 12449 18884
rect 12400 18844 12406 18856
rect 12437 18853 12449 18856
rect 12483 18884 12495 18887
rect 12526 18884 12532 18896
rect 12483 18856 12532 18884
rect 12483 18853 12495 18856
rect 12437 18847 12495 18853
rect 12526 18844 12532 18856
rect 12584 18844 12590 18896
rect 14001 18887 14059 18893
rect 14001 18853 14013 18887
rect 14047 18884 14059 18887
rect 14642 18884 14648 18896
rect 14047 18856 14648 18884
rect 14047 18853 14059 18856
rect 14001 18847 14059 18853
rect 14642 18844 14648 18856
rect 14700 18844 14706 18896
rect 16206 18884 16212 18896
rect 16167 18856 16212 18884
rect 16206 18844 16212 18856
rect 16264 18844 16270 18896
rect 17488 18887 17546 18893
rect 17488 18853 17500 18887
rect 17534 18884 17546 18887
rect 17862 18884 17868 18896
rect 17534 18856 17868 18884
rect 17534 18853 17546 18856
rect 17488 18847 17546 18853
rect 17862 18844 17868 18856
rect 17920 18844 17926 18896
rect 21358 18844 21364 18896
rect 21416 18884 21422 18896
rect 22640 18887 22698 18893
rect 22640 18884 22652 18887
rect 21416 18856 22652 18884
rect 21416 18844 21422 18856
rect 22640 18853 22652 18856
rect 22686 18884 22698 18887
rect 23382 18884 23388 18896
rect 22686 18856 23388 18884
rect 22686 18853 22698 18856
rect 22640 18847 22698 18853
rect 23382 18844 23388 18856
rect 23440 18844 23446 18896
rect 25038 18844 25044 18896
rect 25096 18884 25102 18896
rect 25409 18887 25467 18893
rect 25409 18884 25421 18887
rect 25096 18856 25421 18884
rect 25096 18844 25102 18856
rect 25409 18853 25421 18856
rect 25455 18853 25467 18887
rect 25409 18847 25467 18853
rect 3142 18816 3148 18828
rect 2884 18788 3148 18816
rect 3142 18776 3148 18788
rect 3200 18816 3206 18828
rect 3602 18816 3608 18828
rect 3200 18788 3608 18816
rect 3200 18776 3206 18788
rect 3602 18776 3608 18788
rect 3660 18776 3666 18828
rect 4154 18776 4160 18828
rect 4212 18816 4218 18828
rect 5353 18819 5411 18825
rect 5353 18816 5365 18819
rect 4212 18788 5365 18816
rect 4212 18776 4218 18788
rect 5353 18785 5365 18788
rect 5399 18816 5411 18819
rect 5442 18816 5448 18828
rect 5399 18788 5448 18816
rect 5399 18785 5411 18788
rect 5353 18779 5411 18785
rect 5442 18776 5448 18788
rect 5500 18776 5506 18828
rect 6540 18819 6598 18825
rect 6540 18785 6552 18819
rect 6586 18816 6598 18819
rect 7006 18816 7012 18828
rect 6586 18788 7012 18816
rect 6586 18785 6598 18788
rect 6540 18779 6598 18785
rect 7006 18776 7012 18788
rect 7064 18776 7070 18828
rect 9858 18776 9864 18828
rect 9916 18816 9922 18828
rect 10689 18819 10747 18825
rect 10689 18816 10701 18819
rect 9916 18788 10701 18816
rect 9916 18776 9922 18788
rect 10689 18785 10701 18788
rect 10735 18785 10747 18819
rect 10689 18779 10747 18785
rect 12802 18776 12808 18828
rect 12860 18816 12866 18828
rect 13722 18816 13728 18828
rect 12860 18788 13728 18816
rect 12860 18776 12866 18788
rect 13722 18776 13728 18788
rect 13780 18816 13786 18828
rect 14093 18819 14151 18825
rect 14093 18816 14105 18819
rect 13780 18788 14105 18816
rect 13780 18776 13786 18788
rect 14093 18785 14105 18788
rect 14139 18785 14151 18819
rect 16022 18816 16028 18828
rect 15983 18788 16028 18816
rect 14093 18779 14151 18785
rect 16022 18776 16028 18788
rect 16080 18776 16086 18828
rect 21174 18776 21180 18828
rect 21232 18816 21238 18828
rect 21269 18819 21327 18825
rect 21269 18816 21281 18819
rect 21232 18788 21281 18816
rect 21232 18776 21238 18788
rect 21269 18785 21281 18788
rect 21315 18785 21327 18819
rect 22370 18816 22376 18828
rect 22331 18788 22376 18816
rect 21269 18779 21327 18785
rect 22370 18776 22376 18788
rect 22428 18776 22434 18828
rect 25222 18816 25228 18828
rect 25135 18788 25228 18816
rect 25222 18776 25228 18788
rect 25280 18816 25286 18828
rect 25774 18816 25780 18828
rect 25280 18788 25780 18816
rect 25280 18776 25286 18788
rect 25774 18776 25780 18788
rect 25832 18776 25838 18828
rect 2774 18708 2780 18760
rect 2832 18748 2838 18760
rect 5258 18748 5264 18760
rect 2832 18720 2877 18748
rect 5219 18720 5264 18748
rect 2832 18708 2838 18720
rect 5258 18708 5264 18720
rect 5316 18708 5322 18760
rect 6178 18708 6184 18760
rect 6236 18748 6242 18760
rect 6273 18751 6331 18757
rect 6273 18748 6285 18751
rect 6236 18720 6285 18748
rect 6236 18708 6242 18720
rect 6273 18717 6285 18720
rect 6319 18717 6331 18751
rect 10962 18748 10968 18760
rect 10923 18720 10968 18748
rect 6273 18711 6331 18717
rect 10962 18708 10968 18720
rect 11020 18748 11026 18760
rect 12066 18748 12072 18760
rect 11020 18720 12072 18748
rect 11020 18708 11026 18720
rect 12066 18708 12072 18720
rect 12124 18708 12130 18760
rect 12345 18751 12403 18757
rect 12345 18717 12357 18751
rect 12391 18717 12403 18751
rect 12526 18748 12532 18760
rect 12487 18720 12532 18748
rect 12345 18711 12403 18717
rect 2409 18683 2467 18689
rect 2409 18649 2421 18683
rect 2455 18680 2467 18683
rect 2682 18680 2688 18692
rect 2455 18652 2688 18680
rect 2455 18649 2467 18652
rect 2409 18643 2467 18649
rect 2682 18640 2688 18652
rect 2740 18640 2746 18692
rect 4798 18680 4804 18692
rect 4759 18652 4804 18680
rect 4798 18640 4804 18652
rect 4856 18640 4862 18692
rect 10413 18683 10471 18689
rect 10413 18649 10425 18683
rect 10459 18680 10471 18683
rect 12250 18680 12256 18692
rect 10459 18652 12256 18680
rect 10459 18649 10471 18652
rect 10413 18643 10471 18649
rect 12250 18640 12256 18652
rect 12308 18680 12314 18692
rect 12360 18680 12388 18711
rect 12526 18708 12532 18720
rect 12584 18708 12590 18760
rect 13998 18748 14004 18760
rect 13911 18720 14004 18748
rect 13998 18708 14004 18720
rect 14056 18748 14062 18760
rect 14458 18748 14464 18760
rect 14056 18720 14464 18748
rect 14056 18708 14062 18720
rect 14458 18708 14464 18720
rect 14516 18708 14522 18760
rect 16114 18708 16120 18760
rect 16172 18748 16178 18760
rect 16301 18751 16359 18757
rect 16301 18748 16313 18751
rect 16172 18720 16313 18748
rect 16172 18708 16178 18720
rect 16301 18717 16313 18720
rect 16347 18748 16359 18751
rect 16347 18720 16804 18748
rect 16347 18717 16359 18720
rect 16301 18711 16359 18717
rect 12308 18652 12388 18680
rect 12308 18640 12314 18652
rect 13078 18640 13084 18692
rect 13136 18680 13142 18692
rect 14918 18680 14924 18692
rect 13136 18652 14924 18680
rect 13136 18640 13142 18652
rect 14918 18640 14924 18652
rect 14976 18640 14982 18692
rect 15746 18680 15752 18692
rect 15707 18652 15752 18680
rect 15746 18640 15752 18652
rect 15804 18640 15810 18692
rect 1578 18612 1584 18624
rect 1539 18584 1584 18612
rect 1578 18572 1584 18584
rect 1636 18572 1642 18624
rect 1854 18572 1860 18624
rect 1912 18612 1918 18624
rect 1949 18615 2007 18621
rect 1949 18612 1961 18615
rect 1912 18584 1961 18612
rect 1912 18572 1918 18584
rect 1949 18581 1961 18584
rect 1995 18612 2007 18615
rect 2498 18612 2504 18624
rect 1995 18584 2504 18612
rect 1995 18581 2007 18584
rect 1949 18575 2007 18581
rect 2498 18572 2504 18584
rect 2556 18572 2562 18624
rect 5534 18572 5540 18624
rect 5592 18612 5598 18624
rect 5721 18615 5779 18621
rect 5721 18612 5733 18615
rect 5592 18584 5733 18612
rect 5592 18572 5598 18584
rect 5721 18581 5733 18584
rect 5767 18581 5779 18615
rect 6086 18612 6092 18624
rect 6047 18584 6092 18612
rect 5721 18575 5779 18581
rect 6086 18572 6092 18584
rect 6144 18572 6150 18624
rect 8662 18612 8668 18624
rect 8623 18584 8668 18612
rect 8662 18572 8668 18584
rect 8720 18572 8726 18624
rect 9030 18612 9036 18624
rect 8991 18584 9036 18612
rect 9030 18572 9036 18584
rect 9088 18572 9094 18624
rect 11974 18612 11980 18624
rect 11935 18584 11980 18612
rect 11974 18572 11980 18584
rect 12032 18572 12038 18624
rect 13538 18612 13544 18624
rect 13499 18584 13544 18612
rect 13538 18572 13544 18584
rect 13596 18572 13602 18624
rect 13722 18572 13728 18624
rect 13780 18612 13786 18624
rect 14829 18615 14887 18621
rect 14829 18612 14841 18615
rect 13780 18584 14841 18612
rect 13780 18572 13786 18584
rect 14829 18581 14841 18584
rect 14875 18612 14887 18615
rect 15378 18612 15384 18624
rect 14875 18584 15384 18612
rect 14875 18581 14887 18584
rect 14829 18575 14887 18581
rect 15378 18572 15384 18584
rect 15436 18572 15442 18624
rect 16776 18621 16804 18720
rect 17126 18708 17132 18760
rect 17184 18748 17190 18760
rect 17221 18751 17279 18757
rect 17221 18748 17233 18751
rect 17184 18720 17233 18748
rect 17184 18708 17190 18720
rect 17221 18717 17233 18720
rect 17267 18717 17279 18751
rect 17221 18711 17279 18717
rect 19334 18708 19340 18760
rect 19392 18748 19398 18760
rect 19797 18751 19855 18757
rect 19797 18748 19809 18751
rect 19392 18720 19809 18748
rect 19392 18708 19398 18720
rect 19797 18717 19809 18720
rect 19843 18717 19855 18751
rect 19797 18711 19855 18717
rect 25130 18708 25136 18760
rect 25188 18748 25194 18760
rect 25498 18748 25504 18760
rect 25188 18720 25504 18748
rect 25188 18708 25194 18720
rect 25498 18708 25504 18720
rect 25556 18708 25562 18760
rect 23382 18640 23388 18692
rect 23440 18680 23446 18692
rect 23842 18680 23848 18692
rect 23440 18652 23848 18680
rect 23440 18640 23446 18652
rect 23842 18640 23848 18652
rect 23900 18640 23906 18692
rect 24397 18683 24455 18689
rect 24397 18649 24409 18683
rect 24443 18680 24455 18683
rect 24762 18680 24768 18692
rect 24443 18652 24768 18680
rect 24443 18649 24455 18652
rect 24397 18643 24455 18649
rect 24762 18640 24768 18652
rect 24820 18680 24826 18692
rect 24949 18683 25007 18689
rect 24949 18680 24961 18683
rect 24820 18652 24961 18680
rect 24820 18640 24826 18652
rect 24949 18649 24961 18652
rect 24995 18649 25007 18683
rect 24949 18643 25007 18649
rect 16761 18615 16819 18621
rect 16761 18581 16773 18615
rect 16807 18612 16819 18615
rect 17034 18612 17040 18624
rect 16807 18584 17040 18612
rect 16807 18581 16819 18584
rect 16761 18575 16819 18581
rect 17034 18572 17040 18584
rect 17092 18572 17098 18624
rect 19518 18612 19524 18624
rect 19479 18584 19524 18612
rect 19518 18572 19524 18584
rect 19576 18572 19582 18624
rect 22094 18572 22100 18624
rect 22152 18612 22158 18624
rect 22152 18584 22197 18612
rect 22152 18572 22158 18584
rect 23566 18572 23572 18624
rect 23624 18612 23630 18624
rect 23753 18615 23811 18621
rect 23753 18612 23765 18615
rect 23624 18584 23765 18612
rect 23624 18572 23630 18584
rect 23753 18581 23765 18584
rect 23799 18581 23811 18615
rect 23753 18575 23811 18581
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 2866 18368 2872 18420
rect 2924 18408 2930 18420
rect 2961 18411 3019 18417
rect 2961 18408 2973 18411
rect 2924 18380 2973 18408
rect 2924 18368 2930 18380
rect 2961 18377 2973 18380
rect 3007 18408 3019 18411
rect 5350 18408 5356 18420
rect 3007 18380 5356 18408
rect 3007 18377 3019 18380
rect 2961 18371 3019 18377
rect 5350 18368 5356 18380
rect 5408 18368 5414 18420
rect 6638 18368 6644 18420
rect 6696 18408 6702 18420
rect 7006 18408 7012 18420
rect 6696 18380 7012 18408
rect 6696 18368 6702 18380
rect 7006 18368 7012 18380
rect 7064 18368 7070 18420
rect 8662 18368 8668 18420
rect 8720 18408 8726 18420
rect 10229 18411 10287 18417
rect 10229 18408 10241 18411
rect 8720 18380 10241 18408
rect 8720 18368 8726 18380
rect 10229 18377 10241 18380
rect 10275 18377 10287 18411
rect 10229 18371 10287 18377
rect 10778 18368 10784 18420
rect 10836 18408 10842 18420
rect 11149 18411 11207 18417
rect 11149 18408 11161 18411
rect 10836 18380 11161 18408
rect 10836 18368 10842 18380
rect 11149 18377 11161 18380
rect 11195 18377 11207 18411
rect 11149 18371 11207 18377
rect 11609 18411 11667 18417
rect 11609 18377 11621 18411
rect 11655 18408 11667 18411
rect 12158 18408 12164 18420
rect 11655 18380 12164 18408
rect 11655 18377 11667 18380
rect 11609 18371 11667 18377
rect 9858 18300 9864 18352
rect 9916 18340 9922 18352
rect 9953 18343 10011 18349
rect 9953 18340 9965 18343
rect 9916 18312 9965 18340
rect 9916 18300 9922 18312
rect 9953 18309 9965 18312
rect 9999 18309 10011 18343
rect 9953 18303 10011 18309
rect 10689 18275 10747 18281
rect 10689 18241 10701 18275
rect 10735 18272 10747 18275
rect 11624 18272 11652 18371
rect 12158 18368 12164 18380
rect 12216 18368 12222 18420
rect 12802 18408 12808 18420
rect 12763 18380 12808 18408
rect 12802 18368 12808 18380
rect 12860 18368 12866 18420
rect 13173 18411 13231 18417
rect 13173 18377 13185 18411
rect 13219 18408 13231 18411
rect 13998 18408 14004 18420
rect 13219 18380 14004 18408
rect 13219 18377 13231 18380
rect 13173 18371 13231 18377
rect 13998 18368 14004 18380
rect 14056 18368 14062 18420
rect 14369 18411 14427 18417
rect 14369 18377 14381 18411
rect 14415 18408 14427 18411
rect 14642 18408 14648 18420
rect 14415 18380 14648 18408
rect 14415 18377 14427 18380
rect 14369 18371 14427 18377
rect 14642 18368 14648 18380
rect 14700 18368 14706 18420
rect 14826 18368 14832 18420
rect 14884 18408 14890 18420
rect 14921 18411 14979 18417
rect 14921 18408 14933 18411
rect 14884 18380 14933 18408
rect 14884 18368 14890 18380
rect 14921 18377 14933 18380
rect 14967 18377 14979 18411
rect 14921 18371 14979 18377
rect 15470 18368 15476 18420
rect 15528 18408 15534 18420
rect 16117 18411 16175 18417
rect 16117 18408 16129 18411
rect 15528 18380 16129 18408
rect 15528 18368 15534 18380
rect 16117 18377 16129 18380
rect 16163 18408 16175 18411
rect 16209 18411 16267 18417
rect 16209 18408 16221 18411
rect 16163 18380 16221 18408
rect 16163 18377 16175 18380
rect 16117 18371 16175 18377
rect 16209 18377 16221 18380
rect 16255 18377 16267 18411
rect 16209 18371 16267 18377
rect 16390 18368 16396 18420
rect 16448 18408 16454 18420
rect 16485 18411 16543 18417
rect 16485 18408 16497 18411
rect 16448 18380 16497 18408
rect 16448 18368 16454 18380
rect 16485 18377 16497 18380
rect 16531 18377 16543 18411
rect 17862 18408 17868 18420
rect 17823 18380 17868 18408
rect 16485 18371 16543 18377
rect 17862 18368 17868 18380
rect 17920 18368 17926 18420
rect 19426 18408 19432 18420
rect 19387 18380 19432 18408
rect 19426 18368 19432 18380
rect 19484 18368 19490 18420
rect 20162 18368 20168 18420
rect 20220 18408 20226 18420
rect 20901 18411 20959 18417
rect 20901 18408 20913 18411
rect 20220 18380 20913 18408
rect 20220 18368 20226 18380
rect 20901 18377 20913 18380
rect 20947 18377 20959 18411
rect 20901 18371 20959 18377
rect 21358 18368 21364 18420
rect 21416 18408 21422 18420
rect 21453 18411 21511 18417
rect 21453 18408 21465 18411
rect 21416 18380 21465 18408
rect 21416 18368 21422 18380
rect 21453 18377 21465 18380
rect 21499 18377 21511 18411
rect 21453 18371 21511 18377
rect 22097 18411 22155 18417
rect 22097 18377 22109 18411
rect 22143 18408 22155 18411
rect 23474 18408 23480 18420
rect 22143 18380 23480 18408
rect 22143 18377 22155 18380
rect 22097 18371 22155 18377
rect 23474 18368 23480 18380
rect 23532 18368 23538 18420
rect 25038 18408 25044 18420
rect 24044 18380 24716 18408
rect 24999 18380 25044 18408
rect 11698 18300 11704 18352
rect 11756 18340 11762 18352
rect 12820 18340 12848 18368
rect 11756 18312 12848 18340
rect 13357 18343 13415 18349
rect 11756 18300 11762 18312
rect 13357 18309 13369 18343
rect 13403 18340 13415 18343
rect 13630 18340 13636 18352
rect 13403 18312 13636 18340
rect 13403 18309 13415 18312
rect 13357 18303 13415 18309
rect 13630 18300 13636 18312
rect 13688 18300 13694 18352
rect 14734 18300 14740 18352
rect 14792 18340 14798 18352
rect 18233 18343 18291 18349
rect 18233 18340 18245 18343
rect 14792 18312 18245 18340
rect 14792 18300 14798 18312
rect 13906 18272 13912 18284
rect 10735 18244 11652 18272
rect 13867 18244 13912 18272
rect 10735 18241 10747 18244
rect 10689 18235 10747 18241
rect 13906 18232 13912 18244
rect 13964 18232 13970 18284
rect 15396 18281 15424 18312
rect 18233 18309 18245 18312
rect 18279 18309 18291 18343
rect 18233 18303 18291 18309
rect 15381 18275 15439 18281
rect 15381 18241 15393 18275
rect 15427 18241 15439 18275
rect 15381 18235 15439 18241
rect 16574 18232 16580 18284
rect 16632 18272 16638 18284
rect 16945 18275 17003 18281
rect 16945 18272 16957 18275
rect 16632 18244 16957 18272
rect 16632 18232 16638 18244
rect 16945 18241 16957 18244
rect 16991 18272 17003 18275
rect 19334 18272 19340 18284
rect 16991 18244 19340 18272
rect 16991 18241 17003 18244
rect 16945 18235 17003 18241
rect 19334 18232 19340 18244
rect 19392 18232 19398 18284
rect 19444 18272 19472 18368
rect 22186 18300 22192 18352
rect 22244 18340 22250 18352
rect 22370 18340 22376 18352
rect 22244 18312 22376 18340
rect 22244 18300 22250 18312
rect 22370 18300 22376 18312
rect 22428 18340 22434 18352
rect 23017 18343 23075 18349
rect 23017 18340 23029 18343
rect 22428 18312 23029 18340
rect 22428 18300 22434 18312
rect 23017 18309 23029 18312
rect 23063 18309 23075 18343
rect 24044 18340 24072 18380
rect 23017 18303 23075 18309
rect 23492 18312 24072 18340
rect 24121 18343 24179 18349
rect 19521 18275 19579 18281
rect 19521 18272 19533 18275
rect 19444 18244 19533 18272
rect 19521 18241 19533 18244
rect 19567 18241 19579 18275
rect 19521 18235 19579 18241
rect 21913 18275 21971 18281
rect 21913 18241 21925 18275
rect 21959 18272 21971 18275
rect 22554 18272 22560 18284
rect 21959 18244 22560 18272
rect 21959 18241 21971 18244
rect 21913 18235 21971 18241
rect 22554 18232 22560 18244
rect 22612 18232 22618 18284
rect 23492 18281 23520 18312
rect 24121 18309 24133 18343
rect 24167 18309 24179 18343
rect 24121 18303 24179 18309
rect 23477 18275 23535 18281
rect 23477 18241 23489 18275
rect 23523 18241 23535 18275
rect 23842 18272 23848 18284
rect 23803 18244 23848 18272
rect 23477 18235 23535 18241
rect 23842 18232 23848 18244
rect 23900 18232 23906 18284
rect 1578 18204 1584 18216
rect 1539 18176 1584 18204
rect 1578 18164 1584 18176
rect 1636 18164 1642 18216
rect 1854 18213 1860 18216
rect 1848 18167 1860 18213
rect 1912 18204 1918 18216
rect 4157 18207 4215 18213
rect 1912 18176 1948 18204
rect 1854 18164 1860 18167
rect 1912 18164 1918 18176
rect 4157 18173 4169 18207
rect 4203 18204 4215 18207
rect 4246 18204 4252 18216
rect 4203 18176 4252 18204
rect 4203 18173 4215 18176
rect 4157 18167 4215 18173
rect 4246 18164 4252 18176
rect 4304 18204 4310 18216
rect 6178 18204 6184 18216
rect 4304 18176 6184 18204
rect 4304 18164 4310 18176
rect 6178 18164 6184 18176
rect 6236 18164 6242 18216
rect 7653 18207 7711 18213
rect 7653 18204 7665 18207
rect 7484 18176 7665 18204
rect 3694 18096 3700 18148
rect 3752 18136 3758 18148
rect 4338 18136 4344 18148
rect 3752 18108 4344 18136
rect 3752 18096 3758 18108
rect 4338 18096 4344 18108
rect 4396 18136 4402 18148
rect 4494 18139 4552 18145
rect 4494 18136 4506 18139
rect 4396 18108 4506 18136
rect 4396 18096 4402 18108
rect 4494 18105 4506 18108
rect 4540 18105 4552 18139
rect 4494 18099 4552 18105
rect 3602 18068 3608 18080
rect 3563 18040 3608 18068
rect 3602 18028 3608 18040
rect 3660 18028 3666 18080
rect 5534 18028 5540 18080
rect 5592 18068 5598 18080
rect 5629 18071 5687 18077
rect 5629 18068 5641 18071
rect 5592 18040 5641 18068
rect 5592 18028 5598 18040
rect 5629 18037 5641 18040
rect 5675 18037 5687 18071
rect 5629 18031 5687 18037
rect 6178 18028 6184 18080
rect 6236 18068 6242 18080
rect 7484 18077 7512 18176
rect 7653 18173 7665 18176
rect 7699 18173 7711 18207
rect 7653 18167 7711 18173
rect 9677 18207 9735 18213
rect 9677 18173 9689 18207
rect 9723 18204 9735 18207
rect 9723 18176 10732 18204
rect 9723 18173 9735 18176
rect 9677 18167 9735 18173
rect 10704 18148 10732 18176
rect 12986 18164 12992 18216
rect 13044 18204 13050 18216
rect 13633 18207 13691 18213
rect 13633 18204 13645 18207
rect 13044 18176 13645 18204
rect 13044 18164 13050 18176
rect 13633 18173 13645 18176
rect 13679 18173 13691 18207
rect 13633 18167 13691 18173
rect 14737 18207 14795 18213
rect 14737 18173 14749 18207
rect 14783 18204 14795 18207
rect 15473 18207 15531 18213
rect 15473 18204 15485 18207
rect 14783 18176 15485 18204
rect 14783 18173 14795 18176
rect 14737 18167 14795 18173
rect 15473 18173 15485 18176
rect 15519 18204 15531 18207
rect 16390 18204 16396 18216
rect 15519 18176 16396 18204
rect 15519 18173 15531 18176
rect 15473 18167 15531 18173
rect 16390 18164 16396 18176
rect 16448 18164 16454 18216
rect 17034 18204 17040 18216
rect 16995 18176 17040 18204
rect 17034 18164 17040 18176
rect 17092 18164 17098 18216
rect 22094 18164 22100 18216
rect 22152 18204 22158 18216
rect 24136 18204 24164 18303
rect 22152 18176 24164 18204
rect 22152 18164 22158 18176
rect 7834 18096 7840 18148
rect 7892 18145 7898 18148
rect 7892 18139 7956 18145
rect 7892 18105 7910 18139
rect 7944 18105 7956 18139
rect 10686 18136 10692 18148
rect 10647 18108 10692 18136
rect 7892 18099 7956 18105
rect 7892 18096 7898 18099
rect 10686 18096 10692 18108
rect 10744 18096 10750 18148
rect 10778 18096 10784 18148
rect 10836 18136 10842 18148
rect 12158 18136 12164 18148
rect 10836 18108 10881 18136
rect 10980 18108 12164 18136
rect 10836 18096 10842 18108
rect 6273 18071 6331 18077
rect 6273 18068 6285 18071
rect 6236 18040 6285 18068
rect 6236 18028 6242 18040
rect 6273 18037 6285 18040
rect 6319 18068 6331 18071
rect 7469 18071 7527 18077
rect 7469 18068 7481 18071
rect 6319 18040 7481 18068
rect 6319 18037 6331 18040
rect 6273 18031 6331 18037
rect 7469 18037 7481 18040
rect 7515 18037 7527 18071
rect 7469 18031 7527 18037
rect 9033 18071 9091 18077
rect 9033 18037 9045 18071
rect 9079 18068 9091 18071
rect 9306 18068 9312 18080
rect 9079 18040 9312 18068
rect 9079 18037 9091 18040
rect 9033 18031 9091 18037
rect 9306 18028 9312 18040
rect 9364 18028 9370 18080
rect 9766 18028 9772 18080
rect 9824 18068 9830 18080
rect 10980 18068 11008 18108
rect 12158 18096 12164 18108
rect 12216 18096 12222 18148
rect 13354 18096 13360 18148
rect 13412 18136 13418 18148
rect 13817 18139 13875 18145
rect 13817 18136 13829 18139
rect 13412 18108 13829 18136
rect 13412 18096 13418 18108
rect 13817 18105 13829 18108
rect 13863 18105 13875 18139
rect 15378 18136 15384 18148
rect 15339 18108 15384 18136
rect 13817 18099 13875 18105
rect 15378 18096 15384 18108
rect 15436 18096 15442 18148
rect 16117 18139 16175 18145
rect 16117 18105 16129 18139
rect 16163 18136 16175 18139
rect 16942 18136 16948 18148
rect 16163 18108 16948 18136
rect 16163 18105 16175 18108
rect 16117 18099 16175 18105
rect 16942 18096 16948 18108
rect 17000 18096 17006 18148
rect 19426 18096 19432 18148
rect 19484 18136 19490 18148
rect 22572 18145 22600 18176
rect 19766 18139 19824 18145
rect 19766 18136 19778 18139
rect 19484 18108 19778 18136
rect 19484 18096 19490 18108
rect 19766 18105 19778 18108
rect 19812 18105 19824 18139
rect 19766 18099 19824 18105
rect 22557 18139 22615 18145
rect 22557 18105 22569 18139
rect 22603 18105 22615 18139
rect 22557 18099 22615 18105
rect 22649 18139 22707 18145
rect 22649 18105 22661 18139
rect 22695 18136 22707 18139
rect 24026 18136 24032 18148
rect 22695 18108 24032 18136
rect 22695 18105 22707 18108
rect 22649 18099 22707 18105
rect 9824 18040 11008 18068
rect 11977 18071 12035 18077
rect 9824 18028 9830 18040
rect 11977 18037 11989 18071
rect 12023 18068 12035 18071
rect 12526 18068 12532 18080
rect 12023 18040 12532 18068
rect 12023 18037 12035 18040
rect 11977 18031 12035 18037
rect 12526 18028 12532 18040
rect 12584 18028 12590 18080
rect 15933 18071 15991 18077
rect 15933 18037 15945 18071
rect 15979 18068 15991 18071
rect 16022 18068 16028 18080
rect 15979 18040 16028 18068
rect 15979 18037 15991 18040
rect 15933 18031 15991 18037
rect 16022 18028 16028 18040
rect 16080 18028 16086 18080
rect 16666 18028 16672 18080
rect 16724 18068 16730 18080
rect 17126 18068 17132 18080
rect 16724 18040 17132 18068
rect 16724 18028 16730 18040
rect 17126 18028 17132 18040
rect 17184 18068 17190 18080
rect 17405 18071 17463 18077
rect 17405 18068 17417 18071
rect 17184 18040 17417 18068
rect 17184 18028 17190 18040
rect 17405 18037 17417 18040
rect 17451 18037 17463 18071
rect 18598 18068 18604 18080
rect 18559 18040 18604 18068
rect 17405 18031 17463 18037
rect 18598 18028 18604 18040
rect 18656 18028 18662 18080
rect 22094 18028 22100 18080
rect 22152 18068 22158 18080
rect 22664 18068 22692 18099
rect 24026 18096 24032 18108
rect 24084 18096 24090 18148
rect 24688 18145 24716 18380
rect 25038 18368 25044 18380
rect 25096 18368 25102 18420
rect 25501 18411 25559 18417
rect 25501 18377 25513 18411
rect 25547 18408 25559 18411
rect 25774 18408 25780 18420
rect 25547 18380 25780 18408
rect 25547 18377 25559 18380
rect 25501 18371 25559 18377
rect 25774 18368 25780 18380
rect 25832 18368 25838 18420
rect 24397 18139 24455 18145
rect 24397 18105 24409 18139
rect 24443 18105 24455 18139
rect 24397 18099 24455 18105
rect 24673 18139 24731 18145
rect 24673 18105 24685 18139
rect 24719 18105 24731 18139
rect 24673 18099 24731 18105
rect 22152 18040 22692 18068
rect 22152 18028 22158 18040
rect 23842 18028 23848 18080
rect 23900 18068 23906 18080
rect 24412 18068 24440 18099
rect 24578 18068 24584 18080
rect 23900 18040 24440 18068
rect 24539 18040 24584 18068
rect 23900 18028 23906 18040
rect 24578 18028 24584 18040
rect 24636 18028 24642 18080
rect 24688 18068 24716 18099
rect 25498 18068 25504 18080
rect 24688 18040 25504 18068
rect 25498 18028 25504 18040
rect 25556 18068 25562 18080
rect 25777 18071 25835 18077
rect 25777 18068 25789 18071
rect 25556 18040 25789 18068
rect 25556 18028 25562 18040
rect 25777 18037 25789 18040
rect 25823 18037 25835 18071
rect 25777 18031 25835 18037
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 2774 17824 2780 17876
rect 2832 17864 2838 17876
rect 2832 17836 2877 17864
rect 2832 17824 2838 17836
rect 2958 17824 2964 17876
rect 3016 17864 3022 17876
rect 3421 17867 3479 17873
rect 3421 17864 3433 17867
rect 3016 17836 3433 17864
rect 3016 17824 3022 17836
rect 3421 17833 3433 17836
rect 3467 17833 3479 17867
rect 3421 17827 3479 17833
rect 3881 17867 3939 17873
rect 3881 17833 3893 17867
rect 3927 17864 3939 17867
rect 4154 17864 4160 17876
rect 3927 17836 4160 17864
rect 3927 17833 3939 17836
rect 3881 17827 3939 17833
rect 4154 17824 4160 17836
rect 4212 17824 4218 17876
rect 4338 17864 4344 17876
rect 4299 17836 4344 17864
rect 4338 17824 4344 17836
rect 4396 17824 4402 17876
rect 4433 17867 4491 17873
rect 4433 17833 4445 17867
rect 4479 17864 4491 17867
rect 5258 17864 5264 17876
rect 4479 17836 5264 17864
rect 4479 17833 4491 17836
rect 4433 17827 4491 17833
rect 5258 17824 5264 17836
rect 5316 17824 5322 17876
rect 5442 17824 5448 17876
rect 5500 17864 5506 17876
rect 6825 17867 6883 17873
rect 6825 17864 6837 17867
rect 5500 17836 6837 17864
rect 5500 17824 5506 17836
rect 6825 17833 6837 17836
rect 6871 17864 6883 17867
rect 6914 17864 6920 17876
rect 6871 17836 6920 17864
rect 6871 17833 6883 17836
rect 6825 17827 6883 17833
rect 6914 17824 6920 17836
rect 6972 17824 6978 17876
rect 8573 17867 8631 17873
rect 8573 17833 8585 17867
rect 8619 17864 8631 17867
rect 8662 17864 8668 17876
rect 8619 17836 8668 17864
rect 8619 17833 8631 17836
rect 8573 17827 8631 17833
rect 8662 17824 8668 17836
rect 8720 17824 8726 17876
rect 9306 17864 9312 17876
rect 9267 17836 9312 17864
rect 9306 17824 9312 17836
rect 9364 17864 9370 17876
rect 10137 17867 10195 17873
rect 10137 17864 10149 17867
rect 9364 17836 10149 17864
rect 9364 17824 9370 17836
rect 10137 17833 10149 17836
rect 10183 17864 10195 17867
rect 10778 17864 10784 17876
rect 10183 17836 10784 17864
rect 10183 17833 10195 17836
rect 10137 17827 10195 17833
rect 10778 17824 10784 17836
rect 10836 17824 10842 17876
rect 13354 17864 13360 17876
rect 13315 17836 13360 17864
rect 13354 17824 13360 17836
rect 13412 17824 13418 17876
rect 14185 17867 14243 17873
rect 14185 17833 14197 17867
rect 14231 17864 14243 17867
rect 14550 17864 14556 17876
rect 14231 17836 14556 17864
rect 14231 17833 14243 17836
rect 14185 17827 14243 17833
rect 14550 17824 14556 17836
rect 14608 17824 14614 17876
rect 16114 17864 16120 17876
rect 16075 17836 16120 17864
rect 16114 17824 16120 17836
rect 16172 17824 16178 17876
rect 16482 17864 16488 17876
rect 16443 17836 16488 17864
rect 16482 17824 16488 17836
rect 16540 17824 16546 17876
rect 18966 17824 18972 17876
rect 19024 17864 19030 17876
rect 19518 17864 19524 17876
rect 19024 17836 19524 17864
rect 19024 17824 19030 17836
rect 19518 17824 19524 17836
rect 19576 17864 19582 17876
rect 19576 17836 19932 17864
rect 19576 17824 19582 17836
rect 2225 17799 2283 17805
rect 2225 17765 2237 17799
rect 2271 17796 2283 17799
rect 3234 17796 3240 17808
rect 2271 17768 3240 17796
rect 2271 17765 2283 17768
rect 2225 17759 2283 17765
rect 3234 17756 3240 17768
rect 3292 17796 3298 17808
rect 4522 17796 4528 17808
rect 3292 17768 4528 17796
rect 3292 17756 3298 17768
rect 4522 17756 4528 17768
rect 4580 17756 4586 17808
rect 4798 17756 4804 17808
rect 4856 17796 4862 17808
rect 4893 17799 4951 17805
rect 4893 17796 4905 17799
rect 4856 17768 4905 17796
rect 4856 17756 4862 17768
rect 4893 17765 4905 17768
rect 4939 17765 4951 17799
rect 4893 17759 4951 17765
rect 7745 17799 7803 17805
rect 7745 17765 7757 17799
rect 7791 17796 7803 17799
rect 7834 17796 7840 17808
rect 7791 17768 7840 17796
rect 7791 17765 7803 17768
rect 7745 17759 7803 17765
rect 7834 17756 7840 17768
rect 7892 17756 7898 17808
rect 15565 17799 15623 17805
rect 15565 17765 15577 17799
rect 15611 17796 15623 17799
rect 15654 17796 15660 17808
rect 15611 17768 15660 17796
rect 15611 17765 15623 17768
rect 15565 17759 15623 17765
rect 15654 17756 15660 17768
rect 15712 17756 15718 17808
rect 19610 17756 19616 17808
rect 19668 17796 19674 17808
rect 19904 17805 19932 17836
rect 21174 17824 21180 17876
rect 21232 17864 21238 17876
rect 21269 17867 21327 17873
rect 21269 17864 21281 17867
rect 21232 17836 21281 17864
rect 21232 17824 21238 17836
rect 21269 17833 21281 17836
rect 21315 17833 21327 17867
rect 21269 17827 21327 17833
rect 22094 17824 22100 17876
rect 22152 17864 22158 17876
rect 22152 17836 22197 17864
rect 22152 17824 22158 17836
rect 19797 17799 19855 17805
rect 19797 17796 19809 17799
rect 19668 17768 19809 17796
rect 19668 17756 19674 17768
rect 19797 17765 19809 17768
rect 19843 17765 19855 17799
rect 19797 17759 19855 17765
rect 19889 17799 19947 17805
rect 19889 17765 19901 17799
rect 19935 17765 19947 17799
rect 19889 17759 19947 17765
rect 23474 17756 23480 17808
rect 23532 17796 23538 17808
rect 24121 17799 24179 17805
rect 24121 17796 24133 17799
rect 23532 17768 24133 17796
rect 23532 17756 23538 17768
rect 24121 17765 24133 17768
rect 24167 17796 24179 17799
rect 24578 17796 24584 17808
rect 24167 17768 24584 17796
rect 24167 17765 24179 17768
rect 24121 17759 24179 17765
rect 24578 17756 24584 17768
rect 24636 17796 24642 17808
rect 24946 17796 24952 17808
rect 24636 17768 24952 17796
rect 24636 17756 24642 17768
rect 24946 17756 24952 17768
rect 25004 17756 25010 17808
rect 25038 17756 25044 17808
rect 25096 17796 25102 17808
rect 25225 17799 25283 17805
rect 25225 17796 25237 17799
rect 25096 17768 25237 17796
rect 25096 17756 25102 17768
rect 25225 17765 25237 17768
rect 25271 17765 25283 17799
rect 25225 17759 25283 17765
rect 5534 17688 5540 17740
rect 5592 17728 5598 17740
rect 11054 17737 11060 17740
rect 5701 17731 5759 17737
rect 5701 17728 5713 17731
rect 5592 17700 5713 17728
rect 5592 17688 5598 17700
rect 5701 17697 5713 17700
rect 5747 17697 5759 17731
rect 11048 17728 11060 17737
rect 11015 17700 11060 17728
rect 5701 17691 5759 17697
rect 11048 17691 11060 17700
rect 11054 17688 11060 17691
rect 11112 17688 11118 17740
rect 13906 17688 13912 17740
rect 13964 17728 13970 17740
rect 14277 17731 14335 17737
rect 14277 17728 14289 17731
rect 13964 17700 14289 17728
rect 13964 17688 13970 17700
rect 14277 17697 14289 17700
rect 14323 17697 14335 17731
rect 15286 17728 15292 17740
rect 15247 17700 15292 17728
rect 14277 17691 14335 17697
rect 15286 17688 15292 17700
rect 15344 17688 15350 17740
rect 16942 17737 16948 17740
rect 16936 17728 16948 17737
rect 16903 17700 16948 17728
rect 16936 17691 16948 17700
rect 16942 17688 16948 17691
rect 17000 17688 17006 17740
rect 21450 17688 21456 17740
rect 21508 17728 21514 17740
rect 22445 17731 22503 17737
rect 22445 17728 22457 17731
rect 21508 17700 22457 17728
rect 21508 17688 21514 17700
rect 22445 17697 22457 17700
rect 22491 17728 22503 17731
rect 23566 17728 23572 17740
rect 22491 17700 23572 17728
rect 22491 17697 22503 17700
rect 22445 17691 22503 17697
rect 23566 17688 23572 17700
rect 23624 17688 23630 17740
rect 2222 17660 2228 17672
rect 2183 17632 2228 17660
rect 2222 17620 2228 17632
rect 2280 17620 2286 17672
rect 2317 17663 2375 17669
rect 2317 17629 2329 17663
rect 2363 17660 2375 17663
rect 2682 17660 2688 17672
rect 2363 17632 2688 17660
rect 2363 17629 2375 17632
rect 2317 17623 2375 17629
rect 2682 17620 2688 17632
rect 2740 17660 2746 17672
rect 3053 17663 3111 17669
rect 3053 17660 3065 17663
rect 2740 17632 3065 17660
rect 2740 17620 2746 17632
rect 3053 17629 3065 17632
rect 3099 17629 3111 17663
rect 3053 17623 3111 17629
rect 5445 17663 5503 17669
rect 5445 17629 5457 17663
rect 5491 17629 5503 17663
rect 5445 17623 5503 17629
rect 8481 17663 8539 17669
rect 8481 17629 8493 17663
rect 8527 17629 8539 17663
rect 8662 17660 8668 17672
rect 8623 17632 8668 17660
rect 8481 17623 8539 17629
rect 1762 17592 1768 17604
rect 1723 17564 1768 17592
rect 1762 17552 1768 17564
rect 1820 17552 1826 17604
rect 5460 17524 5488 17623
rect 8113 17595 8171 17601
rect 8113 17561 8125 17595
rect 8159 17592 8171 17595
rect 8202 17592 8208 17604
rect 8159 17564 8208 17592
rect 8159 17561 8171 17564
rect 8113 17555 8171 17561
rect 8202 17552 8208 17564
rect 8260 17552 8266 17604
rect 8496 17592 8524 17623
rect 8662 17620 8668 17632
rect 8720 17620 8726 17672
rect 9674 17660 9680 17672
rect 9635 17632 9680 17660
rect 9674 17620 9680 17632
rect 9732 17620 9738 17672
rect 10778 17660 10784 17672
rect 10739 17632 10784 17660
rect 10778 17620 10784 17632
rect 10836 17620 10842 17672
rect 13630 17620 13636 17672
rect 13688 17660 13694 17672
rect 14182 17660 14188 17672
rect 13688 17632 14188 17660
rect 13688 17620 13694 17632
rect 14182 17620 14188 17632
rect 14240 17620 14246 17672
rect 16666 17660 16672 17672
rect 16627 17632 16672 17660
rect 16666 17620 16672 17632
rect 16724 17620 16730 17672
rect 19797 17663 19855 17669
rect 19797 17629 19809 17663
rect 19843 17660 19855 17663
rect 19978 17660 19984 17672
rect 19843 17632 19984 17660
rect 19843 17629 19855 17632
rect 19797 17623 19855 17629
rect 19978 17620 19984 17632
rect 20036 17620 20042 17672
rect 22186 17660 22192 17672
rect 22147 17632 22192 17660
rect 22186 17620 22192 17632
rect 22244 17620 22250 17672
rect 25130 17660 25136 17672
rect 25091 17632 25136 17660
rect 25130 17620 25136 17632
rect 25188 17620 25194 17672
rect 25317 17663 25375 17669
rect 25317 17629 25329 17663
rect 25363 17660 25375 17663
rect 25498 17660 25504 17672
rect 25363 17632 25504 17660
rect 25363 17629 25375 17632
rect 25317 17623 25375 17629
rect 25498 17620 25504 17632
rect 25556 17620 25562 17672
rect 9030 17592 9036 17604
rect 8496 17564 9036 17592
rect 9030 17552 9036 17564
rect 9088 17592 9094 17604
rect 9582 17592 9588 17604
rect 9088 17564 9588 17592
rect 9088 17552 9094 17564
rect 9582 17552 9588 17564
rect 9640 17552 9646 17604
rect 13722 17592 13728 17604
rect 13683 17564 13728 17592
rect 13722 17552 13728 17564
rect 13780 17552 13786 17604
rect 24026 17552 24032 17604
rect 24084 17592 24090 17604
rect 24489 17595 24547 17601
rect 24489 17592 24501 17595
rect 24084 17564 24501 17592
rect 24084 17552 24090 17564
rect 24489 17561 24501 17564
rect 24535 17561 24547 17595
rect 24489 17555 24547 17561
rect 24670 17552 24676 17604
rect 24728 17592 24734 17604
rect 24765 17595 24823 17601
rect 24765 17592 24777 17595
rect 24728 17564 24777 17592
rect 24728 17552 24734 17564
rect 24765 17561 24777 17564
rect 24811 17561 24823 17595
rect 24765 17555 24823 17561
rect 6178 17524 6184 17536
rect 5460 17496 6184 17524
rect 6178 17484 6184 17496
rect 6236 17484 6242 17536
rect 10597 17527 10655 17533
rect 10597 17493 10609 17527
rect 10643 17524 10655 17527
rect 10962 17524 10968 17536
rect 10643 17496 10968 17524
rect 10643 17493 10655 17496
rect 10597 17487 10655 17493
rect 10962 17484 10968 17496
rect 11020 17524 11026 17536
rect 12158 17524 12164 17536
rect 11020 17496 12164 17524
rect 11020 17484 11026 17496
rect 12158 17484 12164 17496
rect 12216 17484 12222 17536
rect 12526 17484 12532 17536
rect 12584 17524 12590 17536
rect 12713 17527 12771 17533
rect 12713 17524 12725 17527
rect 12584 17496 12725 17524
rect 12584 17484 12590 17496
rect 12713 17493 12725 17496
rect 12759 17493 12771 17527
rect 14826 17524 14832 17536
rect 14787 17496 14832 17524
rect 12713 17487 12771 17493
rect 14826 17484 14832 17496
rect 14884 17484 14890 17536
rect 18046 17524 18052 17536
rect 18007 17496 18052 17524
rect 18046 17484 18052 17496
rect 18104 17484 18110 17536
rect 19337 17527 19395 17533
rect 19337 17493 19349 17527
rect 19383 17524 19395 17527
rect 20162 17524 20168 17536
rect 19383 17496 20168 17524
rect 19383 17493 19395 17496
rect 19337 17487 19395 17493
rect 20162 17484 20168 17496
rect 20220 17484 20226 17536
rect 23382 17484 23388 17536
rect 23440 17524 23446 17536
rect 23569 17527 23627 17533
rect 23569 17524 23581 17527
rect 23440 17496 23581 17524
rect 23440 17484 23446 17496
rect 23569 17493 23581 17496
rect 23615 17493 23627 17527
rect 23569 17487 23627 17493
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 4985 17323 5043 17329
rect 4985 17289 4997 17323
rect 5031 17320 5043 17323
rect 5166 17320 5172 17332
rect 5031 17292 5172 17320
rect 5031 17289 5043 17292
rect 4985 17283 5043 17289
rect 5166 17280 5172 17292
rect 5224 17280 5230 17332
rect 7190 17280 7196 17332
rect 7248 17320 7254 17332
rect 8018 17320 8024 17332
rect 7248 17292 8024 17320
rect 7248 17280 7254 17292
rect 8018 17280 8024 17292
rect 8076 17280 8082 17332
rect 8662 17280 8668 17332
rect 8720 17320 8726 17332
rect 8757 17323 8815 17329
rect 8757 17320 8769 17323
rect 8720 17292 8769 17320
rect 8720 17280 8726 17292
rect 8757 17289 8769 17292
rect 8803 17320 8815 17323
rect 10689 17323 10747 17329
rect 10689 17320 10701 17323
rect 8803 17292 10701 17320
rect 8803 17289 8815 17292
rect 8757 17283 8815 17289
rect 10689 17289 10701 17292
rect 10735 17320 10747 17323
rect 11054 17320 11060 17332
rect 10735 17292 11060 17320
rect 10735 17289 10747 17292
rect 10689 17283 10747 17289
rect 11054 17280 11060 17292
rect 11112 17320 11118 17332
rect 11609 17323 11667 17329
rect 11609 17320 11621 17323
rect 11112 17292 11621 17320
rect 11112 17280 11118 17292
rect 11609 17289 11621 17292
rect 11655 17289 11667 17323
rect 11609 17283 11667 17289
rect 15838 17280 15844 17332
rect 15896 17320 15902 17332
rect 16485 17323 16543 17329
rect 16485 17320 16497 17323
rect 15896 17292 16497 17320
rect 15896 17280 15902 17292
rect 16485 17289 16497 17292
rect 16531 17289 16543 17323
rect 16485 17283 16543 17289
rect 16574 17280 16580 17332
rect 16632 17320 16638 17332
rect 17405 17323 17463 17329
rect 17405 17320 17417 17323
rect 16632 17292 17417 17320
rect 16632 17280 16638 17292
rect 17405 17289 17417 17292
rect 17451 17320 17463 17323
rect 18046 17320 18052 17332
rect 17451 17292 18052 17320
rect 17451 17289 17463 17292
rect 17405 17283 17463 17289
rect 18046 17280 18052 17292
rect 18104 17280 18110 17332
rect 19518 17280 19524 17332
rect 19576 17320 19582 17332
rect 21450 17320 21456 17332
rect 19576 17292 21456 17320
rect 19576 17280 19582 17292
rect 21450 17280 21456 17292
rect 21508 17280 21514 17332
rect 22186 17280 22192 17332
rect 22244 17320 22250 17332
rect 23014 17320 23020 17332
rect 22244 17292 23020 17320
rect 22244 17280 22250 17292
rect 23014 17280 23020 17292
rect 23072 17280 23078 17332
rect 4433 17255 4491 17261
rect 4433 17221 4445 17255
rect 4479 17252 4491 17255
rect 5534 17252 5540 17264
rect 4479 17224 5540 17252
rect 4479 17221 4491 17224
rect 4433 17215 4491 17221
rect 5534 17212 5540 17224
rect 5592 17212 5598 17264
rect 4798 17144 4804 17196
rect 4856 17184 4862 17196
rect 18064 17184 18092 17280
rect 19610 17212 19616 17264
rect 19668 17252 19674 17264
rect 19981 17255 20039 17261
rect 19981 17252 19993 17255
rect 19668 17224 19993 17252
rect 19668 17212 19674 17224
rect 19981 17221 19993 17224
rect 20027 17252 20039 17255
rect 20346 17252 20352 17264
rect 20027 17224 20352 17252
rect 20027 17221 20039 17224
rect 19981 17215 20039 17221
rect 20346 17212 20352 17224
rect 20404 17212 20410 17264
rect 22097 17255 22155 17261
rect 22097 17221 22109 17255
rect 22143 17252 22155 17255
rect 22830 17252 22836 17264
rect 22143 17224 22836 17252
rect 22143 17221 22155 17224
rect 22097 17215 22155 17221
rect 22830 17212 22836 17224
rect 22888 17212 22894 17264
rect 23753 17255 23811 17261
rect 23753 17221 23765 17255
rect 23799 17252 23811 17255
rect 23934 17252 23940 17264
rect 23799 17224 23940 17252
rect 23799 17221 23811 17224
rect 23753 17215 23811 17221
rect 23934 17212 23940 17224
rect 23992 17212 23998 17264
rect 22554 17184 22560 17196
rect 4856 17156 5396 17184
rect 18064 17156 18184 17184
rect 22515 17156 22560 17184
rect 4856 17144 4862 17156
rect 2406 17116 2412 17128
rect 2367 17088 2412 17116
rect 2406 17076 2412 17088
rect 2464 17076 2470 17128
rect 2682 17125 2688 17128
rect 2676 17116 2688 17125
rect 2516 17088 2688 17116
rect 1670 17008 1676 17060
rect 1728 17048 1734 17060
rect 1765 17051 1823 17057
rect 1765 17048 1777 17051
rect 1728 17020 1777 17048
rect 1728 17008 1734 17020
rect 1765 17017 1777 17020
rect 1811 17048 1823 17051
rect 2516 17048 2544 17088
rect 2676 17079 2688 17088
rect 2682 17076 2688 17079
rect 2740 17076 2746 17128
rect 1811 17020 2544 17048
rect 5261 17051 5319 17057
rect 1811 17017 1823 17020
rect 1765 17011 1823 17017
rect 5261 17017 5273 17051
rect 5307 17017 5319 17051
rect 5261 17011 5319 17017
rect 1578 16940 1584 16992
rect 1636 16980 1642 16992
rect 2225 16983 2283 16989
rect 2225 16980 2237 16983
rect 1636 16952 2237 16980
rect 1636 16940 1642 16952
rect 2225 16949 2237 16952
rect 2271 16980 2283 16983
rect 2406 16980 2412 16992
rect 2271 16952 2412 16980
rect 2271 16949 2283 16952
rect 2225 16943 2283 16949
rect 2406 16940 2412 16952
rect 2464 16940 2470 16992
rect 3418 16940 3424 16992
rect 3476 16980 3482 16992
rect 3789 16983 3847 16989
rect 3789 16980 3801 16983
rect 3476 16952 3801 16980
rect 3476 16940 3482 16952
rect 3789 16949 3801 16952
rect 3835 16949 3847 16983
rect 3789 16943 3847 16949
rect 4154 16940 4160 16992
rect 4212 16980 4218 16992
rect 4709 16983 4767 16989
rect 4709 16980 4721 16983
rect 4212 16952 4721 16980
rect 4212 16940 4218 16952
rect 4709 16949 4721 16952
rect 4755 16980 4767 16983
rect 5276 16980 5304 17011
rect 4755 16952 5304 16980
rect 5368 16980 5396 17156
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17085 6883 17119
rect 6825 17079 6883 17085
rect 5534 17048 5540 17060
rect 5495 17020 5540 17048
rect 5534 17008 5540 17020
rect 5592 17008 5598 17060
rect 5997 17051 6055 17057
rect 5997 17017 6009 17051
rect 6043 17048 6055 17051
rect 6178 17048 6184 17060
rect 6043 17020 6184 17048
rect 6043 17017 6055 17020
rect 5997 17011 6055 17017
rect 6178 17008 6184 17020
rect 6236 17048 6242 17060
rect 6641 17051 6699 17057
rect 6641 17048 6653 17051
rect 6236 17020 6653 17048
rect 6236 17008 6242 17020
rect 6641 17017 6653 17020
rect 6687 17048 6699 17051
rect 6840 17048 6868 17079
rect 6914 17076 6920 17128
rect 6972 17116 6978 17128
rect 7081 17119 7139 17125
rect 7081 17116 7093 17119
rect 6972 17088 7093 17116
rect 6972 17076 6978 17088
rect 7081 17085 7093 17088
rect 7127 17085 7139 17119
rect 7081 17079 7139 17085
rect 9309 17119 9367 17125
rect 9309 17085 9321 17119
rect 9355 17085 9367 17119
rect 9309 17079 9367 17085
rect 6687 17020 9076 17048
rect 6687 17017 6699 17020
rect 6641 17011 6699 17017
rect 9048 16992 9076 17020
rect 5445 16983 5503 16989
rect 5445 16980 5457 16983
rect 5368 16952 5457 16980
rect 4755 16949 4767 16952
rect 4709 16943 4767 16949
rect 5445 16949 5457 16952
rect 5491 16949 5503 16983
rect 8202 16980 8208 16992
rect 8163 16952 8208 16980
rect 5445 16943 5503 16949
rect 8202 16940 8208 16952
rect 8260 16940 8266 16992
rect 9030 16940 9036 16992
rect 9088 16980 9094 16992
rect 9125 16983 9183 16989
rect 9125 16980 9137 16983
rect 9088 16952 9137 16980
rect 9088 16940 9094 16952
rect 9125 16949 9137 16952
rect 9171 16980 9183 16983
rect 9324 16980 9352 17079
rect 9398 17076 9404 17128
rect 9456 17116 9462 17128
rect 9565 17119 9623 17125
rect 9565 17116 9577 17119
rect 9456 17088 9577 17116
rect 9456 17076 9462 17088
rect 9565 17085 9577 17088
rect 9611 17116 9623 17119
rect 10134 17116 10140 17128
rect 9611 17088 10140 17116
rect 9611 17085 9623 17088
rect 9565 17079 9623 17085
rect 10134 17076 10140 17088
rect 10192 17076 10198 17128
rect 12621 17119 12679 17125
rect 12621 17116 12633 17119
rect 12176 17088 12633 17116
rect 10778 16980 10784 16992
rect 9171 16952 10784 16980
rect 9171 16949 9183 16952
rect 9125 16943 9183 16949
rect 10778 16940 10784 16952
rect 10836 16980 10842 16992
rect 12176 16989 12204 17088
rect 12621 17085 12633 17088
rect 12667 17085 12679 17119
rect 12621 17079 12679 17085
rect 15105 17119 15163 17125
rect 15105 17085 15117 17119
rect 15151 17116 15163 17119
rect 15194 17116 15200 17128
rect 15151 17088 15200 17116
rect 15151 17085 15163 17088
rect 15105 17079 15163 17085
rect 15194 17076 15200 17088
rect 15252 17076 15258 17128
rect 18049 17119 18107 17125
rect 18049 17116 18061 17119
rect 17788 17088 18061 17116
rect 12526 17008 12532 17060
rect 12584 17048 12590 17060
rect 12888 17051 12946 17057
rect 12888 17048 12900 17051
rect 12584 17020 12900 17048
rect 12584 17008 12590 17020
rect 12888 17017 12900 17020
rect 12934 17048 12946 17051
rect 13538 17048 13544 17060
rect 12934 17020 13544 17048
rect 12934 17017 12946 17020
rect 12888 17011 12946 17017
rect 13538 17008 13544 17020
rect 13596 17008 13602 17060
rect 15350 17051 15408 17057
rect 15350 17048 15362 17051
rect 14568 17020 15362 17048
rect 11241 16983 11299 16989
rect 11241 16980 11253 16983
rect 10836 16952 11253 16980
rect 10836 16940 10842 16952
rect 11241 16949 11253 16952
rect 11287 16980 11299 16983
rect 12161 16983 12219 16989
rect 12161 16980 12173 16983
rect 11287 16952 12173 16980
rect 11287 16949 11299 16952
rect 11241 16943 11299 16949
rect 12161 16949 12173 16952
rect 12207 16949 12219 16983
rect 12161 16943 12219 16949
rect 13354 16940 13360 16992
rect 13412 16980 13418 16992
rect 14568 16989 14596 17020
rect 15350 17017 15362 17020
rect 15396 17017 15408 17051
rect 15350 17011 15408 17017
rect 14001 16983 14059 16989
rect 14001 16980 14013 16983
rect 13412 16952 14013 16980
rect 13412 16940 13418 16952
rect 14001 16949 14013 16952
rect 14047 16980 14059 16983
rect 14553 16983 14611 16989
rect 14553 16980 14565 16983
rect 14047 16952 14565 16980
rect 14047 16949 14059 16952
rect 14001 16943 14059 16949
rect 14553 16949 14565 16952
rect 14599 16949 14611 16983
rect 14553 16943 14611 16949
rect 15013 16983 15071 16989
rect 15013 16949 15025 16983
rect 15059 16980 15071 16983
rect 15194 16980 15200 16992
rect 15059 16952 15200 16980
rect 15059 16949 15071 16952
rect 15013 16943 15071 16949
rect 15194 16940 15200 16952
rect 15252 16980 15258 16992
rect 16666 16980 16672 16992
rect 15252 16952 16672 16980
rect 15252 16940 15258 16952
rect 16666 16940 16672 16952
rect 16724 16980 16730 16992
rect 17788 16989 17816 17088
rect 18049 17085 18061 17088
rect 18095 17085 18107 17119
rect 18156 17116 18184 17156
rect 22554 17144 22560 17156
rect 22612 17144 22618 17196
rect 25222 17184 25228 17196
rect 25183 17156 25228 17184
rect 25222 17144 25228 17156
rect 25280 17144 25286 17196
rect 18305 17119 18363 17125
rect 18305 17116 18317 17119
rect 18156 17088 18317 17116
rect 18049 17079 18107 17085
rect 18305 17085 18317 17088
rect 18351 17085 18363 17119
rect 18305 17079 18363 17085
rect 20990 17008 20996 17060
rect 21048 17048 21054 17060
rect 21085 17051 21143 17057
rect 21085 17048 21097 17051
rect 21048 17020 21097 17048
rect 21048 17008 21054 17020
rect 21085 17017 21097 17020
rect 21131 17048 21143 17051
rect 22557 17051 22615 17057
rect 22557 17048 22569 17051
rect 21131 17020 22569 17048
rect 21131 17017 21143 17020
rect 21085 17011 21143 17017
rect 22557 17017 22569 17020
rect 22603 17017 22615 17051
rect 22557 17011 22615 17017
rect 22649 17051 22707 17057
rect 22649 17017 22661 17051
rect 22695 17048 22707 17051
rect 22738 17048 22744 17060
rect 22695 17020 22744 17048
rect 22695 17017 22707 17020
rect 22649 17011 22707 17017
rect 22738 17008 22744 17020
rect 22796 17008 22802 17060
rect 24026 17048 24032 17060
rect 23987 17020 24032 17048
rect 24026 17008 24032 17020
rect 24084 17008 24090 17060
rect 24118 17008 24124 17060
rect 24176 17048 24182 17060
rect 24213 17051 24271 17057
rect 24213 17048 24225 17051
rect 24176 17020 24225 17048
rect 24176 17008 24182 17020
rect 24213 17017 24225 17020
rect 24259 17017 24271 17051
rect 24213 17011 24271 17017
rect 24305 17051 24363 17057
rect 24305 17017 24317 17051
rect 24351 17017 24363 17051
rect 24305 17011 24363 17017
rect 24765 17051 24823 17057
rect 24765 17017 24777 17051
rect 24811 17048 24823 17051
rect 25130 17048 25136 17060
rect 24811 17020 25136 17048
rect 24811 17017 24823 17020
rect 24765 17011 24823 17017
rect 17037 16983 17095 16989
rect 17037 16980 17049 16983
rect 16724 16952 17049 16980
rect 16724 16940 16730 16952
rect 17037 16949 17049 16952
rect 17083 16980 17095 16983
rect 17773 16983 17831 16989
rect 17773 16980 17785 16983
rect 17083 16952 17785 16980
rect 17083 16949 17095 16952
rect 17037 16943 17095 16949
rect 17773 16949 17785 16952
rect 17819 16949 17831 16983
rect 19426 16980 19432 16992
rect 19387 16952 19432 16980
rect 17773 16943 17831 16949
rect 19426 16940 19432 16952
rect 19484 16940 19490 16992
rect 21818 16980 21824 16992
rect 21779 16952 21824 16980
rect 21818 16940 21824 16952
rect 21876 16940 21882 16992
rect 23382 16980 23388 16992
rect 23343 16952 23388 16980
rect 23382 16940 23388 16952
rect 23440 16980 23446 16992
rect 24320 16980 24348 17011
rect 25130 17008 25136 17020
rect 25188 17008 25194 17060
rect 25038 16980 25044 16992
rect 23440 16952 24348 16980
rect 24999 16952 25044 16980
rect 23440 16940 23446 16952
rect 25038 16940 25044 16952
rect 25096 16940 25102 16992
rect 25498 16940 25504 16992
rect 25556 16980 25562 16992
rect 25685 16983 25743 16989
rect 25685 16980 25697 16983
rect 25556 16952 25697 16980
rect 25556 16940 25562 16952
rect 25685 16949 25697 16952
rect 25731 16949 25743 16983
rect 25685 16943 25743 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1670 16776 1676 16788
rect 1631 16748 1676 16776
rect 1670 16736 1676 16748
rect 1728 16736 1734 16788
rect 1762 16736 1768 16788
rect 1820 16736 1826 16788
rect 2222 16736 2228 16788
rect 2280 16776 2286 16788
rect 3513 16779 3571 16785
rect 3513 16776 3525 16779
rect 2280 16748 3525 16776
rect 2280 16736 2286 16748
rect 3513 16745 3525 16748
rect 3559 16745 3571 16779
rect 5442 16776 5448 16788
rect 5403 16748 5448 16776
rect 3513 16739 3571 16745
rect 5442 16736 5448 16748
rect 5500 16736 5506 16788
rect 5534 16736 5540 16788
rect 5592 16776 5598 16788
rect 5997 16779 6055 16785
rect 5997 16776 6009 16779
rect 5592 16748 6009 16776
rect 5592 16736 5598 16748
rect 5997 16745 6009 16748
rect 6043 16745 6055 16779
rect 6914 16776 6920 16788
rect 6875 16748 6920 16776
rect 5997 16739 6055 16745
rect 6914 16736 6920 16748
rect 6972 16736 6978 16788
rect 8573 16779 8631 16785
rect 8573 16745 8585 16779
rect 8619 16776 8631 16779
rect 8754 16776 8760 16788
rect 8619 16748 8760 16776
rect 8619 16745 8631 16748
rect 8573 16739 8631 16745
rect 8754 16736 8760 16748
rect 8812 16736 8818 16788
rect 9122 16776 9128 16788
rect 9083 16748 9128 16776
rect 9122 16736 9128 16748
rect 9180 16776 9186 16788
rect 9858 16776 9864 16788
rect 9180 16748 9864 16776
rect 9180 16736 9186 16748
rect 9858 16736 9864 16748
rect 9916 16736 9922 16788
rect 11977 16779 12035 16785
rect 11977 16745 11989 16779
rect 12023 16776 12035 16779
rect 12342 16776 12348 16788
rect 12023 16748 12348 16776
rect 12023 16745 12035 16748
rect 11977 16739 12035 16745
rect 12342 16736 12348 16748
rect 12400 16736 12406 16788
rect 12611 16779 12669 16785
rect 12611 16745 12623 16779
rect 12657 16776 12669 16779
rect 12657 16748 14136 16776
rect 12657 16745 12669 16748
rect 12611 16739 12669 16745
rect 1780 16708 1808 16736
rect 2317 16711 2375 16717
rect 2317 16708 2329 16711
rect 1780 16680 2329 16708
rect 2317 16677 2329 16680
rect 2363 16677 2375 16711
rect 2317 16671 2375 16677
rect 2409 16711 2467 16717
rect 2409 16677 2421 16711
rect 2455 16708 2467 16711
rect 3418 16708 3424 16720
rect 2455 16680 3424 16708
rect 2455 16677 2467 16680
rect 2409 16671 2467 16677
rect 3418 16668 3424 16680
rect 3476 16708 3482 16720
rect 4310 16711 4368 16717
rect 4310 16708 4322 16711
rect 3476 16680 4322 16708
rect 3476 16668 3482 16680
rect 4310 16677 4322 16680
rect 4356 16677 4368 16711
rect 4310 16671 4368 16677
rect 7929 16711 7987 16717
rect 7929 16677 7941 16711
rect 7975 16708 7987 16711
rect 8202 16708 8208 16720
rect 7975 16680 8208 16708
rect 7975 16677 7987 16680
rect 7929 16671 7987 16677
rect 8202 16668 8208 16680
rect 8260 16708 8266 16720
rect 8260 16680 8524 16708
rect 8260 16668 8266 16680
rect 1839 16643 1897 16649
rect 1839 16609 1851 16643
rect 1885 16640 1897 16643
rect 1946 16640 1952 16652
rect 1885 16612 1952 16640
rect 1885 16609 1897 16612
rect 1839 16603 1897 16609
rect 1946 16600 1952 16612
rect 2004 16600 2010 16652
rect 2130 16640 2136 16652
rect 2091 16612 2136 16640
rect 2130 16600 2136 16612
rect 2188 16600 2194 16652
rect 2866 16640 2872 16652
rect 2827 16612 2872 16640
rect 2866 16600 2872 16612
rect 2924 16600 2930 16652
rect 3234 16640 3240 16652
rect 3195 16612 3240 16640
rect 3234 16600 3240 16612
rect 3292 16600 3298 16652
rect 4065 16643 4123 16649
rect 4065 16609 4077 16643
rect 4111 16640 4123 16643
rect 4798 16640 4804 16652
rect 4111 16612 4804 16640
rect 4111 16609 4123 16612
rect 4065 16603 4123 16609
rect 4798 16600 4804 16612
rect 4856 16600 4862 16652
rect 8386 16640 8392 16652
rect 8347 16612 8392 16640
rect 8386 16600 8392 16612
rect 8444 16600 8450 16652
rect 8496 16640 8524 16680
rect 9766 16668 9772 16720
rect 9824 16708 9830 16720
rect 10229 16711 10287 16717
rect 10229 16708 10241 16711
rect 9824 16680 10241 16708
rect 9824 16668 9830 16680
rect 10229 16677 10241 16680
rect 10275 16708 10287 16711
rect 10689 16711 10747 16717
rect 10689 16708 10701 16711
rect 10275 16680 10701 16708
rect 10275 16677 10287 16680
rect 10229 16671 10287 16677
rect 10689 16677 10701 16680
rect 10735 16677 10747 16711
rect 12250 16708 12256 16720
rect 12211 16680 12256 16708
rect 10689 16671 10747 16677
rect 12250 16668 12256 16680
rect 12308 16668 12314 16720
rect 13078 16668 13084 16720
rect 13136 16708 13142 16720
rect 13722 16708 13728 16720
rect 13136 16680 13728 16708
rect 13136 16668 13142 16680
rect 13722 16668 13728 16680
rect 13780 16668 13786 16720
rect 13906 16708 13912 16720
rect 13867 16680 13912 16708
rect 13906 16668 13912 16680
rect 13964 16668 13970 16720
rect 14108 16708 14136 16748
rect 14182 16736 14188 16788
rect 14240 16776 14246 16788
rect 14645 16779 14703 16785
rect 14645 16776 14657 16779
rect 14240 16748 14657 16776
rect 14240 16736 14246 16748
rect 14645 16745 14657 16748
rect 14691 16745 14703 16779
rect 14645 16739 14703 16745
rect 18877 16779 18935 16785
rect 18877 16745 18889 16779
rect 18923 16776 18935 16779
rect 19150 16776 19156 16788
rect 18923 16748 19156 16776
rect 18923 16745 18935 16748
rect 18877 16739 18935 16745
rect 19150 16736 19156 16748
rect 19208 16736 19214 16788
rect 19518 16736 19524 16788
rect 19576 16776 19582 16788
rect 19613 16779 19671 16785
rect 19613 16776 19625 16779
rect 19576 16748 19625 16776
rect 19576 16736 19582 16748
rect 19613 16745 19625 16748
rect 19659 16745 19671 16779
rect 19613 16739 19671 16745
rect 21637 16779 21695 16785
rect 21637 16745 21649 16779
rect 21683 16776 21695 16779
rect 21818 16776 21824 16788
rect 21683 16748 21824 16776
rect 21683 16745 21695 16748
rect 21637 16739 21695 16745
rect 21818 16736 21824 16748
rect 21876 16776 21882 16788
rect 21876 16748 22140 16776
rect 21876 16736 21882 16748
rect 15013 16711 15071 16717
rect 15013 16708 15025 16711
rect 14108 16680 15025 16708
rect 15013 16677 15025 16680
rect 15059 16708 15071 16711
rect 15286 16708 15292 16720
rect 15059 16680 15292 16708
rect 15059 16677 15071 16680
rect 15013 16671 15071 16677
rect 15286 16668 15292 16680
rect 15344 16668 15350 16720
rect 15556 16711 15614 16717
rect 15556 16708 15568 16711
rect 15396 16680 15568 16708
rect 8665 16643 8723 16649
rect 8665 16640 8677 16643
rect 8496 16612 8677 16640
rect 8665 16609 8677 16612
rect 8711 16640 8723 16643
rect 9490 16640 9496 16652
rect 8711 16612 9496 16640
rect 8711 16609 8723 16612
rect 8665 16603 8723 16609
rect 9490 16600 9496 16612
rect 9548 16600 9554 16652
rect 10045 16643 10103 16649
rect 10045 16640 10057 16643
rect 9600 16612 10057 16640
rect 9214 16532 9220 16584
rect 9272 16572 9278 16584
rect 9600 16572 9628 16612
rect 10045 16609 10057 16612
rect 10091 16640 10103 16643
rect 10962 16640 10968 16652
rect 10091 16612 10968 16640
rect 10091 16609 10103 16612
rect 10045 16603 10103 16609
rect 10962 16600 10968 16612
rect 11020 16600 11026 16652
rect 14369 16643 14427 16649
rect 14369 16609 14381 16643
rect 14415 16640 14427 16643
rect 14550 16640 14556 16652
rect 14415 16612 14556 16640
rect 14415 16609 14427 16612
rect 14369 16603 14427 16609
rect 14550 16600 14556 16612
rect 14608 16600 14614 16652
rect 15396 16640 15424 16680
rect 15556 16677 15568 16680
rect 15602 16708 15614 16711
rect 15838 16708 15844 16720
rect 15602 16680 15844 16708
rect 15602 16677 15614 16680
rect 15556 16671 15614 16677
rect 15838 16668 15844 16680
rect 15896 16668 15902 16720
rect 18138 16708 18144 16720
rect 18099 16680 18144 16708
rect 18138 16668 18144 16680
rect 18196 16668 18202 16720
rect 18322 16708 18328 16720
rect 18283 16680 18328 16708
rect 18322 16668 18328 16680
rect 18380 16668 18386 16720
rect 19337 16711 19395 16717
rect 19337 16677 19349 16711
rect 19383 16708 19395 16711
rect 19978 16708 19984 16720
rect 19383 16680 19984 16708
rect 19383 16677 19395 16680
rect 19337 16671 19395 16677
rect 19978 16668 19984 16680
rect 20036 16668 20042 16720
rect 16942 16640 16948 16652
rect 15120 16612 15424 16640
rect 16684 16612 16948 16640
rect 9272 16544 9628 16572
rect 9272 16532 9278 16544
rect 10134 16532 10140 16584
rect 10192 16572 10198 16584
rect 10321 16575 10379 16581
rect 10321 16572 10333 16575
rect 10192 16544 10333 16572
rect 10192 16532 10198 16544
rect 10321 16541 10333 16544
rect 10367 16541 10379 16575
rect 10321 16535 10379 16541
rect 12989 16575 13047 16581
rect 12989 16541 13001 16575
rect 13035 16541 13047 16575
rect 12989 16535 13047 16541
rect 9582 16464 9588 16516
rect 9640 16504 9646 16516
rect 9769 16507 9827 16513
rect 9769 16504 9781 16507
rect 9640 16476 9781 16504
rect 9640 16464 9646 16476
rect 9769 16473 9781 16476
rect 9815 16473 9827 16507
rect 9769 16467 9827 16473
rect 11974 16464 11980 16516
rect 12032 16504 12038 16516
rect 13004 16504 13032 16535
rect 13078 16532 13084 16584
rect 13136 16572 13142 16584
rect 13173 16575 13231 16581
rect 13173 16572 13185 16575
rect 13136 16544 13185 16572
rect 13136 16532 13142 16544
rect 13173 16541 13185 16544
rect 13219 16572 13231 16575
rect 13354 16572 13360 16584
rect 13219 16544 13360 16572
rect 13219 16541 13231 16544
rect 13173 16535 13231 16541
rect 13354 16532 13360 16544
rect 13412 16532 13418 16584
rect 13633 16575 13691 16581
rect 13633 16541 13645 16575
rect 13679 16572 13691 16575
rect 14642 16572 14648 16584
rect 13679 16544 14648 16572
rect 13679 16541 13691 16544
rect 13633 16535 13691 16541
rect 14642 16532 14648 16544
rect 14700 16572 14706 16584
rect 15120 16572 15148 16612
rect 15286 16572 15292 16584
rect 14700 16544 15148 16572
rect 15247 16544 15292 16572
rect 14700 16532 14706 16544
rect 15286 16532 15292 16544
rect 15344 16532 15350 16584
rect 12032 16476 13032 16504
rect 12032 16464 12038 16476
rect 6457 16439 6515 16445
rect 6457 16405 6469 16439
rect 6503 16436 6515 16439
rect 6730 16436 6736 16448
rect 6503 16408 6736 16436
rect 6503 16405 6515 16408
rect 6457 16399 6515 16405
rect 6730 16396 6736 16408
rect 6788 16396 6794 16448
rect 7098 16396 7104 16448
rect 7156 16436 7162 16448
rect 7285 16439 7343 16445
rect 7285 16436 7297 16439
rect 7156 16408 7297 16436
rect 7156 16396 7162 16408
rect 7285 16405 7297 16408
rect 7331 16405 7343 16439
rect 8110 16436 8116 16448
rect 8071 16408 8116 16436
rect 7285 16399 7343 16405
rect 8110 16396 8116 16408
rect 8168 16396 8174 16448
rect 11149 16439 11207 16445
rect 11149 16405 11161 16439
rect 11195 16436 11207 16439
rect 11330 16436 11336 16448
rect 11195 16408 11336 16436
rect 11195 16405 11207 16408
rect 11149 16399 11207 16405
rect 11330 16396 11336 16408
rect 11388 16396 11394 16448
rect 15470 16396 15476 16448
rect 15528 16436 15534 16448
rect 16684 16445 16712 16612
rect 16942 16600 16948 16612
rect 17000 16640 17006 16652
rect 17221 16643 17279 16649
rect 17221 16640 17233 16643
rect 17000 16612 17233 16640
rect 17000 16600 17006 16612
rect 17221 16609 17233 16612
rect 17267 16609 17279 16643
rect 18417 16643 18475 16649
rect 18417 16640 18429 16643
rect 17221 16603 17279 16609
rect 17880 16612 18429 16640
rect 17494 16532 17500 16584
rect 17552 16572 17558 16584
rect 17880 16572 17908 16612
rect 18417 16609 18429 16612
rect 18463 16640 18475 16643
rect 18690 16640 18696 16652
rect 18463 16612 18696 16640
rect 18463 16609 18475 16612
rect 18417 16603 18475 16609
rect 18690 16600 18696 16612
rect 18748 16600 18754 16652
rect 22112 16640 22140 16748
rect 22370 16736 22376 16788
rect 22428 16776 22434 16788
rect 23109 16779 23167 16785
rect 23109 16776 23121 16779
rect 22428 16748 23121 16776
rect 22428 16736 22434 16748
rect 23109 16745 23121 16748
rect 23155 16776 23167 16779
rect 23382 16776 23388 16788
rect 23155 16748 23388 16776
rect 23155 16745 23167 16748
rect 23109 16739 23167 16745
rect 23382 16736 23388 16748
rect 23440 16736 23446 16788
rect 23658 16736 23664 16788
rect 23716 16776 23722 16788
rect 24673 16779 24731 16785
rect 24673 16776 24685 16779
rect 23716 16748 24685 16776
rect 23716 16736 23722 16748
rect 24673 16745 24685 16748
rect 24719 16745 24731 16779
rect 24673 16739 24731 16745
rect 22278 16708 22284 16720
rect 22239 16680 22284 16708
rect 22278 16668 22284 16680
rect 22336 16668 22342 16720
rect 22554 16668 22560 16720
rect 22612 16708 22618 16720
rect 22833 16711 22891 16717
rect 22833 16708 22845 16711
rect 22612 16680 22845 16708
rect 22612 16668 22618 16680
rect 22833 16677 22845 16680
rect 22879 16708 22891 16711
rect 23290 16708 23296 16720
rect 22879 16680 23296 16708
rect 22879 16677 22891 16680
rect 22833 16671 22891 16677
rect 23290 16668 23296 16680
rect 23348 16668 23354 16720
rect 23400 16708 23428 16736
rect 23538 16711 23596 16717
rect 23538 16708 23550 16711
rect 23400 16680 23550 16708
rect 23538 16677 23550 16680
rect 23584 16677 23596 16711
rect 23538 16671 23596 16677
rect 22373 16643 22431 16649
rect 22373 16640 22385 16643
rect 22112 16612 22385 16640
rect 22373 16609 22385 16612
rect 22419 16640 22431 16643
rect 22738 16640 22744 16652
rect 22419 16612 22744 16640
rect 22419 16609 22431 16612
rect 22373 16603 22431 16609
rect 22738 16600 22744 16612
rect 22796 16600 22802 16652
rect 24026 16600 24032 16652
rect 24084 16640 24090 16652
rect 25225 16643 25283 16649
rect 25225 16640 25237 16643
rect 24084 16612 25237 16640
rect 24084 16600 24090 16612
rect 25225 16609 25237 16612
rect 25271 16609 25283 16643
rect 25225 16603 25283 16609
rect 17552 16544 17908 16572
rect 22281 16575 22339 16581
rect 17552 16532 17558 16544
rect 22281 16541 22293 16575
rect 22327 16572 22339 16575
rect 22462 16572 22468 16584
rect 22327 16544 22468 16572
rect 22327 16541 22339 16544
rect 22281 16535 22339 16541
rect 22462 16532 22468 16544
rect 22520 16532 22526 16584
rect 23014 16532 23020 16584
rect 23072 16572 23078 16584
rect 23293 16575 23351 16581
rect 23293 16572 23305 16575
rect 23072 16544 23305 16572
rect 23072 16532 23078 16544
rect 23293 16541 23305 16544
rect 23339 16541 23351 16575
rect 23293 16535 23351 16541
rect 16669 16439 16727 16445
rect 16669 16436 16681 16439
rect 15528 16408 16681 16436
rect 15528 16396 15534 16408
rect 16669 16405 16681 16408
rect 16715 16405 16727 16439
rect 17862 16436 17868 16448
rect 17823 16408 17868 16436
rect 16669 16399 16727 16405
rect 17862 16396 17868 16408
rect 17920 16396 17926 16448
rect 21818 16436 21824 16448
rect 21779 16408 21824 16436
rect 21818 16396 21824 16408
rect 21876 16396 21882 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2222 16192 2228 16244
rect 2280 16232 2286 16244
rect 2501 16235 2559 16241
rect 2501 16232 2513 16235
rect 2280 16204 2513 16232
rect 2280 16192 2286 16204
rect 2501 16201 2513 16204
rect 2547 16201 2559 16235
rect 3418 16232 3424 16244
rect 3379 16204 3424 16232
rect 2501 16195 2559 16201
rect 3418 16192 3424 16204
rect 3476 16232 3482 16244
rect 4433 16235 4491 16241
rect 4433 16232 4445 16235
rect 3476 16204 4445 16232
rect 3476 16192 3482 16204
rect 4433 16201 4445 16204
rect 4479 16201 4491 16235
rect 8938 16232 8944 16244
rect 8899 16204 8944 16232
rect 4433 16195 4491 16201
rect 8938 16192 8944 16204
rect 8996 16192 9002 16244
rect 9214 16232 9220 16244
rect 9175 16204 9220 16232
rect 9214 16192 9220 16204
rect 9272 16192 9278 16244
rect 10134 16232 10140 16244
rect 10095 16204 10140 16232
rect 10134 16192 10140 16204
rect 10192 16192 10198 16244
rect 12253 16235 12311 16241
rect 12253 16201 12265 16235
rect 12299 16232 12311 16235
rect 13078 16232 13084 16244
rect 12299 16204 13084 16232
rect 12299 16201 12311 16204
rect 12253 16195 12311 16201
rect 13078 16192 13084 16204
rect 13136 16192 13142 16244
rect 13814 16192 13820 16244
rect 13872 16232 13878 16244
rect 14277 16235 14335 16241
rect 14277 16232 14289 16235
rect 13872 16204 14289 16232
rect 13872 16192 13878 16204
rect 14277 16201 14289 16204
rect 14323 16201 14335 16235
rect 14642 16232 14648 16244
rect 14603 16204 14648 16232
rect 14277 16195 14335 16201
rect 14642 16192 14648 16204
rect 14700 16192 14706 16244
rect 14734 16192 14740 16244
rect 14792 16232 14798 16244
rect 14921 16235 14979 16241
rect 14921 16232 14933 16235
rect 14792 16204 14933 16232
rect 14792 16192 14798 16204
rect 14921 16201 14933 16204
rect 14967 16201 14979 16235
rect 14921 16195 14979 16201
rect 15286 16192 15292 16244
rect 15344 16232 15350 16244
rect 15838 16232 15844 16244
rect 15344 16204 15844 16232
rect 15344 16192 15350 16204
rect 15838 16192 15844 16204
rect 15896 16192 15902 16244
rect 16206 16192 16212 16244
rect 16264 16232 16270 16244
rect 16485 16235 16543 16241
rect 16485 16232 16497 16235
rect 16264 16204 16497 16232
rect 16264 16192 16270 16204
rect 16485 16201 16497 16204
rect 16531 16201 16543 16235
rect 17494 16232 17500 16244
rect 17455 16204 17500 16232
rect 16485 16195 16543 16201
rect 17494 16192 17500 16204
rect 17552 16192 17558 16244
rect 17865 16235 17923 16241
rect 17865 16201 17877 16235
rect 17911 16232 17923 16235
rect 18138 16232 18144 16244
rect 17911 16204 18144 16232
rect 17911 16201 17923 16204
rect 17865 16195 17923 16201
rect 18138 16192 18144 16204
rect 18196 16192 18202 16244
rect 18322 16232 18328 16244
rect 18283 16204 18328 16232
rect 18322 16192 18328 16204
rect 18380 16192 18386 16244
rect 23014 16192 23020 16244
rect 23072 16232 23078 16244
rect 23293 16235 23351 16241
rect 23293 16232 23305 16235
rect 23072 16204 23305 16232
rect 23072 16192 23078 16204
rect 23293 16201 23305 16204
rect 23339 16201 23351 16235
rect 23293 16195 23351 16201
rect 23845 16235 23903 16241
rect 23845 16201 23857 16235
rect 23891 16232 23903 16235
rect 24026 16232 24032 16244
rect 23891 16204 24032 16232
rect 23891 16201 23903 16204
rect 23845 16195 23903 16201
rect 24026 16192 24032 16204
rect 24084 16192 24090 16244
rect 2317 16167 2375 16173
rect 2317 16133 2329 16167
rect 2363 16164 2375 16167
rect 4246 16164 4252 16176
rect 2363 16136 4252 16164
rect 2363 16133 2375 16136
rect 2317 16127 2375 16133
rect 2976 16105 3004 16136
rect 4246 16124 4252 16136
rect 4304 16124 4310 16176
rect 4614 16124 4620 16176
rect 4672 16164 4678 16176
rect 5261 16167 5319 16173
rect 5261 16164 5273 16167
rect 4672 16136 5273 16164
rect 4672 16124 4678 16136
rect 5261 16133 5273 16136
rect 5307 16133 5319 16167
rect 5261 16127 5319 16133
rect 6641 16167 6699 16173
rect 6641 16133 6653 16167
rect 6687 16164 6699 16167
rect 7374 16164 7380 16176
rect 6687 16136 7380 16164
rect 6687 16133 6699 16136
rect 6641 16127 6699 16133
rect 7374 16124 7380 16136
rect 7432 16124 7438 16176
rect 10873 16167 10931 16173
rect 10873 16133 10885 16167
rect 10919 16164 10931 16167
rect 11974 16164 11980 16176
rect 10919 16136 11980 16164
rect 10919 16133 10931 16136
rect 10873 16127 10931 16133
rect 11974 16124 11980 16136
rect 12032 16124 12038 16176
rect 13357 16167 13415 16173
rect 13357 16133 13369 16167
rect 13403 16133 13415 16167
rect 18874 16164 18880 16176
rect 18835 16136 18880 16164
rect 13357 16127 13415 16133
rect 2961 16099 3019 16105
rect 2961 16065 2973 16099
rect 3007 16065 3019 16099
rect 2961 16059 3019 16065
rect 3050 16056 3056 16108
rect 3108 16096 3114 16108
rect 5721 16099 5779 16105
rect 3108 16068 3153 16096
rect 3108 16056 3114 16068
rect 5721 16065 5733 16099
rect 5767 16096 5779 16099
rect 6730 16096 6736 16108
rect 5767 16068 6736 16096
rect 5767 16065 5779 16068
rect 5721 16059 5779 16065
rect 6730 16056 6736 16068
rect 6788 16056 6794 16108
rect 7193 16099 7251 16105
rect 7193 16065 7205 16099
rect 7239 16096 7251 16099
rect 7837 16099 7895 16105
rect 7837 16096 7849 16099
rect 7239 16068 7849 16096
rect 7239 16065 7251 16068
rect 7193 16059 7251 16065
rect 7837 16065 7849 16068
rect 7883 16096 7895 16099
rect 9398 16096 9404 16108
rect 7883 16068 9404 16096
rect 7883 16065 7895 16068
rect 7837 16059 7895 16065
rect 9398 16056 9404 16068
rect 9456 16056 9462 16108
rect 9582 16096 9588 16108
rect 9543 16068 9588 16096
rect 9582 16056 9588 16068
rect 9640 16056 9646 16108
rect 9769 16099 9827 16105
rect 9769 16065 9781 16099
rect 9815 16096 9827 16099
rect 9858 16096 9864 16108
rect 9815 16068 9864 16096
rect 9815 16065 9827 16068
rect 9769 16059 9827 16065
rect 9858 16056 9864 16068
rect 9916 16056 9922 16108
rect 10689 16099 10747 16105
rect 10689 16065 10701 16099
rect 10735 16096 10747 16099
rect 11425 16099 11483 16105
rect 11425 16096 11437 16099
rect 10735 16068 11437 16096
rect 10735 16065 10747 16068
rect 10689 16059 10747 16065
rect 11425 16065 11437 16068
rect 11471 16096 11483 16099
rect 12342 16096 12348 16108
rect 11471 16068 12348 16096
rect 11471 16065 11483 16068
rect 11425 16059 11483 16065
rect 12342 16056 12348 16068
rect 12400 16056 12406 16108
rect 13372 16096 13400 16127
rect 18874 16124 18880 16136
rect 18932 16124 18938 16176
rect 14826 16096 14832 16108
rect 13372 16068 14832 16096
rect 14826 16056 14832 16068
rect 14884 16096 14890 16108
rect 15289 16099 15347 16105
rect 15289 16096 15301 16099
rect 14884 16068 15301 16096
rect 14884 16056 14890 16068
rect 15289 16065 15301 16068
rect 15335 16065 15347 16099
rect 15289 16059 15347 16065
rect 16301 16099 16359 16105
rect 16301 16065 16313 16099
rect 16347 16096 16359 16099
rect 16942 16096 16948 16108
rect 16347 16068 16948 16096
rect 16347 16065 16359 16068
rect 16301 16059 16359 16065
rect 16942 16056 16948 16068
rect 17000 16056 17006 16108
rect 23566 16056 23572 16108
rect 23624 16096 23630 16108
rect 24397 16099 24455 16105
rect 24397 16096 24409 16099
rect 23624 16068 24409 16096
rect 23624 16056 23630 16068
rect 24397 16065 24409 16068
rect 24443 16096 24455 16099
rect 24765 16099 24823 16105
rect 24765 16096 24777 16099
rect 24443 16068 24777 16096
rect 24443 16065 24455 16068
rect 24397 16059 24455 16065
rect 24765 16065 24777 16068
rect 24811 16096 24823 16099
rect 24854 16096 24860 16108
rect 24811 16068 24860 16096
rect 24811 16065 24823 16068
rect 24765 16059 24823 16065
rect 24854 16056 24860 16068
rect 24912 16056 24918 16108
rect 1949 16031 2007 16037
rect 1949 15997 1961 16031
rect 1995 16028 2007 16031
rect 3326 16028 3332 16040
rect 1995 16000 3332 16028
rect 1995 15997 2007 16000
rect 1949 15991 2007 15997
rect 3326 15988 3332 16000
rect 3384 15988 3390 16040
rect 5077 16031 5135 16037
rect 5077 15997 5089 16031
rect 5123 16028 5135 16031
rect 5813 16031 5871 16037
rect 5813 16028 5825 16031
rect 5123 16000 5825 16028
rect 5123 15997 5135 16000
rect 5077 15991 5135 15997
rect 5813 15997 5825 16000
rect 5859 16028 5871 16031
rect 6638 16028 6644 16040
rect 5859 16000 6644 16028
rect 5859 15997 5871 16000
rect 5813 15991 5871 15997
rect 6638 15988 6644 16000
rect 6696 15988 6702 16040
rect 13170 16028 13176 16040
rect 13083 16000 13176 16028
rect 13170 15988 13176 16000
rect 13228 16028 13234 16040
rect 13909 16031 13967 16037
rect 13228 16000 13860 16028
rect 13228 15988 13234 16000
rect 13832 15972 13860 16000
rect 13909 15997 13921 16031
rect 13955 16028 13967 16031
rect 14642 16028 14648 16040
rect 13955 16000 14648 16028
rect 13955 15997 13967 16000
rect 13909 15991 13967 15997
rect 14642 15988 14648 16000
rect 14700 15988 14706 16040
rect 19150 16028 19156 16040
rect 19111 16000 19156 16028
rect 19150 15988 19156 16000
rect 19208 15988 19214 16040
rect 20809 16031 20867 16037
rect 20809 15997 20821 16031
rect 20855 16028 20867 16031
rect 20898 16028 20904 16040
rect 20855 16000 20904 16028
rect 20855 15997 20867 16000
rect 20809 15991 20867 15997
rect 20898 15988 20904 16000
rect 20956 16028 20962 16040
rect 23014 16028 23020 16040
rect 20956 16000 23020 16028
rect 20956 15988 20962 16000
rect 23014 15988 23020 16000
rect 23072 15988 23078 16040
rect 24121 16031 24179 16037
rect 24121 15997 24133 16031
rect 24167 16028 24179 16031
rect 24210 16028 24216 16040
rect 24167 16000 24216 16028
rect 24167 15997 24179 16000
rect 24121 15991 24179 15997
rect 7929 15963 7987 15969
rect 7929 15929 7941 15963
rect 7975 15960 7987 15963
rect 8018 15960 8024 15972
rect 7975 15932 8024 15960
rect 7975 15929 7987 15932
rect 7929 15923 7987 15929
rect 8018 15920 8024 15932
rect 8076 15920 8082 15972
rect 8938 15920 8944 15972
rect 8996 15960 9002 15972
rect 9677 15963 9735 15969
rect 9677 15960 9689 15963
rect 8996 15932 9689 15960
rect 8996 15920 9002 15932
rect 9677 15929 9689 15932
rect 9723 15960 9735 15963
rect 10778 15960 10784 15972
rect 9723 15932 10784 15960
rect 9723 15929 9735 15932
rect 9677 15923 9735 15929
rect 10778 15920 10784 15932
rect 10836 15920 10842 15972
rect 11149 15963 11207 15969
rect 11149 15929 11161 15963
rect 11195 15960 11207 15963
rect 12805 15963 12863 15969
rect 11195 15932 11928 15960
rect 11195 15929 11207 15932
rect 11149 15923 11207 15929
rect 1394 15892 1400 15904
rect 1355 15864 1400 15892
rect 1394 15852 1400 15864
rect 1452 15852 1458 15904
rect 2961 15895 3019 15901
rect 2961 15861 2973 15895
rect 3007 15892 3019 15895
rect 3326 15892 3332 15904
rect 3007 15864 3332 15892
rect 3007 15861 3019 15864
rect 2961 15855 3019 15861
rect 3326 15852 3332 15864
rect 3384 15852 3390 15904
rect 4157 15895 4215 15901
rect 4157 15861 4169 15895
rect 4203 15892 4215 15895
rect 4798 15892 4804 15904
rect 4203 15864 4804 15892
rect 4203 15861 4215 15864
rect 4157 15855 4215 15861
rect 4798 15852 4804 15864
rect 4856 15852 4862 15904
rect 5721 15895 5779 15901
rect 5721 15861 5733 15895
rect 5767 15892 5779 15895
rect 6273 15895 6331 15901
rect 6273 15892 6285 15895
rect 5767 15864 6285 15892
rect 5767 15861 5779 15864
rect 5721 15855 5779 15861
rect 6273 15861 6285 15864
rect 6319 15892 6331 15895
rect 6822 15892 6828 15904
rect 6319 15864 6828 15892
rect 6319 15861 6331 15864
rect 6273 15855 6331 15861
rect 6822 15852 6828 15864
rect 6880 15852 6886 15904
rect 7006 15852 7012 15904
rect 7064 15892 7070 15904
rect 7837 15895 7895 15901
rect 7837 15892 7849 15895
rect 7064 15864 7849 15892
rect 7064 15852 7070 15864
rect 7837 15861 7849 15864
rect 7883 15892 7895 15895
rect 8202 15892 8208 15904
rect 7883 15864 8208 15892
rect 7883 15861 7895 15864
rect 7837 15855 7895 15861
rect 8202 15852 8208 15864
rect 8260 15852 8266 15904
rect 8386 15892 8392 15904
rect 8347 15864 8392 15892
rect 8386 15852 8392 15864
rect 8444 15852 8450 15904
rect 11330 15892 11336 15904
rect 11291 15864 11336 15892
rect 11330 15852 11336 15864
rect 11388 15852 11394 15904
rect 11900 15901 11928 15932
rect 12805 15929 12817 15963
rect 12851 15960 12863 15963
rect 13630 15960 13636 15972
rect 12851 15932 13636 15960
rect 12851 15929 12863 15932
rect 12805 15923 12863 15929
rect 13630 15920 13636 15932
rect 13688 15920 13694 15972
rect 13814 15960 13820 15972
rect 13775 15932 13820 15960
rect 13814 15920 13820 15932
rect 13872 15920 13878 15972
rect 15470 15960 15476 15972
rect 15431 15932 15476 15960
rect 15470 15920 15476 15932
rect 15528 15920 15534 15972
rect 15654 15920 15660 15972
rect 15712 15960 15718 15972
rect 17034 15960 17040 15972
rect 15712 15932 17040 15960
rect 15712 15920 15718 15932
rect 17034 15920 17040 15932
rect 17092 15920 17098 15972
rect 18138 15920 18144 15972
rect 18196 15960 18202 15972
rect 19429 15963 19487 15969
rect 19429 15960 19441 15963
rect 18196 15932 19441 15960
rect 18196 15920 18202 15932
rect 19429 15929 19441 15932
rect 19475 15960 19487 15963
rect 19797 15963 19855 15969
rect 19797 15960 19809 15963
rect 19475 15932 19809 15960
rect 19475 15929 19487 15932
rect 19429 15923 19487 15929
rect 19797 15929 19809 15932
rect 19843 15960 19855 15963
rect 19978 15960 19984 15972
rect 19843 15932 19984 15960
rect 19843 15929 19855 15932
rect 19797 15923 19855 15929
rect 19978 15920 19984 15932
rect 20036 15920 20042 15972
rect 21082 15969 21088 15972
rect 20349 15963 20407 15969
rect 20349 15929 20361 15963
rect 20395 15960 20407 15963
rect 21076 15960 21088 15969
rect 20395 15932 21088 15960
rect 20395 15929 20407 15932
rect 20349 15923 20407 15929
rect 21076 15923 21088 15932
rect 21082 15920 21088 15923
rect 21140 15920 21146 15972
rect 22278 15920 22284 15972
rect 22336 15960 22342 15972
rect 22925 15963 22983 15969
rect 22925 15960 22937 15963
rect 22336 15932 22937 15960
rect 22336 15920 22342 15932
rect 22925 15929 22937 15932
rect 22971 15960 22983 15963
rect 24136 15960 24164 15991
rect 24210 15988 24216 16000
rect 24268 15988 24274 16040
rect 24670 15988 24676 16040
rect 24728 16028 24734 16040
rect 25317 16031 25375 16037
rect 25317 16028 25329 16031
rect 24728 16000 25329 16028
rect 24728 15988 24734 16000
rect 25317 15997 25329 16000
rect 25363 16028 25375 16031
rect 25869 16031 25927 16037
rect 25869 16028 25881 16031
rect 25363 16000 25881 16028
rect 25363 15997 25375 16000
rect 25317 15991 25375 15997
rect 25869 15997 25881 16000
rect 25915 15997 25927 16031
rect 25869 15991 25927 15997
rect 22971 15932 24164 15960
rect 22971 15929 22983 15932
rect 22925 15923 22983 15929
rect 11885 15895 11943 15901
rect 11885 15861 11897 15895
rect 11931 15892 11943 15895
rect 12342 15892 12348 15904
rect 11931 15864 12348 15892
rect 11931 15861 11943 15864
rect 11885 15855 11943 15861
rect 12342 15852 12348 15864
rect 12400 15852 12406 15904
rect 15381 15895 15439 15901
rect 15381 15861 15393 15895
rect 15427 15892 15439 15895
rect 15562 15892 15568 15904
rect 15427 15864 15568 15892
rect 15427 15861 15439 15864
rect 15381 15855 15439 15861
rect 15562 15852 15568 15864
rect 15620 15852 15626 15904
rect 15838 15892 15844 15904
rect 15799 15864 15844 15892
rect 15838 15852 15844 15864
rect 15896 15852 15902 15904
rect 16390 15852 16396 15904
rect 16448 15892 16454 15904
rect 16945 15895 17003 15901
rect 16945 15892 16957 15895
rect 16448 15864 16957 15892
rect 16448 15852 16454 15864
rect 16945 15861 16957 15864
rect 16991 15861 17003 15895
rect 18598 15892 18604 15904
rect 18559 15864 18604 15892
rect 16945 15855 17003 15861
rect 18598 15852 18604 15864
rect 18656 15892 18662 15904
rect 19337 15895 19395 15901
rect 19337 15892 19349 15895
rect 18656 15864 19349 15892
rect 18656 15852 18662 15864
rect 19337 15861 19349 15864
rect 19383 15861 19395 15895
rect 19337 15855 19395 15861
rect 20717 15895 20775 15901
rect 20717 15861 20729 15895
rect 20763 15892 20775 15895
rect 20898 15892 20904 15904
rect 20763 15864 20904 15892
rect 20763 15861 20775 15864
rect 20717 15855 20775 15861
rect 20898 15852 20904 15864
rect 20956 15852 20962 15904
rect 21910 15852 21916 15904
rect 21968 15892 21974 15904
rect 22189 15895 22247 15901
rect 22189 15892 22201 15895
rect 21968 15864 22201 15892
rect 21968 15852 21974 15864
rect 22189 15861 22201 15864
rect 22235 15861 22247 15895
rect 22189 15855 22247 15861
rect 23474 15852 23480 15904
rect 23532 15892 23538 15904
rect 24305 15895 24363 15901
rect 24305 15892 24317 15895
rect 23532 15864 24317 15892
rect 23532 15852 23538 15864
rect 24305 15861 24317 15864
rect 24351 15861 24363 15895
rect 24305 15855 24363 15861
rect 25501 15895 25559 15901
rect 25501 15861 25513 15895
rect 25547 15892 25559 15895
rect 25682 15892 25688 15904
rect 25547 15864 25688 15892
rect 25547 15861 25559 15864
rect 25501 15855 25559 15861
rect 25682 15852 25688 15864
rect 25740 15852 25746 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 2774 15648 2780 15700
rect 2832 15688 2838 15700
rect 2869 15691 2927 15697
rect 2869 15688 2881 15691
rect 2832 15660 2881 15688
rect 2832 15648 2838 15660
rect 2869 15657 2881 15660
rect 2915 15657 2927 15691
rect 6638 15688 6644 15700
rect 6599 15660 6644 15688
rect 2869 15651 2927 15657
rect 6638 15648 6644 15660
rect 6696 15648 6702 15700
rect 7006 15648 7012 15700
rect 7064 15688 7070 15700
rect 7285 15691 7343 15697
rect 7285 15688 7297 15691
rect 7064 15660 7297 15688
rect 7064 15648 7070 15660
rect 7285 15657 7297 15660
rect 7331 15657 7343 15691
rect 8294 15688 8300 15700
rect 8255 15660 8300 15688
rect 7285 15651 7343 15657
rect 8294 15648 8300 15660
rect 8352 15648 8358 15700
rect 8754 15688 8760 15700
rect 8715 15660 8760 15688
rect 8754 15648 8760 15660
rect 8812 15648 8818 15700
rect 9217 15691 9275 15697
rect 9217 15657 9229 15691
rect 9263 15688 9275 15691
rect 9582 15688 9588 15700
rect 9263 15660 9588 15688
rect 9263 15657 9275 15660
rect 9217 15651 9275 15657
rect 9582 15648 9588 15660
rect 9640 15648 9646 15700
rect 10962 15648 10968 15700
rect 11020 15688 11026 15700
rect 11057 15691 11115 15697
rect 11057 15688 11069 15691
rect 11020 15660 11069 15688
rect 11020 15648 11026 15660
rect 11057 15657 11069 15660
rect 11103 15657 11115 15691
rect 11974 15688 11980 15700
rect 11935 15660 11980 15688
rect 11057 15651 11115 15657
rect 11974 15648 11980 15660
rect 12032 15648 12038 15700
rect 13538 15648 13544 15700
rect 13596 15688 13602 15700
rect 13817 15691 13875 15697
rect 13817 15688 13829 15691
rect 13596 15660 13829 15688
rect 13596 15648 13602 15660
rect 13817 15657 13829 15660
rect 13863 15657 13875 15691
rect 13817 15651 13875 15657
rect 14553 15691 14611 15697
rect 14553 15657 14565 15691
rect 14599 15688 14611 15691
rect 15562 15688 15568 15700
rect 14599 15660 15568 15688
rect 14599 15657 14611 15660
rect 14553 15651 14611 15657
rect 15562 15648 15568 15660
rect 15620 15648 15626 15700
rect 15746 15688 15752 15700
rect 15707 15660 15752 15688
rect 15746 15648 15752 15660
rect 15804 15648 15810 15700
rect 16850 15648 16856 15700
rect 16908 15688 16914 15700
rect 17313 15691 17371 15697
rect 17313 15688 17325 15691
rect 16908 15660 17325 15688
rect 16908 15648 16914 15660
rect 17313 15657 17325 15660
rect 17359 15688 17371 15691
rect 17402 15688 17408 15700
rect 17359 15660 17408 15688
rect 17359 15657 17371 15660
rect 17313 15651 17371 15657
rect 17402 15648 17408 15660
rect 17460 15648 17466 15700
rect 19521 15691 19579 15697
rect 19521 15688 19533 15691
rect 18892 15660 19533 15688
rect 18892 15632 18920 15660
rect 19521 15657 19533 15660
rect 19567 15657 19579 15691
rect 19521 15651 19579 15657
rect 21266 15648 21272 15700
rect 21324 15688 21330 15700
rect 21453 15691 21511 15697
rect 21453 15688 21465 15691
rect 21324 15660 21465 15688
rect 21324 15648 21330 15660
rect 21453 15657 21465 15660
rect 21499 15657 21511 15691
rect 21453 15651 21511 15657
rect 22005 15691 22063 15697
rect 22005 15657 22017 15691
rect 22051 15688 22063 15691
rect 22278 15688 22284 15700
rect 22051 15660 22284 15688
rect 22051 15657 22063 15660
rect 22005 15651 22063 15657
rect 22278 15648 22284 15660
rect 22336 15648 22342 15700
rect 22373 15691 22431 15697
rect 22373 15657 22385 15691
rect 22419 15688 22431 15691
rect 22462 15688 22468 15700
rect 22419 15660 22468 15688
rect 22419 15657 22431 15660
rect 22373 15651 22431 15657
rect 22462 15648 22468 15660
rect 22520 15648 22526 15700
rect 23474 15648 23480 15700
rect 23532 15688 23538 15700
rect 23753 15691 23811 15697
rect 23753 15688 23765 15691
rect 23532 15660 23765 15688
rect 23532 15648 23538 15660
rect 23753 15657 23765 15660
rect 23799 15657 23811 15691
rect 23753 15651 23811 15657
rect 4709 15623 4767 15629
rect 4709 15589 4721 15623
rect 4755 15620 4767 15623
rect 4798 15620 4804 15632
rect 4755 15592 4804 15620
rect 4755 15589 4767 15592
rect 4709 15583 4767 15589
rect 4798 15580 4804 15592
rect 4856 15620 4862 15632
rect 6086 15620 6092 15632
rect 4856 15592 6092 15620
rect 4856 15580 4862 15592
rect 1489 15555 1547 15561
rect 1489 15521 1501 15555
rect 1535 15552 1547 15555
rect 1578 15552 1584 15564
rect 1535 15524 1584 15552
rect 1535 15521 1547 15524
rect 1489 15515 1547 15521
rect 1578 15512 1584 15524
rect 1636 15512 1642 15564
rect 1756 15555 1814 15561
rect 1756 15521 1768 15555
rect 1802 15552 1814 15555
rect 2866 15552 2872 15564
rect 1802 15524 2872 15552
rect 1802 15521 1814 15524
rect 1756 15515 1814 15521
rect 2866 15512 2872 15524
rect 2924 15512 2930 15564
rect 4062 15552 4068 15564
rect 4023 15524 4068 15552
rect 4062 15512 4068 15524
rect 4120 15512 4126 15564
rect 5276 15561 5304 15592
rect 6086 15580 6092 15592
rect 6144 15580 6150 15632
rect 9950 15580 9956 15632
rect 10008 15620 10014 15632
rect 10229 15623 10287 15629
rect 10229 15620 10241 15623
rect 10008 15592 10241 15620
rect 10008 15580 10014 15592
rect 10229 15589 10241 15592
rect 10275 15589 10287 15623
rect 10229 15583 10287 15589
rect 13906 15580 13912 15632
rect 13964 15620 13970 15632
rect 14829 15623 14887 15629
rect 14829 15620 14841 15623
rect 13964 15592 14841 15620
rect 13964 15580 13970 15592
rect 14829 15589 14841 15592
rect 14875 15620 14887 15623
rect 15470 15620 15476 15632
rect 14875 15592 15476 15620
rect 14875 15589 14887 15592
rect 14829 15583 14887 15589
rect 15470 15580 15476 15592
rect 15528 15580 15534 15632
rect 15654 15620 15660 15632
rect 15615 15592 15660 15620
rect 15654 15580 15660 15592
rect 15712 15580 15718 15632
rect 18874 15620 18880 15632
rect 18835 15592 18880 15620
rect 18874 15580 18880 15592
rect 18932 15580 18938 15632
rect 19061 15623 19119 15629
rect 19061 15620 19073 15623
rect 18984 15592 19073 15620
rect 5534 15561 5540 15564
rect 5261 15555 5319 15561
rect 5261 15521 5273 15555
rect 5307 15521 5319 15555
rect 5261 15515 5319 15521
rect 5528 15515 5540 15561
rect 5592 15552 5598 15564
rect 5592 15524 5628 15552
rect 5534 15512 5540 15515
rect 5592 15512 5598 15524
rect 7098 15512 7104 15564
rect 7156 15552 7162 15564
rect 8018 15552 8024 15564
rect 7156 15524 8024 15552
rect 7156 15512 7162 15524
rect 8018 15512 8024 15524
rect 8076 15552 8082 15564
rect 8389 15555 8447 15561
rect 8389 15552 8401 15555
rect 8076 15524 8401 15552
rect 8076 15512 8082 15524
rect 8389 15521 8401 15524
rect 8435 15521 8447 15555
rect 8389 15515 8447 15521
rect 9674 15512 9680 15564
rect 9732 15552 9738 15564
rect 10045 15555 10103 15561
rect 10045 15552 10057 15555
rect 9732 15524 10057 15552
rect 9732 15512 9738 15524
rect 10045 15521 10057 15524
rect 10091 15521 10103 15555
rect 10045 15515 10103 15521
rect 12158 15512 12164 15564
rect 12216 15552 12222 15564
rect 12345 15555 12403 15561
rect 12345 15552 12357 15555
rect 12216 15524 12357 15552
rect 12216 15512 12222 15524
rect 12345 15521 12357 15524
rect 12391 15552 12403 15555
rect 12704 15555 12762 15561
rect 12704 15552 12716 15555
rect 12391 15524 12716 15552
rect 12391 15521 12403 15524
rect 12345 15515 12403 15521
rect 12704 15521 12716 15524
rect 12750 15552 12762 15555
rect 12986 15552 12992 15564
rect 12750 15524 12992 15552
rect 12750 15521 12762 15524
rect 12704 15515 12762 15521
rect 12986 15512 12992 15524
rect 13044 15512 13050 15564
rect 15378 15512 15384 15564
rect 15436 15552 15442 15564
rect 16390 15552 16396 15564
rect 15436 15524 16396 15552
rect 15436 15512 15442 15524
rect 16390 15512 16396 15524
rect 16448 15512 16454 15564
rect 16666 15552 16672 15564
rect 16500 15524 16672 15552
rect 8202 15484 8208 15496
rect 8163 15456 8208 15484
rect 8202 15444 8208 15456
rect 8260 15444 8266 15496
rect 9398 15444 9404 15496
rect 9456 15484 9462 15496
rect 9858 15484 9864 15496
rect 9456 15456 9864 15484
rect 9456 15444 9462 15456
rect 9858 15444 9864 15456
rect 9916 15484 9922 15496
rect 10321 15487 10379 15493
rect 10321 15484 10333 15487
rect 9916 15456 10333 15484
rect 9916 15444 9922 15456
rect 10321 15453 10333 15456
rect 10367 15453 10379 15487
rect 10321 15447 10379 15453
rect 11698 15444 11704 15496
rect 11756 15484 11762 15496
rect 12434 15484 12440 15496
rect 11756 15456 12440 15484
rect 11756 15444 11762 15456
rect 12434 15444 12440 15456
rect 12492 15444 12498 15496
rect 14550 15444 14556 15496
rect 14608 15484 14614 15496
rect 16500 15484 16528 15524
rect 16666 15512 16672 15524
rect 16724 15552 16730 15564
rect 17129 15555 17187 15561
rect 17129 15552 17141 15555
rect 16724 15524 17141 15552
rect 16724 15512 16730 15524
rect 17129 15521 17141 15524
rect 17175 15521 17187 15555
rect 17129 15515 17187 15521
rect 14608 15456 16528 15484
rect 14608 15444 14614 15456
rect 16574 15444 16580 15496
rect 16632 15484 16638 15496
rect 17405 15487 17463 15493
rect 17405 15484 17417 15487
rect 16632 15456 17417 15484
rect 16632 15444 16638 15456
rect 17405 15453 17417 15456
rect 17451 15484 17463 15487
rect 18049 15487 18107 15493
rect 18049 15484 18061 15487
rect 17451 15456 18061 15484
rect 17451 15453 17463 15456
rect 17405 15447 17463 15453
rect 18049 15453 18061 15456
rect 18095 15484 18107 15487
rect 18138 15484 18144 15496
rect 18095 15456 18144 15484
rect 18095 15453 18107 15456
rect 18049 15447 18107 15453
rect 18138 15444 18144 15456
rect 18196 15444 18202 15496
rect 2498 15376 2504 15428
rect 2556 15416 2562 15428
rect 3881 15419 3939 15425
rect 3881 15416 3893 15419
rect 2556 15388 3893 15416
rect 2556 15376 2562 15388
rect 3881 15385 3893 15388
rect 3927 15385 3939 15419
rect 9766 15416 9772 15428
rect 9727 15388 9772 15416
rect 3881 15379 3939 15385
rect 9766 15376 9772 15388
rect 9824 15376 9830 15428
rect 16853 15419 16911 15425
rect 16853 15385 16865 15419
rect 16899 15416 16911 15419
rect 18874 15416 18880 15428
rect 16899 15388 18880 15416
rect 16899 15385 16911 15388
rect 16853 15379 16911 15385
rect 18874 15376 18880 15388
rect 18932 15416 18938 15428
rect 18984 15416 19012 15592
rect 19061 15589 19073 15592
rect 19107 15589 19119 15623
rect 19061 15583 19119 15589
rect 22646 15580 22652 15632
rect 22704 15620 22710 15632
rect 22833 15623 22891 15629
rect 22833 15620 22845 15623
rect 22704 15592 22845 15620
rect 22704 15580 22710 15592
rect 22833 15589 22845 15592
rect 22879 15589 22891 15623
rect 23014 15620 23020 15632
rect 22975 15592 23020 15620
rect 22833 15583 22891 15589
rect 23014 15580 23020 15592
rect 23072 15620 23078 15632
rect 23198 15620 23204 15632
rect 23072 15592 23204 15620
rect 23072 15580 23078 15592
rect 23198 15580 23204 15592
rect 23256 15580 23262 15632
rect 24394 15620 24400 15632
rect 24355 15592 24400 15620
rect 24394 15580 24400 15592
rect 24452 15580 24458 15632
rect 24581 15623 24639 15629
rect 24581 15589 24593 15623
rect 24627 15620 24639 15623
rect 25130 15620 25136 15632
rect 24627 15592 25136 15620
rect 24627 15589 24639 15592
rect 24581 15583 24639 15589
rect 20806 15512 20812 15564
rect 20864 15552 20870 15564
rect 21269 15555 21327 15561
rect 21269 15552 21281 15555
rect 20864 15524 21281 15552
rect 20864 15512 20870 15524
rect 21269 15521 21281 15524
rect 21315 15552 21327 15555
rect 22002 15552 22008 15564
rect 21315 15524 22008 15552
rect 21315 15521 21327 15524
rect 21269 15515 21327 15521
rect 22002 15512 22008 15524
rect 22060 15512 22066 15564
rect 23109 15555 23167 15561
rect 23109 15552 23121 15555
rect 22572 15524 23121 15552
rect 19150 15484 19156 15496
rect 19111 15456 19156 15484
rect 19150 15444 19156 15456
rect 19208 15444 19214 15496
rect 19978 15444 19984 15496
rect 20036 15484 20042 15496
rect 21545 15487 21603 15493
rect 21545 15484 21557 15487
rect 20036 15456 21557 15484
rect 20036 15444 20042 15456
rect 21545 15453 21557 15456
rect 21591 15484 21603 15487
rect 21910 15484 21916 15496
rect 21591 15456 21916 15484
rect 21591 15453 21603 15456
rect 21545 15447 21603 15453
rect 21910 15444 21916 15456
rect 21968 15484 21974 15496
rect 22572 15484 22600 15524
rect 23109 15521 23121 15524
rect 23155 15521 23167 15555
rect 23109 15515 23167 15521
rect 23474 15512 23480 15564
rect 23532 15552 23538 15564
rect 24596 15552 24624 15583
rect 25130 15580 25136 15592
rect 25188 15580 25194 15632
rect 23532 15524 24624 15552
rect 24673 15555 24731 15561
rect 23532 15512 23538 15524
rect 24673 15521 24685 15555
rect 24719 15552 24731 15555
rect 24854 15552 24860 15564
rect 24719 15524 24860 15552
rect 24719 15521 24731 15524
rect 24673 15515 24731 15521
rect 24854 15512 24860 15524
rect 24912 15552 24918 15564
rect 25041 15555 25099 15561
rect 25041 15552 25053 15555
rect 24912 15524 25053 15552
rect 24912 15512 24918 15524
rect 25041 15521 25053 15524
rect 25087 15521 25099 15555
rect 25041 15515 25099 15521
rect 21968 15456 22600 15484
rect 21968 15444 21974 15456
rect 18932 15388 19012 15416
rect 20257 15419 20315 15425
rect 18932 15376 18938 15388
rect 20257 15385 20269 15419
rect 20303 15416 20315 15419
rect 20990 15416 20996 15428
rect 20303 15388 20996 15416
rect 20303 15385 20315 15388
rect 20257 15379 20315 15385
rect 20990 15376 20996 15388
rect 21048 15376 21054 15428
rect 2590 15308 2596 15360
rect 2648 15348 2654 15360
rect 3421 15351 3479 15357
rect 3421 15348 3433 15351
rect 2648 15320 3433 15348
rect 2648 15308 2654 15320
rect 3421 15317 3433 15320
rect 3467 15317 3479 15351
rect 3421 15311 3479 15317
rect 3786 15308 3792 15360
rect 3844 15348 3850 15360
rect 4249 15351 4307 15357
rect 4249 15348 4261 15351
rect 3844 15320 4261 15348
rect 3844 15308 3850 15320
rect 4249 15317 4261 15320
rect 4295 15317 4307 15351
rect 5074 15348 5080 15360
rect 5035 15320 5080 15348
rect 4249 15311 4307 15317
rect 5074 15308 5080 15320
rect 5132 15308 5138 15360
rect 7834 15348 7840 15360
rect 7795 15320 7840 15348
rect 7834 15308 7840 15320
rect 7892 15308 7898 15360
rect 10686 15348 10692 15360
rect 10647 15320 10692 15348
rect 10686 15308 10692 15320
rect 10744 15308 10750 15360
rect 18601 15351 18659 15357
rect 18601 15317 18613 15351
rect 18647 15348 18659 15351
rect 19242 15348 19248 15360
rect 18647 15320 19248 15348
rect 18647 15317 18659 15320
rect 18601 15311 18659 15317
rect 19242 15308 19248 15320
rect 19300 15308 19306 15360
rect 20625 15351 20683 15357
rect 20625 15317 20637 15351
rect 20671 15348 20683 15351
rect 20714 15348 20720 15360
rect 20671 15320 20720 15348
rect 20671 15317 20683 15320
rect 20625 15311 20683 15317
rect 20714 15308 20720 15320
rect 20772 15348 20778 15360
rect 22557 15351 22615 15357
rect 22557 15348 22569 15351
rect 20772 15320 22569 15348
rect 20772 15308 20778 15320
rect 22557 15317 22569 15320
rect 22603 15317 22615 15351
rect 22557 15311 22615 15317
rect 24121 15351 24179 15357
rect 24121 15317 24133 15351
rect 24167 15348 24179 15351
rect 24762 15348 24768 15360
rect 24167 15320 24768 15348
rect 24167 15317 24179 15320
rect 24121 15311 24179 15317
rect 24762 15308 24768 15320
rect 24820 15308 24826 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1489 15147 1547 15153
rect 1489 15113 1501 15147
rect 1535 15144 1547 15147
rect 2130 15144 2136 15156
rect 1535 15116 2136 15144
rect 1535 15113 1547 15116
rect 1489 15107 1547 15113
rect 2130 15104 2136 15116
rect 2188 15104 2194 15156
rect 2866 15144 2872 15156
rect 2827 15116 2872 15144
rect 2866 15104 2872 15116
rect 2924 15104 2930 15156
rect 3602 15144 3608 15156
rect 3563 15116 3608 15144
rect 3602 15104 3608 15116
rect 3660 15104 3666 15156
rect 4154 15144 4160 15156
rect 4115 15116 4160 15144
rect 4154 15104 4160 15116
rect 4212 15104 4218 15156
rect 5534 15104 5540 15156
rect 5592 15144 5598 15156
rect 5629 15147 5687 15153
rect 5629 15144 5641 15147
rect 5592 15116 5641 15144
rect 5592 15104 5598 15116
rect 5629 15113 5641 15116
rect 5675 15113 5687 15147
rect 6178 15144 6184 15156
rect 6139 15116 6184 15144
rect 5629 15107 5687 15113
rect 6178 15104 6184 15116
rect 6236 15104 6242 15156
rect 6914 15144 6920 15156
rect 6875 15116 6920 15144
rect 6914 15104 6920 15116
rect 6972 15104 6978 15156
rect 7006 15104 7012 15156
rect 7064 15144 7070 15156
rect 7929 15147 7987 15153
rect 7929 15144 7941 15147
rect 7064 15116 7941 15144
rect 7064 15104 7070 15116
rect 7929 15113 7941 15116
rect 7975 15144 7987 15147
rect 8294 15144 8300 15156
rect 7975 15116 8300 15144
rect 7975 15113 7987 15116
rect 7929 15107 7987 15113
rect 8294 15104 8300 15116
rect 8352 15104 8358 15156
rect 10134 15104 10140 15156
rect 10192 15144 10198 15156
rect 10192 15116 11192 15144
rect 10192 15104 10198 15116
rect 2498 15076 2504 15088
rect 1964 15048 2504 15076
rect 1762 14968 1768 15020
rect 1820 15008 1826 15020
rect 1964 15017 1992 15048
rect 2498 15036 2504 15048
rect 2556 15036 2562 15088
rect 11164 15076 11192 15116
rect 11422 15104 11428 15156
rect 11480 15144 11486 15156
rect 12161 15147 12219 15153
rect 12161 15144 12173 15147
rect 11480 15116 12173 15144
rect 11480 15104 11486 15116
rect 12161 15113 12173 15116
rect 12207 15113 12219 15147
rect 12161 15107 12219 15113
rect 11793 15079 11851 15085
rect 11793 15076 11805 15079
rect 11164 15048 11805 15076
rect 11793 15045 11805 15048
rect 11839 15076 11851 15079
rect 11839 15048 12112 15076
rect 11839 15045 11851 15048
rect 11793 15039 11851 15045
rect 1949 15011 2007 15017
rect 1949 15008 1961 15011
rect 1820 14980 1961 15008
rect 1820 14968 1826 14980
rect 1949 14977 1961 14980
rect 1995 14977 2007 15011
rect 1949 14971 2007 14977
rect 2041 15011 2099 15017
rect 2041 14977 2053 15011
rect 2087 15008 2099 15011
rect 2682 15008 2688 15020
rect 2087 14980 2688 15008
rect 2087 14977 2099 14980
rect 2041 14971 2099 14977
rect 2682 14968 2688 14980
rect 2740 14968 2746 15020
rect 2961 14943 3019 14949
rect 2961 14909 2973 14943
rect 3007 14940 3019 14943
rect 3050 14940 3056 14952
rect 3007 14912 3056 14940
rect 3007 14909 3019 14912
rect 2961 14903 3019 14909
rect 3050 14900 3056 14912
rect 3108 14940 3114 14952
rect 3602 14940 3608 14952
rect 3108 14912 3608 14940
rect 3108 14900 3114 14912
rect 3602 14900 3608 14912
rect 3660 14900 3666 14952
rect 4062 14900 4068 14952
rect 4120 14940 4126 14952
rect 4249 14943 4307 14949
rect 4249 14940 4261 14943
rect 4120 14912 4261 14940
rect 4120 14900 4126 14912
rect 4249 14909 4261 14912
rect 4295 14940 4307 14943
rect 4798 14940 4804 14952
rect 4295 14912 4804 14940
rect 4295 14909 4307 14912
rect 4249 14903 4307 14909
rect 4798 14900 4804 14912
rect 4856 14900 4862 14952
rect 6730 14900 6736 14952
rect 6788 14940 6794 14952
rect 7193 14943 7251 14949
rect 7193 14940 7205 14943
rect 6788 14912 7205 14940
rect 6788 14900 6794 14912
rect 7193 14909 7205 14912
rect 7239 14909 7251 14943
rect 9030 14940 9036 14952
rect 8943 14912 9036 14940
rect 7193 14903 7251 14909
rect 9030 14900 9036 14912
rect 9088 14940 9094 14952
rect 9861 14943 9919 14949
rect 9861 14940 9873 14943
rect 9088 14912 9873 14940
rect 9088 14900 9094 14912
rect 9861 14909 9873 14912
rect 9907 14940 9919 14943
rect 11698 14940 11704 14952
rect 9907 14912 11704 14940
rect 9907 14909 9919 14912
rect 9861 14903 9919 14909
rect 11698 14900 11704 14912
rect 11756 14900 11762 14952
rect 12084 14940 12112 15048
rect 12176 15008 12204 15107
rect 12434 15104 12440 15156
rect 12492 15144 12498 15156
rect 13449 15147 13507 15153
rect 13449 15144 13461 15147
rect 12492 15116 13461 15144
rect 12492 15104 12498 15116
rect 13449 15113 13461 15116
rect 13495 15113 13507 15147
rect 16482 15144 16488 15156
rect 16443 15116 16488 15144
rect 13449 15107 13507 15113
rect 16482 15104 16488 15116
rect 16540 15104 16546 15156
rect 16666 15104 16672 15156
rect 16724 15144 16730 15156
rect 16761 15147 16819 15153
rect 16761 15144 16773 15147
rect 16724 15116 16773 15144
rect 16724 15104 16730 15116
rect 16761 15113 16773 15116
rect 16807 15113 16819 15147
rect 17402 15144 17408 15156
rect 17363 15116 17408 15144
rect 16761 15107 16819 15113
rect 17402 15104 17408 15116
rect 17460 15104 17466 15156
rect 19978 15144 19984 15156
rect 19939 15116 19984 15144
rect 19978 15104 19984 15116
rect 20036 15104 20042 15156
rect 20441 15147 20499 15153
rect 20441 15113 20453 15147
rect 20487 15144 20499 15147
rect 20806 15144 20812 15156
rect 20487 15116 20812 15144
rect 20487 15113 20499 15116
rect 20441 15107 20499 15113
rect 20806 15104 20812 15116
rect 20864 15104 20870 15156
rect 21266 15104 21272 15156
rect 21324 15144 21330 15156
rect 21545 15147 21603 15153
rect 21545 15144 21557 15147
rect 21324 15116 21557 15144
rect 21324 15104 21330 15116
rect 21545 15113 21557 15116
rect 21591 15144 21603 15147
rect 21634 15144 21640 15156
rect 21591 15116 21640 15144
rect 21591 15113 21603 15116
rect 21545 15107 21603 15113
rect 21634 15104 21640 15116
rect 21692 15104 21698 15156
rect 21910 15144 21916 15156
rect 21871 15116 21916 15144
rect 21910 15104 21916 15116
rect 21968 15104 21974 15156
rect 22646 15144 22652 15156
rect 22607 15116 22652 15144
rect 22646 15104 22652 15116
rect 22704 15104 22710 15156
rect 23474 15144 23480 15156
rect 23435 15116 23480 15144
rect 23474 15104 23480 15116
rect 23532 15104 23538 15156
rect 24670 15144 24676 15156
rect 24631 15116 24676 15144
rect 24670 15104 24676 15116
rect 24728 15104 24734 15156
rect 12529 15079 12587 15085
rect 12529 15045 12541 15079
rect 12575 15076 12587 15079
rect 13262 15076 13268 15088
rect 12575 15048 13268 15076
rect 12575 15045 12587 15048
rect 12529 15039 12587 15045
rect 13262 15036 13268 15048
rect 13320 15036 13326 15088
rect 15102 15076 15108 15088
rect 15063 15048 15108 15076
rect 15102 15036 15108 15048
rect 15160 15036 15166 15088
rect 20622 15076 20628 15088
rect 20583 15048 20628 15076
rect 20622 15036 20628 15048
rect 20680 15036 20686 15088
rect 23750 15076 23756 15088
rect 23711 15048 23756 15076
rect 23750 15036 23756 15048
rect 23808 15036 23814 15088
rect 12897 15011 12955 15017
rect 12897 15008 12909 15011
rect 12176 14980 12909 15008
rect 12897 14977 12909 14980
rect 12943 14977 12955 15011
rect 13078 15008 13084 15020
rect 12991 14980 13084 15008
rect 12897 14971 12955 14977
rect 13078 14968 13084 14980
rect 13136 15008 13142 15020
rect 13906 15008 13912 15020
rect 13136 14980 13912 15008
rect 13136 14968 13142 14980
rect 13906 14968 13912 14980
rect 13964 14968 13970 15020
rect 15378 14968 15384 15020
rect 15436 15008 15442 15020
rect 15565 15011 15623 15017
rect 15565 15008 15577 15011
rect 15436 14980 15577 15008
rect 15436 14968 15442 14980
rect 15565 14977 15577 14980
rect 15611 15008 15623 15011
rect 16025 15011 16083 15017
rect 16025 15008 16037 15011
rect 15611 14980 16037 15008
rect 15611 14977 15623 14980
rect 15565 14971 15623 14977
rect 16025 14977 16037 14980
rect 16071 14977 16083 15011
rect 20990 15008 20996 15020
rect 20951 14980 20996 15008
rect 16025 14971 16083 14977
rect 20990 14968 20996 14980
rect 21048 14968 21054 15020
rect 22094 14968 22100 15020
rect 22152 15008 22158 15020
rect 22152 14980 22197 15008
rect 22152 14968 22158 14980
rect 12084 14912 13032 14940
rect 1946 14872 1952 14884
rect 1859 14844 1952 14872
rect 1946 14832 1952 14844
rect 2004 14872 2010 14884
rect 2590 14872 2596 14884
rect 2004 14844 2596 14872
rect 2004 14832 2010 14844
rect 2590 14832 2596 14844
rect 2648 14832 2654 14884
rect 4338 14832 4344 14884
rect 4396 14872 4402 14884
rect 4494 14875 4552 14881
rect 4494 14872 4506 14875
rect 4396 14844 4506 14872
rect 4396 14832 4402 14844
rect 4494 14841 4506 14844
rect 4540 14841 4552 14875
rect 4494 14835 4552 14841
rect 5074 14832 5080 14884
rect 5132 14872 5138 14884
rect 6549 14875 6607 14881
rect 6549 14872 6561 14875
rect 5132 14844 6561 14872
rect 5132 14832 5138 14844
rect 6549 14841 6561 14844
rect 6595 14872 6607 14875
rect 7098 14872 7104 14884
rect 6595 14844 7104 14872
rect 6595 14841 6607 14844
rect 6549 14835 6607 14841
rect 7098 14832 7104 14844
rect 7156 14832 7162 14884
rect 7374 14872 7380 14884
rect 7335 14844 7380 14872
rect 7374 14832 7380 14844
rect 7432 14832 7438 14884
rect 7466 14832 7472 14884
rect 7524 14872 7530 14884
rect 8294 14872 8300 14884
rect 7524 14844 7569 14872
rect 8255 14844 8300 14872
rect 7524 14832 7530 14844
rect 8294 14832 8300 14844
rect 8352 14832 8358 14884
rect 9490 14832 9496 14884
rect 9548 14872 9554 14884
rect 10106 14875 10164 14881
rect 10106 14872 10118 14875
rect 9548 14844 10118 14872
rect 9548 14832 9554 14844
rect 10106 14841 10118 14844
rect 10152 14872 10164 14875
rect 10686 14872 10692 14884
rect 10152 14844 10692 14872
rect 10152 14841 10164 14844
rect 10106 14835 10164 14841
rect 10686 14832 10692 14844
rect 10744 14832 10750 14884
rect 13004 14881 13032 14912
rect 13814 14900 13820 14952
rect 13872 14940 13878 14952
rect 14001 14943 14059 14949
rect 14001 14940 14013 14943
rect 13872 14912 14013 14940
rect 13872 14900 13878 14912
rect 14001 14909 14013 14912
rect 14047 14909 14059 14943
rect 14001 14903 14059 14909
rect 14921 14943 14979 14949
rect 14921 14909 14933 14943
rect 14967 14940 14979 14943
rect 15657 14943 15715 14949
rect 15657 14940 15669 14943
rect 14967 14912 15669 14940
rect 14967 14909 14979 14912
rect 14921 14903 14979 14909
rect 15657 14909 15669 14912
rect 15703 14940 15715 14943
rect 16390 14940 16396 14952
rect 15703 14912 16396 14940
rect 15703 14909 15715 14912
rect 15657 14903 15715 14909
rect 16390 14900 16396 14912
rect 16448 14900 16454 14952
rect 18049 14943 18107 14949
rect 18049 14909 18061 14943
rect 18095 14909 18107 14943
rect 18049 14903 18107 14909
rect 12989 14875 13047 14881
rect 12989 14841 13001 14875
rect 13035 14841 13047 14875
rect 15565 14875 15623 14881
rect 15565 14872 15577 14875
rect 12989 14835 13047 14841
rect 14476 14844 15577 14872
rect 14476 14816 14504 14844
rect 15565 14841 15577 14844
rect 15611 14841 15623 14875
rect 15565 14835 15623 14841
rect 15838 14832 15844 14884
rect 15896 14872 15902 14884
rect 17773 14875 17831 14881
rect 17773 14872 17785 14875
rect 15896 14844 17785 14872
rect 15896 14832 15902 14844
rect 17773 14841 17785 14844
rect 17819 14872 17831 14875
rect 18064 14872 18092 14903
rect 18138 14900 18144 14952
rect 18196 14940 18202 14952
rect 18305 14943 18363 14949
rect 18305 14940 18317 14943
rect 18196 14912 18317 14940
rect 18196 14900 18202 14912
rect 18305 14909 18317 14912
rect 18351 14909 18363 14943
rect 19978 14940 19984 14952
rect 19891 14912 19984 14940
rect 18305 14903 18363 14909
rect 19518 14872 19524 14884
rect 17819 14844 19524 14872
rect 17819 14841 17831 14844
rect 17773 14835 17831 14841
rect 19518 14832 19524 14844
rect 19576 14832 19582 14884
rect 1578 14764 1584 14816
rect 1636 14804 1642 14816
rect 2130 14804 2136 14816
rect 1636 14776 2136 14804
rect 1636 14764 1642 14776
rect 2130 14764 2136 14776
rect 2188 14804 2194 14816
rect 2409 14807 2467 14813
rect 2409 14804 2421 14807
rect 2188 14776 2421 14804
rect 2188 14764 2194 14776
rect 2409 14773 2421 14776
rect 2455 14773 2467 14807
rect 3142 14804 3148 14816
rect 3103 14776 3148 14804
rect 2409 14767 2467 14773
rect 3142 14764 3148 14776
rect 3200 14764 3206 14816
rect 8478 14804 8484 14816
rect 8439 14776 8484 14804
rect 8478 14764 8484 14776
rect 8536 14764 8542 14816
rect 9401 14807 9459 14813
rect 9401 14773 9413 14807
rect 9447 14804 9459 14807
rect 9582 14804 9588 14816
rect 9447 14776 9588 14804
rect 9447 14773 9459 14776
rect 9401 14767 9459 14773
rect 9582 14764 9588 14776
rect 9640 14764 9646 14816
rect 9766 14804 9772 14816
rect 9727 14776 9772 14804
rect 9766 14764 9772 14776
rect 9824 14804 9830 14816
rect 9950 14804 9956 14816
rect 9824 14776 9956 14804
rect 9824 14764 9830 14776
rect 9950 14764 9956 14776
rect 10008 14764 10014 14816
rect 11238 14804 11244 14816
rect 11199 14776 11244 14804
rect 11238 14764 11244 14776
rect 11296 14764 11302 14816
rect 14458 14804 14464 14816
rect 14419 14776 14464 14804
rect 14458 14764 14464 14776
rect 14516 14764 14522 14816
rect 16942 14804 16948 14816
rect 16903 14776 16948 14804
rect 16942 14764 16948 14776
rect 17000 14764 17006 14816
rect 19150 14764 19156 14816
rect 19208 14804 19214 14816
rect 19429 14807 19487 14813
rect 19429 14804 19441 14807
rect 19208 14776 19441 14804
rect 19208 14764 19214 14776
rect 19429 14773 19441 14776
rect 19475 14804 19487 14807
rect 19904 14804 19932 14912
rect 19978 14900 19984 14912
rect 20036 14940 20042 14952
rect 24026 14940 24032 14952
rect 20036 14912 21220 14940
rect 23987 14912 24032 14940
rect 20036 14900 20042 14912
rect 21192 14884 21220 14912
rect 24026 14900 24032 14912
rect 24084 14900 24090 14952
rect 24946 14900 24952 14952
rect 25004 14940 25010 14952
rect 25225 14943 25283 14949
rect 25225 14940 25237 14943
rect 25004 14912 25237 14940
rect 25004 14900 25010 14912
rect 25225 14909 25237 14912
rect 25271 14940 25283 14943
rect 25777 14943 25835 14949
rect 25777 14940 25789 14943
rect 25271 14912 25789 14940
rect 25271 14909 25283 14912
rect 25225 14903 25283 14909
rect 25777 14909 25789 14912
rect 25823 14909 25835 14943
rect 25777 14903 25835 14909
rect 20714 14832 20720 14884
rect 20772 14872 20778 14884
rect 21085 14875 21143 14881
rect 21085 14872 21097 14875
rect 20772 14844 21097 14872
rect 20772 14832 20778 14844
rect 21085 14841 21097 14844
rect 21131 14841 21143 14875
rect 21085 14835 21143 14841
rect 21174 14832 21180 14884
rect 21232 14872 21238 14884
rect 21232 14844 21277 14872
rect 21232 14832 21238 14844
rect 22830 14832 22836 14884
rect 22888 14872 22894 14884
rect 24213 14875 24271 14881
rect 24213 14872 24225 14875
rect 22888 14844 24225 14872
rect 22888 14832 22894 14844
rect 24213 14841 24225 14844
rect 24259 14841 24271 14875
rect 24213 14835 24271 14841
rect 24305 14875 24363 14881
rect 24305 14841 24317 14875
rect 24351 14872 24363 14875
rect 25038 14872 25044 14884
rect 24351 14844 25044 14872
rect 24351 14841 24363 14844
rect 24305 14835 24363 14841
rect 25038 14832 25044 14844
rect 25096 14832 25102 14884
rect 19475 14776 19932 14804
rect 19475 14773 19487 14776
rect 19429 14767 19487 14773
rect 22094 14764 22100 14816
rect 22152 14804 22158 14816
rect 22925 14807 22983 14813
rect 22925 14804 22937 14807
rect 22152 14776 22937 14804
rect 22152 14764 22158 14776
rect 22925 14773 22937 14776
rect 22971 14804 22983 14807
rect 23014 14804 23020 14816
rect 22971 14776 23020 14804
rect 22971 14773 22983 14776
rect 22925 14767 22983 14773
rect 23014 14764 23020 14776
rect 23072 14764 23078 14816
rect 25409 14807 25467 14813
rect 25409 14773 25421 14807
rect 25455 14804 25467 14807
rect 25590 14804 25596 14816
rect 25455 14776 25596 14804
rect 25455 14773 25467 14776
rect 25409 14767 25467 14773
rect 25590 14764 25596 14776
rect 25648 14764 25654 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 2777 14603 2835 14609
rect 2777 14569 2789 14603
rect 2823 14600 2835 14603
rect 2866 14600 2872 14612
rect 2823 14572 2872 14600
rect 2823 14569 2835 14572
rect 2777 14563 2835 14569
rect 1394 14492 1400 14544
rect 1452 14532 1458 14544
rect 2038 14532 2044 14544
rect 1452 14504 2044 14532
rect 1452 14492 1458 14504
rect 2038 14492 2044 14504
rect 2096 14492 2102 14544
rect 2222 14532 2228 14544
rect 2135 14504 2228 14532
rect 2222 14492 2228 14504
rect 2280 14492 2286 14544
rect 2314 14492 2320 14544
rect 2372 14532 2378 14544
rect 2792 14532 2820 14563
rect 2866 14560 2872 14572
rect 2924 14600 2930 14612
rect 3053 14603 3111 14609
rect 3053 14600 3065 14603
rect 2924 14572 3065 14600
rect 2924 14560 2930 14572
rect 3053 14569 3065 14572
rect 3099 14569 3111 14603
rect 3053 14563 3111 14569
rect 4338 14560 4344 14612
rect 4396 14600 4402 14612
rect 5074 14600 5080 14612
rect 4396 14572 5080 14600
rect 4396 14560 4402 14572
rect 5074 14560 5080 14572
rect 5132 14600 5138 14612
rect 5445 14603 5503 14609
rect 5445 14600 5457 14603
rect 5132 14572 5457 14600
rect 5132 14560 5138 14572
rect 5445 14569 5457 14572
rect 5491 14569 5503 14603
rect 5445 14563 5503 14569
rect 5534 14560 5540 14612
rect 5592 14600 5598 14612
rect 5997 14603 6055 14609
rect 5997 14600 6009 14603
rect 5592 14572 6009 14600
rect 5592 14560 5598 14572
rect 5997 14569 6009 14572
rect 6043 14600 6055 14603
rect 6457 14603 6515 14609
rect 6457 14600 6469 14603
rect 6043 14572 6469 14600
rect 6043 14569 6055 14572
rect 5997 14563 6055 14569
rect 6457 14569 6469 14572
rect 6503 14600 6515 14603
rect 6825 14603 6883 14609
rect 6825 14600 6837 14603
rect 6503 14572 6837 14600
rect 6503 14569 6515 14572
rect 6457 14563 6515 14569
rect 6825 14569 6837 14572
rect 6871 14600 6883 14603
rect 7466 14600 7472 14612
rect 6871 14572 7472 14600
rect 6871 14569 6883 14572
rect 6825 14563 6883 14569
rect 7466 14560 7472 14572
rect 7524 14560 7530 14612
rect 8386 14600 8392 14612
rect 8347 14572 8392 14600
rect 8386 14560 8392 14572
rect 8444 14600 8450 14612
rect 8938 14600 8944 14612
rect 8444 14572 8944 14600
rect 8444 14560 8450 14572
rect 8938 14560 8944 14572
rect 8996 14560 9002 14612
rect 9398 14600 9404 14612
rect 9359 14572 9404 14600
rect 9398 14560 9404 14572
rect 9456 14560 9462 14612
rect 9858 14560 9864 14612
rect 9916 14600 9922 14612
rect 10413 14603 10471 14609
rect 10413 14600 10425 14603
rect 9916 14572 10425 14600
rect 9916 14560 9922 14572
rect 10413 14569 10425 14572
rect 10459 14569 10471 14603
rect 10413 14563 10471 14569
rect 12805 14603 12863 14609
rect 12805 14569 12817 14603
rect 12851 14600 12863 14603
rect 13078 14600 13084 14612
rect 12851 14572 13084 14600
rect 12851 14569 12863 14572
rect 12805 14563 12863 14569
rect 13078 14560 13084 14572
rect 13136 14560 13142 14612
rect 14274 14560 14280 14612
rect 14332 14600 14338 14612
rect 15841 14603 15899 14609
rect 15841 14600 15853 14603
rect 14332 14572 15853 14600
rect 14332 14560 14338 14572
rect 15841 14569 15853 14572
rect 15887 14569 15899 14603
rect 15841 14563 15899 14569
rect 16942 14560 16948 14612
rect 17000 14600 17006 14612
rect 18049 14603 18107 14609
rect 18049 14600 18061 14603
rect 17000 14572 18061 14600
rect 17000 14560 17006 14572
rect 18049 14569 18061 14572
rect 18095 14600 18107 14603
rect 18414 14600 18420 14612
rect 18095 14572 18420 14600
rect 18095 14569 18107 14572
rect 18049 14563 18107 14569
rect 18414 14560 18420 14572
rect 18472 14560 18478 14612
rect 18874 14600 18880 14612
rect 18835 14572 18880 14600
rect 18874 14560 18880 14572
rect 18932 14560 18938 14612
rect 19334 14560 19340 14612
rect 19392 14600 19398 14612
rect 19797 14603 19855 14609
rect 19797 14600 19809 14603
rect 19392 14572 19809 14600
rect 19392 14560 19398 14572
rect 19797 14569 19809 14572
rect 19843 14569 19855 14603
rect 19797 14563 19855 14569
rect 20625 14603 20683 14609
rect 20625 14569 20637 14603
rect 20671 14600 20683 14603
rect 21174 14600 21180 14612
rect 20671 14572 21180 14600
rect 20671 14569 20683 14572
rect 20625 14563 20683 14569
rect 21174 14560 21180 14572
rect 21232 14560 21238 14612
rect 22830 14600 22836 14612
rect 22791 14572 22836 14600
rect 22830 14560 22836 14572
rect 22888 14560 22894 14612
rect 24026 14560 24032 14612
rect 24084 14600 24090 14612
rect 25317 14603 25375 14609
rect 25317 14600 25329 14603
rect 24084 14572 25329 14600
rect 24084 14560 24090 14572
rect 25317 14569 25329 14572
rect 25363 14569 25375 14603
rect 25317 14563 25375 14569
rect 2372 14504 2820 14532
rect 7745 14535 7803 14541
rect 2372 14492 2378 14504
rect 7745 14501 7757 14535
rect 7791 14532 7803 14535
rect 8110 14532 8116 14544
rect 7791 14504 8116 14532
rect 7791 14501 7803 14504
rect 7745 14495 7803 14501
rect 8110 14492 8116 14504
rect 8168 14492 8174 14544
rect 11241 14535 11299 14541
rect 11241 14532 11253 14535
rect 10520 14504 11253 14532
rect 2240 14464 2268 14492
rect 2498 14464 2504 14476
rect 2240 14436 2504 14464
rect 2498 14424 2504 14436
rect 2556 14424 2562 14476
rect 3326 14424 3332 14476
rect 3384 14464 3390 14476
rect 4321 14467 4379 14473
rect 4321 14464 4333 14467
rect 3384 14436 4333 14464
rect 3384 14424 3390 14436
rect 4321 14433 4333 14436
rect 4367 14433 4379 14467
rect 4321 14427 4379 14433
rect 7098 14424 7104 14476
rect 7156 14464 7162 14476
rect 7837 14467 7895 14473
rect 7837 14464 7849 14467
rect 7156 14436 7849 14464
rect 7156 14424 7162 14436
rect 7837 14433 7849 14436
rect 7883 14433 7895 14467
rect 10226 14464 10232 14476
rect 10187 14436 10232 14464
rect 7837 14427 7895 14433
rect 10226 14424 10232 14436
rect 10284 14464 10290 14476
rect 10520 14464 10548 14504
rect 11241 14501 11253 14504
rect 11287 14501 11299 14535
rect 11241 14495 11299 14501
rect 17310 14492 17316 14544
rect 17368 14532 17374 14544
rect 17405 14535 17463 14541
rect 17405 14532 17417 14535
rect 17368 14504 17417 14532
rect 17368 14492 17374 14504
rect 17405 14501 17417 14504
rect 17451 14532 17463 14535
rect 17862 14532 17868 14544
rect 17451 14504 17868 14532
rect 17451 14501 17463 14504
rect 17405 14495 17463 14501
rect 17862 14492 17868 14504
rect 17920 14492 17926 14544
rect 18601 14535 18659 14541
rect 18601 14501 18613 14535
rect 18647 14532 18659 14535
rect 19150 14532 19156 14544
rect 18647 14504 19156 14532
rect 18647 14501 18659 14504
rect 18601 14495 18659 14501
rect 19150 14492 19156 14504
rect 19208 14492 19214 14544
rect 23382 14492 23388 14544
rect 23440 14532 23446 14544
rect 23630 14535 23688 14541
rect 23630 14532 23642 14535
rect 23440 14504 23642 14532
rect 23440 14492 23446 14504
rect 23630 14501 23642 14504
rect 23676 14501 23688 14535
rect 23630 14495 23688 14501
rect 11681 14467 11739 14473
rect 11681 14464 11693 14467
rect 10284 14436 10548 14464
rect 11256 14436 11693 14464
rect 10284 14424 10290 14436
rect 11256 14408 11284 14436
rect 11681 14433 11693 14436
rect 11727 14464 11739 14467
rect 12158 14464 12164 14476
rect 11727 14436 12164 14464
rect 11727 14433 11739 14436
rect 11681 14427 11739 14433
rect 12158 14424 12164 14436
rect 12216 14424 12222 14476
rect 13446 14464 13452 14476
rect 13407 14436 13452 14464
rect 13446 14424 13452 14436
rect 13504 14424 13510 14476
rect 15562 14424 15568 14476
rect 15620 14464 15626 14476
rect 15657 14467 15715 14473
rect 15657 14464 15669 14467
rect 15620 14436 15669 14464
rect 15620 14424 15626 14436
rect 15657 14433 15669 14436
rect 15703 14433 15715 14467
rect 15657 14427 15715 14433
rect 16390 14424 16396 14476
rect 16448 14464 16454 14476
rect 17497 14467 17555 14473
rect 17497 14464 17509 14467
rect 16448 14436 17509 14464
rect 16448 14424 16454 14436
rect 17497 14433 17509 14436
rect 17543 14433 17555 14467
rect 17497 14427 17555 14433
rect 19334 14424 19340 14476
rect 19392 14464 19398 14476
rect 19613 14467 19671 14473
rect 19613 14464 19625 14467
rect 19392 14436 19625 14464
rect 19392 14424 19398 14436
rect 19613 14433 19625 14436
rect 19659 14464 19671 14467
rect 20622 14464 20628 14476
rect 19659 14436 20628 14464
rect 19659 14433 19671 14436
rect 19613 14427 19671 14433
rect 20622 14424 20628 14436
rect 20680 14424 20686 14476
rect 20990 14424 20996 14476
rect 21048 14464 21054 14476
rect 21157 14467 21215 14473
rect 21157 14464 21169 14467
rect 21048 14436 21169 14464
rect 21048 14424 21054 14436
rect 21157 14433 21169 14436
rect 21203 14433 21215 14467
rect 21157 14427 21215 14433
rect 4062 14396 4068 14408
rect 4023 14368 4068 14396
rect 4062 14356 4068 14368
rect 4120 14356 4126 14408
rect 7745 14399 7803 14405
rect 7745 14365 7757 14399
rect 7791 14365 7803 14399
rect 10502 14396 10508 14408
rect 10463 14368 10508 14396
rect 7745 14359 7803 14365
rect 1762 14328 1768 14340
rect 1723 14300 1768 14328
rect 1762 14288 1768 14300
rect 1820 14288 1826 14340
rect 6638 14288 6644 14340
rect 6696 14328 6702 14340
rect 7760 14328 7788 14359
rect 10502 14356 10508 14368
rect 10560 14396 10566 14408
rect 11238 14396 11244 14408
rect 10560 14368 11244 14396
rect 10560 14356 10566 14368
rect 11238 14356 11244 14368
rect 11296 14356 11302 14408
rect 11425 14399 11483 14405
rect 11425 14365 11437 14399
rect 11471 14365 11483 14399
rect 11425 14359 11483 14365
rect 15105 14399 15163 14405
rect 15105 14365 15117 14399
rect 15151 14396 15163 14399
rect 15933 14399 15991 14405
rect 15933 14396 15945 14399
rect 15151 14368 15945 14396
rect 15151 14365 15163 14368
rect 15105 14359 15163 14365
rect 15933 14365 15945 14368
rect 15979 14396 15991 14399
rect 16022 14396 16028 14408
rect 15979 14368 16028 14396
rect 15979 14365 15991 14368
rect 15933 14359 15991 14365
rect 8202 14328 8208 14340
rect 6696 14300 8208 14328
rect 6696 14288 6702 14300
rect 8202 14288 8208 14300
rect 8260 14288 8266 14340
rect 9953 14331 10011 14337
rect 9953 14297 9965 14331
rect 9999 14328 10011 14331
rect 10962 14328 10968 14340
rect 9999 14300 10968 14328
rect 9999 14297 10011 14300
rect 9953 14291 10011 14297
rect 10962 14288 10968 14300
rect 11020 14288 11026 14340
rect 3513 14263 3571 14269
rect 3513 14229 3525 14263
rect 3559 14260 3571 14263
rect 3602 14260 3608 14272
rect 3559 14232 3608 14260
rect 3559 14229 3571 14232
rect 3513 14223 3571 14229
rect 3602 14220 3608 14232
rect 3660 14220 3666 14272
rect 3881 14263 3939 14269
rect 3881 14229 3893 14263
rect 3927 14260 3939 14263
rect 4062 14260 4068 14272
rect 3927 14232 4068 14260
rect 3927 14229 3939 14232
rect 3881 14223 3939 14229
rect 4062 14220 4068 14232
rect 4120 14220 4126 14272
rect 7282 14260 7288 14272
rect 7243 14232 7288 14260
rect 7282 14220 7288 14232
rect 7340 14220 7346 14272
rect 8849 14263 8907 14269
rect 8849 14229 8861 14263
rect 8895 14260 8907 14263
rect 9030 14260 9036 14272
rect 8895 14232 9036 14260
rect 8895 14229 8907 14232
rect 8849 14223 8907 14229
rect 9030 14220 9036 14232
rect 9088 14220 9094 14272
rect 10873 14263 10931 14269
rect 10873 14229 10885 14263
rect 10919 14260 10931 14263
rect 11146 14260 11152 14272
rect 10919 14232 11152 14260
rect 10919 14229 10931 14232
rect 10873 14223 10931 14229
rect 11146 14220 11152 14232
rect 11204 14220 11210 14272
rect 11440 14260 11468 14359
rect 16022 14356 16028 14368
rect 16080 14356 16086 14408
rect 16761 14399 16819 14405
rect 16761 14365 16773 14399
rect 16807 14396 16819 14399
rect 17402 14396 17408 14408
rect 16807 14368 17408 14396
rect 16807 14365 16819 14368
rect 16761 14359 16819 14365
rect 17402 14356 17408 14368
rect 17460 14356 17466 14408
rect 19886 14396 19892 14408
rect 19847 14368 19892 14396
rect 19886 14356 19892 14368
rect 19944 14356 19950 14408
rect 20898 14396 20904 14408
rect 20859 14368 20904 14396
rect 20898 14356 20904 14368
rect 20956 14356 20962 14408
rect 23382 14396 23388 14408
rect 23343 14368 23388 14396
rect 23382 14356 23388 14368
rect 23440 14356 23446 14408
rect 15378 14328 15384 14340
rect 15339 14300 15384 14328
rect 15378 14288 15384 14300
rect 15436 14288 15442 14340
rect 11698 14260 11704 14272
rect 11440 14232 11704 14260
rect 11698 14220 11704 14232
rect 11756 14220 11762 14272
rect 16942 14260 16948 14272
rect 16903 14232 16948 14260
rect 16942 14220 16948 14232
rect 17000 14220 17006 14272
rect 19337 14263 19395 14269
rect 19337 14229 19349 14263
rect 19383 14260 19395 14263
rect 20530 14260 20536 14272
rect 19383 14232 20536 14260
rect 19383 14229 19395 14232
rect 19337 14223 19395 14229
rect 20530 14220 20536 14232
rect 20588 14220 20594 14272
rect 22278 14260 22284 14272
rect 22239 14232 22284 14260
rect 22278 14220 22284 14232
rect 22336 14220 22342 14272
rect 22830 14220 22836 14272
rect 22888 14260 22894 14272
rect 23293 14263 23351 14269
rect 23293 14260 23305 14263
rect 22888 14232 23305 14260
rect 22888 14220 22894 14232
rect 23293 14229 23305 14232
rect 23339 14260 23351 14263
rect 24765 14263 24823 14269
rect 24765 14260 24777 14263
rect 23339 14232 24777 14260
rect 23339 14229 23351 14232
rect 23293 14223 23351 14229
rect 24765 14229 24777 14232
rect 24811 14260 24823 14263
rect 24946 14260 24952 14272
rect 24811 14232 24952 14260
rect 24811 14229 24823 14232
rect 24765 14223 24823 14229
rect 24946 14220 24952 14232
rect 25004 14220 25010 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1489 14059 1547 14065
rect 1489 14025 1501 14059
rect 1535 14056 1547 14059
rect 1946 14056 1952 14068
rect 1535 14028 1952 14056
rect 1535 14025 1547 14028
rect 1489 14019 1547 14025
rect 1946 14016 1952 14028
rect 2004 14016 2010 14068
rect 2038 14016 2044 14068
rect 2096 14056 2102 14068
rect 2777 14059 2835 14065
rect 2777 14056 2789 14059
rect 2096 14028 2789 14056
rect 2096 14016 2102 14028
rect 2777 14025 2789 14028
rect 2823 14025 2835 14059
rect 3326 14056 3332 14068
rect 3287 14028 3332 14056
rect 2777 14019 2835 14025
rect 3326 14016 3332 14028
rect 3384 14016 3390 14068
rect 4154 14016 4160 14068
rect 4212 14056 4218 14068
rect 4433 14059 4491 14065
rect 4433 14056 4445 14059
rect 4212 14028 4445 14056
rect 4212 14016 4218 14028
rect 4433 14025 4445 14028
rect 4479 14025 4491 14059
rect 6638 14056 6644 14068
rect 6599 14028 6644 14056
rect 4433 14019 4491 14025
rect 6638 14016 6644 14028
rect 6696 14016 6702 14068
rect 6914 14056 6920 14068
rect 6875 14028 6920 14056
rect 6914 14016 6920 14028
rect 6972 14016 6978 14068
rect 9953 14059 10011 14065
rect 9953 14025 9965 14059
rect 9999 14056 10011 14059
rect 10502 14056 10508 14068
rect 9999 14028 10508 14056
rect 9999 14025 10011 14028
rect 9953 14019 10011 14025
rect 10502 14016 10508 14028
rect 10560 14016 10566 14068
rect 12158 14056 12164 14068
rect 12119 14028 12164 14056
rect 12158 14016 12164 14028
rect 12216 14016 12222 14068
rect 13173 14059 13231 14065
rect 13173 14056 13185 14059
rect 12268 14028 13185 14056
rect 2498 13988 2504 14000
rect 2459 13960 2504 13988
rect 2498 13948 2504 13960
rect 2556 13948 2562 14000
rect 3513 13991 3571 13997
rect 3513 13988 3525 13991
rect 2792 13960 3525 13988
rect 2792 13932 2820 13960
rect 3513 13957 3525 13960
rect 3559 13957 3571 13991
rect 3513 13951 3571 13957
rect 3602 13948 3608 14000
rect 3660 13988 3666 14000
rect 5169 13991 5227 13997
rect 5169 13988 5181 13991
rect 3660 13960 5181 13988
rect 3660 13948 3666 13960
rect 5169 13957 5181 13960
rect 5215 13957 5227 13991
rect 5169 13951 5227 13957
rect 8386 13948 8392 14000
rect 8444 13988 8450 14000
rect 8481 13991 8539 13997
rect 8481 13988 8493 13991
rect 8444 13960 8493 13988
rect 8444 13948 8450 13960
rect 8481 13957 8493 13960
rect 8527 13957 8539 13991
rect 8481 13951 8539 13957
rect 10134 13948 10140 14000
rect 10192 13988 10198 14000
rect 10229 13991 10287 13997
rect 10229 13988 10241 13991
rect 10192 13960 10241 13988
rect 10192 13948 10198 13960
rect 10229 13957 10241 13960
rect 10275 13957 10287 13991
rect 10229 13951 10287 13957
rect 10873 13991 10931 13997
rect 10873 13957 10885 13991
rect 10919 13988 10931 13991
rect 10962 13988 10968 14000
rect 10919 13960 10968 13988
rect 10919 13957 10931 13960
rect 10873 13951 10931 13957
rect 10962 13948 10968 13960
rect 11020 13948 11026 14000
rect 11054 13948 11060 14000
rect 11112 13988 11118 14000
rect 12268 13988 12296 14028
rect 13173 14025 13185 14028
rect 13219 14056 13231 14059
rect 13265 14059 13323 14065
rect 13265 14056 13277 14059
rect 13219 14028 13277 14056
rect 13219 14025 13231 14028
rect 13173 14019 13231 14025
rect 13265 14025 13277 14028
rect 13311 14025 13323 14059
rect 13265 14019 13323 14025
rect 13541 14059 13599 14065
rect 13541 14025 13553 14059
rect 13587 14056 13599 14059
rect 14458 14056 14464 14068
rect 13587 14028 14464 14056
rect 13587 14025 13599 14028
rect 13541 14019 13599 14025
rect 14458 14016 14464 14028
rect 14516 14016 14522 14068
rect 16390 14056 16396 14068
rect 16351 14028 16396 14056
rect 16390 14016 16396 14028
rect 16448 14056 16454 14068
rect 16945 14059 17003 14065
rect 16945 14056 16957 14059
rect 16448 14028 16957 14056
rect 16448 14016 16454 14028
rect 16945 14025 16957 14028
rect 16991 14025 17003 14059
rect 17310 14056 17316 14068
rect 17271 14028 17316 14056
rect 16945 14019 17003 14025
rect 17310 14016 17316 14028
rect 17368 14016 17374 14068
rect 17402 14016 17408 14068
rect 17460 14056 17466 14068
rect 18141 14059 18199 14065
rect 18141 14056 18153 14059
rect 17460 14028 18153 14056
rect 17460 14016 17466 14028
rect 18141 14025 18153 14028
rect 18187 14025 18199 14059
rect 18141 14019 18199 14025
rect 19153 14059 19211 14065
rect 19153 14025 19165 14059
rect 19199 14056 19211 14059
rect 19886 14056 19892 14068
rect 19199 14028 19892 14056
rect 19199 14025 19211 14028
rect 19153 14019 19211 14025
rect 19886 14016 19892 14028
rect 19944 14056 19950 14068
rect 20990 14056 20996 14068
rect 19944 14028 20996 14056
rect 19944 14016 19950 14028
rect 20990 14016 20996 14028
rect 21048 14016 21054 14068
rect 25038 14056 25044 14068
rect 24999 14028 25044 14056
rect 25038 14016 25044 14028
rect 25096 14016 25102 14068
rect 11112 13960 12296 13988
rect 12989 13991 13047 13997
rect 11112 13948 11118 13960
rect 12989 13957 13001 13991
rect 13035 13988 13047 13991
rect 13035 13960 14136 13988
rect 13035 13957 13047 13960
rect 12989 13951 13047 13957
rect 2041 13923 2099 13929
rect 2041 13889 2053 13923
rect 2087 13920 2099 13923
rect 2314 13920 2320 13932
rect 2087 13892 2320 13920
rect 2087 13889 2099 13892
rect 2041 13883 2099 13889
rect 2314 13880 2320 13892
rect 2372 13880 2378 13932
rect 2774 13880 2780 13932
rect 2832 13880 2838 13932
rect 3881 13923 3939 13929
rect 3881 13889 3893 13923
rect 3927 13920 3939 13923
rect 4062 13920 4068 13932
rect 3927 13892 4068 13920
rect 3927 13889 3939 13892
rect 3881 13883 3939 13889
rect 4062 13880 4068 13892
rect 4120 13880 4126 13932
rect 4985 13923 5043 13929
rect 4985 13889 4997 13923
rect 5031 13920 5043 13923
rect 5626 13920 5632 13932
rect 5031 13892 5632 13920
rect 5031 13889 5043 13892
rect 4985 13883 5043 13889
rect 5626 13880 5632 13892
rect 5684 13880 5690 13932
rect 7282 13880 7288 13932
rect 7340 13920 7346 13932
rect 7377 13923 7435 13929
rect 7377 13920 7389 13923
rect 7340 13892 7389 13920
rect 7340 13880 7346 13892
rect 7377 13889 7389 13892
rect 7423 13920 7435 13923
rect 9401 13923 9459 13929
rect 9401 13920 9413 13923
rect 7423 13892 9413 13920
rect 7423 13889 7435 13892
rect 7377 13883 7435 13889
rect 9401 13889 9413 13892
rect 9447 13889 9459 13923
rect 9401 13883 9459 13889
rect 11146 13880 11152 13932
rect 11204 13920 11210 13932
rect 14108 13929 14136 13960
rect 14274 13948 14280 14000
rect 14332 13988 14338 14000
rect 14829 13991 14887 13997
rect 14829 13988 14841 13991
rect 14332 13960 14841 13988
rect 14332 13948 14338 13960
rect 14829 13957 14841 13960
rect 14875 13957 14887 13991
rect 17770 13988 17776 14000
rect 17731 13960 17776 13988
rect 14829 13951 14887 13957
rect 17770 13948 17776 13960
rect 17828 13988 17834 14000
rect 19518 13988 19524 14000
rect 17828 13960 17908 13988
rect 19431 13960 19524 13988
rect 17828 13948 17834 13960
rect 11425 13923 11483 13929
rect 11425 13920 11437 13923
rect 11204 13892 11437 13920
rect 11204 13880 11210 13892
rect 11425 13889 11437 13892
rect 11471 13889 11483 13923
rect 11425 13883 11483 13889
rect 13173 13923 13231 13929
rect 13173 13889 13185 13923
rect 13219 13920 13231 13923
rect 13909 13923 13967 13929
rect 13909 13920 13921 13923
rect 13219 13892 13921 13920
rect 13219 13889 13231 13892
rect 13173 13883 13231 13889
rect 13909 13889 13921 13892
rect 13955 13889 13967 13923
rect 13909 13883 13967 13889
rect 14093 13923 14151 13929
rect 14093 13889 14105 13923
rect 14139 13920 14151 13923
rect 14553 13923 14611 13929
rect 14553 13920 14565 13923
rect 14139 13892 14565 13920
rect 14139 13889 14151 13892
rect 14093 13883 14151 13889
rect 14553 13889 14565 13892
rect 14599 13920 14611 13923
rect 14599 13892 15148 13920
rect 14599 13889 14611 13892
rect 14553 13883 14611 13889
rect 1762 13852 1768 13864
rect 1723 13824 1768 13852
rect 1762 13812 1768 13824
rect 1820 13812 1826 13864
rect 5534 13812 5540 13864
rect 5592 13852 5598 13864
rect 5721 13855 5779 13861
rect 5721 13852 5733 13855
rect 5592 13824 5733 13852
rect 5592 13812 5598 13824
rect 5721 13821 5733 13824
rect 5767 13852 5779 13855
rect 6822 13852 6828 13864
rect 5767 13824 6828 13852
rect 5767 13821 5779 13824
rect 5721 13815 5779 13821
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 7466 13852 7472 13864
rect 7427 13824 7472 13852
rect 7466 13812 7472 13824
rect 7524 13812 7530 13864
rect 7929 13855 7987 13861
rect 7929 13821 7941 13855
rect 7975 13852 7987 13855
rect 8110 13852 8116 13864
rect 7975 13824 8116 13852
rect 7975 13821 7987 13824
rect 7929 13815 7987 13821
rect 8110 13812 8116 13824
rect 8168 13812 8174 13864
rect 8297 13855 8355 13861
rect 8297 13821 8309 13855
rect 8343 13852 8355 13855
rect 8754 13852 8760 13864
rect 8343 13824 8760 13852
rect 8343 13821 8355 13824
rect 8297 13815 8355 13821
rect 8754 13812 8760 13824
rect 8812 13812 8818 13864
rect 9030 13852 9036 13864
rect 8991 13824 9036 13852
rect 9030 13812 9036 13824
rect 9088 13812 9094 13864
rect 10689 13855 10747 13861
rect 10689 13821 10701 13855
rect 10735 13852 10747 13855
rect 11330 13852 11336 13864
rect 10735 13824 11336 13852
rect 10735 13821 10747 13824
rect 10689 13815 10747 13821
rect 4062 13784 4068 13796
rect 4023 13756 4068 13784
rect 4062 13744 4068 13756
rect 4120 13744 4126 13796
rect 4522 13744 4528 13796
rect 4580 13784 4586 13796
rect 6181 13787 6239 13793
rect 6181 13784 6193 13787
rect 4580 13756 6193 13784
rect 4580 13744 4586 13756
rect 6181 13753 6193 13756
rect 6227 13784 6239 13787
rect 6730 13784 6736 13796
rect 6227 13756 6736 13784
rect 6227 13753 6239 13756
rect 6181 13747 6239 13753
rect 6730 13744 6736 13756
rect 6788 13744 6794 13796
rect 8938 13784 8944 13796
rect 8899 13756 8944 13784
rect 8938 13744 8944 13756
rect 8996 13744 9002 13796
rect 11164 13793 11192 13824
rect 11330 13812 11336 13824
rect 11388 13812 11394 13864
rect 13446 13812 13452 13864
rect 13504 13852 13510 13864
rect 15010 13852 15016 13864
rect 13504 13824 13768 13852
rect 14971 13824 15016 13852
rect 13504 13812 13510 13824
rect 11149 13787 11207 13793
rect 11149 13753 11161 13787
rect 11195 13753 11207 13787
rect 13740 13784 13768 13824
rect 15010 13812 15016 13824
rect 15068 13812 15074 13864
rect 15120 13852 15148 13892
rect 15280 13855 15338 13861
rect 15280 13852 15292 13855
rect 15120 13824 15292 13852
rect 15280 13821 15292 13824
rect 15326 13852 15338 13855
rect 16022 13852 16028 13864
rect 15326 13824 16028 13852
rect 15326 13821 15338 13824
rect 15280 13815 15338 13821
rect 16022 13812 16028 13824
rect 16080 13812 16086 13864
rect 14001 13787 14059 13793
rect 14001 13784 14013 13787
rect 13740 13756 14013 13784
rect 11149 13747 11207 13753
rect 14001 13753 14013 13756
rect 14047 13753 14059 13787
rect 17880 13784 17908 13960
rect 19518 13948 19524 13960
rect 19576 13988 19582 14000
rect 19576 13960 19656 13988
rect 19576 13948 19582 13960
rect 18690 13920 18696 13932
rect 18651 13892 18696 13920
rect 18690 13880 18696 13892
rect 18748 13880 18754 13932
rect 18414 13852 18420 13864
rect 18375 13824 18420 13852
rect 18414 13812 18420 13824
rect 18472 13812 18478 13864
rect 19628 13861 19656 13960
rect 19613 13855 19671 13861
rect 19613 13821 19625 13855
rect 19659 13852 19671 13855
rect 20898 13852 20904 13864
rect 19659 13824 20904 13852
rect 19659 13821 19671 13824
rect 19613 13815 19671 13821
rect 20898 13812 20904 13824
rect 20956 13852 20962 13864
rect 21545 13855 21603 13861
rect 21545 13852 21557 13855
rect 20956 13824 21557 13852
rect 20956 13812 20962 13824
rect 21545 13821 21557 13824
rect 21591 13852 21603 13855
rect 23017 13855 23075 13861
rect 23017 13852 23029 13855
rect 21591 13824 23029 13852
rect 21591 13821 21603 13824
rect 21545 13815 21603 13821
rect 23017 13821 23029 13824
rect 23063 13852 23075 13855
rect 23382 13852 23388 13864
rect 23063 13824 23388 13852
rect 23063 13821 23075 13824
rect 23017 13815 23075 13821
rect 23382 13812 23388 13824
rect 23440 13852 23446 13864
rect 23661 13855 23719 13861
rect 23661 13852 23673 13855
rect 23440 13824 23673 13852
rect 23440 13812 23446 13824
rect 23661 13821 23673 13824
rect 23707 13821 23719 13855
rect 23661 13815 23719 13821
rect 23928 13855 23986 13861
rect 23928 13821 23940 13855
rect 23974 13852 23986 13855
rect 24946 13852 24952 13864
rect 23974 13824 24952 13852
rect 23974 13821 23986 13824
rect 23928 13815 23986 13821
rect 24946 13812 24952 13824
rect 25004 13812 25010 13864
rect 18601 13787 18659 13793
rect 18601 13784 18613 13787
rect 17880 13756 18613 13784
rect 14001 13747 14059 13753
rect 18601 13753 18613 13756
rect 18647 13784 18659 13787
rect 18874 13784 18880 13796
rect 18647 13756 18880 13784
rect 18647 13753 18659 13756
rect 18601 13747 18659 13753
rect 18874 13744 18880 13756
rect 18932 13744 18938 13796
rect 19880 13787 19938 13793
rect 19880 13753 19892 13787
rect 19926 13784 19938 13787
rect 19978 13784 19984 13796
rect 19926 13756 19984 13784
rect 19926 13753 19938 13756
rect 19880 13747 19938 13753
rect 19978 13744 19984 13756
rect 20036 13744 20042 13796
rect 1946 13716 1952 13728
rect 1907 13688 1952 13716
rect 1946 13676 1952 13688
rect 2004 13676 2010 13728
rect 3602 13676 3608 13728
rect 3660 13716 3666 13728
rect 3973 13719 4031 13725
rect 3973 13716 3985 13719
rect 3660 13688 3985 13716
rect 3660 13676 3666 13688
rect 3973 13685 3985 13688
rect 4019 13685 4031 13719
rect 5626 13716 5632 13728
rect 5587 13688 5632 13716
rect 3973 13679 4031 13685
rect 5626 13676 5632 13688
rect 5684 13676 5690 13728
rect 7377 13719 7435 13725
rect 7377 13685 7389 13719
rect 7423 13716 7435 13719
rect 7834 13716 7840 13728
rect 7423 13688 7840 13716
rect 7423 13685 7435 13688
rect 7377 13679 7435 13685
rect 7834 13676 7840 13688
rect 7892 13676 7898 13728
rect 10134 13676 10140 13728
rect 10192 13716 10198 13728
rect 11333 13719 11391 13725
rect 11333 13716 11345 13719
rect 10192 13688 11345 13716
rect 10192 13676 10198 13688
rect 11333 13685 11345 13688
rect 11379 13685 11391 13719
rect 11333 13679 11391 13685
rect 11698 13676 11704 13728
rect 11756 13716 11762 13728
rect 11793 13719 11851 13725
rect 11793 13716 11805 13719
rect 11756 13688 11805 13716
rect 11756 13676 11762 13688
rect 11793 13685 11805 13688
rect 11839 13685 11851 13719
rect 11793 13679 11851 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1673 13515 1731 13521
rect 1673 13481 1685 13515
rect 1719 13512 1731 13515
rect 1762 13512 1768 13524
rect 1719 13484 1768 13512
rect 1719 13481 1731 13484
rect 1673 13475 1731 13481
rect 1762 13472 1768 13484
rect 1820 13472 1826 13524
rect 3050 13512 3056 13524
rect 2792 13484 3056 13512
rect 2038 13404 2044 13456
rect 2096 13444 2102 13456
rect 2792 13453 2820 13484
rect 3050 13472 3056 13484
rect 3108 13472 3114 13524
rect 3513 13515 3571 13521
rect 3513 13481 3525 13515
rect 3559 13512 3571 13515
rect 3878 13512 3884 13524
rect 3559 13484 3884 13512
rect 3559 13481 3571 13484
rect 3513 13475 3571 13481
rect 3878 13472 3884 13484
rect 3936 13512 3942 13524
rect 4062 13512 4068 13524
rect 3936 13484 4068 13512
rect 3936 13472 3942 13484
rect 4062 13472 4068 13484
rect 4120 13472 4126 13524
rect 5077 13515 5135 13521
rect 5077 13481 5089 13515
rect 5123 13512 5135 13515
rect 5442 13512 5448 13524
rect 5123 13484 5448 13512
rect 5123 13481 5135 13484
rect 5077 13475 5135 13481
rect 5442 13472 5448 13484
rect 5500 13472 5506 13524
rect 6822 13472 6828 13524
rect 6880 13512 6886 13524
rect 6917 13515 6975 13521
rect 6917 13512 6929 13515
rect 6880 13484 6929 13512
rect 6880 13472 6886 13484
rect 6917 13481 6929 13484
rect 6963 13481 6975 13515
rect 6917 13475 6975 13481
rect 7098 13472 7104 13524
rect 7156 13512 7162 13524
rect 7469 13515 7527 13521
rect 7469 13512 7481 13515
rect 7156 13484 7481 13512
rect 7156 13472 7162 13484
rect 7469 13481 7481 13484
rect 7515 13481 7527 13515
rect 7834 13512 7840 13524
rect 7795 13484 7840 13512
rect 7469 13475 7527 13481
rect 7834 13472 7840 13484
rect 7892 13472 7898 13524
rect 8018 13472 8024 13524
rect 8076 13512 8082 13524
rect 8573 13515 8631 13521
rect 8573 13512 8585 13515
rect 8076 13484 8585 13512
rect 8076 13472 8082 13484
rect 8573 13481 8585 13484
rect 8619 13481 8631 13515
rect 8573 13475 8631 13481
rect 9858 13472 9864 13524
rect 9916 13512 9922 13524
rect 10505 13515 10563 13521
rect 10505 13512 10517 13515
rect 9916 13484 10517 13512
rect 9916 13472 9922 13484
rect 10505 13481 10517 13484
rect 10551 13481 10563 13515
rect 10505 13475 10563 13481
rect 11146 13472 11152 13524
rect 11204 13512 11210 13524
rect 12069 13515 12127 13521
rect 12069 13512 12081 13515
rect 11204 13484 12081 13512
rect 11204 13472 11210 13484
rect 12069 13481 12081 13484
rect 12115 13512 12127 13515
rect 12342 13512 12348 13524
rect 12115 13484 12348 13512
rect 12115 13481 12127 13484
rect 12069 13475 12127 13481
rect 12342 13472 12348 13484
rect 12400 13472 12406 13524
rect 18233 13515 18291 13521
rect 18233 13481 18245 13515
rect 18279 13512 18291 13515
rect 18690 13512 18696 13524
rect 18279 13484 18696 13512
rect 18279 13481 18291 13484
rect 18233 13475 18291 13481
rect 18690 13472 18696 13484
rect 18748 13472 18754 13524
rect 19153 13515 19211 13521
rect 19153 13481 19165 13515
rect 19199 13512 19211 13515
rect 19242 13512 19248 13524
rect 19199 13484 19248 13512
rect 19199 13481 19211 13484
rect 19153 13475 19211 13481
rect 19242 13472 19248 13484
rect 19300 13472 19306 13524
rect 19978 13472 19984 13524
rect 20036 13512 20042 13524
rect 20257 13515 20315 13521
rect 20257 13512 20269 13515
rect 20036 13484 20269 13512
rect 20036 13472 20042 13484
rect 20257 13481 20269 13484
rect 20303 13481 20315 13515
rect 20257 13475 20315 13481
rect 20990 13472 20996 13524
rect 21048 13512 21054 13524
rect 21085 13515 21143 13521
rect 21085 13512 21097 13515
rect 21048 13484 21097 13512
rect 21048 13472 21054 13484
rect 21085 13481 21097 13484
rect 21131 13481 21143 13515
rect 21085 13475 21143 13481
rect 23290 13472 23296 13524
rect 23348 13512 23354 13524
rect 23385 13515 23443 13521
rect 23385 13512 23397 13515
rect 23348 13484 23397 13512
rect 23348 13472 23354 13484
rect 23385 13481 23397 13484
rect 23431 13512 23443 13515
rect 23566 13512 23572 13524
rect 23431 13484 23572 13512
rect 23431 13481 23443 13484
rect 23385 13475 23443 13481
rect 23566 13472 23572 13484
rect 23624 13472 23630 13524
rect 2777 13447 2835 13453
rect 2777 13444 2789 13447
rect 2096 13416 2789 13444
rect 2096 13404 2102 13416
rect 2777 13413 2789 13416
rect 2823 13413 2835 13447
rect 2958 13444 2964 13456
rect 2919 13416 2964 13444
rect 2777 13407 2835 13413
rect 2958 13404 2964 13416
rect 3016 13404 3022 13456
rect 3789 13447 3847 13453
rect 3789 13413 3801 13447
rect 3835 13444 3847 13447
rect 3970 13444 3976 13456
rect 3835 13416 3976 13444
rect 3835 13413 3847 13416
rect 3789 13407 3847 13413
rect 3970 13404 3976 13416
rect 4028 13404 4034 13456
rect 4430 13404 4436 13456
rect 4488 13444 4494 13456
rect 5534 13444 5540 13456
rect 4488 13416 5540 13444
rect 4488 13404 4494 13416
rect 5534 13404 5540 13416
rect 5592 13404 5598 13456
rect 5810 13453 5816 13456
rect 5804 13444 5816 13453
rect 5771 13416 5816 13444
rect 5804 13407 5816 13416
rect 5810 13404 5816 13407
rect 5868 13404 5874 13456
rect 8389 13447 8447 13453
rect 8389 13413 8401 13447
rect 8435 13444 8447 13447
rect 8478 13444 8484 13456
rect 8435 13416 8484 13444
rect 8435 13413 8447 13416
rect 8389 13407 8447 13413
rect 8478 13404 8484 13416
rect 8536 13404 8542 13456
rect 10686 13404 10692 13456
rect 10744 13444 10750 13456
rect 10934 13447 10992 13453
rect 10934 13444 10946 13447
rect 10744 13416 10946 13444
rect 10744 13404 10750 13416
rect 10934 13413 10946 13416
rect 10980 13413 10992 13447
rect 10934 13407 10992 13413
rect 12802 13404 12808 13456
rect 12860 13444 12866 13456
rect 13725 13447 13783 13453
rect 13725 13444 13737 13447
rect 12860 13416 13737 13444
rect 12860 13404 12866 13416
rect 13725 13413 13737 13416
rect 13771 13413 13783 13447
rect 15562 13444 15568 13456
rect 15523 13416 15568 13444
rect 13725 13407 13783 13413
rect 15562 13404 15568 13416
rect 15620 13404 15626 13456
rect 16390 13404 16396 13456
rect 16448 13453 16454 13456
rect 16448 13447 16512 13453
rect 16448 13413 16466 13447
rect 16500 13413 16512 13447
rect 16448 13407 16512 13413
rect 18785 13447 18843 13453
rect 18785 13413 18797 13447
rect 18831 13444 18843 13447
rect 19334 13444 19340 13456
rect 18831 13416 19340 13444
rect 18831 13413 18843 13416
rect 18785 13407 18843 13413
rect 16448 13404 16454 13407
rect 19334 13404 19340 13416
rect 19392 13404 19398 13456
rect 19702 13404 19708 13456
rect 19760 13444 19766 13456
rect 19797 13447 19855 13453
rect 19797 13444 19809 13447
rect 19760 13416 19809 13444
rect 19760 13404 19766 13416
rect 19797 13413 19809 13416
rect 19843 13413 19855 13447
rect 22554 13444 22560 13456
rect 22515 13416 22560 13444
rect 19797 13407 19855 13413
rect 22554 13404 22560 13416
rect 22612 13404 22618 13456
rect 22649 13447 22707 13453
rect 22649 13413 22661 13447
rect 22695 13444 22707 13447
rect 22830 13444 22836 13456
rect 22695 13416 22836 13444
rect 22695 13413 22707 13416
rect 22649 13407 22707 13413
rect 22830 13404 22836 13416
rect 22888 13404 22894 13456
rect 24118 13444 24124 13456
rect 24079 13416 24124 13444
rect 24118 13404 24124 13416
rect 24176 13404 24182 13456
rect 24213 13447 24271 13453
rect 24213 13413 24225 13447
rect 24259 13444 24271 13447
rect 24854 13444 24860 13456
rect 24259 13416 24860 13444
rect 24259 13413 24271 13416
rect 24213 13407 24271 13413
rect 24854 13404 24860 13416
rect 24912 13444 24918 13456
rect 25038 13444 25044 13456
rect 24912 13416 25044 13444
rect 24912 13404 24918 13416
rect 25038 13404 25044 13416
rect 25096 13404 25102 13456
rect 4062 13376 4068 13388
rect 4023 13348 4068 13376
rect 4062 13336 4068 13348
rect 4120 13336 4126 13388
rect 11698 13376 11704 13388
rect 10704 13348 11704 13376
rect 3053 13311 3111 13317
rect 3053 13277 3065 13311
rect 3099 13308 3111 13311
rect 3234 13308 3240 13320
rect 3099 13280 3240 13308
rect 3099 13277 3111 13280
rect 3053 13271 3111 13277
rect 3234 13268 3240 13280
rect 3292 13268 3298 13320
rect 5350 13268 5356 13320
rect 5408 13308 5414 13320
rect 5537 13311 5595 13317
rect 5537 13308 5549 13311
rect 5408 13280 5549 13308
rect 5408 13268 5414 13280
rect 5537 13277 5549 13280
rect 5583 13277 5595 13311
rect 5537 13271 5595 13277
rect 8665 13311 8723 13317
rect 8665 13277 8677 13311
rect 8711 13308 8723 13311
rect 8754 13308 8760 13320
rect 8711 13280 8760 13308
rect 8711 13277 8723 13280
rect 8665 13271 8723 13277
rect 8754 13268 8760 13280
rect 8812 13308 8818 13320
rect 9490 13308 9496 13320
rect 8812 13280 9496 13308
rect 8812 13268 8818 13280
rect 9490 13268 9496 13280
rect 9548 13268 9554 13320
rect 9677 13311 9735 13317
rect 9677 13277 9689 13311
rect 9723 13308 9735 13311
rect 9858 13308 9864 13320
rect 9723 13280 9864 13308
rect 9723 13277 9735 13280
rect 9677 13271 9735 13277
rect 9858 13268 9864 13280
rect 9916 13268 9922 13320
rect 10594 13268 10600 13320
rect 10652 13308 10658 13320
rect 10704 13317 10732 13348
rect 11698 13336 11704 13348
rect 11756 13336 11762 13388
rect 12986 13336 12992 13388
rect 13044 13376 13050 13388
rect 13081 13379 13139 13385
rect 13081 13376 13093 13379
rect 13044 13348 13093 13376
rect 13044 13336 13050 13348
rect 13081 13345 13093 13348
rect 13127 13376 13139 13379
rect 13127 13348 13860 13376
rect 13127 13345 13139 13348
rect 13081 13339 13139 13345
rect 10689 13311 10747 13317
rect 10689 13308 10701 13311
rect 10652 13280 10701 13308
rect 10652 13268 10658 13280
rect 10689 13277 10701 13280
rect 10735 13277 10747 13311
rect 13722 13308 13728 13320
rect 13683 13280 13728 13308
rect 10689 13271 10747 13277
rect 13722 13268 13728 13280
rect 13780 13268 13786 13320
rect 13832 13317 13860 13348
rect 19426 13336 19432 13388
rect 19484 13376 19490 13388
rect 19889 13379 19947 13385
rect 19889 13376 19901 13379
rect 19484 13348 19901 13376
rect 19484 13336 19490 13348
rect 19889 13345 19901 13348
rect 19935 13345 19947 13379
rect 19889 13339 19947 13345
rect 22373 13379 22431 13385
rect 22373 13345 22385 13379
rect 22419 13376 22431 13379
rect 22462 13376 22468 13388
rect 22419 13348 22468 13376
rect 22419 13345 22431 13348
rect 22373 13339 22431 13345
rect 22462 13336 22468 13348
rect 22520 13376 22526 13388
rect 25133 13379 25191 13385
rect 25133 13376 25145 13379
rect 22520 13348 25145 13376
rect 22520 13336 22526 13348
rect 25133 13345 25145 13348
rect 25179 13345 25191 13379
rect 25133 13339 25191 13345
rect 13817 13311 13875 13317
rect 13817 13277 13829 13311
rect 13863 13308 13875 13311
rect 13906 13308 13912 13320
rect 13863 13280 13912 13308
rect 13863 13277 13875 13280
rect 13817 13271 13875 13277
rect 13906 13268 13912 13280
rect 13964 13268 13970 13320
rect 14274 13268 14280 13320
rect 14332 13308 14338 13320
rect 15010 13308 15016 13320
rect 14332 13280 15016 13308
rect 14332 13268 14338 13280
rect 15010 13268 15016 13280
rect 15068 13308 15074 13320
rect 15838 13308 15844 13320
rect 15068 13280 15844 13308
rect 15068 13268 15074 13280
rect 15838 13268 15844 13280
rect 15896 13308 15902 13320
rect 16022 13308 16028 13320
rect 15896 13280 16028 13308
rect 15896 13268 15902 13280
rect 16022 13268 16028 13280
rect 16080 13308 16086 13320
rect 16209 13311 16267 13317
rect 16209 13308 16221 13311
rect 16080 13280 16221 13308
rect 16080 13268 16086 13280
rect 16209 13277 16221 13280
rect 16255 13277 16267 13311
rect 16209 13271 16267 13277
rect 19058 13268 19064 13320
rect 19116 13308 19122 13320
rect 19705 13311 19763 13317
rect 19705 13308 19717 13311
rect 19116 13280 19717 13308
rect 19116 13268 19122 13280
rect 19705 13277 19717 13280
rect 19751 13277 19763 13311
rect 24029 13311 24087 13317
rect 24029 13308 24041 13311
rect 19705 13271 19763 13277
rect 23032 13280 24041 13308
rect 2501 13243 2559 13249
rect 2501 13209 2513 13243
rect 2547 13240 2559 13243
rect 4522 13240 4528 13252
rect 2547 13212 4528 13240
rect 2547 13209 2559 13212
rect 2501 13203 2559 13209
rect 4522 13200 4528 13212
rect 4580 13200 4586 13252
rect 4706 13240 4712 13252
rect 4667 13212 4712 13240
rect 4706 13200 4712 13212
rect 4764 13200 4770 13252
rect 8113 13243 8171 13249
rect 8113 13209 8125 13243
rect 8159 13240 8171 13243
rect 8202 13240 8208 13252
rect 8159 13212 8208 13240
rect 8159 13209 8171 13212
rect 8113 13203 8171 13209
rect 8202 13200 8208 13212
rect 8260 13200 8266 13252
rect 12526 13200 12532 13252
rect 12584 13240 12590 13252
rect 13265 13243 13323 13249
rect 13265 13240 13277 13243
rect 12584 13212 13277 13240
rect 12584 13200 12590 13212
rect 13265 13209 13277 13212
rect 13311 13209 13323 13243
rect 13265 13203 13323 13209
rect 22097 13243 22155 13249
rect 22097 13209 22109 13243
rect 22143 13240 22155 13243
rect 23032 13240 23060 13280
rect 24029 13277 24041 13280
rect 24075 13308 24087 13311
rect 25038 13308 25044 13320
rect 24075 13280 25044 13308
rect 24075 13277 24087 13280
rect 24029 13271 24087 13277
rect 25038 13268 25044 13280
rect 25096 13268 25102 13320
rect 22143 13212 23060 13240
rect 23109 13243 23167 13249
rect 22143 13209 22155 13212
rect 22097 13203 22155 13209
rect 23109 13209 23121 13243
rect 23155 13240 23167 13243
rect 23658 13240 23664 13252
rect 23155 13212 23664 13240
rect 23155 13209 23167 13212
rect 23109 13203 23167 13209
rect 23658 13200 23664 13212
rect 23716 13200 23722 13252
rect 1946 13172 1952 13184
rect 1907 13144 1952 13172
rect 1946 13132 1952 13144
rect 2004 13132 2010 13184
rect 3970 13132 3976 13184
rect 4028 13172 4034 13184
rect 4249 13175 4307 13181
rect 4249 13172 4261 13175
rect 4028 13144 4261 13172
rect 4028 13132 4034 13144
rect 4249 13141 4261 13144
rect 4295 13141 4307 13175
rect 4249 13135 4307 13141
rect 9217 13175 9275 13181
rect 9217 13141 9229 13175
rect 9263 13172 9275 13175
rect 9582 13172 9588 13184
rect 9263 13144 9588 13172
rect 9263 13141 9275 13144
rect 9217 13135 9275 13141
rect 9582 13132 9588 13144
rect 9640 13132 9646 13184
rect 10134 13172 10140 13184
rect 10095 13144 10140 13172
rect 10134 13132 10140 13144
rect 10192 13132 10198 13184
rect 17586 13172 17592 13184
rect 17547 13144 17592 13172
rect 17586 13132 17592 13144
rect 17644 13132 17650 13184
rect 19337 13175 19395 13181
rect 19337 13141 19349 13175
rect 19383 13172 19395 13175
rect 19794 13172 19800 13184
rect 19383 13144 19800 13172
rect 19383 13141 19395 13144
rect 19337 13135 19395 13141
rect 19794 13132 19800 13144
rect 19852 13132 19858 13184
rect 21450 13172 21456 13184
rect 21411 13144 21456 13172
rect 21450 13132 21456 13144
rect 21508 13132 21514 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1673 12971 1731 12977
rect 1673 12937 1685 12971
rect 1719 12968 1731 12971
rect 2866 12968 2872 12980
rect 1719 12940 2872 12968
rect 1719 12937 1731 12940
rect 1673 12931 1731 12937
rect 2866 12928 2872 12940
rect 2924 12928 2930 12980
rect 3326 12928 3332 12980
rect 3384 12968 3390 12980
rect 3513 12971 3571 12977
rect 3513 12968 3525 12971
rect 3384 12940 3525 12968
rect 3384 12928 3390 12940
rect 3513 12937 3525 12940
rect 3559 12937 3571 12971
rect 3513 12931 3571 12937
rect 4154 12928 4160 12980
rect 4212 12968 4218 12980
rect 4709 12971 4767 12977
rect 4709 12968 4721 12971
rect 4212 12940 4721 12968
rect 4212 12928 4218 12940
rect 4709 12937 4721 12940
rect 4755 12937 4767 12971
rect 5994 12968 6000 12980
rect 5955 12940 6000 12968
rect 4709 12931 4767 12937
rect 5994 12928 6000 12940
rect 6052 12928 6058 12980
rect 12802 12928 12808 12980
rect 12860 12968 12866 12980
rect 13081 12971 13139 12977
rect 13081 12968 13093 12971
rect 12860 12940 13093 12968
rect 12860 12928 12866 12940
rect 13081 12937 13093 12940
rect 13127 12937 13139 12971
rect 13354 12968 13360 12980
rect 13315 12940 13360 12968
rect 13081 12931 13139 12937
rect 13354 12928 13360 12940
rect 13412 12928 13418 12980
rect 14369 12971 14427 12977
rect 14369 12937 14381 12971
rect 14415 12968 14427 12971
rect 14550 12968 14556 12980
rect 14415 12940 14556 12968
rect 14415 12937 14427 12940
rect 14369 12931 14427 12937
rect 2038 12900 2044 12912
rect 1999 12872 2044 12900
rect 2038 12860 2044 12872
rect 2096 12860 2102 12912
rect 6822 12860 6828 12912
rect 6880 12900 6886 12912
rect 7009 12903 7067 12909
rect 7009 12900 7021 12903
rect 6880 12872 7021 12900
rect 6880 12860 6886 12872
rect 7009 12869 7021 12872
rect 7055 12869 7067 12903
rect 8018 12900 8024 12912
rect 7979 12872 8024 12900
rect 7009 12863 7067 12869
rect 8018 12860 8024 12872
rect 8076 12860 8082 12912
rect 14384 12900 14412 12931
rect 14550 12928 14556 12940
rect 14608 12928 14614 12980
rect 15381 12971 15439 12977
rect 15381 12937 15393 12971
rect 15427 12968 15439 12971
rect 16390 12968 16396 12980
rect 15427 12940 16396 12968
rect 15427 12937 15439 12940
rect 15381 12931 15439 12937
rect 16390 12928 16396 12940
rect 16448 12928 16454 12980
rect 16942 12928 16948 12980
rect 17000 12968 17006 12980
rect 17221 12971 17279 12977
rect 17221 12968 17233 12971
rect 17000 12940 17233 12968
rect 17000 12928 17006 12940
rect 17221 12937 17233 12940
rect 17267 12937 17279 12971
rect 17221 12931 17279 12937
rect 18969 12971 19027 12977
rect 18969 12937 18981 12971
rect 19015 12968 19027 12971
rect 19058 12968 19064 12980
rect 19015 12940 19064 12968
rect 19015 12937 19027 12940
rect 18969 12931 19027 12937
rect 19058 12928 19064 12940
rect 19116 12928 19122 12980
rect 19334 12968 19340 12980
rect 19295 12940 19340 12968
rect 19334 12928 19340 12940
rect 19392 12968 19398 12980
rect 19702 12968 19708 12980
rect 19392 12940 19708 12968
rect 19392 12928 19398 12940
rect 19702 12928 19708 12940
rect 19760 12928 19766 12980
rect 22097 12971 22155 12977
rect 22097 12937 22109 12971
rect 22143 12968 22155 12971
rect 22186 12968 22192 12980
rect 22143 12940 22192 12968
rect 22143 12937 22155 12940
rect 22097 12931 22155 12937
rect 22186 12928 22192 12940
rect 22244 12968 22250 12980
rect 22554 12968 22560 12980
rect 22244 12940 22560 12968
rect 22244 12928 22250 12940
rect 22554 12928 22560 12940
rect 22612 12928 22618 12980
rect 22830 12968 22836 12980
rect 22791 12940 22836 12968
rect 22830 12928 22836 12940
rect 22888 12928 22894 12980
rect 24118 12928 24124 12980
rect 24176 12968 24182 12980
rect 24673 12971 24731 12977
rect 24673 12968 24685 12971
rect 24176 12940 24685 12968
rect 24176 12928 24182 12940
rect 24673 12937 24685 12940
rect 24719 12937 24731 12971
rect 25038 12968 25044 12980
rect 24999 12940 25044 12968
rect 24673 12931 24731 12937
rect 25038 12928 25044 12940
rect 25096 12928 25102 12980
rect 16022 12900 16028 12912
rect 13740 12872 14412 12900
rect 15983 12872 16028 12900
rect 4062 12792 4068 12844
rect 4120 12832 4126 12844
rect 4157 12835 4215 12841
rect 4157 12832 4169 12835
rect 4120 12804 4169 12832
rect 4120 12792 4126 12804
rect 4157 12801 4169 12804
rect 4203 12832 4215 12835
rect 4525 12835 4583 12841
rect 4525 12832 4537 12835
rect 4203 12804 4537 12832
rect 4203 12801 4215 12804
rect 4157 12795 4215 12801
rect 4525 12801 4537 12804
rect 4571 12832 4583 12835
rect 5166 12832 5172 12844
rect 4571 12804 5172 12832
rect 4571 12801 4583 12804
rect 4525 12795 4583 12801
rect 5166 12792 5172 12804
rect 5224 12792 5230 12844
rect 5261 12835 5319 12841
rect 5261 12801 5273 12835
rect 5307 12832 5319 12835
rect 5442 12832 5448 12844
rect 5307 12804 5448 12832
rect 5307 12801 5319 12804
rect 5261 12795 5319 12801
rect 5442 12792 5448 12804
rect 5500 12792 5506 12844
rect 7466 12832 7472 12844
rect 7427 12804 7472 12832
rect 7466 12792 7472 12804
rect 7524 12792 7530 12844
rect 8294 12792 8300 12844
rect 8352 12832 8358 12844
rect 13740 12841 13768 12872
rect 16022 12860 16028 12872
rect 16080 12860 16086 12912
rect 16301 12903 16359 12909
rect 16301 12869 16313 12903
rect 16347 12900 16359 12903
rect 16482 12900 16488 12912
rect 16347 12872 16488 12900
rect 16347 12869 16359 12872
rect 16301 12863 16359 12869
rect 16482 12860 16488 12872
rect 16540 12860 16546 12912
rect 8481 12835 8539 12841
rect 8481 12832 8493 12835
rect 8352 12804 8493 12832
rect 8352 12792 8358 12804
rect 8481 12801 8493 12804
rect 8527 12801 8539 12835
rect 8481 12795 8539 12801
rect 13725 12835 13783 12841
rect 13725 12801 13737 12835
rect 13771 12801 13783 12835
rect 13906 12832 13912 12844
rect 13819 12804 13912 12832
rect 13725 12795 13783 12801
rect 13906 12792 13912 12804
rect 13964 12832 13970 12844
rect 14645 12835 14703 12841
rect 14645 12832 14657 12835
rect 13964 12804 14657 12832
rect 13964 12792 13970 12804
rect 14645 12801 14657 12804
rect 14691 12801 14703 12835
rect 14645 12795 14703 12801
rect 16761 12835 16819 12841
rect 16761 12801 16773 12835
rect 16807 12832 16819 12835
rect 16960 12832 16988 12928
rect 19518 12900 19524 12912
rect 19479 12872 19524 12900
rect 19518 12860 19524 12872
rect 19576 12860 19582 12912
rect 21082 12900 21088 12912
rect 21043 12872 21088 12900
rect 21082 12860 21088 12872
rect 21140 12860 21146 12912
rect 22462 12900 22468 12912
rect 22423 12872 22468 12900
rect 22462 12860 22468 12872
rect 22520 12860 22526 12912
rect 23753 12903 23811 12909
rect 23753 12900 23765 12903
rect 23400 12872 23765 12900
rect 21450 12832 21456 12844
rect 16807 12804 16988 12832
rect 20088 12804 21456 12832
rect 16807 12801 16819 12804
rect 16761 12795 16819 12801
rect 2130 12764 2136 12776
rect 2091 12736 2136 12764
rect 2130 12724 2136 12736
rect 2188 12724 2194 12776
rect 9401 12767 9459 12773
rect 9401 12764 9413 12767
rect 6104 12736 9413 12764
rect 2400 12699 2458 12705
rect 2400 12665 2412 12699
rect 2446 12696 2458 12699
rect 3878 12696 3884 12708
rect 2446 12668 3884 12696
rect 2446 12665 2458 12668
rect 2400 12659 2458 12665
rect 3878 12656 3884 12668
rect 3936 12656 3942 12708
rect 4062 12656 4068 12708
rect 4120 12696 4126 12708
rect 4706 12696 4712 12708
rect 4120 12668 4712 12696
rect 4120 12656 4126 12668
rect 4706 12656 4712 12668
rect 4764 12696 4770 12708
rect 5169 12699 5227 12705
rect 5169 12696 5181 12699
rect 4764 12668 5181 12696
rect 4764 12656 4770 12668
rect 5169 12665 5181 12668
rect 5215 12665 5227 12699
rect 5169 12659 5227 12665
rect 6104 12640 6132 12736
rect 9401 12733 9413 12736
rect 9447 12764 9459 12767
rect 9585 12767 9643 12773
rect 9585 12764 9597 12767
rect 9447 12736 9597 12764
rect 9447 12733 9459 12736
rect 9401 12727 9459 12733
rect 9585 12733 9597 12736
rect 9631 12764 9643 12767
rect 10594 12764 10600 12776
rect 9631 12736 10600 12764
rect 9631 12733 9643 12736
rect 9585 12727 9643 12733
rect 10594 12724 10600 12736
rect 10652 12724 10658 12776
rect 10778 12724 10784 12776
rect 10836 12764 10842 12776
rect 15749 12767 15807 12773
rect 10836 12736 12848 12764
rect 10836 12724 10842 12736
rect 6641 12699 6699 12705
rect 6641 12665 6653 12699
rect 6687 12696 6699 12699
rect 7561 12699 7619 12705
rect 7561 12696 7573 12699
rect 6687 12668 7573 12696
rect 6687 12665 6699 12668
rect 6641 12659 6699 12665
rect 7561 12665 7573 12668
rect 7607 12696 7619 12699
rect 8294 12696 8300 12708
rect 7607 12668 8300 12696
rect 7607 12665 7619 12668
rect 7561 12659 7619 12665
rect 8294 12656 8300 12668
rect 8352 12656 8358 12708
rect 9125 12699 9183 12705
rect 9125 12665 9137 12699
rect 9171 12696 9183 12699
rect 9852 12699 9910 12705
rect 9852 12696 9864 12699
rect 9171 12668 9864 12696
rect 9171 12665 9183 12668
rect 9125 12659 9183 12665
rect 9852 12665 9864 12668
rect 9898 12696 9910 12699
rect 10870 12696 10876 12708
rect 9898 12668 10876 12696
rect 9898 12665 9910 12668
rect 9852 12659 9910 12665
rect 10870 12656 10876 12668
rect 10928 12656 10934 12708
rect 12820 12705 12848 12736
rect 15749 12733 15761 12767
rect 15795 12764 15807 12767
rect 16853 12767 16911 12773
rect 16853 12764 16865 12767
rect 15795 12736 16865 12764
rect 15795 12733 15807 12736
rect 15749 12727 15807 12733
rect 16853 12733 16865 12736
rect 16899 12764 16911 12767
rect 17586 12764 17592 12776
rect 16899 12736 17592 12764
rect 16899 12733 16911 12736
rect 16853 12727 16911 12733
rect 17586 12724 17592 12736
rect 17644 12724 17650 12776
rect 19794 12764 19800 12776
rect 19755 12736 19800 12764
rect 19794 12724 19800 12736
rect 19852 12724 19858 12776
rect 20088 12708 20116 12804
rect 21450 12792 21456 12804
rect 21508 12832 21514 12844
rect 21637 12835 21695 12841
rect 21637 12832 21649 12835
rect 21508 12804 21649 12832
rect 21508 12792 21514 12804
rect 21637 12801 21649 12804
rect 21683 12832 21695 12835
rect 22002 12832 22008 12844
rect 21683 12804 22008 12832
rect 21683 12801 21695 12804
rect 21637 12795 21695 12801
rect 22002 12792 22008 12804
rect 22060 12792 22066 12844
rect 22094 12764 22100 12776
rect 21376 12736 22100 12764
rect 12805 12699 12863 12705
rect 12805 12665 12817 12699
rect 12851 12696 12863 12699
rect 13817 12699 13875 12705
rect 13817 12696 13829 12699
rect 12851 12668 13829 12696
rect 12851 12665 12863 12668
rect 12805 12659 12863 12665
rect 13817 12665 13829 12668
rect 13863 12696 13875 12699
rect 13998 12696 14004 12708
rect 13863 12668 14004 12696
rect 13863 12665 13875 12668
rect 13817 12659 13875 12665
rect 13998 12656 14004 12668
rect 14056 12656 14062 12708
rect 16758 12696 16764 12708
rect 16719 12668 16764 12696
rect 16758 12656 16764 12668
rect 16816 12656 16822 12708
rect 18598 12696 18604 12708
rect 18511 12668 18604 12696
rect 18598 12656 18604 12668
rect 18656 12696 18662 12708
rect 19981 12699 20039 12705
rect 19981 12696 19993 12699
rect 18656 12668 19993 12696
rect 18656 12656 18662 12668
rect 19981 12665 19993 12668
rect 20027 12665 20039 12699
rect 19981 12659 20039 12665
rect 20070 12656 20076 12708
rect 20128 12696 20134 12708
rect 21376 12705 21404 12736
rect 22094 12724 22100 12736
rect 22152 12724 22158 12776
rect 22646 12724 22652 12776
rect 22704 12764 22710 12776
rect 23106 12764 23112 12776
rect 22704 12736 23112 12764
rect 22704 12724 22710 12736
rect 23106 12724 23112 12736
rect 23164 12724 23170 12776
rect 20533 12699 20591 12705
rect 20128 12668 20173 12696
rect 20128 12656 20134 12668
rect 20533 12665 20545 12699
rect 20579 12696 20591 12699
rect 21361 12699 21419 12705
rect 21361 12696 21373 12699
rect 20579 12668 21373 12696
rect 20579 12665 20591 12668
rect 20533 12659 20591 12665
rect 21361 12665 21373 12668
rect 21407 12665 21419 12699
rect 21542 12696 21548 12708
rect 21503 12668 21548 12696
rect 21361 12659 21419 12665
rect 21542 12656 21548 12668
rect 21600 12656 21606 12708
rect 5350 12588 5356 12640
rect 5408 12628 5414 12640
rect 5721 12631 5779 12637
rect 5721 12628 5733 12631
rect 5408 12600 5733 12628
rect 5408 12588 5414 12600
rect 5721 12597 5733 12600
rect 5767 12628 5779 12631
rect 6086 12628 6092 12640
rect 5767 12600 6092 12628
rect 5767 12597 5779 12600
rect 5721 12591 5779 12597
rect 6086 12588 6092 12600
rect 6144 12588 6150 12640
rect 7006 12588 7012 12640
rect 7064 12628 7070 12640
rect 7469 12631 7527 12637
rect 7469 12628 7481 12631
rect 7064 12600 7481 12628
rect 7064 12588 7070 12600
rect 7469 12597 7481 12600
rect 7515 12597 7527 12631
rect 7469 12591 7527 12597
rect 7742 12588 7748 12640
rect 7800 12628 7806 12640
rect 8662 12628 8668 12640
rect 7800 12600 8668 12628
rect 7800 12588 7806 12600
rect 8662 12588 8668 12600
rect 8720 12588 8726 12640
rect 10686 12588 10692 12640
rect 10744 12628 10750 12640
rect 10965 12631 11023 12637
rect 10965 12628 10977 12631
rect 10744 12600 10977 12628
rect 10744 12588 10750 12600
rect 10965 12597 10977 12600
rect 11011 12597 11023 12631
rect 10965 12591 11023 12597
rect 11609 12631 11667 12637
rect 11609 12597 11621 12631
rect 11655 12628 11667 12631
rect 11698 12628 11704 12640
rect 11655 12600 11704 12628
rect 11655 12597 11667 12600
rect 11609 12591 11667 12597
rect 11698 12588 11704 12600
rect 11756 12588 11762 12640
rect 20806 12588 20812 12640
rect 20864 12628 20870 12640
rect 20901 12631 20959 12637
rect 20901 12628 20913 12631
rect 20864 12600 20913 12628
rect 20864 12588 20870 12600
rect 20901 12597 20913 12600
rect 20947 12628 20959 12631
rect 21560 12628 21588 12656
rect 23400 12640 23428 12872
rect 23753 12869 23765 12872
rect 23799 12869 23811 12903
rect 23753 12863 23811 12869
rect 23658 12724 23664 12776
rect 23716 12764 23722 12776
rect 24029 12767 24087 12773
rect 24029 12764 24041 12767
rect 23716 12736 24041 12764
rect 23716 12724 23722 12736
rect 24029 12733 24041 12736
rect 24075 12733 24087 12767
rect 24029 12727 24087 12733
rect 24210 12724 24216 12776
rect 24268 12724 24274 12776
rect 24670 12724 24676 12776
rect 24728 12764 24734 12776
rect 25225 12767 25283 12773
rect 25225 12764 25237 12767
rect 24728 12736 25237 12764
rect 24728 12724 24734 12736
rect 25225 12733 25237 12736
rect 25271 12764 25283 12767
rect 25777 12767 25835 12773
rect 25777 12764 25789 12767
rect 25271 12736 25789 12764
rect 25271 12733 25283 12736
rect 25225 12727 25283 12733
rect 25777 12733 25789 12736
rect 25823 12733 25835 12767
rect 25777 12727 25835 12733
rect 23477 12699 23535 12705
rect 23477 12665 23489 12699
rect 23523 12696 23535 12699
rect 24228 12696 24256 12724
rect 24305 12699 24363 12705
rect 24305 12696 24317 12699
rect 23523 12668 24317 12696
rect 23523 12665 23535 12668
rect 23477 12659 23535 12665
rect 24305 12665 24317 12668
rect 24351 12665 24363 12699
rect 24305 12659 24363 12665
rect 20947 12600 21588 12628
rect 20947 12597 20959 12600
rect 20901 12591 20959 12597
rect 23382 12588 23388 12640
rect 23440 12588 23446 12640
rect 23750 12588 23756 12640
rect 23808 12628 23814 12640
rect 24213 12631 24271 12637
rect 24213 12628 24225 12631
rect 23808 12600 24225 12628
rect 23808 12588 23814 12600
rect 24213 12597 24225 12600
rect 24259 12597 24271 12631
rect 25406 12628 25412 12640
rect 25367 12600 25412 12628
rect 24213 12591 24271 12597
rect 25406 12588 25412 12600
rect 25464 12588 25470 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 2961 12427 3019 12433
rect 2961 12424 2973 12427
rect 2832 12396 2973 12424
rect 2832 12384 2838 12396
rect 2961 12393 2973 12396
rect 3007 12393 3019 12427
rect 2961 12387 3019 12393
rect 3234 12384 3240 12436
rect 3292 12424 3298 12436
rect 3421 12427 3479 12433
rect 3421 12424 3433 12427
rect 3292 12396 3433 12424
rect 3292 12384 3298 12396
rect 3421 12393 3433 12396
rect 3467 12393 3479 12427
rect 8478 12424 8484 12436
rect 8439 12396 8484 12424
rect 3421 12387 3479 12393
rect 8478 12384 8484 12396
rect 8536 12384 8542 12436
rect 8754 12424 8760 12436
rect 8715 12396 8760 12424
rect 8754 12384 8760 12396
rect 8812 12384 8818 12436
rect 11149 12427 11207 12433
rect 11149 12393 11161 12427
rect 11195 12424 11207 12427
rect 11238 12424 11244 12436
rect 11195 12396 11244 12424
rect 11195 12393 11207 12396
rect 11149 12387 11207 12393
rect 11238 12384 11244 12396
rect 11296 12384 11302 12436
rect 13814 12424 13820 12436
rect 13775 12396 13820 12424
rect 13814 12384 13820 12396
rect 13872 12384 13878 12436
rect 16758 12424 16764 12436
rect 16719 12396 16764 12424
rect 16758 12384 16764 12396
rect 16816 12384 16822 12436
rect 19978 12424 19984 12436
rect 19939 12396 19984 12424
rect 19978 12384 19984 12396
rect 20036 12384 20042 12436
rect 22094 12384 22100 12436
rect 22152 12424 22158 12436
rect 22281 12427 22339 12433
rect 22281 12424 22293 12427
rect 22152 12396 22293 12424
rect 22152 12384 22158 12396
rect 22281 12393 22293 12396
rect 22327 12393 22339 12427
rect 22281 12387 22339 12393
rect 23293 12427 23351 12433
rect 23293 12393 23305 12427
rect 23339 12424 23351 12427
rect 23750 12424 23756 12436
rect 23339 12396 23756 12424
rect 23339 12393 23351 12396
rect 23293 12387 23351 12393
rect 23750 12384 23756 12396
rect 23808 12384 23814 12436
rect 23934 12384 23940 12436
rect 23992 12424 23998 12436
rect 24670 12424 24676 12436
rect 23992 12396 24676 12424
rect 23992 12384 23998 12396
rect 24670 12384 24676 12396
rect 24728 12384 24734 12436
rect 3050 12356 3056 12368
rect 2963 12328 3056 12356
rect 3050 12316 3056 12328
rect 3108 12356 3114 12368
rect 3326 12356 3332 12368
rect 3108 12328 3332 12356
rect 3108 12316 3114 12328
rect 3326 12316 3332 12328
rect 3384 12316 3390 12368
rect 7282 12316 7288 12368
rect 7340 12356 7346 12368
rect 7929 12359 7987 12365
rect 7929 12356 7941 12359
rect 7340 12328 7941 12356
rect 7340 12316 7346 12328
rect 7929 12325 7941 12328
rect 7975 12325 7987 12359
rect 7929 12319 7987 12325
rect 8938 12316 8944 12368
rect 8996 12356 9002 12368
rect 10229 12359 10287 12365
rect 10229 12356 10241 12359
rect 8996 12328 10241 12356
rect 8996 12316 9002 12328
rect 10229 12325 10241 12328
rect 10275 12325 10287 12359
rect 10229 12319 10287 12325
rect 14366 12316 14372 12368
rect 14424 12356 14430 12368
rect 16206 12356 16212 12368
rect 14424 12328 16212 12356
rect 14424 12316 14430 12328
rect 16206 12316 16212 12328
rect 16264 12316 16270 12368
rect 17488 12359 17546 12365
rect 17488 12325 17500 12359
rect 17534 12356 17546 12359
rect 17586 12356 17592 12368
rect 17534 12328 17592 12356
rect 17534 12325 17546 12328
rect 17488 12319 17546 12325
rect 17586 12316 17592 12328
rect 17644 12316 17650 12368
rect 23106 12316 23112 12368
rect 23164 12356 23170 12368
rect 23661 12359 23719 12365
rect 23661 12356 23673 12359
rect 23164 12328 23673 12356
rect 23164 12316 23170 12328
rect 23661 12325 23673 12328
rect 23707 12356 23719 12359
rect 24112 12359 24170 12365
rect 24112 12356 24124 12359
rect 23707 12328 24124 12356
rect 23707 12325 23719 12328
rect 23661 12319 23719 12325
rect 24112 12325 24124 12328
rect 24158 12356 24170 12359
rect 24854 12356 24860 12368
rect 24158 12328 24860 12356
rect 24158 12325 24170 12328
rect 24112 12319 24170 12325
rect 24854 12316 24860 12328
rect 24912 12316 24918 12368
rect 2130 12248 2136 12300
rect 2188 12288 2194 12300
rect 2225 12291 2283 12297
rect 2225 12288 2237 12291
rect 2188 12260 2237 12288
rect 2188 12248 2194 12260
rect 2225 12257 2237 12260
rect 2271 12288 2283 12291
rect 4065 12291 4123 12297
rect 4065 12288 4077 12291
rect 2271 12260 4077 12288
rect 2271 12257 2283 12260
rect 2225 12251 2283 12257
rect 4065 12257 4077 12260
rect 4111 12257 4123 12291
rect 4065 12251 4123 12257
rect 4332 12291 4390 12297
rect 4332 12257 4344 12291
rect 4378 12288 4390 12291
rect 5442 12288 5448 12300
rect 4378 12260 5448 12288
rect 4378 12257 4390 12260
rect 4332 12251 4390 12257
rect 5442 12248 5448 12260
rect 5500 12248 5506 12300
rect 7374 12248 7380 12300
rect 7432 12288 7438 12300
rect 7742 12288 7748 12300
rect 7432 12260 7748 12288
rect 7432 12248 7438 12260
rect 7742 12248 7748 12260
rect 7800 12248 7806 12300
rect 10042 12288 10048 12300
rect 10003 12260 10048 12288
rect 10042 12248 10048 12260
rect 10100 12248 10106 12300
rect 12158 12297 12164 12300
rect 12152 12288 12164 12297
rect 12071 12260 12164 12288
rect 12152 12251 12164 12260
rect 12216 12288 12222 12300
rect 15654 12288 15660 12300
rect 12216 12260 15660 12288
rect 12158 12248 12164 12251
rect 12216 12248 12222 12260
rect 15654 12248 15660 12260
rect 15712 12248 15718 12300
rect 19337 12291 19395 12297
rect 19337 12257 19349 12291
rect 19383 12288 19395 12291
rect 19426 12288 19432 12300
rect 19383 12260 19432 12288
rect 19383 12257 19395 12260
rect 19337 12251 19395 12257
rect 19426 12248 19432 12260
rect 19484 12288 19490 12300
rect 21174 12297 21180 12300
rect 21168 12288 21180 12297
rect 19484 12260 21180 12288
rect 19484 12248 19490 12260
rect 21168 12251 21180 12260
rect 21174 12248 21180 12251
rect 21232 12248 21238 12300
rect 1394 12220 1400 12232
rect 1355 12192 1400 12220
rect 1394 12180 1400 12192
rect 1452 12180 1458 12232
rect 2961 12223 3019 12229
rect 2961 12189 2973 12223
rect 3007 12189 3019 12223
rect 5994 12220 6000 12232
rect 5955 12192 6000 12220
rect 2961 12183 3019 12189
rect 2976 12152 3004 12183
rect 5994 12180 6000 12192
rect 6052 12180 6058 12232
rect 7466 12180 7472 12232
rect 7524 12180 7530 12232
rect 8018 12220 8024 12232
rect 7979 12192 8024 12220
rect 8018 12180 8024 12192
rect 8076 12180 8082 12232
rect 9674 12180 9680 12232
rect 9732 12220 9738 12232
rect 9858 12220 9864 12232
rect 9732 12192 9864 12220
rect 9732 12180 9738 12192
rect 9858 12180 9864 12192
rect 9916 12180 9922 12232
rect 10318 12220 10324 12232
rect 10279 12192 10324 12220
rect 10318 12180 10324 12192
rect 10376 12180 10382 12232
rect 11885 12223 11943 12229
rect 11885 12220 11897 12223
rect 11716 12192 11897 12220
rect 3326 12152 3332 12164
rect 2976 12124 3332 12152
rect 3326 12112 3332 12124
rect 3384 12112 3390 12164
rect 6641 12155 6699 12161
rect 6641 12121 6653 12155
rect 6687 12152 6699 12155
rect 7484 12152 7512 12180
rect 7650 12152 7656 12164
rect 6687 12124 7656 12152
rect 6687 12121 6699 12124
rect 6641 12115 6699 12121
rect 7650 12112 7656 12124
rect 7708 12112 7714 12164
rect 11716 12096 11744 12192
rect 11885 12189 11897 12192
rect 11931 12189 11943 12223
rect 16114 12220 16120 12232
rect 16075 12192 16120 12220
rect 11885 12183 11943 12189
rect 16114 12180 16120 12192
rect 16172 12180 16178 12232
rect 16298 12220 16304 12232
rect 16259 12192 16304 12220
rect 16298 12180 16304 12192
rect 16356 12180 16362 12232
rect 17218 12220 17224 12232
rect 17179 12192 17224 12220
rect 17218 12180 17224 12192
rect 17276 12180 17282 12232
rect 20898 12220 20904 12232
rect 20811 12192 20904 12220
rect 20898 12180 20904 12192
rect 20956 12180 20962 12232
rect 23842 12220 23848 12232
rect 23803 12192 23848 12220
rect 23842 12180 23848 12192
rect 23900 12180 23906 12232
rect 13262 12152 13268 12164
rect 13223 12124 13268 12152
rect 13262 12112 13268 12124
rect 13320 12112 13326 12164
rect 2406 12044 2412 12096
rect 2464 12084 2470 12096
rect 2501 12087 2559 12093
rect 2501 12084 2513 12087
rect 2464 12056 2513 12084
rect 2464 12044 2470 12056
rect 2501 12053 2513 12056
rect 2547 12053 2559 12087
rect 3878 12084 3884 12096
rect 3791 12056 3884 12084
rect 2501 12047 2559 12053
rect 3878 12044 3884 12056
rect 3936 12084 3942 12096
rect 5445 12087 5503 12093
rect 5445 12084 5457 12087
rect 3936 12056 5457 12084
rect 3936 12044 3942 12056
rect 5445 12053 5457 12056
rect 5491 12053 5503 12087
rect 7006 12084 7012 12096
rect 6967 12056 7012 12084
rect 5445 12047 5503 12053
rect 7006 12044 7012 12056
rect 7064 12044 7070 12096
rect 7466 12084 7472 12096
rect 7427 12056 7472 12084
rect 7466 12044 7472 12056
rect 7524 12044 7530 12096
rect 8294 12044 8300 12096
rect 8352 12084 8358 12096
rect 9122 12084 9128 12096
rect 8352 12056 9128 12084
rect 8352 12044 8358 12056
rect 9122 12044 9128 12056
rect 9180 12044 9186 12096
rect 9674 12044 9680 12096
rect 9732 12084 9738 12096
rect 9769 12087 9827 12093
rect 9769 12084 9781 12087
rect 9732 12056 9781 12084
rect 9732 12044 9738 12056
rect 9769 12053 9781 12056
rect 9815 12053 9827 12087
rect 10686 12084 10692 12096
rect 10647 12056 10692 12084
rect 9769 12047 9827 12053
rect 10686 12044 10692 12056
rect 10744 12044 10750 12096
rect 11698 12084 11704 12096
rect 11659 12056 11704 12084
rect 11698 12044 11704 12056
rect 11756 12044 11762 12096
rect 15746 12084 15752 12096
rect 15707 12056 15752 12084
rect 15746 12044 15752 12056
rect 15804 12044 15810 12096
rect 17954 12044 17960 12096
rect 18012 12084 18018 12096
rect 18601 12087 18659 12093
rect 18601 12084 18613 12087
rect 18012 12056 18613 12084
rect 18012 12044 18018 12056
rect 18601 12053 18613 12056
rect 18647 12053 18659 12087
rect 18601 12047 18659 12053
rect 19705 12087 19763 12093
rect 19705 12053 19717 12087
rect 19751 12084 19763 12087
rect 20070 12084 20076 12096
rect 19751 12056 20076 12084
rect 19751 12053 19763 12056
rect 19705 12047 19763 12053
rect 20070 12044 20076 12056
rect 20128 12044 20134 12096
rect 20916 12084 20944 12180
rect 21818 12084 21824 12096
rect 20916 12056 21824 12084
rect 21818 12044 21824 12056
rect 21876 12044 21882 12096
rect 25222 12084 25228 12096
rect 25183 12056 25228 12084
rect 25222 12044 25228 12056
rect 25280 12044 25286 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 2777 11883 2835 11889
rect 2777 11849 2789 11883
rect 2823 11880 2835 11883
rect 3050 11880 3056 11892
rect 2823 11852 3056 11880
rect 2823 11849 2835 11852
rect 2777 11843 2835 11849
rect 3050 11840 3056 11852
rect 3108 11840 3114 11892
rect 3326 11880 3332 11892
rect 3287 11852 3332 11880
rect 3326 11840 3332 11852
rect 3384 11840 3390 11892
rect 5905 11883 5963 11889
rect 5905 11849 5917 11883
rect 5951 11880 5963 11883
rect 6086 11880 6092 11892
rect 5951 11852 6092 11880
rect 5951 11849 5963 11852
rect 5905 11843 5963 11849
rect 6086 11840 6092 11852
rect 6144 11840 6150 11892
rect 6273 11883 6331 11889
rect 6273 11849 6285 11883
rect 6319 11880 6331 11883
rect 6454 11880 6460 11892
rect 6319 11852 6460 11880
rect 6319 11849 6331 11852
rect 6273 11843 6331 11849
rect 6454 11840 6460 11852
rect 6512 11880 6518 11892
rect 6822 11880 6828 11892
rect 6512 11852 6828 11880
rect 6512 11840 6518 11852
rect 6822 11840 6828 11852
rect 6880 11840 6886 11892
rect 7282 11840 7288 11892
rect 7340 11880 7346 11892
rect 7377 11883 7435 11889
rect 7377 11880 7389 11883
rect 7340 11852 7389 11880
rect 7340 11840 7346 11852
rect 7377 11849 7389 11852
rect 7423 11849 7435 11883
rect 7650 11880 7656 11892
rect 7611 11852 7656 11880
rect 7377 11843 7435 11849
rect 7650 11840 7656 11852
rect 7708 11840 7714 11892
rect 11790 11880 11796 11892
rect 11751 11852 11796 11880
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 15654 11880 15660 11892
rect 15615 11852 15660 11880
rect 15654 11840 15660 11852
rect 15712 11840 15718 11892
rect 16206 11880 16212 11892
rect 16167 11852 16212 11880
rect 16206 11840 16212 11852
rect 16264 11840 16270 11892
rect 17586 11880 17592 11892
rect 17547 11852 17592 11880
rect 17586 11840 17592 11852
rect 17644 11840 17650 11892
rect 18598 11840 18604 11892
rect 18656 11880 18662 11892
rect 18877 11883 18935 11889
rect 18877 11880 18889 11883
rect 18656 11852 18889 11880
rect 18656 11840 18662 11852
rect 18877 11849 18889 11852
rect 18923 11849 18935 11883
rect 18877 11843 18935 11849
rect 20625 11883 20683 11889
rect 20625 11849 20637 11883
rect 20671 11880 20683 11883
rect 21174 11880 21180 11892
rect 20671 11852 21180 11880
rect 20671 11849 20683 11852
rect 20625 11843 20683 11849
rect 21174 11840 21180 11852
rect 21232 11840 21238 11892
rect 23106 11880 23112 11892
rect 23067 11852 23112 11880
rect 23106 11840 23112 11852
rect 23164 11840 23170 11892
rect 24854 11840 24860 11892
rect 24912 11880 24918 11892
rect 25501 11883 25559 11889
rect 25501 11880 25513 11883
rect 24912 11852 25513 11880
rect 24912 11840 24918 11852
rect 25501 11849 25513 11852
rect 25547 11849 25559 11883
rect 25501 11843 25559 11849
rect 1765 11815 1823 11821
rect 1765 11781 1777 11815
rect 1811 11812 1823 11815
rect 1854 11812 1860 11824
rect 1811 11784 1860 11812
rect 1811 11781 1823 11784
rect 1765 11775 1823 11781
rect 1854 11772 1860 11784
rect 1912 11772 1918 11824
rect 9214 11812 9220 11824
rect 9175 11784 9220 11812
rect 9214 11772 9220 11784
rect 9272 11772 9278 11824
rect 10870 11812 10876 11824
rect 10831 11784 10876 11812
rect 10870 11772 10876 11784
rect 10928 11772 10934 11824
rect 3789 11747 3847 11753
rect 3789 11713 3801 11747
rect 3835 11744 3847 11747
rect 4062 11744 4068 11756
rect 3835 11716 4068 11744
rect 3835 11713 3847 11716
rect 3789 11707 3847 11713
rect 4062 11704 4068 11716
rect 4120 11704 4126 11756
rect 5442 11744 5448 11756
rect 5403 11716 5448 11744
rect 5442 11704 5448 11716
rect 5500 11704 5506 11756
rect 7926 11704 7932 11756
rect 7984 11744 7990 11756
rect 8113 11747 8171 11753
rect 8113 11744 8125 11747
rect 7984 11716 8125 11744
rect 7984 11704 7990 11716
rect 8113 11713 8125 11716
rect 8159 11744 8171 11747
rect 8294 11744 8300 11756
rect 8159 11716 8300 11744
rect 8159 11713 8171 11716
rect 8113 11707 8171 11713
rect 8294 11704 8300 11716
rect 8352 11744 8358 11756
rect 8573 11747 8631 11753
rect 8573 11744 8585 11747
rect 8352 11716 8585 11744
rect 8352 11704 8358 11716
rect 8573 11713 8585 11716
rect 8619 11713 8631 11747
rect 8573 11707 8631 11713
rect 11146 11704 11152 11756
rect 11204 11744 11210 11756
rect 11425 11747 11483 11753
rect 11425 11744 11437 11747
rect 11204 11716 11437 11744
rect 11204 11704 11210 11716
rect 11425 11713 11437 11716
rect 11471 11713 11483 11747
rect 11808 11744 11836 11840
rect 12805 11815 12863 11821
rect 12805 11781 12817 11815
rect 12851 11812 12863 11815
rect 13906 11812 13912 11824
rect 12851 11784 13912 11812
rect 12851 11781 12863 11784
rect 12805 11775 12863 11781
rect 13906 11772 13912 11784
rect 13964 11772 13970 11824
rect 20806 11812 20812 11824
rect 20767 11784 20812 11812
rect 20806 11772 20812 11784
rect 20864 11772 20870 11824
rect 21818 11772 21824 11824
rect 21876 11812 21882 11824
rect 23477 11815 23535 11821
rect 23477 11812 23489 11815
rect 21876 11784 23489 11812
rect 21876 11772 21882 11784
rect 23477 11781 23489 11784
rect 23523 11812 23535 11815
rect 23842 11812 23848 11824
rect 23523 11784 23848 11812
rect 23523 11781 23535 11784
rect 23477 11775 23535 11781
rect 23842 11772 23848 11784
rect 23900 11812 23906 11824
rect 23937 11815 23995 11821
rect 23937 11812 23949 11815
rect 23900 11784 23949 11812
rect 23900 11772 23906 11784
rect 23937 11781 23949 11784
rect 23983 11812 23995 11815
rect 23983 11784 24164 11812
rect 23983 11781 23995 11784
rect 23937 11775 23995 11781
rect 13170 11744 13176 11756
rect 11808 11716 13176 11744
rect 11425 11707 11483 11713
rect 13170 11704 13176 11716
rect 13228 11704 13234 11756
rect 18325 11747 18383 11753
rect 18325 11713 18337 11747
rect 18371 11744 18383 11747
rect 19426 11744 19432 11756
rect 18371 11716 19432 11744
rect 18371 11713 18383 11716
rect 18325 11707 18383 11713
rect 19426 11704 19432 11716
rect 19484 11704 19490 11756
rect 19889 11747 19947 11753
rect 19889 11713 19901 11747
rect 19935 11744 19947 11747
rect 21082 11744 21088 11756
rect 19935 11716 21088 11744
rect 19935 11713 19947 11716
rect 19889 11707 19947 11713
rect 21082 11704 21088 11716
rect 21140 11744 21146 11756
rect 24136 11753 24164 11784
rect 21177 11747 21235 11753
rect 21177 11744 21189 11747
rect 21140 11716 21189 11744
rect 21140 11704 21146 11716
rect 21177 11713 21189 11716
rect 21223 11713 21235 11747
rect 21177 11707 21235 11713
rect 24121 11747 24179 11753
rect 24121 11713 24133 11747
rect 24167 11713 24179 11747
rect 24121 11707 24179 11713
rect 3145 11679 3203 11685
rect 3145 11645 3157 11679
rect 3191 11676 3203 11679
rect 3878 11676 3884 11688
rect 3191 11648 3884 11676
rect 3191 11645 3203 11648
rect 3145 11639 3203 11645
rect 3878 11636 3884 11648
rect 3936 11636 3942 11688
rect 4341 11679 4399 11685
rect 4341 11645 4353 11679
rect 4387 11676 4399 11679
rect 4982 11676 4988 11688
rect 4387 11648 4988 11676
rect 4387 11645 4399 11648
rect 4341 11639 4399 11645
rect 4982 11636 4988 11648
rect 5040 11676 5046 11688
rect 5169 11679 5227 11685
rect 5169 11676 5181 11679
rect 5040 11648 5181 11676
rect 5040 11636 5046 11648
rect 5169 11645 5181 11648
rect 5215 11645 5227 11679
rect 5169 11639 5227 11645
rect 7466 11636 7472 11688
rect 7524 11676 7530 11688
rect 8846 11676 8852 11688
rect 7524 11648 8852 11676
rect 7524 11636 7530 11648
rect 8846 11636 8852 11648
rect 8904 11676 8910 11688
rect 9493 11679 9551 11685
rect 9493 11676 9505 11679
rect 8904 11648 9505 11676
rect 8904 11636 8910 11648
rect 9493 11645 9505 11648
rect 9539 11645 9551 11679
rect 9493 11639 9551 11645
rect 11698 11636 11704 11688
rect 11756 11676 11762 11688
rect 14093 11679 14151 11685
rect 14093 11676 14105 11679
rect 11756 11648 14105 11676
rect 11756 11636 11762 11648
rect 14093 11645 14105 11648
rect 14139 11676 14151 11679
rect 14274 11676 14280 11688
rect 14139 11648 14280 11676
rect 14139 11645 14151 11648
rect 14093 11639 14151 11645
rect 14274 11636 14280 11648
rect 14332 11636 14338 11688
rect 24210 11636 24216 11688
rect 24268 11676 24274 11688
rect 24388 11679 24446 11685
rect 24388 11676 24400 11679
rect 24268 11648 24400 11676
rect 24268 11636 24274 11648
rect 24388 11645 24400 11648
rect 24434 11676 24446 11679
rect 25222 11676 25228 11688
rect 24434 11648 25228 11676
rect 24434 11645 24446 11648
rect 24388 11639 24446 11645
rect 25222 11636 25228 11648
rect 25280 11636 25286 11688
rect 2041 11611 2099 11617
rect 2041 11577 2053 11611
rect 2087 11608 2099 11611
rect 2130 11608 2136 11620
rect 2087 11580 2136 11608
rect 2087 11577 2099 11580
rect 2041 11571 2099 11577
rect 2130 11568 2136 11580
rect 2188 11568 2194 11620
rect 2314 11608 2320 11620
rect 2227 11580 2320 11608
rect 2314 11568 2320 11580
rect 2372 11608 2378 11620
rect 2866 11608 2872 11620
rect 2372 11580 2872 11608
rect 2372 11568 2378 11580
rect 2866 11568 2872 11580
rect 2924 11568 2930 11620
rect 4875 11611 4933 11617
rect 4875 11608 4887 11611
rect 3988 11580 4887 11608
rect 2222 11540 2228 11552
rect 2183 11512 2228 11540
rect 2222 11500 2228 11512
rect 2280 11500 2286 11552
rect 3326 11500 3332 11552
rect 3384 11540 3390 11552
rect 3789 11543 3847 11549
rect 3789 11540 3801 11543
rect 3384 11512 3801 11540
rect 3384 11500 3390 11512
rect 3789 11509 3801 11512
rect 3835 11540 3847 11543
rect 3988 11540 4016 11580
rect 4875 11577 4887 11580
rect 4921 11577 4933 11611
rect 4875 11571 4933 11577
rect 7101 11611 7159 11617
rect 7101 11577 7113 11611
rect 7147 11608 7159 11611
rect 7742 11608 7748 11620
rect 7147 11580 7748 11608
rect 7147 11577 7159 11580
rect 7101 11571 7159 11577
rect 7742 11568 7748 11580
rect 7800 11568 7806 11620
rect 8018 11568 8024 11620
rect 8076 11608 8082 11620
rect 8205 11611 8263 11617
rect 8205 11608 8217 11611
rect 8076 11580 8217 11608
rect 8076 11568 8082 11580
rect 8205 11577 8217 11580
rect 8251 11577 8263 11611
rect 8205 11571 8263 11577
rect 3835 11512 4016 11540
rect 4709 11543 4767 11549
rect 3835 11509 3847 11512
rect 3789 11503 3847 11509
rect 4709 11509 4721 11543
rect 4755 11540 4767 11543
rect 5350 11540 5356 11552
rect 4755 11512 5356 11540
rect 4755 11509 4767 11512
rect 4709 11503 4767 11509
rect 5350 11500 5356 11512
rect 5408 11500 5414 11552
rect 6638 11540 6644 11552
rect 6599 11512 6644 11540
rect 6638 11500 6644 11512
rect 6696 11500 6702 11552
rect 7650 11500 7656 11552
rect 7708 11540 7714 11552
rect 8110 11540 8116 11552
rect 7708 11512 8116 11540
rect 7708 11500 7714 11512
rect 8110 11500 8116 11512
rect 8168 11500 8174 11552
rect 8220 11540 8248 11571
rect 9122 11568 9128 11620
rect 9180 11608 9186 11620
rect 9769 11611 9827 11617
rect 9769 11608 9781 11611
rect 9180 11580 9781 11608
rect 9180 11568 9186 11580
rect 9769 11577 9781 11580
rect 9815 11608 9827 11611
rect 10137 11611 10195 11617
rect 10137 11608 10149 11611
rect 9815 11580 10149 11608
rect 9815 11577 9827 11580
rect 9769 11571 9827 11577
rect 10137 11577 10149 11580
rect 10183 11608 10195 11611
rect 10318 11608 10324 11620
rect 10183 11580 10324 11608
rect 10183 11577 10195 11580
rect 10137 11571 10195 11577
rect 10318 11568 10324 11580
rect 10376 11568 10382 11620
rect 11149 11611 11207 11617
rect 11149 11577 11161 11611
rect 11195 11577 11207 11611
rect 11149 11571 11207 11577
rect 9030 11540 9036 11552
rect 8220 11512 9036 11540
rect 9030 11500 9036 11512
rect 9088 11500 9094 11552
rect 9674 11540 9680 11552
rect 9635 11512 9680 11540
rect 9674 11500 9680 11512
rect 9732 11500 9738 11552
rect 9858 11500 9864 11552
rect 9916 11540 9922 11552
rect 10597 11543 10655 11549
rect 10597 11540 10609 11543
rect 9916 11512 10609 11540
rect 9916 11500 9922 11512
rect 10597 11509 10609 11512
rect 10643 11540 10655 11543
rect 11164 11540 11192 11571
rect 11238 11568 11244 11620
rect 11296 11608 11302 11620
rect 11333 11611 11391 11617
rect 11333 11608 11345 11611
rect 11296 11580 11345 11608
rect 11296 11568 11302 11580
rect 11333 11577 11345 11580
rect 11379 11577 11391 11611
rect 11333 11571 11391 11577
rect 11606 11568 11612 11620
rect 11664 11608 11670 11620
rect 12161 11611 12219 11617
rect 12161 11608 12173 11611
rect 11664 11580 12173 11608
rect 11664 11568 11670 11580
rect 12161 11577 12173 11580
rect 12207 11577 12219 11611
rect 12161 11571 12219 11577
rect 13357 11611 13415 11617
rect 13357 11577 13369 11611
rect 13403 11608 13415 11611
rect 13725 11611 13783 11617
rect 13725 11608 13737 11611
rect 13403 11580 13737 11608
rect 13403 11577 13415 11580
rect 13357 11571 13415 11577
rect 13725 11577 13737 11580
rect 13771 11608 13783 11611
rect 14458 11608 14464 11620
rect 13771 11580 14464 11608
rect 13771 11577 13783 11580
rect 13725 11571 13783 11577
rect 12066 11540 12072 11552
rect 10643 11512 12072 11540
rect 10643 11509 10655 11512
rect 10597 11503 10655 11509
rect 12066 11500 12072 11512
rect 12124 11500 12130 11552
rect 12176 11540 12204 11571
rect 14458 11568 14464 11580
rect 14516 11617 14522 11620
rect 14516 11611 14580 11617
rect 14516 11577 14534 11611
rect 14568 11577 14580 11611
rect 14516 11571 14580 11577
rect 14516 11568 14522 11571
rect 18782 11568 18788 11620
rect 18840 11608 18846 11620
rect 19153 11611 19211 11617
rect 19153 11608 19165 11611
rect 18840 11580 19165 11608
rect 18840 11568 18846 11580
rect 19153 11577 19165 11580
rect 19199 11577 19211 11611
rect 19153 11571 19211 11577
rect 20257 11611 20315 11617
rect 20257 11577 20269 11611
rect 20303 11608 20315 11611
rect 21358 11608 21364 11620
rect 20303 11580 21364 11608
rect 20303 11577 20315 11580
rect 20257 11571 20315 11577
rect 21358 11568 21364 11580
rect 21416 11568 21422 11620
rect 13262 11540 13268 11552
rect 12176 11512 13268 11540
rect 13262 11500 13268 11512
rect 13320 11500 13326 11552
rect 16666 11500 16672 11552
rect 16724 11540 16730 11552
rect 17218 11540 17224 11552
rect 16724 11512 17224 11540
rect 16724 11500 16730 11512
rect 17218 11500 17224 11512
rect 17276 11500 17282 11552
rect 18598 11540 18604 11552
rect 18559 11512 18604 11540
rect 18598 11500 18604 11512
rect 18656 11540 18662 11552
rect 19337 11543 19395 11549
rect 19337 11540 19349 11543
rect 18656 11512 19349 11540
rect 18656 11500 18662 11512
rect 19337 11509 19349 11512
rect 19383 11509 19395 11543
rect 19337 11503 19395 11509
rect 19518 11500 19524 11552
rect 19576 11540 19582 11552
rect 21082 11540 21088 11552
rect 19576 11512 21088 11540
rect 19576 11500 19582 11512
rect 21082 11500 21088 11512
rect 21140 11540 21146 11552
rect 21269 11543 21327 11549
rect 21269 11540 21281 11543
rect 21140 11512 21281 11540
rect 21140 11500 21146 11512
rect 21269 11509 21281 11512
rect 21315 11509 21327 11543
rect 21818 11540 21824 11552
rect 21779 11512 21824 11540
rect 21269 11503 21327 11509
rect 21818 11500 21824 11512
rect 21876 11500 21882 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 2225 11339 2283 11345
rect 2225 11305 2237 11339
rect 2271 11336 2283 11339
rect 2314 11336 2320 11348
rect 2271 11308 2320 11336
rect 2271 11305 2283 11308
rect 2225 11299 2283 11305
rect 2314 11296 2320 11308
rect 2372 11296 2378 11348
rect 2869 11339 2927 11345
rect 2869 11305 2881 11339
rect 2915 11336 2927 11339
rect 2958 11336 2964 11348
rect 2915 11308 2964 11336
rect 2915 11305 2927 11308
rect 2869 11299 2927 11305
rect 2958 11296 2964 11308
rect 3016 11296 3022 11348
rect 3881 11339 3939 11345
rect 3881 11305 3893 11339
rect 3927 11336 3939 11339
rect 4338 11336 4344 11348
rect 3927 11308 4344 11336
rect 3927 11305 3939 11308
rect 3881 11299 3939 11305
rect 4338 11296 4344 11308
rect 4396 11336 4402 11348
rect 5442 11336 5448 11348
rect 4396 11308 5448 11336
rect 4396 11296 4402 11308
rect 4430 11268 4436 11280
rect 4391 11240 4436 11268
rect 4430 11228 4436 11240
rect 4488 11228 4494 11280
rect 4522 11228 4528 11280
rect 4580 11268 4586 11280
rect 4724 11277 4752 11308
rect 5442 11296 5448 11308
rect 5500 11296 5506 11348
rect 6454 11336 6460 11348
rect 6415 11308 6460 11336
rect 6454 11296 6460 11308
rect 6512 11296 6518 11348
rect 8297 11339 8355 11345
rect 8297 11305 8309 11339
rect 8343 11336 8355 11339
rect 8386 11336 8392 11348
rect 8343 11308 8392 11336
rect 8343 11305 8355 11308
rect 8297 11299 8355 11305
rect 8386 11296 8392 11308
rect 8444 11296 8450 11348
rect 8938 11336 8944 11348
rect 8899 11308 8944 11336
rect 8938 11296 8944 11308
rect 8996 11296 9002 11348
rect 10778 11336 10784 11348
rect 10060 11308 10784 11336
rect 4617 11271 4675 11277
rect 4617 11268 4629 11271
rect 4580 11240 4629 11268
rect 4580 11228 4586 11240
rect 4617 11237 4629 11240
rect 4663 11237 4675 11271
rect 4617 11231 4675 11237
rect 4709 11271 4767 11277
rect 4709 11237 4721 11271
rect 4755 11237 4767 11271
rect 4709 11231 4767 11237
rect 4982 11228 4988 11280
rect 5040 11268 5046 11280
rect 8113 11271 8171 11277
rect 8113 11268 8125 11271
rect 5040 11240 8125 11268
rect 5040 11228 5046 11240
rect 8113 11237 8125 11240
rect 8159 11268 8171 11271
rect 8202 11268 8208 11280
rect 8159 11240 8208 11268
rect 8159 11237 8171 11240
rect 8113 11231 8171 11237
rect 8202 11228 8208 11240
rect 8260 11228 8266 11280
rect 10060 11277 10088 11308
rect 10778 11296 10784 11308
rect 10836 11296 10842 11348
rect 10870 11296 10876 11348
rect 10928 11336 10934 11348
rect 11149 11339 11207 11345
rect 11149 11336 11161 11339
rect 10928 11308 11161 11336
rect 10928 11296 10934 11308
rect 11149 11305 11161 11308
rect 11195 11336 11207 11339
rect 11330 11336 11336 11348
rect 11195 11308 11336 11336
rect 11195 11305 11207 11308
rect 11149 11299 11207 11305
rect 11330 11296 11336 11308
rect 11388 11296 11394 11348
rect 11609 11339 11667 11345
rect 11609 11305 11621 11339
rect 11655 11336 11667 11339
rect 11790 11336 11796 11348
rect 11655 11308 11796 11336
rect 11655 11305 11667 11308
rect 11609 11299 11667 11305
rect 11790 11296 11796 11308
rect 11848 11336 11854 11348
rect 12158 11336 12164 11348
rect 11848 11308 12164 11336
rect 11848 11296 11854 11308
rect 12158 11296 12164 11308
rect 12216 11296 12222 11348
rect 14369 11339 14427 11345
rect 14369 11305 14381 11339
rect 14415 11336 14427 11339
rect 14458 11336 14464 11348
rect 14415 11308 14464 11336
rect 14415 11305 14427 11308
rect 14369 11299 14427 11305
rect 14458 11296 14464 11308
rect 14516 11296 14522 11348
rect 15749 11339 15807 11345
rect 15749 11305 15761 11339
rect 15795 11336 15807 11339
rect 16114 11336 16120 11348
rect 15795 11308 16120 11336
rect 15795 11305 15807 11308
rect 15749 11299 15807 11305
rect 16114 11296 16120 11308
rect 16172 11296 16178 11348
rect 18782 11336 18788 11348
rect 18743 11308 18788 11336
rect 18782 11296 18788 11308
rect 18840 11296 18846 11348
rect 21082 11336 21088 11348
rect 21043 11308 21088 11336
rect 21082 11296 21088 11308
rect 21140 11296 21146 11348
rect 22094 11296 22100 11348
rect 22152 11336 22158 11348
rect 23201 11339 23259 11345
rect 23201 11336 23213 11339
rect 22152 11308 23213 11336
rect 22152 11296 22158 11308
rect 23201 11305 23213 11308
rect 23247 11336 23259 11339
rect 23750 11336 23756 11348
rect 23247 11308 23756 11336
rect 23247 11305 23259 11308
rect 23201 11299 23259 11305
rect 23750 11296 23756 11308
rect 23808 11296 23814 11348
rect 24210 11336 24216 11348
rect 24171 11308 24216 11336
rect 24210 11296 24216 11308
rect 24268 11296 24274 11348
rect 25130 11336 25136 11348
rect 24872 11308 25136 11336
rect 24872 11280 24900 11308
rect 25130 11296 25136 11308
rect 25188 11296 25194 11348
rect 10045 11271 10103 11277
rect 10045 11237 10057 11271
rect 10091 11237 10103 11271
rect 10226 11268 10232 11280
rect 10187 11240 10232 11268
rect 10045 11231 10103 11237
rect 10226 11228 10232 11240
rect 10284 11228 10290 11280
rect 11968 11271 12026 11277
rect 11968 11237 11980 11271
rect 12014 11268 12026 11271
rect 12342 11268 12348 11280
rect 12014 11240 12348 11268
rect 12014 11237 12026 11240
rect 11968 11231 12026 11237
rect 12342 11228 12348 11240
rect 12400 11228 12406 11280
rect 19334 11228 19340 11280
rect 19392 11268 19398 11280
rect 19705 11271 19763 11277
rect 19705 11268 19717 11271
rect 19392 11240 19717 11268
rect 19392 11228 19398 11240
rect 19705 11237 19717 11240
rect 19751 11237 19763 11271
rect 24670 11268 24676 11280
rect 24631 11240 24676 11268
rect 19705 11231 19763 11237
rect 24670 11228 24676 11240
rect 24728 11228 24734 11280
rect 24854 11268 24860 11280
rect 24815 11240 24860 11268
rect 24854 11228 24860 11240
rect 24912 11228 24918 11280
rect 24946 11228 24952 11280
rect 25004 11268 25010 11280
rect 25004 11240 25049 11268
rect 25004 11228 25010 11240
rect 1394 11200 1400 11212
rect 1355 11172 1400 11200
rect 1394 11160 1400 11172
rect 1452 11160 1458 11212
rect 2685 11203 2743 11209
rect 2685 11169 2697 11203
rect 2731 11200 2743 11203
rect 2774 11200 2780 11212
rect 2731 11172 2780 11200
rect 2731 11169 2743 11172
rect 2685 11163 2743 11169
rect 2774 11160 2780 11172
rect 2832 11160 2838 11212
rect 6270 11200 6276 11212
rect 6231 11172 6276 11200
rect 6270 11160 6276 11172
rect 6328 11160 6334 11212
rect 6638 11160 6644 11212
rect 6696 11200 6702 11212
rect 7009 11203 7067 11209
rect 7009 11200 7021 11203
rect 6696 11172 7021 11200
rect 6696 11160 6702 11172
rect 7009 11169 7021 11172
rect 7055 11200 7067 11203
rect 8389 11203 8447 11209
rect 8389 11200 8401 11203
rect 7055 11172 8401 11200
rect 7055 11169 7067 11172
rect 7009 11163 7067 11169
rect 8389 11169 8401 11172
rect 8435 11200 8447 11203
rect 9030 11200 9036 11212
rect 8435 11172 9036 11200
rect 8435 11169 8447 11172
rect 8389 11163 8447 11169
rect 9030 11160 9036 11172
rect 9088 11200 9094 11212
rect 9309 11203 9367 11209
rect 9309 11200 9321 11203
rect 9088 11172 9321 11200
rect 9088 11160 9094 11172
rect 9309 11169 9321 11172
rect 9355 11200 9367 11203
rect 16117 11203 16175 11209
rect 9355 11172 10364 11200
rect 9355 11169 9367 11172
rect 9309 11163 9367 11169
rect 10336 11144 10364 11172
rect 16117 11169 16129 11203
rect 16163 11200 16175 11203
rect 16298 11200 16304 11212
rect 16163 11172 16304 11200
rect 16163 11169 16175 11172
rect 16117 11163 16175 11169
rect 16298 11160 16304 11172
rect 16356 11200 16362 11212
rect 16942 11209 16948 11212
rect 16936 11200 16948 11209
rect 16356 11172 16948 11200
rect 16356 11160 16362 11172
rect 16936 11163 16948 11172
rect 16942 11160 16948 11163
rect 17000 11160 17006 11212
rect 19518 11160 19524 11212
rect 19576 11200 19582 11212
rect 19797 11203 19855 11209
rect 19797 11200 19809 11203
rect 19576 11172 19809 11200
rect 19576 11160 19582 11172
rect 19797 11169 19809 11172
rect 19843 11169 19855 11203
rect 19797 11163 19855 11169
rect 21358 11160 21364 11212
rect 21416 11200 21422 11212
rect 22094 11209 22100 11212
rect 22088 11200 22100 11209
rect 21416 11172 22100 11200
rect 21416 11160 21422 11172
rect 22088 11163 22100 11172
rect 22152 11200 22158 11212
rect 22152 11172 22236 11200
rect 22094 11160 22100 11163
rect 22152 11160 22158 11172
rect 23382 11160 23388 11212
rect 23440 11200 23446 11212
rect 24210 11200 24216 11212
rect 23440 11172 24216 11200
rect 23440 11160 23446 11172
rect 24210 11160 24216 11172
rect 24268 11160 24274 11212
rect 1673 11135 1731 11141
rect 1673 11101 1685 11135
rect 1719 11132 1731 11135
rect 2866 11132 2872 11144
rect 1719 11104 2872 11132
rect 1719 11101 1731 11104
rect 1673 11095 1731 11101
rect 2866 11092 2872 11104
rect 2924 11092 2930 11144
rect 3513 11135 3571 11141
rect 3513 11101 3525 11135
rect 3559 11132 3571 11135
rect 4154 11132 4160 11144
rect 3559 11104 4160 11132
rect 3559 11101 3571 11104
rect 3513 11095 3571 11101
rect 4154 11092 4160 11104
rect 4212 11092 4218 11144
rect 6546 11132 6552 11144
rect 6507 11104 6552 11132
rect 6546 11092 6552 11104
rect 6604 11092 6610 11144
rect 7650 11132 7656 11144
rect 7611 11104 7656 11132
rect 7650 11092 7656 11104
rect 7708 11092 7714 11144
rect 10318 11132 10324 11144
rect 10279 11104 10324 11132
rect 10318 11092 10324 11104
rect 10376 11092 10382 11144
rect 11698 11132 11704 11144
rect 11659 11104 11704 11132
rect 11698 11092 11704 11104
rect 11756 11092 11762 11144
rect 16666 11132 16672 11144
rect 16627 11104 16672 11132
rect 16666 11092 16672 11104
rect 16724 11092 16730 11144
rect 19426 11092 19432 11144
rect 19484 11132 19490 11144
rect 19613 11135 19671 11141
rect 19613 11132 19625 11135
rect 19484 11104 19625 11132
rect 19484 11092 19490 11104
rect 19613 11101 19625 11104
rect 19659 11101 19671 11135
rect 21818 11132 21824 11144
rect 21779 11104 21824 11132
rect 19613 11095 19671 11101
rect 21818 11092 21824 11104
rect 21876 11092 21882 11144
rect 24118 11092 24124 11144
rect 24176 11132 24182 11144
rect 24176 11104 24440 11132
rect 24176 11092 24182 11104
rect 2314 11024 2320 11076
rect 2372 11064 2378 11076
rect 2501 11067 2559 11073
rect 2501 11064 2513 11067
rect 2372 11036 2513 11064
rect 2372 11024 2378 11036
rect 2501 11033 2513 11036
rect 2547 11033 2559 11067
rect 2501 11027 2559 11033
rect 4062 11024 4068 11076
rect 4120 11064 4126 11076
rect 4120 11036 4200 11064
rect 4120 11024 4126 11036
rect 4172 11005 4200 11036
rect 5534 11024 5540 11076
rect 5592 11064 5598 11076
rect 5997 11067 6055 11073
rect 5997 11064 6009 11067
rect 5592 11036 6009 11064
rect 5592 11024 5598 11036
rect 5997 11033 6009 11036
rect 6043 11033 6055 11067
rect 5997 11027 6055 11033
rect 7006 11024 7012 11076
rect 7064 11064 7070 11076
rect 7837 11067 7895 11073
rect 7837 11064 7849 11067
rect 7064 11036 7849 11064
rect 7064 11024 7070 11036
rect 7837 11033 7849 11036
rect 7883 11033 7895 11067
rect 7837 11027 7895 11033
rect 9769 11067 9827 11073
rect 9769 11033 9781 11067
rect 9815 11064 9827 11067
rect 10042 11064 10048 11076
rect 9815 11036 10048 11064
rect 9815 11033 9827 11036
rect 9769 11027 9827 11033
rect 10042 11024 10048 11036
rect 10100 11024 10106 11076
rect 10873 11067 10931 11073
rect 10873 11033 10885 11067
rect 10919 11064 10931 11067
rect 11146 11064 11152 11076
rect 10919 11036 11152 11064
rect 10919 11033 10931 11036
rect 10873 11027 10931 11033
rect 11146 11024 11152 11036
rect 11204 11024 11210 11076
rect 18874 11024 18880 11076
rect 18932 11064 18938 11076
rect 24412 11073 24440 11104
rect 19245 11067 19303 11073
rect 19245 11064 19257 11067
rect 18932 11036 19257 11064
rect 18932 11024 18938 11036
rect 19245 11033 19257 11036
rect 19291 11033 19303 11067
rect 19245 11027 19303 11033
rect 24397 11067 24455 11073
rect 24397 11033 24409 11067
rect 24443 11033 24455 11067
rect 24397 11027 24455 11033
rect 4157 10999 4215 11005
rect 4157 10965 4169 10999
rect 4203 10965 4215 10999
rect 5166 10996 5172 11008
rect 5127 10968 5172 10996
rect 4157 10959 4215 10965
rect 5166 10956 5172 10968
rect 5224 10956 5230 11008
rect 7190 10956 7196 11008
rect 7248 10996 7254 11008
rect 8570 10996 8576 11008
rect 7248 10968 8576 10996
rect 7248 10956 7254 10968
rect 8570 10956 8576 10968
rect 8628 10956 8634 11008
rect 13078 10996 13084 11008
rect 13039 10968 13084 10996
rect 13078 10956 13084 10968
rect 13136 10956 13142 11008
rect 18049 10999 18107 11005
rect 18049 10965 18061 10999
rect 18095 10996 18107 10999
rect 19518 10996 19524 11008
rect 18095 10968 19524 10996
rect 18095 10965 18107 10968
rect 18049 10959 18107 10965
rect 19518 10956 19524 10968
rect 19576 10956 19582 11008
rect 21450 10996 21456 11008
rect 21411 10968 21456 10996
rect 21450 10956 21456 10968
rect 21508 10956 21514 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 3786 10792 3792 10804
rect 3747 10764 3792 10792
rect 3786 10752 3792 10764
rect 3844 10752 3850 10804
rect 4430 10752 4436 10804
rect 4488 10792 4494 10804
rect 4525 10795 4583 10801
rect 4525 10792 4537 10795
rect 4488 10764 4537 10792
rect 4488 10752 4494 10764
rect 4525 10761 4537 10764
rect 4571 10761 4583 10795
rect 4525 10755 4583 10761
rect 5997 10795 6055 10801
rect 5997 10761 6009 10795
rect 6043 10792 6055 10795
rect 6546 10792 6552 10804
rect 6043 10764 6552 10792
rect 6043 10761 6055 10764
rect 5997 10755 6055 10761
rect 6546 10752 6552 10764
rect 6604 10792 6610 10804
rect 6822 10792 6828 10804
rect 6604 10764 6828 10792
rect 6604 10752 6610 10764
rect 6822 10752 6828 10764
rect 6880 10752 6886 10804
rect 7006 10792 7012 10804
rect 6967 10764 7012 10792
rect 7006 10752 7012 10764
rect 7064 10752 7070 10804
rect 8021 10795 8079 10801
rect 8021 10761 8033 10795
rect 8067 10792 8079 10795
rect 8386 10792 8392 10804
rect 8067 10764 8392 10792
rect 8067 10761 8079 10764
rect 8021 10755 8079 10761
rect 8386 10752 8392 10764
rect 8444 10752 8450 10804
rect 8938 10752 8944 10804
rect 8996 10792 9002 10804
rect 9309 10795 9367 10801
rect 9309 10792 9321 10795
rect 8996 10764 9321 10792
rect 8996 10752 9002 10764
rect 9309 10761 9321 10764
rect 9355 10761 9367 10795
rect 9309 10755 9367 10761
rect 10321 10795 10379 10801
rect 10321 10761 10333 10795
rect 10367 10792 10379 10795
rect 10778 10792 10784 10804
rect 10367 10764 10784 10792
rect 10367 10761 10379 10764
rect 10321 10755 10379 10761
rect 10778 10752 10784 10764
rect 10836 10752 10842 10804
rect 11054 10752 11060 10804
rect 11112 10792 11118 10804
rect 12069 10795 12127 10801
rect 12069 10792 12081 10795
rect 11112 10764 12081 10792
rect 11112 10752 11118 10764
rect 12069 10761 12081 10764
rect 12115 10792 12127 10795
rect 12161 10795 12219 10801
rect 12161 10792 12173 10795
rect 12115 10764 12173 10792
rect 12115 10761 12127 10764
rect 12069 10755 12127 10761
rect 12161 10761 12173 10764
rect 12207 10761 12219 10795
rect 12161 10755 12219 10761
rect 14274 10752 14280 10804
rect 14332 10792 14338 10804
rect 14369 10795 14427 10801
rect 14369 10792 14381 10795
rect 14332 10764 14381 10792
rect 14332 10752 14338 10764
rect 14369 10761 14381 10764
rect 14415 10792 14427 10795
rect 16666 10792 16672 10804
rect 14415 10764 16672 10792
rect 14415 10761 14427 10764
rect 14369 10755 14427 10761
rect 2682 10724 2688 10736
rect 2643 10696 2688 10724
rect 2682 10684 2688 10696
rect 2740 10684 2746 10736
rect 2774 10684 2780 10736
rect 2832 10724 2838 10736
rect 3513 10727 3571 10733
rect 3513 10724 3525 10727
rect 2832 10696 3525 10724
rect 2832 10684 2838 10696
rect 3513 10693 3525 10696
rect 3559 10724 3571 10727
rect 3970 10724 3976 10736
rect 3559 10696 3976 10724
rect 3559 10693 3571 10696
rect 3513 10687 3571 10693
rect 3970 10684 3976 10696
rect 4028 10684 4034 10736
rect 4614 10684 4620 10736
rect 4672 10724 4678 10736
rect 4801 10727 4859 10733
rect 4801 10724 4813 10727
rect 4672 10696 4813 10724
rect 4672 10684 4678 10696
rect 4801 10693 4813 10696
rect 4847 10693 4859 10727
rect 4801 10687 4859 10693
rect 8202 10684 8208 10736
rect 8260 10724 8266 10736
rect 8297 10727 8355 10733
rect 8297 10724 8309 10727
rect 8260 10696 8309 10724
rect 8260 10684 8266 10696
rect 8297 10693 8309 10696
rect 8343 10724 8355 10727
rect 8478 10724 8484 10736
rect 8343 10696 8484 10724
rect 8343 10693 8355 10696
rect 8297 10687 8355 10693
rect 8478 10684 8484 10696
rect 8536 10684 8542 10736
rect 10870 10724 10876 10736
rect 10831 10696 10876 10724
rect 10870 10684 10876 10696
rect 10928 10684 10934 10736
rect 12526 10724 12532 10736
rect 12487 10696 12532 10724
rect 12526 10684 12532 10696
rect 12584 10684 12590 10736
rect 5166 10616 5172 10668
rect 5224 10656 5230 10668
rect 5353 10659 5411 10665
rect 5353 10656 5365 10659
rect 5224 10628 5365 10656
rect 5224 10616 5230 10628
rect 5353 10625 5365 10628
rect 5399 10625 5411 10659
rect 5353 10619 5411 10625
rect 7098 10616 7104 10668
rect 7156 10656 7162 10668
rect 7469 10659 7527 10665
rect 7469 10656 7481 10659
rect 7156 10628 7481 10656
rect 7156 10616 7162 10628
rect 7469 10625 7481 10628
rect 7515 10656 7527 10659
rect 7558 10656 7564 10668
rect 7515 10628 7564 10656
rect 7515 10625 7527 10628
rect 7469 10619 7527 10625
rect 7558 10616 7564 10628
rect 7616 10616 7622 10668
rect 9125 10659 9183 10665
rect 9125 10625 9137 10659
rect 9171 10656 9183 10659
rect 9769 10659 9827 10665
rect 9769 10656 9781 10659
rect 9171 10628 9781 10656
rect 9171 10625 9183 10628
rect 9125 10619 9183 10625
rect 9769 10625 9781 10628
rect 9815 10656 9827 10659
rect 9950 10656 9956 10668
rect 9815 10628 9956 10656
rect 9815 10625 9827 10628
rect 9769 10619 9827 10625
rect 9950 10616 9956 10628
rect 10008 10656 10014 10668
rect 11333 10659 11391 10665
rect 10008 10628 11284 10656
rect 10008 10616 10014 10628
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10588 1455 10591
rect 1946 10588 1952 10600
rect 1443 10560 1952 10588
rect 1443 10557 1455 10560
rect 1397 10551 1455 10557
rect 1946 10548 1952 10560
rect 2004 10588 2010 10600
rect 2501 10591 2559 10597
rect 2004 10560 2084 10588
rect 2004 10548 2010 10560
rect 2056 10464 2084 10560
rect 2501 10557 2513 10591
rect 2547 10557 2559 10591
rect 2501 10551 2559 10557
rect 2516 10520 2544 10551
rect 2866 10548 2872 10600
rect 2924 10588 2930 10600
rect 3602 10588 3608 10600
rect 2924 10560 3608 10588
rect 2924 10548 2930 10560
rect 3602 10548 3608 10560
rect 3660 10548 3666 10600
rect 4154 10548 4160 10600
rect 4212 10588 4218 10600
rect 5077 10591 5135 10597
rect 5077 10588 5089 10591
rect 4212 10560 5089 10588
rect 4212 10548 4218 10560
rect 5077 10557 5089 10560
rect 5123 10588 5135 10591
rect 5442 10588 5448 10600
rect 5123 10560 5448 10588
rect 5123 10557 5135 10560
rect 5077 10551 5135 10557
rect 5442 10548 5448 10560
rect 5500 10548 5506 10600
rect 11256 10588 11284 10628
rect 11333 10625 11345 10659
rect 11379 10656 11391 10659
rect 13170 10656 13176 10668
rect 11379 10628 13176 10656
rect 11379 10625 11391 10628
rect 11333 10619 11391 10625
rect 13170 10616 13176 10628
rect 13228 10656 13234 10668
rect 13817 10659 13875 10665
rect 13817 10656 13829 10659
rect 13228 10628 13829 10656
rect 13228 10616 13234 10628
rect 13817 10625 13829 10628
rect 13863 10625 13875 10659
rect 14384 10656 14412 10755
rect 16666 10752 16672 10764
rect 16724 10752 16730 10804
rect 19610 10792 19616 10804
rect 19571 10764 19616 10792
rect 19610 10752 19616 10764
rect 19668 10752 19674 10804
rect 20806 10792 20812 10804
rect 20767 10764 20812 10792
rect 20806 10752 20812 10764
rect 20864 10752 20870 10804
rect 21818 10792 21824 10804
rect 21376 10764 21824 10792
rect 18046 10684 18052 10736
rect 18104 10724 18110 10736
rect 18141 10727 18199 10733
rect 18141 10724 18153 10727
rect 18104 10696 18153 10724
rect 18104 10684 18110 10696
rect 18141 10693 18153 10696
rect 18187 10693 18199 10727
rect 18141 10687 18199 10693
rect 19889 10727 19947 10733
rect 19889 10693 19901 10727
rect 19935 10724 19947 10727
rect 20622 10724 20628 10736
rect 19935 10696 20628 10724
rect 19935 10693 19947 10696
rect 19889 10687 19947 10693
rect 20622 10684 20628 10696
rect 20680 10684 20686 10736
rect 20714 10684 20720 10736
rect 20772 10724 20778 10736
rect 21376 10724 21404 10764
rect 21818 10752 21824 10764
rect 21876 10792 21882 10804
rect 22373 10795 22431 10801
rect 22373 10792 22385 10795
rect 21876 10764 22385 10792
rect 21876 10752 21882 10764
rect 22373 10761 22385 10764
rect 22419 10792 22431 10795
rect 23385 10795 23443 10801
rect 23385 10792 23397 10795
rect 22419 10764 23397 10792
rect 22419 10761 22431 10764
rect 22373 10755 22431 10761
rect 23385 10761 23397 10764
rect 23431 10761 23443 10795
rect 23385 10755 23443 10761
rect 25041 10795 25099 10801
rect 25041 10761 25053 10795
rect 25087 10792 25099 10795
rect 25498 10792 25504 10804
rect 25087 10764 25504 10792
rect 25087 10761 25099 10764
rect 25041 10755 25099 10761
rect 20772 10696 21404 10724
rect 21453 10727 21511 10733
rect 20772 10684 20778 10696
rect 21453 10693 21465 10727
rect 21499 10724 21511 10727
rect 21910 10724 21916 10736
rect 21499 10696 21916 10724
rect 21499 10693 21511 10696
rect 21453 10687 21511 10693
rect 21910 10684 21916 10696
rect 21968 10684 21974 10736
rect 14553 10659 14611 10665
rect 14553 10656 14565 10659
rect 14384 10628 14565 10656
rect 13817 10619 13875 10625
rect 14553 10625 14565 10628
rect 14599 10625 14611 10659
rect 14553 10619 14611 10625
rect 21269 10659 21327 10665
rect 21269 10625 21281 10659
rect 21315 10656 21327 10659
rect 22002 10656 22008 10668
rect 21315 10628 22008 10656
rect 21315 10625 21327 10628
rect 21269 10619 21327 10625
rect 22002 10616 22008 10628
rect 22060 10616 22066 10668
rect 23400 10656 23428 10755
rect 25498 10752 25504 10764
rect 25556 10752 25562 10804
rect 24946 10684 24952 10736
rect 25004 10724 25010 10736
rect 25593 10727 25651 10733
rect 25593 10724 25605 10727
rect 25004 10696 25605 10724
rect 25004 10684 25010 10696
rect 25593 10693 25605 10696
rect 25639 10693 25651 10727
rect 25593 10687 25651 10693
rect 23661 10659 23719 10665
rect 23661 10656 23673 10659
rect 23400 10628 23673 10656
rect 23661 10625 23673 10628
rect 23707 10625 23719 10659
rect 23661 10619 23719 10625
rect 11882 10588 11888 10600
rect 11256 10560 11744 10588
rect 11795 10560 11888 10588
rect 3145 10523 3203 10529
rect 3145 10520 3157 10523
rect 2516 10492 3157 10520
rect 3145 10489 3157 10492
rect 3191 10520 3203 10523
rect 6641 10523 6699 10529
rect 6641 10520 6653 10523
rect 3191 10492 6653 10520
rect 3191 10489 3203 10492
rect 3145 10483 3203 10489
rect 6641 10489 6653 10492
rect 6687 10520 6699 10523
rect 7466 10520 7472 10532
rect 6687 10492 7472 10520
rect 6687 10489 6699 10492
rect 6641 10483 6699 10489
rect 7466 10480 7472 10492
rect 7524 10480 7530 10532
rect 7561 10523 7619 10529
rect 7561 10489 7573 10523
rect 7607 10520 7619 10523
rect 8386 10520 8392 10532
rect 7607 10492 8392 10520
rect 7607 10489 7619 10492
rect 7561 10483 7619 10489
rect 8386 10480 8392 10492
rect 8444 10520 8450 10532
rect 8757 10523 8815 10529
rect 8757 10520 8769 10523
rect 8444 10492 8769 10520
rect 8444 10480 8450 10492
rect 8757 10489 8769 10492
rect 8803 10520 8815 10523
rect 9861 10523 9919 10529
rect 9861 10520 9873 10523
rect 8803 10492 9873 10520
rect 8803 10489 8815 10492
rect 8757 10483 8815 10489
rect 9861 10489 9873 10492
rect 9907 10520 9919 10523
rect 10042 10520 10048 10532
rect 9907 10492 10048 10520
rect 9907 10489 9919 10492
rect 9861 10483 9919 10489
rect 10042 10480 10048 10492
rect 10100 10520 10106 10532
rect 10318 10520 10324 10532
rect 10100 10492 10324 10520
rect 10100 10480 10106 10492
rect 10318 10480 10324 10492
rect 10376 10480 10382 10532
rect 11330 10520 11336 10532
rect 11291 10492 11336 10520
rect 11330 10480 11336 10492
rect 11388 10480 11394 10532
rect 11425 10523 11483 10529
rect 11425 10489 11437 10523
rect 11471 10489 11483 10523
rect 11716 10520 11744 10560
rect 11882 10548 11888 10560
rect 11940 10588 11946 10600
rect 12805 10591 12863 10597
rect 12805 10588 12817 10591
rect 11940 10560 12817 10588
rect 11940 10548 11946 10560
rect 12805 10557 12817 10560
rect 12851 10588 12863 10591
rect 13722 10588 13728 10600
rect 12851 10560 13728 10588
rect 12851 10557 12863 10560
rect 12805 10551 12863 10557
rect 13722 10548 13728 10560
rect 13780 10548 13786 10600
rect 17497 10591 17555 10597
rect 17497 10557 17509 10591
rect 17543 10588 17555 10591
rect 17678 10588 17684 10600
rect 17543 10560 17684 10588
rect 17543 10557 17555 10560
rect 17497 10551 17555 10557
rect 17678 10548 17684 10560
rect 17736 10588 17742 10600
rect 19337 10591 19395 10597
rect 17736 10560 18736 10588
rect 17736 10548 17742 10560
rect 12710 10520 12716 10532
rect 11716 10492 12716 10520
rect 11425 10483 11483 10489
rect 1581 10455 1639 10461
rect 1581 10421 1593 10455
rect 1627 10452 1639 10455
rect 1762 10452 1768 10464
rect 1627 10424 1768 10452
rect 1627 10421 1639 10424
rect 1581 10415 1639 10421
rect 1762 10412 1768 10424
rect 1820 10412 1826 10464
rect 2038 10452 2044 10464
rect 1999 10424 2044 10452
rect 2038 10412 2044 10424
rect 2096 10412 2102 10464
rect 2222 10412 2228 10464
rect 2280 10452 2286 10464
rect 2317 10455 2375 10461
rect 2317 10452 2329 10455
rect 2280 10424 2329 10452
rect 2280 10412 2286 10424
rect 2317 10421 2329 10424
rect 2363 10421 2375 10455
rect 2317 10415 2375 10421
rect 3510 10412 3516 10464
rect 3568 10452 3574 10464
rect 4157 10455 4215 10461
rect 4157 10452 4169 10455
rect 3568 10424 4169 10452
rect 3568 10412 3574 10424
rect 4157 10421 4169 10424
rect 4203 10452 4215 10455
rect 4522 10452 4528 10464
rect 4203 10424 4528 10452
rect 4203 10421 4215 10424
rect 4157 10415 4215 10421
rect 4522 10412 4528 10424
rect 4580 10412 4586 10464
rect 5261 10455 5319 10461
rect 5261 10421 5273 10455
rect 5307 10452 5319 10455
rect 5442 10452 5448 10464
rect 5307 10424 5448 10452
rect 5307 10421 5319 10424
rect 5261 10415 5319 10421
rect 5442 10412 5448 10424
rect 5500 10412 5506 10464
rect 9769 10455 9827 10461
rect 9769 10421 9781 10455
rect 9815 10452 9827 10455
rect 9950 10452 9956 10464
rect 9815 10424 9956 10452
rect 9815 10421 9827 10424
rect 9769 10415 9827 10421
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 10689 10455 10747 10461
rect 10689 10421 10701 10455
rect 10735 10452 10747 10455
rect 10778 10452 10784 10464
rect 10735 10424 10784 10452
rect 10735 10421 10747 10424
rect 10689 10415 10747 10421
rect 10778 10412 10784 10424
rect 10836 10452 10842 10464
rect 11440 10452 11468 10483
rect 12710 10480 12716 10492
rect 12768 10480 12774 10532
rect 13078 10520 13084 10532
rect 12991 10492 13084 10520
rect 13078 10480 13084 10492
rect 13136 10480 13142 10532
rect 14642 10480 14648 10532
rect 14700 10520 14706 10532
rect 14798 10523 14856 10529
rect 14798 10520 14810 10523
rect 14700 10492 14810 10520
rect 14700 10480 14706 10492
rect 14798 10489 14810 10492
rect 14844 10489 14856 10523
rect 14798 10483 14856 10489
rect 16942 10480 16948 10532
rect 17000 10520 17006 10532
rect 17129 10523 17187 10529
rect 17129 10520 17141 10523
rect 17000 10492 17141 10520
rect 17000 10480 17006 10492
rect 17129 10489 17141 10492
rect 17175 10520 17187 10523
rect 17862 10520 17868 10532
rect 17175 10492 17868 10520
rect 17175 10489 17187 10492
rect 17129 10483 17187 10489
rect 17862 10480 17868 10492
rect 17920 10480 17926 10532
rect 18708 10529 18736 10560
rect 19337 10557 19349 10591
rect 19383 10588 19395 10591
rect 20070 10588 20076 10600
rect 19383 10560 20076 10588
rect 19383 10557 19395 10560
rect 19337 10551 19395 10557
rect 20070 10548 20076 10560
rect 20128 10588 20134 10600
rect 20128 10560 20484 10588
rect 20128 10548 20134 10560
rect 20456 10532 20484 10560
rect 23750 10548 23756 10600
rect 23808 10588 23814 10600
rect 23917 10591 23975 10597
rect 23917 10588 23929 10591
rect 23808 10560 23929 10588
rect 23808 10548 23814 10560
rect 23917 10557 23929 10560
rect 23963 10557 23975 10591
rect 23917 10551 23975 10557
rect 18417 10523 18475 10529
rect 18417 10489 18429 10523
rect 18463 10489 18475 10523
rect 18417 10483 18475 10489
rect 18693 10523 18751 10529
rect 18693 10489 18705 10523
rect 18739 10520 18751 10523
rect 19518 10520 19524 10532
rect 18739 10492 19524 10520
rect 18739 10489 18751 10492
rect 18693 10483 18751 10489
rect 10836 10424 11468 10452
rect 12069 10455 12127 10461
rect 10836 10412 10842 10424
rect 12069 10421 12081 10455
rect 12115 10452 12127 10455
rect 12989 10455 13047 10461
rect 12989 10452 13001 10455
rect 12115 10424 13001 10452
rect 12115 10421 12127 10424
rect 12069 10415 12127 10421
rect 12989 10421 13001 10424
rect 13035 10421 13047 10455
rect 13096 10452 13124 10480
rect 13446 10452 13452 10464
rect 13096 10424 13452 10452
rect 12989 10415 13047 10421
rect 13446 10412 13452 10424
rect 13504 10412 13510 10464
rect 14458 10412 14464 10464
rect 14516 10452 14522 10464
rect 15562 10452 15568 10464
rect 14516 10424 15568 10452
rect 14516 10412 14522 10424
rect 15562 10412 15568 10424
rect 15620 10452 15626 10464
rect 15933 10455 15991 10461
rect 15933 10452 15945 10455
rect 15620 10424 15945 10452
rect 15620 10412 15626 10424
rect 15933 10421 15945 10424
rect 15979 10421 15991 10455
rect 17770 10452 17776 10464
rect 17731 10424 17776 10452
rect 15933 10415 15991 10421
rect 17770 10412 17776 10424
rect 17828 10452 17834 10464
rect 18432 10452 18460 10483
rect 19518 10480 19524 10492
rect 19576 10480 19582 10532
rect 19610 10480 19616 10532
rect 19668 10480 19674 10532
rect 19978 10480 19984 10532
rect 20036 10520 20042 10532
rect 20165 10523 20223 10529
rect 20165 10520 20177 10523
rect 20036 10492 20177 10520
rect 20036 10480 20042 10492
rect 20165 10489 20177 10492
rect 20211 10489 20223 10523
rect 20438 10520 20444 10532
rect 20399 10492 20444 10520
rect 20165 10483 20223 10489
rect 20438 10480 20444 10492
rect 20496 10480 20502 10532
rect 20898 10480 20904 10532
rect 20956 10520 20962 10532
rect 21450 10520 21456 10532
rect 20956 10492 21456 10520
rect 20956 10480 20962 10492
rect 21450 10480 21456 10492
rect 21508 10520 21514 10532
rect 21729 10523 21787 10529
rect 21729 10520 21741 10523
rect 21508 10492 21741 10520
rect 21508 10480 21514 10492
rect 21729 10489 21741 10492
rect 21775 10489 21787 10523
rect 21729 10483 21787 10489
rect 18598 10452 18604 10464
rect 17828 10424 18460 10452
rect 18559 10424 18604 10452
rect 17828 10412 17834 10424
rect 18598 10412 18604 10424
rect 18656 10412 18662 10464
rect 19628 10452 19656 10480
rect 20254 10452 20260 10464
rect 19628 10424 20260 10452
rect 20254 10412 20260 10424
rect 20312 10452 20318 10464
rect 20349 10455 20407 10461
rect 20349 10452 20361 10455
rect 20312 10424 20361 10452
rect 20312 10412 20318 10424
rect 20349 10421 20361 10424
rect 20395 10421 20407 10455
rect 20349 10415 20407 10421
rect 20806 10412 20812 10464
rect 20864 10452 20870 10464
rect 21913 10455 21971 10461
rect 21913 10452 21925 10455
rect 20864 10424 21925 10452
rect 20864 10412 20870 10424
rect 21913 10421 21925 10424
rect 21959 10421 21971 10455
rect 21913 10415 21971 10421
rect 22094 10412 22100 10464
rect 22152 10452 22158 10464
rect 22741 10455 22799 10461
rect 22741 10452 22753 10455
rect 22152 10424 22753 10452
rect 22152 10412 22158 10424
rect 22741 10421 22753 10424
rect 22787 10421 22799 10455
rect 22741 10415 22799 10421
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1394 10208 1400 10260
rect 1452 10248 1458 10260
rect 1949 10251 2007 10257
rect 1949 10248 1961 10251
rect 1452 10220 1961 10248
rect 1452 10208 1458 10220
rect 1949 10217 1961 10220
rect 1995 10217 2007 10251
rect 1949 10211 2007 10217
rect 2409 10251 2467 10257
rect 2409 10217 2421 10251
rect 2455 10248 2467 10251
rect 2590 10248 2596 10260
rect 2455 10220 2596 10248
rect 2455 10217 2467 10220
rect 2409 10211 2467 10217
rect 2590 10208 2596 10220
rect 2648 10208 2654 10260
rect 3326 10248 3332 10260
rect 3287 10220 3332 10248
rect 3326 10208 3332 10220
rect 3384 10208 3390 10260
rect 3602 10248 3608 10260
rect 3563 10220 3608 10248
rect 3602 10208 3608 10220
rect 3660 10208 3666 10260
rect 4338 10248 4344 10260
rect 4299 10220 4344 10248
rect 4338 10208 4344 10220
rect 4396 10208 4402 10260
rect 6178 10248 6184 10260
rect 6139 10220 6184 10248
rect 6178 10208 6184 10220
rect 6236 10208 6242 10260
rect 7009 10251 7067 10257
rect 7009 10217 7021 10251
rect 7055 10248 7067 10251
rect 7558 10248 7564 10260
rect 7055 10220 7564 10248
rect 7055 10217 7067 10220
rect 7009 10211 7067 10217
rect 7558 10208 7564 10220
rect 7616 10208 7622 10260
rect 7653 10251 7711 10257
rect 7653 10217 7665 10251
rect 7699 10248 7711 10251
rect 8846 10248 8852 10260
rect 7699 10220 8432 10248
rect 8807 10220 8852 10248
rect 7699 10217 7711 10220
rect 7653 10211 7711 10217
rect 8404 10192 8432 10220
rect 8846 10208 8852 10220
rect 8904 10208 8910 10260
rect 9953 10251 10011 10257
rect 9953 10217 9965 10251
rect 9999 10248 10011 10251
rect 10134 10248 10140 10260
rect 9999 10220 10140 10248
rect 9999 10217 10011 10220
rect 9953 10211 10011 10217
rect 10134 10208 10140 10220
rect 10192 10208 10198 10260
rect 12434 10208 12440 10260
rect 12492 10248 12498 10260
rect 13078 10248 13084 10260
rect 12492 10220 12537 10248
rect 13039 10220 13084 10248
rect 12492 10208 12498 10220
rect 13078 10208 13084 10220
rect 13136 10208 13142 10260
rect 14642 10248 14648 10260
rect 14603 10220 14648 10248
rect 14642 10208 14648 10220
rect 14700 10208 14706 10260
rect 15838 10248 15844 10260
rect 15799 10220 15844 10248
rect 15838 10208 15844 10220
rect 15896 10208 15902 10260
rect 17405 10251 17463 10257
rect 17405 10217 17417 10251
rect 17451 10248 17463 10251
rect 18598 10248 18604 10260
rect 17451 10220 18604 10248
rect 17451 10217 17463 10220
rect 17405 10211 17463 10217
rect 18598 10208 18604 10220
rect 18656 10208 18662 10260
rect 18782 10208 18788 10260
rect 18840 10248 18846 10260
rect 18877 10251 18935 10257
rect 18877 10248 18889 10251
rect 18840 10220 18889 10248
rect 18840 10208 18846 10220
rect 18877 10217 18889 10220
rect 18923 10217 18935 10251
rect 19518 10248 19524 10260
rect 19479 10220 19524 10248
rect 18877 10211 18935 10217
rect 19518 10208 19524 10220
rect 19576 10208 19582 10260
rect 23290 10248 23296 10260
rect 23251 10220 23296 10248
rect 23290 10208 23296 10220
rect 23348 10208 23354 10260
rect 23566 10208 23572 10260
rect 23624 10248 23630 10260
rect 23842 10248 23848 10260
rect 23624 10220 23848 10248
rect 23624 10208 23630 10220
rect 23842 10208 23848 10220
rect 23900 10248 23906 10260
rect 23937 10251 23995 10257
rect 23937 10248 23949 10251
rect 23900 10220 23949 10248
rect 23900 10208 23906 10220
rect 23937 10217 23949 10220
rect 23983 10217 23995 10251
rect 23937 10211 23995 10217
rect 24489 10251 24547 10257
rect 24489 10217 24501 10251
rect 24535 10248 24547 10251
rect 24670 10248 24676 10260
rect 24535 10220 24676 10248
rect 24535 10217 24547 10220
rect 24489 10211 24547 10217
rect 24670 10208 24676 10220
rect 24728 10208 24734 10260
rect 25130 10248 25136 10260
rect 25091 10220 25136 10248
rect 25130 10208 25136 10220
rect 25188 10208 25194 10260
rect 5068 10183 5126 10189
rect 5068 10149 5080 10183
rect 5114 10180 5126 10183
rect 5166 10180 5172 10192
rect 5114 10152 5172 10180
rect 5114 10149 5126 10152
rect 5068 10143 5126 10149
rect 5166 10140 5172 10152
rect 5224 10140 5230 10192
rect 8202 10140 8208 10192
rect 8260 10180 8266 10192
rect 8297 10183 8355 10189
rect 8297 10180 8309 10183
rect 8260 10152 8309 10180
rect 8260 10140 8266 10152
rect 8297 10149 8309 10152
rect 8343 10149 8355 10183
rect 8297 10143 8355 10149
rect 8386 10140 8392 10192
rect 8444 10180 8450 10192
rect 11517 10183 11575 10189
rect 11517 10180 11529 10183
rect 8444 10152 8489 10180
rect 10704 10152 11529 10180
rect 8444 10140 8450 10152
rect 10704 10124 10732 10152
rect 11517 10149 11529 10152
rect 11563 10180 11575 10183
rect 12526 10180 12532 10192
rect 11563 10152 12532 10180
rect 11563 10149 11575 10152
rect 11517 10143 11575 10149
rect 12526 10140 12532 10152
rect 12584 10140 12590 10192
rect 12710 10140 12716 10192
rect 12768 10180 12774 10192
rect 12768 10152 14228 10180
rect 12768 10140 12774 10152
rect 1394 10112 1400 10124
rect 1355 10084 1400 10112
rect 1394 10072 1400 10084
rect 1452 10072 1458 10124
rect 2501 10115 2559 10121
rect 2501 10081 2513 10115
rect 2547 10112 2559 10115
rect 2682 10112 2688 10124
rect 2547 10084 2688 10112
rect 2547 10081 2559 10084
rect 2501 10075 2559 10081
rect 2682 10072 2688 10084
rect 2740 10072 2746 10124
rect 7650 10072 7656 10124
rect 7708 10112 7714 10124
rect 8113 10115 8171 10121
rect 8113 10112 8125 10115
rect 7708 10084 8125 10112
rect 7708 10072 7714 10084
rect 8113 10081 8125 10084
rect 8159 10081 8171 10115
rect 8113 10075 8171 10081
rect 8662 10072 8668 10124
rect 8720 10112 8726 10124
rect 9309 10115 9367 10121
rect 9309 10112 9321 10115
rect 8720 10084 9321 10112
rect 8720 10072 8726 10084
rect 9309 10081 9321 10084
rect 9355 10112 9367 10115
rect 9950 10112 9956 10124
rect 9355 10084 9956 10112
rect 9355 10081 9367 10084
rect 9309 10075 9367 10081
rect 9950 10072 9956 10084
rect 10008 10072 10014 10124
rect 10686 10072 10692 10124
rect 10744 10072 10750 10124
rect 11330 10072 11336 10124
rect 11388 10112 11394 10124
rect 11388 10084 11433 10112
rect 11388 10072 11394 10084
rect 11882 10072 11888 10124
rect 11940 10112 11946 10124
rect 12897 10115 12955 10121
rect 12897 10112 12909 10115
rect 11940 10084 12909 10112
rect 11940 10072 11946 10084
rect 12897 10081 12909 10084
rect 12943 10112 12955 10115
rect 14093 10115 14151 10121
rect 14093 10112 14105 10115
rect 12943 10084 14105 10112
rect 12943 10081 12955 10084
rect 12897 10075 12955 10081
rect 14093 10081 14105 10084
rect 14139 10081 14151 10115
rect 14200 10112 14228 10152
rect 14458 10140 14464 10192
rect 14516 10180 14522 10192
rect 14921 10183 14979 10189
rect 14921 10180 14933 10183
rect 14516 10152 14933 10180
rect 14516 10140 14522 10152
rect 14921 10149 14933 10152
rect 14967 10149 14979 10183
rect 15654 10180 15660 10192
rect 14921 10143 14979 10149
rect 15028 10152 15660 10180
rect 15028 10112 15056 10152
rect 15654 10140 15660 10152
rect 15712 10140 15718 10192
rect 15933 10183 15991 10189
rect 15933 10149 15945 10183
rect 15979 10180 15991 10183
rect 16942 10180 16948 10192
rect 15979 10152 16948 10180
rect 15979 10149 15991 10152
rect 15933 10143 15991 10149
rect 14200 10084 15056 10112
rect 14093 10075 14151 10081
rect 15286 10072 15292 10124
rect 15344 10112 15350 10124
rect 15948 10112 15976 10143
rect 16942 10140 16948 10152
rect 17000 10140 17006 10192
rect 17678 10140 17684 10192
rect 17736 10189 17742 10192
rect 17736 10183 17800 10189
rect 17736 10149 17754 10183
rect 17788 10149 17800 10183
rect 17736 10143 17800 10149
rect 17736 10140 17742 10143
rect 23014 10140 23020 10192
rect 23072 10180 23078 10192
rect 23753 10183 23811 10189
rect 23753 10180 23765 10183
rect 23072 10152 23765 10180
rect 23072 10140 23078 10152
rect 23753 10149 23765 10152
rect 23799 10149 23811 10183
rect 23753 10143 23811 10149
rect 15344 10084 15976 10112
rect 21168 10115 21226 10121
rect 15344 10072 15350 10084
rect 21168 10081 21180 10115
rect 21214 10112 21226 10115
rect 21726 10112 21732 10124
rect 21214 10084 21732 10112
rect 21214 10081 21226 10084
rect 21168 10075 21226 10081
rect 21726 10072 21732 10084
rect 21784 10072 21790 10124
rect 23658 10072 23664 10124
rect 23716 10112 23722 10124
rect 24029 10115 24087 10121
rect 24029 10112 24041 10115
rect 23716 10084 24041 10112
rect 23716 10072 23722 10084
rect 24029 10081 24041 10084
rect 24075 10112 24087 10115
rect 24118 10112 24124 10124
rect 24075 10084 24124 10112
rect 24075 10081 24087 10084
rect 24029 10075 24087 10081
rect 24118 10072 24124 10084
rect 24176 10072 24182 10124
rect 24946 10112 24952 10124
rect 24907 10084 24952 10112
rect 24946 10072 24952 10084
rect 25004 10072 25010 10124
rect 4798 10044 4804 10056
rect 4759 10016 4804 10044
rect 4798 10004 4804 10016
rect 4856 10004 4862 10056
rect 10778 10004 10784 10056
rect 10836 10044 10842 10056
rect 11606 10044 11612 10056
rect 10836 10016 11612 10044
rect 10836 10004 10842 10016
rect 11606 10004 11612 10016
rect 11664 10004 11670 10056
rect 13078 10004 13084 10056
rect 13136 10044 13142 10056
rect 13173 10047 13231 10053
rect 13173 10044 13185 10047
rect 13136 10016 13185 10044
rect 13136 10004 13142 10016
rect 13173 10013 13185 10016
rect 13219 10044 13231 10047
rect 13446 10044 13452 10056
rect 13219 10016 13452 10044
rect 13219 10013 13231 10016
rect 13173 10007 13231 10013
rect 13446 10004 13452 10016
rect 13504 10004 13510 10056
rect 17494 10044 17500 10056
rect 17455 10016 17500 10044
rect 17494 10004 17500 10016
rect 17552 10004 17558 10056
rect 20714 10004 20720 10056
rect 20772 10044 20778 10056
rect 20901 10047 20959 10053
rect 20901 10044 20913 10047
rect 20772 10016 20913 10044
rect 20772 10004 20778 10016
rect 20901 10013 20913 10016
rect 20947 10013 20959 10047
rect 20901 10007 20959 10013
rect 2682 9976 2688 9988
rect 2643 9948 2688 9976
rect 2682 9936 2688 9948
rect 2740 9936 2746 9988
rect 10962 9936 10968 9988
rect 11020 9976 11026 9988
rect 11020 9948 11376 9976
rect 11020 9936 11026 9948
rect 11348 9920 11376 9948
rect 11698 9936 11704 9988
rect 11756 9976 11762 9988
rect 11977 9979 12035 9985
rect 11977 9976 11989 9979
rect 11756 9948 11989 9976
rect 11756 9936 11762 9948
rect 11977 9945 11989 9948
rect 12023 9945 12035 9979
rect 23474 9976 23480 9988
rect 23435 9948 23480 9976
rect 11977 9939 12035 9945
rect 23474 9936 23480 9948
rect 23532 9936 23538 9988
rect 23842 9936 23848 9988
rect 23900 9976 23906 9988
rect 24026 9976 24032 9988
rect 23900 9948 24032 9976
rect 23900 9936 23906 9948
rect 24026 9936 24032 9948
rect 24084 9936 24090 9988
rect 1581 9911 1639 9917
rect 1581 9877 1593 9911
rect 1627 9908 1639 9911
rect 1670 9908 1676 9920
rect 1627 9880 1676 9908
rect 1627 9877 1639 9880
rect 1581 9871 1639 9877
rect 1670 9868 1676 9880
rect 1728 9868 1734 9920
rect 4709 9911 4767 9917
rect 4709 9877 4721 9911
rect 4755 9908 4767 9911
rect 5442 9908 5448 9920
rect 4755 9880 5448 9908
rect 4755 9877 4767 9880
rect 4709 9871 4767 9877
rect 5442 9868 5448 9880
rect 5500 9868 5506 9920
rect 7834 9908 7840 9920
rect 7795 9880 7840 9908
rect 7834 9868 7840 9880
rect 7892 9868 7898 9920
rect 10042 9868 10048 9920
rect 10100 9908 10106 9920
rect 10229 9911 10287 9917
rect 10229 9908 10241 9911
rect 10100 9880 10241 9908
rect 10100 9868 10106 9880
rect 10229 9877 10241 9880
rect 10275 9877 10287 9911
rect 10778 9908 10784 9920
rect 10739 9880 10784 9908
rect 10229 9871 10287 9877
rect 10778 9868 10784 9880
rect 10836 9868 10842 9920
rect 11054 9908 11060 9920
rect 11015 9880 11060 9908
rect 11054 9868 11060 9880
rect 11112 9868 11118 9920
rect 11330 9868 11336 9920
rect 11388 9908 11394 9920
rect 12621 9911 12679 9917
rect 12621 9908 12633 9911
rect 11388 9880 12633 9908
rect 11388 9868 11394 9880
rect 12621 9877 12633 9880
rect 12667 9877 12679 9911
rect 15378 9908 15384 9920
rect 15339 9880 15384 9908
rect 12621 9871 12679 9877
rect 15378 9868 15384 9880
rect 15436 9868 15442 9920
rect 19886 9908 19892 9920
rect 19847 9880 19892 9908
rect 19886 9868 19892 9880
rect 19944 9868 19950 9920
rect 22094 9868 22100 9920
rect 22152 9908 22158 9920
rect 22281 9911 22339 9917
rect 22281 9908 22293 9911
rect 22152 9880 22293 9908
rect 22152 9868 22158 9880
rect 22281 9877 22293 9880
rect 22327 9877 22339 9911
rect 22922 9908 22928 9920
rect 22883 9880 22928 9908
rect 22281 9871 22339 9877
rect 22922 9868 22928 9880
rect 22980 9868 22986 9920
rect 24854 9908 24860 9920
rect 24767 9880 24860 9908
rect 24854 9868 24860 9880
rect 24912 9908 24918 9920
rect 25222 9908 25228 9920
rect 24912 9880 25228 9908
rect 24912 9868 24918 9880
rect 25222 9868 25228 9880
rect 25280 9868 25286 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 5166 9664 5172 9716
rect 5224 9664 5230 9716
rect 6822 9704 6828 9716
rect 5736 9676 6828 9704
rect 2498 9596 2504 9648
rect 2556 9636 2562 9648
rect 2685 9639 2743 9645
rect 2685 9636 2697 9639
rect 2556 9608 2697 9636
rect 2556 9596 2562 9608
rect 2685 9605 2697 9608
rect 2731 9605 2743 9639
rect 2685 9599 2743 9605
rect 3513 9639 3571 9645
rect 3513 9605 3525 9639
rect 3559 9636 3571 9639
rect 4062 9636 4068 9648
rect 3559 9608 4068 9636
rect 3559 9605 3571 9608
rect 3513 9599 3571 9605
rect 4062 9596 4068 9608
rect 4120 9596 4126 9648
rect 5184 9636 5212 9664
rect 5629 9639 5687 9645
rect 5629 9636 5641 9639
rect 5184 9608 5641 9636
rect 5629 9605 5641 9608
rect 5675 9605 5687 9639
rect 5629 9599 5687 9605
rect 2409 9571 2467 9577
rect 2409 9537 2421 9571
rect 2455 9568 2467 9571
rect 2866 9568 2872 9580
rect 2455 9540 2872 9568
rect 2455 9537 2467 9540
rect 2409 9531 2467 9537
rect 2516 9509 2544 9540
rect 2866 9528 2872 9540
rect 2924 9528 2930 9580
rect 5736 9568 5764 9676
rect 6822 9664 6828 9676
rect 6880 9664 6886 9716
rect 7650 9704 7656 9716
rect 7611 9676 7656 9704
rect 7650 9664 7656 9676
rect 7708 9664 7714 9716
rect 11882 9704 11888 9716
rect 11843 9676 11888 9704
rect 11882 9664 11888 9676
rect 11940 9664 11946 9716
rect 15286 9704 15292 9716
rect 15120 9676 15292 9704
rect 9950 9596 9956 9648
rect 10008 9636 10014 9648
rect 10413 9639 10471 9645
rect 10413 9636 10425 9639
rect 10008 9608 10425 9636
rect 10008 9596 10014 9608
rect 10413 9605 10425 9608
rect 10459 9605 10471 9639
rect 13814 9636 13820 9648
rect 13775 9608 13820 9636
rect 10413 9599 10471 9605
rect 13814 9596 13820 9608
rect 13872 9596 13878 9648
rect 13998 9596 14004 9648
rect 14056 9636 14062 9648
rect 15013 9639 15071 9645
rect 15013 9636 15025 9639
rect 14056 9608 15025 9636
rect 14056 9596 14062 9608
rect 15013 9605 15025 9608
rect 15059 9605 15071 9639
rect 15013 9599 15071 9605
rect 5460 9540 5764 9568
rect 9861 9571 9919 9577
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9469 1455 9503
rect 1397 9463 1455 9469
rect 2507 9503 2565 9509
rect 2507 9469 2519 9503
rect 2553 9469 2565 9503
rect 2507 9463 2565 9469
rect 4157 9503 4215 9509
rect 4157 9469 4169 9503
rect 4203 9500 4215 9503
rect 4246 9500 4252 9512
rect 4203 9472 4252 9500
rect 4203 9469 4215 9472
rect 4157 9463 4215 9469
rect 1412 9432 1440 9463
rect 4246 9460 4252 9472
rect 4304 9460 4310 9512
rect 4338 9460 4344 9512
rect 4396 9500 4402 9512
rect 4516 9503 4574 9509
rect 4516 9500 4528 9503
rect 4396 9472 4528 9500
rect 4396 9460 4402 9472
rect 4516 9469 4528 9472
rect 4562 9500 4574 9503
rect 5460 9500 5488 9540
rect 9861 9537 9873 9571
rect 9907 9568 9919 9571
rect 10962 9568 10968 9580
rect 9907 9540 10968 9568
rect 9907 9537 9919 9540
rect 9861 9531 9919 9537
rect 10962 9528 10968 9540
rect 11020 9528 11026 9580
rect 11146 9528 11152 9580
rect 11204 9568 11210 9580
rect 11517 9571 11575 9577
rect 11517 9568 11529 9571
rect 11204 9540 11529 9568
rect 11204 9528 11210 9540
rect 11517 9537 11529 9540
rect 11563 9568 11575 9571
rect 14461 9571 14519 9577
rect 11563 9540 12572 9568
rect 11563 9537 11575 9540
rect 11517 9531 11575 9537
rect 4562 9472 5488 9500
rect 4562 9469 4574 9472
rect 4516 9463 4574 9469
rect 6086 9460 6092 9512
rect 6144 9500 6150 9512
rect 7837 9503 7895 9509
rect 7837 9500 7849 9503
rect 6144 9472 7849 9500
rect 6144 9460 6150 9472
rect 7837 9469 7849 9472
rect 7883 9500 7895 9503
rect 7926 9500 7932 9512
rect 7883 9472 7932 9500
rect 7883 9469 7895 9472
rect 7837 9463 7895 9469
rect 7926 9460 7932 9472
rect 7984 9460 7990 9512
rect 8104 9503 8162 9509
rect 8104 9469 8116 9503
rect 8150 9500 8162 9503
rect 8386 9500 8392 9512
rect 8150 9472 8392 9500
rect 8150 9469 8162 9472
rect 8104 9463 8162 9469
rect 8386 9460 8392 9472
rect 8444 9460 8450 9512
rect 11054 9500 11060 9512
rect 10704 9472 11060 9500
rect 2041 9435 2099 9441
rect 2041 9432 2053 9435
rect 1412 9404 2053 9432
rect 2041 9401 2053 9404
rect 2087 9432 2099 9435
rect 2866 9432 2872 9444
rect 2087 9404 2872 9432
rect 2087 9401 2099 9404
rect 2041 9395 2099 9401
rect 2866 9392 2872 9404
rect 2924 9392 2930 9444
rect 7377 9435 7435 9441
rect 7377 9401 7389 9435
rect 7423 9432 7435 9435
rect 8202 9432 8208 9444
rect 7423 9404 8208 9432
rect 7423 9401 7435 9404
rect 7377 9395 7435 9401
rect 8202 9392 8208 9404
rect 8260 9392 8266 9444
rect 9490 9392 9496 9444
rect 9548 9432 9554 9444
rect 10704 9441 10732 9472
rect 11054 9460 11060 9472
rect 11112 9460 11118 9512
rect 12158 9500 12164 9512
rect 12119 9472 12164 9500
rect 12158 9460 12164 9472
rect 12216 9460 12222 9512
rect 12437 9503 12495 9509
rect 12437 9469 12449 9503
rect 12483 9469 12495 9503
rect 12544 9500 12572 9540
rect 14461 9537 14473 9571
rect 14507 9568 14519 9571
rect 15120 9568 15148 9676
rect 15286 9664 15292 9676
rect 15344 9664 15350 9716
rect 15654 9664 15660 9716
rect 15712 9704 15718 9716
rect 15933 9707 15991 9713
rect 15933 9704 15945 9707
rect 15712 9676 15945 9704
rect 15712 9664 15718 9676
rect 15933 9673 15945 9676
rect 15979 9673 15991 9707
rect 15933 9667 15991 9673
rect 16666 9664 16672 9716
rect 16724 9704 16730 9716
rect 17494 9704 17500 9716
rect 16724 9676 17500 9704
rect 16724 9664 16730 9676
rect 17494 9664 17500 9676
rect 17552 9664 17558 9716
rect 20714 9704 20720 9716
rect 20675 9676 20720 9704
rect 20714 9664 20720 9676
rect 20772 9664 20778 9716
rect 20898 9704 20904 9716
rect 20859 9676 20904 9704
rect 20898 9664 20904 9676
rect 20956 9664 20962 9716
rect 23290 9664 23296 9716
rect 23348 9704 23354 9716
rect 23477 9707 23535 9713
rect 23348 9676 23428 9704
rect 23348 9664 23354 9676
rect 15746 9636 15752 9648
rect 15396 9608 15752 9636
rect 15396 9577 15424 9608
rect 15746 9596 15752 9608
rect 15804 9596 15810 9648
rect 18138 9636 18144 9648
rect 18099 9608 18144 9636
rect 18138 9596 18144 9608
rect 18196 9596 18202 9648
rect 19150 9636 19156 9648
rect 19111 9608 19156 9636
rect 19150 9596 19156 9608
rect 19208 9596 19214 9648
rect 19426 9596 19432 9648
rect 19484 9636 19490 9648
rect 19521 9639 19579 9645
rect 19521 9636 19533 9639
rect 19484 9608 19533 9636
rect 19484 9596 19490 9608
rect 19521 9605 19533 9608
rect 19567 9605 19579 9639
rect 19521 9599 19579 9605
rect 20349 9639 20407 9645
rect 20349 9605 20361 9639
rect 20395 9636 20407 9639
rect 20438 9636 20444 9648
rect 20395 9608 20444 9636
rect 20395 9605 20407 9608
rect 20349 9599 20407 9605
rect 20438 9596 20444 9608
rect 20496 9636 20502 9648
rect 21726 9636 21732 9648
rect 20496 9608 21732 9636
rect 20496 9596 20502 9608
rect 21726 9596 21732 9608
rect 21784 9596 21790 9648
rect 23014 9636 23020 9648
rect 22975 9608 23020 9636
rect 23014 9596 23020 9608
rect 23072 9596 23078 9648
rect 23400 9636 23428 9676
rect 23477 9673 23489 9707
rect 23523 9704 23535 9707
rect 23566 9704 23572 9716
rect 23523 9676 23572 9704
rect 23523 9673 23535 9676
rect 23477 9667 23535 9673
rect 23566 9664 23572 9676
rect 23624 9664 23630 9716
rect 24946 9704 24952 9716
rect 24907 9676 24952 9704
rect 24946 9664 24952 9676
rect 25004 9664 25010 9716
rect 23750 9636 23756 9648
rect 23400 9608 23612 9636
rect 23711 9608 23756 9636
rect 14507 9540 15148 9568
rect 15381 9571 15439 9577
rect 14507 9537 14519 9540
rect 14461 9531 14519 9537
rect 15381 9537 15393 9571
rect 15427 9537 15439 9571
rect 15562 9568 15568 9580
rect 15523 9540 15568 9568
rect 15381 9531 15439 9537
rect 14829 9503 14887 9509
rect 12544 9472 12664 9500
rect 12437 9463 12495 9469
rect 10689 9435 10747 9441
rect 10689 9432 10701 9435
rect 9548 9404 10701 9432
rect 9548 9392 9554 9404
rect 10689 9401 10701 9404
rect 10735 9401 10747 9435
rect 10870 9432 10876 9444
rect 10831 9404 10876 9432
rect 10689 9395 10747 9401
rect 10870 9392 10876 9404
rect 10928 9392 10934 9444
rect 10965 9435 11023 9441
rect 10965 9401 10977 9435
rect 11011 9401 11023 9435
rect 10965 9395 11023 9401
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 2774 9324 2780 9376
rect 2832 9364 2838 9376
rect 3145 9367 3203 9373
rect 3145 9364 3157 9367
rect 2832 9336 3157 9364
rect 2832 9324 2838 9336
rect 3145 9333 3157 9336
rect 3191 9364 3203 9367
rect 3234 9364 3240 9376
rect 3191 9336 3240 9364
rect 3191 9333 3203 9336
rect 3145 9327 3203 9333
rect 3234 9324 3240 9336
rect 3292 9324 3298 9376
rect 6270 9364 6276 9376
rect 6231 9336 6276 9364
rect 6270 9324 6276 9336
rect 6328 9324 6334 9376
rect 6825 9367 6883 9373
rect 6825 9333 6837 9367
rect 6871 9364 6883 9367
rect 7190 9364 7196 9376
rect 6871 9336 7196 9364
rect 6871 9333 6883 9336
rect 6825 9327 6883 9333
rect 7190 9324 7196 9336
rect 7248 9324 7254 9376
rect 9214 9364 9220 9376
rect 9175 9336 9220 9364
rect 9214 9324 9220 9336
rect 9272 9324 9278 9376
rect 10134 9364 10140 9376
rect 10095 9336 10140 9364
rect 10134 9324 10140 9336
rect 10192 9364 10198 9376
rect 10980 9364 11008 9395
rect 11698 9392 11704 9444
rect 11756 9432 11762 9444
rect 12342 9432 12348 9444
rect 11756 9404 12348 9432
rect 11756 9392 11762 9404
rect 12342 9392 12348 9404
rect 12400 9432 12406 9444
rect 12452 9432 12480 9463
rect 12400 9404 12480 9432
rect 12636 9432 12664 9472
rect 14829 9469 14841 9503
rect 14875 9500 14887 9503
rect 15396 9500 15424 9531
rect 15562 9528 15568 9540
rect 15620 9528 15626 9580
rect 16945 9571 17003 9577
rect 16945 9537 16957 9571
rect 16991 9568 17003 9571
rect 17770 9568 17776 9580
rect 16991 9540 17776 9568
rect 16991 9537 17003 9540
rect 16945 9531 17003 9537
rect 17770 9528 17776 9540
rect 17828 9528 17834 9580
rect 18693 9571 18751 9577
rect 18693 9537 18705 9571
rect 18739 9568 18751 9571
rect 18782 9568 18788 9580
rect 18739 9540 18788 9568
rect 18739 9537 18751 9540
rect 18693 9531 18751 9537
rect 18782 9528 18788 9540
rect 18840 9528 18846 9580
rect 19981 9571 20039 9577
rect 19981 9537 19993 9571
rect 20027 9568 20039 9571
rect 21453 9571 21511 9577
rect 21453 9568 21465 9571
rect 20027 9540 21465 9568
rect 20027 9537 20039 9540
rect 19981 9531 20039 9537
rect 21453 9537 21465 9540
rect 21499 9568 21511 9571
rect 22002 9568 22008 9580
rect 21499 9540 22008 9568
rect 21499 9537 21511 9540
rect 21453 9531 21511 9537
rect 22002 9528 22008 9540
rect 22060 9528 22066 9580
rect 22370 9568 22376 9580
rect 22331 9540 22376 9568
rect 22370 9528 22376 9540
rect 22428 9528 22434 9580
rect 23584 9568 23612 9608
rect 23750 9596 23756 9608
rect 23808 9596 23814 9648
rect 25409 9639 25467 9645
rect 25409 9605 25421 9639
rect 25455 9636 25467 9639
rect 25498 9636 25504 9648
rect 25455 9608 25504 9636
rect 25455 9605 25467 9608
rect 25409 9599 25467 9605
rect 25498 9596 25504 9608
rect 25556 9596 25562 9648
rect 24305 9571 24363 9577
rect 24305 9568 24317 9571
rect 23584 9540 24317 9568
rect 24305 9537 24317 9540
rect 24351 9537 24363 9571
rect 24305 9531 24363 9537
rect 14875 9472 15424 9500
rect 16853 9503 16911 9509
rect 14875 9469 14887 9472
rect 14829 9463 14887 9469
rect 16853 9469 16865 9503
rect 16899 9500 16911 9503
rect 16899 9472 18644 9500
rect 16899 9469 16911 9472
rect 16853 9463 16911 9469
rect 12704 9435 12762 9441
rect 12704 9432 12716 9435
rect 12636 9404 12716 9432
rect 12400 9392 12406 9404
rect 12704 9401 12716 9404
rect 12750 9432 12762 9435
rect 13078 9432 13084 9444
rect 12750 9404 13084 9432
rect 12750 9401 12762 9404
rect 12704 9395 12762 9401
rect 13078 9392 13084 9404
rect 13136 9392 13142 9444
rect 15470 9432 15476 9444
rect 15431 9404 15476 9432
rect 15470 9392 15476 9404
rect 15528 9392 15534 9444
rect 17218 9392 17224 9444
rect 17276 9432 17282 9444
rect 18046 9432 18052 9444
rect 17276 9404 18052 9432
rect 17276 9392 17282 9404
rect 18046 9392 18052 9404
rect 18104 9432 18110 9444
rect 18417 9435 18475 9441
rect 18417 9432 18429 9435
rect 18104 9404 18429 9432
rect 18104 9392 18110 9404
rect 18417 9401 18429 9404
rect 18463 9401 18475 9435
rect 18417 9395 18475 9401
rect 11974 9364 11980 9376
rect 10192 9336 11980 9364
rect 10192 9324 10198 9336
rect 11974 9324 11980 9336
rect 12032 9324 12038 9376
rect 18616 9373 18644 9472
rect 20714 9460 20720 9512
rect 20772 9500 20778 9512
rect 21177 9503 21235 9509
rect 21177 9500 21189 9503
rect 20772 9472 21189 9500
rect 20772 9460 20778 9472
rect 21177 9469 21189 9472
rect 21223 9500 21235 9503
rect 22189 9503 22247 9509
rect 22189 9500 22201 9503
rect 21223 9472 22201 9500
rect 21223 9469 21235 9472
rect 21177 9463 21235 9469
rect 22189 9469 22201 9472
rect 22235 9469 22247 9503
rect 22189 9463 22247 9469
rect 25038 9460 25044 9512
rect 25096 9500 25102 9512
rect 25225 9503 25283 9509
rect 25225 9500 25237 9503
rect 25096 9472 25237 9500
rect 25096 9460 25102 9472
rect 25225 9469 25237 9472
rect 25271 9500 25283 9503
rect 25777 9503 25835 9509
rect 25777 9500 25789 9503
rect 25271 9472 25789 9500
rect 25271 9469 25283 9472
rect 25225 9463 25283 9469
rect 25777 9469 25789 9472
rect 25823 9469 25835 9503
rect 25777 9463 25835 9469
rect 22922 9392 22928 9444
rect 22980 9432 22986 9444
rect 24029 9435 24087 9441
rect 24029 9432 24041 9435
rect 22980 9404 24041 9432
rect 22980 9392 22986 9404
rect 24029 9401 24041 9404
rect 24075 9401 24087 9435
rect 24029 9395 24087 9401
rect 24213 9435 24271 9441
rect 24213 9401 24225 9435
rect 24259 9432 24271 9435
rect 24762 9432 24768 9444
rect 24259 9404 24768 9432
rect 24259 9401 24271 9404
rect 24213 9395 24271 9401
rect 18601 9367 18659 9373
rect 18601 9333 18613 9367
rect 18647 9364 18659 9367
rect 18874 9364 18880 9376
rect 18647 9336 18880 9364
rect 18647 9333 18659 9336
rect 18601 9327 18659 9333
rect 18874 9324 18880 9336
rect 18932 9324 18938 9376
rect 21082 9324 21088 9376
rect 21140 9364 21146 9376
rect 21361 9367 21419 9373
rect 21361 9364 21373 9367
rect 21140 9336 21373 9364
rect 21140 9324 21146 9336
rect 21361 9333 21373 9336
rect 21407 9364 21419 9367
rect 21821 9367 21879 9373
rect 21821 9364 21833 9367
rect 21407 9336 21833 9364
rect 21407 9333 21419 9336
rect 21361 9327 21419 9333
rect 21821 9333 21833 9336
rect 21867 9333 21879 9367
rect 21821 9327 21879 9333
rect 23106 9324 23112 9376
rect 23164 9364 23170 9376
rect 24228 9364 24256 9395
rect 24762 9392 24768 9404
rect 24820 9392 24826 9444
rect 23164 9336 24256 9364
rect 23164 9324 23170 9336
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1394 9120 1400 9172
rect 1452 9160 1458 9172
rect 1949 9163 2007 9169
rect 1949 9160 1961 9163
rect 1452 9132 1961 9160
rect 1452 9120 1458 9132
rect 1949 9129 1961 9132
rect 1995 9129 2007 9163
rect 4338 9160 4344 9172
rect 4299 9132 4344 9160
rect 1949 9123 2007 9129
rect 4338 9120 4344 9132
rect 4396 9120 4402 9172
rect 5166 9160 5172 9172
rect 5127 9132 5172 9160
rect 5166 9120 5172 9132
rect 5224 9120 5230 9172
rect 6914 9120 6920 9172
rect 6972 9160 6978 9172
rect 7653 9163 7711 9169
rect 7653 9160 7665 9163
rect 6972 9132 7665 9160
rect 6972 9120 6978 9132
rect 7653 9129 7665 9132
rect 7699 9129 7711 9163
rect 7653 9123 7711 9129
rect 7926 9120 7932 9172
rect 7984 9160 7990 9172
rect 8205 9163 8263 9169
rect 8205 9160 8217 9163
rect 7984 9132 8217 9160
rect 7984 9120 7990 9132
rect 8205 9129 8217 9132
rect 8251 9129 8263 9163
rect 9490 9160 9496 9172
rect 9451 9132 9496 9160
rect 8205 9123 8263 9129
rect 9490 9120 9496 9132
rect 9548 9120 9554 9172
rect 10137 9163 10195 9169
rect 10137 9129 10149 9163
rect 10183 9160 10195 9163
rect 10870 9160 10876 9172
rect 10183 9132 10876 9160
rect 10183 9129 10195 9132
rect 10137 9123 10195 9129
rect 10870 9120 10876 9132
rect 10928 9120 10934 9172
rect 11974 9160 11980 9172
rect 11935 9132 11980 9160
rect 11974 9120 11980 9132
rect 12032 9120 12038 9172
rect 13630 9160 13636 9172
rect 13591 9132 13636 9160
rect 13630 9120 13636 9132
rect 13688 9120 13694 9172
rect 14182 9160 14188 9172
rect 14143 9132 14188 9160
rect 14182 9120 14188 9132
rect 14240 9120 14246 9172
rect 15013 9163 15071 9169
rect 15013 9129 15025 9163
rect 15059 9160 15071 9163
rect 15470 9160 15476 9172
rect 15059 9132 15476 9160
rect 15059 9129 15071 9132
rect 15013 9123 15071 9129
rect 15470 9120 15476 9132
rect 15528 9120 15534 9172
rect 15565 9163 15623 9169
rect 15565 9129 15577 9163
rect 15611 9160 15623 9163
rect 15838 9160 15844 9172
rect 15611 9132 15844 9160
rect 15611 9129 15623 9132
rect 15565 9123 15623 9129
rect 15838 9120 15844 9132
rect 15896 9120 15902 9172
rect 17218 9160 17224 9172
rect 17179 9132 17224 9160
rect 17218 9120 17224 9132
rect 17276 9120 17282 9172
rect 17589 9163 17647 9169
rect 17589 9129 17601 9163
rect 17635 9160 17647 9163
rect 17678 9160 17684 9172
rect 17635 9132 17684 9160
rect 17635 9129 17647 9132
rect 17589 9123 17647 9129
rect 17678 9120 17684 9132
rect 17736 9120 17742 9172
rect 18141 9163 18199 9169
rect 18141 9129 18153 9163
rect 18187 9160 18199 9163
rect 18690 9160 18696 9172
rect 18187 9132 18696 9160
rect 18187 9129 18199 9132
rect 18141 9123 18199 9129
rect 18690 9120 18696 9132
rect 18748 9120 18754 9172
rect 23106 9160 23112 9172
rect 23067 9132 23112 9160
rect 23106 9120 23112 9132
rect 23164 9120 23170 9172
rect 24118 9120 24124 9172
rect 24176 9160 24182 9172
rect 24213 9163 24271 9169
rect 24213 9160 24225 9163
rect 24176 9132 24225 9160
rect 24176 9120 24182 9132
rect 24213 9129 24225 9132
rect 24259 9129 24271 9163
rect 24946 9160 24952 9172
rect 24907 9132 24952 9160
rect 24213 9123 24271 9129
rect 24946 9120 24952 9132
rect 25004 9120 25010 9172
rect 4246 9052 4252 9104
rect 4304 9092 4310 9104
rect 4798 9092 4804 9104
rect 4304 9064 4804 9092
rect 4304 9052 4310 9064
rect 4798 9052 4804 9064
rect 4856 9052 4862 9104
rect 8665 9095 8723 9101
rect 8665 9061 8677 9095
rect 8711 9092 8723 9095
rect 10042 9092 10048 9104
rect 8711 9064 10048 9092
rect 8711 9061 8723 9064
rect 8665 9055 8723 9061
rect 10042 9052 10048 9064
rect 10100 9052 10106 9104
rect 10505 9095 10563 9101
rect 10505 9061 10517 9095
rect 10551 9092 10563 9095
rect 10686 9092 10692 9104
rect 10551 9064 10692 9092
rect 10551 9061 10563 9064
rect 10505 9055 10563 9061
rect 10686 9052 10692 9064
rect 10744 9052 10750 9104
rect 13449 9095 13507 9101
rect 13449 9061 13461 9095
rect 13495 9092 13507 9095
rect 13538 9092 13544 9104
rect 13495 9064 13544 9092
rect 13495 9061 13507 9064
rect 13449 9055 13507 9061
rect 13538 9052 13544 9064
rect 13596 9052 13602 9104
rect 18782 9092 18788 9104
rect 18743 9064 18788 9092
rect 18782 9052 18788 9064
rect 18840 9052 18846 9104
rect 21542 9092 21548 9104
rect 21503 9064 21548 9092
rect 21542 9052 21548 9064
rect 21600 9052 21606 9104
rect 23566 9092 23572 9104
rect 23527 9064 23572 9092
rect 23566 9052 23572 9064
rect 23624 9052 23630 9104
rect 23753 9095 23811 9101
rect 23753 9061 23765 9095
rect 23799 9092 23811 9095
rect 24670 9092 24676 9104
rect 23799 9064 24676 9092
rect 23799 9061 23811 9064
rect 23753 9055 23811 9061
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 2038 9024 2044 9036
rect 1443 8996 2044 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 2038 8984 2044 8996
rect 2096 8984 2102 9036
rect 4816 8956 4844 9052
rect 6178 8984 6184 9036
rect 6236 9024 6242 9036
rect 10870 9033 10876 9036
rect 6529 9027 6587 9033
rect 6529 9024 6541 9027
rect 6236 8996 6541 9024
rect 6236 8984 6242 8996
rect 6529 8993 6541 8996
rect 6575 8993 6587 9027
rect 10864 9024 10876 9033
rect 10831 8996 10876 9024
rect 6529 8987 6587 8993
rect 10864 8987 10876 8996
rect 10870 8984 10876 8987
rect 10928 8984 10934 9036
rect 12342 8984 12348 9036
rect 12400 9024 12406 9036
rect 12529 9027 12587 9033
rect 12529 9024 12541 9027
rect 12400 8996 12541 9024
rect 12400 8984 12406 8996
rect 12529 8993 12541 8996
rect 12575 8993 12587 9027
rect 12529 8987 12587 8993
rect 17954 8984 17960 9036
rect 18012 9024 18018 9036
rect 21358 9024 21364 9036
rect 18012 8996 18920 9024
rect 21319 8996 21364 9024
rect 18012 8984 18018 8996
rect 18892 8968 18920 8996
rect 21358 8984 21364 8996
rect 21416 8984 21422 9036
rect 23014 8984 23020 9036
rect 23072 9024 23078 9036
rect 23768 9024 23796 9055
rect 24670 9052 24676 9064
rect 24728 9052 24734 9104
rect 24762 9024 24768 9036
rect 23072 8996 23796 9024
rect 24723 8996 24768 9024
rect 23072 8984 23078 8996
rect 24762 8984 24768 8996
rect 24820 8984 24826 9036
rect 6086 8956 6092 8968
rect 4816 8928 6092 8956
rect 6086 8916 6092 8928
rect 6144 8956 6150 8968
rect 6273 8959 6331 8965
rect 6273 8956 6285 8959
rect 6144 8928 6285 8956
rect 6144 8916 6150 8928
rect 6273 8925 6285 8928
rect 6319 8925 6331 8959
rect 6273 8919 6331 8925
rect 10597 8959 10655 8965
rect 10597 8925 10609 8959
rect 10643 8925 10655 8959
rect 10597 8919 10655 8925
rect 13725 8959 13783 8965
rect 13725 8925 13737 8959
rect 13771 8925 13783 8959
rect 13725 8919 13783 8925
rect 1486 8780 1492 8832
rect 1544 8820 1550 8832
rect 1581 8823 1639 8829
rect 1581 8820 1593 8823
rect 1544 8792 1593 8820
rect 1544 8780 1550 8792
rect 1581 8789 1593 8792
rect 1627 8789 1639 8823
rect 1581 8783 1639 8789
rect 9306 8780 9312 8832
rect 9364 8820 9370 8832
rect 10612 8820 10640 8919
rect 13170 8888 13176 8900
rect 13131 8860 13176 8888
rect 13170 8848 13176 8860
rect 13228 8848 13234 8900
rect 11698 8820 11704 8832
rect 9364 8792 11704 8820
rect 9364 8780 9370 8792
rect 11698 8780 11704 8792
rect 11756 8780 11762 8832
rect 12989 8823 13047 8829
rect 12989 8789 13001 8823
rect 13035 8820 13047 8823
rect 13078 8820 13084 8832
rect 13035 8792 13084 8820
rect 13035 8789 13047 8792
rect 12989 8783 13047 8789
rect 13078 8780 13084 8792
rect 13136 8820 13142 8832
rect 13740 8820 13768 8919
rect 17310 8916 17316 8968
rect 17368 8956 17374 8968
rect 18693 8959 18751 8965
rect 18693 8956 18705 8959
rect 17368 8928 18705 8956
rect 17368 8916 17374 8928
rect 18693 8925 18705 8928
rect 18739 8925 18751 8959
rect 18874 8956 18880 8968
rect 18835 8928 18880 8956
rect 18693 8919 18751 8925
rect 18325 8891 18383 8897
rect 18325 8857 18337 8891
rect 18371 8888 18383 8891
rect 18598 8888 18604 8900
rect 18371 8860 18604 8888
rect 18371 8857 18383 8860
rect 18325 8851 18383 8857
rect 18598 8848 18604 8860
rect 18656 8848 18662 8900
rect 18708 8888 18736 8919
rect 18874 8916 18880 8928
rect 18932 8916 18938 8968
rect 21637 8959 21695 8965
rect 21637 8925 21649 8959
rect 21683 8956 21695 8959
rect 21726 8956 21732 8968
rect 21683 8928 21732 8956
rect 21683 8925 21695 8928
rect 21637 8919 21695 8925
rect 21726 8916 21732 8928
rect 21784 8916 21790 8968
rect 23842 8956 23848 8968
rect 23803 8928 23848 8956
rect 23842 8916 23848 8928
rect 23900 8916 23906 8968
rect 19150 8888 19156 8900
rect 18708 8860 19156 8888
rect 19150 8848 19156 8860
rect 19208 8848 19214 8900
rect 21082 8888 21088 8900
rect 21043 8860 21088 8888
rect 21082 8848 21088 8860
rect 21140 8848 21146 8900
rect 22922 8848 22928 8900
rect 22980 8888 22986 8900
rect 23293 8891 23351 8897
rect 23293 8888 23305 8891
rect 22980 8860 23305 8888
rect 22980 8848 22986 8860
rect 23293 8857 23305 8860
rect 23339 8857 23351 8891
rect 23293 8851 23351 8857
rect 13136 8792 13768 8820
rect 13136 8780 13142 8792
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1578 8616 1584 8628
rect 1539 8588 1584 8616
rect 1578 8576 1584 8588
rect 1636 8576 1642 8628
rect 2038 8616 2044 8628
rect 1999 8588 2044 8616
rect 2038 8576 2044 8588
rect 2096 8576 2102 8628
rect 5629 8619 5687 8625
rect 5629 8585 5641 8619
rect 5675 8616 5687 8619
rect 5905 8619 5963 8625
rect 5905 8616 5917 8619
rect 5675 8588 5917 8616
rect 5675 8585 5687 8588
rect 5629 8579 5687 8585
rect 5905 8585 5917 8588
rect 5951 8616 5963 8619
rect 6178 8616 6184 8628
rect 5951 8588 6184 8616
rect 5951 8585 5963 8588
rect 5905 8579 5963 8585
rect 6178 8576 6184 8588
rect 6236 8576 6242 8628
rect 6270 8576 6276 8628
rect 6328 8616 6334 8628
rect 6917 8619 6975 8625
rect 6917 8616 6929 8619
rect 6328 8588 6929 8616
rect 6328 8576 6334 8588
rect 6917 8585 6929 8588
rect 6963 8585 6975 8619
rect 6917 8579 6975 8585
rect 7926 8576 7932 8628
rect 7984 8616 7990 8628
rect 9217 8619 9275 8625
rect 9217 8616 9229 8619
rect 7984 8588 9229 8616
rect 7984 8576 7990 8588
rect 9217 8585 9229 8588
rect 9263 8616 9275 8619
rect 9306 8616 9312 8628
rect 9263 8588 9312 8616
rect 9263 8585 9275 8588
rect 9217 8579 9275 8585
rect 9306 8576 9312 8588
rect 9364 8576 9370 8628
rect 10042 8576 10048 8628
rect 10100 8616 10106 8628
rect 10781 8619 10839 8625
rect 10781 8616 10793 8619
rect 10100 8588 10793 8616
rect 10100 8576 10106 8588
rect 10781 8585 10793 8588
rect 10827 8585 10839 8619
rect 11790 8616 11796 8628
rect 11751 8588 11796 8616
rect 10781 8579 10839 8585
rect 11790 8576 11796 8588
rect 11848 8576 11854 8628
rect 13541 8619 13599 8625
rect 13541 8585 13553 8619
rect 13587 8616 13599 8619
rect 13630 8616 13636 8628
rect 13587 8588 13636 8616
rect 13587 8585 13599 8588
rect 13541 8579 13599 8585
rect 13630 8576 13636 8588
rect 13688 8576 13694 8628
rect 17865 8619 17923 8625
rect 17865 8585 17877 8619
rect 17911 8616 17923 8619
rect 18782 8616 18788 8628
rect 17911 8588 18788 8616
rect 17911 8585 17923 8588
rect 17865 8579 17923 8585
rect 18782 8576 18788 8588
rect 18840 8616 18846 8628
rect 21361 8619 21419 8625
rect 21361 8616 21373 8619
rect 18840 8588 21373 8616
rect 18840 8576 18846 8588
rect 21361 8585 21373 8588
rect 21407 8616 21419 8619
rect 21542 8616 21548 8628
rect 21407 8588 21548 8616
rect 21407 8585 21419 8588
rect 21361 8579 21419 8585
rect 21542 8576 21548 8588
rect 21600 8576 21606 8628
rect 21726 8616 21732 8628
rect 21687 8588 21732 8616
rect 21726 8576 21732 8588
rect 21784 8576 21790 8628
rect 22462 8576 22468 8628
rect 22520 8616 22526 8628
rect 23201 8619 23259 8625
rect 23201 8616 23213 8619
rect 22520 8588 23213 8616
rect 22520 8576 22526 8588
rect 23201 8585 23213 8588
rect 23247 8616 23259 8619
rect 23842 8616 23848 8628
rect 23247 8588 23848 8616
rect 23247 8585 23259 8588
rect 23201 8579 23259 8585
rect 23842 8576 23848 8588
rect 23900 8576 23906 8628
rect 24854 8616 24860 8628
rect 24815 8588 24860 8616
rect 24854 8576 24860 8588
rect 24912 8576 24918 8628
rect 25130 8616 25136 8628
rect 25091 8588 25136 8616
rect 25130 8576 25136 8588
rect 25188 8576 25194 8628
rect 6196 8480 6224 8576
rect 7469 8483 7527 8489
rect 7469 8480 7481 8483
rect 6196 8452 7481 8480
rect 7469 8449 7481 8452
rect 7515 8480 7527 8483
rect 9214 8480 9220 8492
rect 7515 8452 9220 8480
rect 7515 8449 7527 8452
rect 7469 8443 7527 8449
rect 9214 8440 9220 8452
rect 9272 8440 9278 8492
rect 1394 8412 1400 8424
rect 1355 8384 1400 8412
rect 1394 8372 1400 8384
rect 1452 8412 1458 8424
rect 2317 8415 2375 8421
rect 2317 8412 2329 8415
rect 1452 8384 2329 8412
rect 1452 8372 1458 8384
rect 2317 8381 2329 8384
rect 2363 8381 2375 8415
rect 2317 8375 2375 8381
rect 6086 8372 6092 8424
rect 6144 8412 6150 8424
rect 6273 8415 6331 8421
rect 6273 8412 6285 8415
rect 6144 8384 6285 8412
rect 6144 8372 6150 8384
rect 6273 8381 6285 8384
rect 6319 8381 6331 8415
rect 7190 8412 7196 8424
rect 7151 8384 7196 8412
rect 6273 8375 6331 8381
rect 7190 8372 7196 8384
rect 7248 8372 7254 8424
rect 9324 8412 9352 8576
rect 11425 8551 11483 8557
rect 11425 8517 11437 8551
rect 11471 8548 11483 8551
rect 11698 8548 11704 8560
rect 11471 8520 11704 8548
rect 11471 8517 11483 8520
rect 11425 8511 11483 8517
rect 11698 8508 11704 8520
rect 11756 8508 11762 8560
rect 11808 8480 11836 8576
rect 12434 8508 12440 8560
rect 12492 8548 12498 8560
rect 12529 8551 12587 8557
rect 12529 8548 12541 8551
rect 12492 8520 12541 8548
rect 12492 8508 12498 8520
rect 12529 8517 12541 8520
rect 12575 8517 12587 8551
rect 12529 8511 12587 8517
rect 14093 8551 14151 8557
rect 14093 8517 14105 8551
rect 14139 8517 14151 8551
rect 14093 8511 14151 8517
rect 22925 8551 22983 8557
rect 22925 8517 22937 8551
rect 22971 8548 22983 8551
rect 23014 8548 23020 8560
rect 22971 8520 23020 8548
rect 22971 8517 22983 8520
rect 22925 8511 22983 8517
rect 13081 8483 13139 8489
rect 13081 8480 13093 8483
rect 11808 8452 13093 8480
rect 13081 8449 13093 8452
rect 13127 8480 13139 8483
rect 13446 8480 13452 8492
rect 13127 8452 13452 8480
rect 13127 8449 13139 8452
rect 13081 8443 13139 8449
rect 13446 8440 13452 8452
rect 13504 8440 13510 8492
rect 9401 8415 9459 8421
rect 9401 8412 9413 8415
rect 9324 8384 9413 8412
rect 9401 8381 9413 8384
rect 9447 8381 9459 8415
rect 12250 8412 12256 8424
rect 12163 8384 12256 8412
rect 9401 8375 9459 8381
rect 12250 8372 12256 8384
rect 12308 8412 12314 8424
rect 12805 8415 12863 8421
rect 12805 8412 12817 8415
rect 12308 8384 12817 8412
rect 12308 8372 12314 8384
rect 12805 8381 12817 8384
rect 12851 8381 12863 8415
rect 14108 8412 14136 8511
rect 23014 8508 23020 8520
rect 23072 8508 23078 8560
rect 14458 8440 14464 8492
rect 14516 8480 14522 8492
rect 14645 8483 14703 8489
rect 14645 8480 14657 8483
rect 14516 8452 14657 8480
rect 14516 8440 14522 8452
rect 14645 8449 14657 8452
rect 14691 8449 14703 8483
rect 14645 8443 14703 8449
rect 21085 8483 21143 8489
rect 21085 8449 21097 8483
rect 21131 8480 21143 8483
rect 21358 8480 21364 8492
rect 21131 8452 21364 8480
rect 21131 8449 21143 8452
rect 21085 8443 21143 8449
rect 21358 8440 21364 8452
rect 21416 8440 21422 8492
rect 12805 8375 12863 8381
rect 13004 8384 14136 8412
rect 7650 8304 7656 8356
rect 7708 8344 7714 8356
rect 8386 8344 8392 8356
rect 7708 8316 8392 8344
rect 7708 8304 7714 8316
rect 8386 8304 8392 8316
rect 8444 8304 8450 8356
rect 9490 8304 9496 8356
rect 9548 8344 9554 8356
rect 9646 8347 9704 8353
rect 9646 8344 9658 8347
rect 9548 8316 9658 8344
rect 9548 8304 9554 8316
rect 9646 8313 9658 8316
rect 9692 8344 9704 8347
rect 10134 8344 10140 8356
rect 9692 8316 10140 8344
rect 9692 8313 9704 8316
rect 9646 8307 9704 8313
rect 10134 8304 10140 8316
rect 10192 8304 10198 8356
rect 12710 8304 12716 8356
rect 12768 8344 12774 8356
rect 13004 8353 13032 8384
rect 14182 8372 14188 8424
rect 14240 8412 14246 8424
rect 14369 8415 14427 8421
rect 14369 8412 14381 8415
rect 14240 8384 14381 8412
rect 14240 8372 14246 8384
rect 14369 8381 14381 8384
rect 14415 8381 14427 8415
rect 14369 8375 14427 8381
rect 17497 8415 17555 8421
rect 17497 8381 17509 8415
rect 17543 8412 17555 8415
rect 18138 8412 18144 8424
rect 17543 8384 18144 8412
rect 17543 8381 17555 8384
rect 17497 8375 17555 8381
rect 18138 8372 18144 8384
rect 18196 8412 18202 8424
rect 18233 8415 18291 8421
rect 18233 8412 18245 8415
rect 18196 8384 18245 8412
rect 18196 8372 18202 8384
rect 18233 8381 18245 8384
rect 18279 8381 18291 8415
rect 23658 8412 23664 8424
rect 23619 8384 23664 8412
rect 18233 8375 18291 8381
rect 23658 8372 23664 8384
rect 23716 8412 23722 8424
rect 24397 8415 24455 8421
rect 24397 8412 24409 8415
rect 23716 8384 24409 8412
rect 23716 8372 23722 8384
rect 24397 8381 24409 8384
rect 24443 8381 24455 8415
rect 24946 8412 24952 8424
rect 24907 8384 24952 8412
rect 24397 8375 24455 8381
rect 24946 8372 24952 8384
rect 25004 8412 25010 8424
rect 25501 8415 25559 8421
rect 25501 8412 25513 8415
rect 25004 8384 25513 8412
rect 25004 8372 25010 8384
rect 25501 8381 25513 8384
rect 25547 8381 25559 8415
rect 25501 8375 25559 8381
rect 12989 8347 13047 8353
rect 12989 8344 13001 8347
rect 12768 8316 13001 8344
rect 12768 8304 12774 8316
rect 12989 8313 13001 8316
rect 13035 8313 13047 8347
rect 12989 8307 13047 8313
rect 13909 8347 13967 8353
rect 13909 8313 13921 8347
rect 13955 8344 13967 8347
rect 14090 8344 14096 8356
rect 13955 8316 14096 8344
rect 13955 8313 13967 8316
rect 13909 8307 13967 8313
rect 14090 8304 14096 8316
rect 14148 8344 14154 8356
rect 14550 8344 14556 8356
rect 14148 8316 14556 8344
rect 14148 8304 14154 8316
rect 14550 8304 14556 8316
rect 14608 8304 14614 8356
rect 18506 8344 18512 8356
rect 18467 8316 18512 8344
rect 18506 8304 18512 8316
rect 18564 8304 18570 8356
rect 19061 8347 19119 8353
rect 19061 8313 19073 8347
rect 19107 8344 19119 8347
rect 19150 8344 19156 8356
rect 19107 8316 19156 8344
rect 19107 8313 19119 8316
rect 19061 8307 19119 8313
rect 19150 8304 19156 8316
rect 19208 8304 19214 8356
rect 23934 8344 23940 8356
rect 23895 8316 23940 8344
rect 23934 8304 23940 8316
rect 23992 8304 23998 8356
rect 7374 8276 7380 8288
rect 7287 8248 7380 8276
rect 7374 8236 7380 8248
rect 7432 8276 7438 8288
rect 7834 8276 7840 8288
rect 7432 8248 7840 8276
rect 7432 8236 7438 8248
rect 7834 8236 7840 8248
rect 7892 8236 7898 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1578 8072 1584 8084
rect 1539 8044 1584 8072
rect 1578 8032 1584 8044
rect 1636 8032 1642 8084
rect 6457 8075 6515 8081
rect 6457 8041 6469 8075
rect 6503 8072 6515 8075
rect 6730 8072 6736 8084
rect 6503 8044 6736 8072
rect 6503 8041 6515 8044
rect 6457 8035 6515 8041
rect 6730 8032 6736 8044
rect 6788 8032 6794 8084
rect 7009 8075 7067 8081
rect 7009 8041 7021 8075
rect 7055 8072 7067 8075
rect 7190 8072 7196 8084
rect 7055 8044 7196 8072
rect 7055 8041 7067 8044
rect 7009 8035 7067 8041
rect 7190 8032 7196 8044
rect 7248 8032 7254 8084
rect 7374 8072 7380 8084
rect 7335 8044 7380 8072
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 8103 8075 8161 8081
rect 8103 8041 8115 8075
rect 8149 8072 8161 8075
rect 9858 8072 9864 8084
rect 8149 8044 9864 8072
rect 8149 8041 8161 8044
rect 8103 8035 8161 8041
rect 9858 8032 9864 8044
rect 9916 8072 9922 8084
rect 10229 8075 10287 8081
rect 10229 8072 10241 8075
rect 9916 8044 10241 8072
rect 9916 8032 9922 8044
rect 10229 8041 10241 8044
rect 10275 8041 10287 8075
rect 10229 8035 10287 8041
rect 10781 8075 10839 8081
rect 10781 8041 10793 8075
rect 10827 8072 10839 8075
rect 10870 8072 10876 8084
rect 10827 8044 10876 8072
rect 10827 8041 10839 8044
rect 10781 8035 10839 8041
rect 10870 8032 10876 8044
rect 10928 8032 10934 8084
rect 13906 8032 13912 8084
rect 13964 8072 13970 8084
rect 14001 8075 14059 8081
rect 14001 8072 14013 8075
rect 13964 8044 14013 8072
rect 13964 8032 13970 8044
rect 14001 8041 14013 8044
rect 14047 8041 14059 8075
rect 14458 8072 14464 8084
rect 14419 8044 14464 8072
rect 14001 8035 14059 8041
rect 14458 8032 14464 8044
rect 14516 8032 14522 8084
rect 18325 8075 18383 8081
rect 18325 8041 18337 8075
rect 18371 8072 18383 8075
rect 18874 8072 18880 8084
rect 18371 8044 18880 8072
rect 18371 8041 18383 8044
rect 18325 8035 18383 8041
rect 18874 8032 18880 8044
rect 18932 8032 18938 8084
rect 23293 8075 23351 8081
rect 23293 8041 23305 8075
rect 23339 8072 23351 8075
rect 23382 8072 23388 8084
rect 23339 8044 23388 8072
rect 23339 8041 23351 8044
rect 23293 8035 23351 8041
rect 23382 8032 23388 8044
rect 23440 8032 23446 8084
rect 24762 8072 24768 8084
rect 24723 8044 24768 8072
rect 24762 8032 24768 8044
rect 24820 8032 24826 8084
rect 6549 8007 6607 8013
rect 6549 7973 6561 8007
rect 6595 8004 6607 8007
rect 6822 8004 6828 8016
rect 6595 7976 6828 8004
rect 6595 7973 6607 7976
rect 6549 7967 6607 7973
rect 6822 7964 6828 7976
rect 6880 7964 6886 8016
rect 7926 7964 7932 8016
rect 7984 8004 7990 8016
rect 8478 8004 8484 8016
rect 7984 7976 8484 8004
rect 7984 7964 7990 7976
rect 8478 7964 8484 7976
rect 8536 8004 8542 8016
rect 8573 8007 8631 8013
rect 8573 8004 8585 8007
rect 8536 7976 8585 8004
rect 8536 7964 8542 7976
rect 8573 7973 8585 7976
rect 8619 7973 8631 8007
rect 9490 8004 9496 8016
rect 9451 7976 9496 8004
rect 8573 7967 8631 7973
rect 9490 7964 9496 7976
rect 9548 7964 9554 8016
rect 11606 7964 11612 8016
rect 11664 8004 11670 8016
rect 12437 8007 12495 8013
rect 12437 8004 12449 8007
rect 11664 7976 12449 8004
rect 11664 7964 11670 7976
rect 12437 7973 12449 7976
rect 12483 8004 12495 8007
rect 13523 8007 13581 8013
rect 13523 8004 13535 8007
rect 12483 7976 13535 8004
rect 12483 7973 12495 7976
rect 12437 7967 12495 7973
rect 13523 7973 13535 7976
rect 13569 7973 13581 8007
rect 13523 7967 13581 7973
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 2038 7936 2044 7948
rect 1443 7908 2044 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 2038 7896 2044 7908
rect 2096 7896 2102 7948
rect 8294 7896 8300 7948
rect 8352 7936 8358 7948
rect 8389 7939 8447 7945
rect 8389 7936 8401 7939
rect 8352 7908 8401 7936
rect 8352 7896 8358 7908
rect 8389 7905 8401 7908
rect 8435 7905 8447 7939
rect 8389 7899 8447 7905
rect 9674 7896 9680 7948
rect 9732 7936 9738 7948
rect 10045 7939 10103 7945
rect 10045 7936 10057 7939
rect 9732 7908 10057 7936
rect 9732 7896 9738 7908
rect 10045 7905 10057 7908
rect 10091 7905 10103 7939
rect 12250 7936 12256 7948
rect 12211 7908 12256 7936
rect 10045 7899 10103 7905
rect 12250 7896 12256 7908
rect 12308 7896 12314 7948
rect 16574 7896 16580 7948
rect 16632 7936 16638 7948
rect 16942 7936 16948 7948
rect 16632 7908 16948 7936
rect 16632 7896 16638 7908
rect 16942 7896 16948 7908
rect 17000 7896 17006 7948
rect 23477 7939 23535 7945
rect 23477 7905 23489 7939
rect 23523 7936 23535 7939
rect 23934 7936 23940 7948
rect 23523 7908 23940 7936
rect 23523 7905 23535 7908
rect 23477 7899 23535 7905
rect 23934 7896 23940 7908
rect 23992 7896 23998 7948
rect 24026 7896 24032 7948
rect 24084 7936 24090 7948
rect 24581 7939 24639 7945
rect 24581 7936 24593 7939
rect 24084 7908 24593 7936
rect 24084 7896 24090 7908
rect 24581 7905 24593 7908
rect 24627 7905 24639 7939
rect 24581 7899 24639 7905
rect 6454 7868 6460 7880
rect 6415 7840 6460 7868
rect 6454 7828 6460 7840
rect 6512 7828 6518 7880
rect 8662 7868 8668 7880
rect 8623 7840 8668 7868
rect 8662 7828 8668 7840
rect 8720 7828 8726 7880
rect 10318 7868 10324 7880
rect 10231 7840 10324 7868
rect 10318 7828 10324 7840
rect 10376 7868 10382 7880
rect 12066 7868 12072 7880
rect 10376 7840 12072 7868
rect 10376 7828 10382 7840
rect 12066 7828 12072 7840
rect 12124 7868 12130 7880
rect 12529 7871 12587 7877
rect 12529 7868 12541 7871
rect 12124 7840 12541 7868
rect 12124 7828 12130 7840
rect 12529 7837 12541 7840
rect 12575 7868 12587 7871
rect 12618 7868 12624 7880
rect 12575 7840 12624 7868
rect 12575 7837 12587 7840
rect 12529 7831 12587 7837
rect 12618 7828 12624 7840
rect 12676 7828 12682 7880
rect 13173 7871 13231 7877
rect 13173 7837 13185 7871
rect 13219 7868 13231 7871
rect 13538 7868 13544 7880
rect 13219 7840 13544 7868
rect 13219 7837 13231 7840
rect 13173 7831 13231 7837
rect 13538 7828 13544 7840
rect 13596 7828 13602 7880
rect 13998 7868 14004 7880
rect 13959 7840 14004 7868
rect 13998 7828 14004 7840
rect 14056 7828 14062 7880
rect 14093 7871 14151 7877
rect 14093 7837 14105 7871
rect 14139 7837 14151 7871
rect 17218 7868 17224 7880
rect 17179 7840 17224 7868
rect 14093 7831 14151 7837
rect 5442 7760 5448 7812
rect 5500 7800 5506 7812
rect 5997 7803 6055 7809
rect 5997 7800 6009 7803
rect 5500 7772 6009 7800
rect 5500 7760 5506 7772
rect 5997 7769 6009 7772
rect 6043 7769 6055 7803
rect 9766 7800 9772 7812
rect 9727 7772 9772 7800
rect 5997 7763 6055 7769
rect 9766 7760 9772 7772
rect 9824 7760 9830 7812
rect 13446 7760 13452 7812
rect 13504 7800 13510 7812
rect 14108 7800 14136 7831
rect 17218 7828 17224 7840
rect 17276 7828 17282 7880
rect 13504 7772 14136 7800
rect 13504 7760 13510 7772
rect 11974 7732 11980 7744
rect 11935 7704 11980 7732
rect 11974 7692 11980 7704
rect 12032 7692 12038 7744
rect 23658 7732 23664 7744
rect 23619 7704 23664 7732
rect 23658 7692 23664 7704
rect 23716 7692 23722 7744
rect 23842 7692 23848 7744
rect 23900 7732 23906 7744
rect 24118 7732 24124 7744
rect 23900 7704 24124 7732
rect 23900 7692 23906 7704
rect 24118 7692 24124 7704
rect 24176 7692 24182 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 2038 7528 2044 7540
rect 1999 7500 2044 7528
rect 2038 7488 2044 7500
rect 2096 7488 2102 7540
rect 5997 7531 6055 7537
rect 5997 7497 6009 7531
rect 6043 7528 6055 7531
rect 6822 7528 6828 7540
rect 6043 7500 6828 7528
rect 6043 7497 6055 7500
rect 5997 7491 6055 7497
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 7926 7528 7932 7540
rect 7887 7500 7932 7528
rect 7926 7488 7932 7500
rect 7984 7488 7990 7540
rect 8297 7531 8355 7537
rect 8297 7497 8309 7531
rect 8343 7528 8355 7531
rect 8386 7528 8392 7540
rect 8343 7500 8392 7528
rect 8343 7497 8355 7500
rect 8297 7491 8355 7497
rect 8386 7488 8392 7500
rect 8444 7488 8450 7540
rect 8481 7531 8539 7537
rect 8481 7497 8493 7531
rect 8527 7528 8539 7531
rect 9674 7528 9680 7540
rect 8527 7500 9680 7528
rect 8527 7497 8539 7500
rect 8481 7491 8539 7497
rect 9674 7488 9680 7500
rect 9732 7488 9738 7540
rect 9769 7531 9827 7537
rect 9769 7497 9781 7531
rect 9815 7528 9827 7531
rect 10318 7528 10324 7540
rect 9815 7500 10324 7528
rect 9815 7497 9827 7500
rect 9769 7491 9827 7497
rect 10318 7488 10324 7500
rect 10376 7488 10382 7540
rect 11606 7528 11612 7540
rect 11567 7500 11612 7528
rect 11606 7488 11612 7500
rect 11664 7488 11670 7540
rect 11977 7531 12035 7537
rect 11977 7497 11989 7531
rect 12023 7528 12035 7531
rect 12066 7528 12072 7540
rect 12023 7500 12072 7528
rect 12023 7497 12035 7500
rect 11977 7491 12035 7497
rect 12066 7488 12072 7500
rect 12124 7488 12130 7540
rect 12710 7528 12716 7540
rect 12671 7500 12716 7528
rect 12710 7488 12716 7500
rect 12768 7488 12774 7540
rect 13078 7528 13084 7540
rect 13039 7500 13084 7528
rect 13078 7488 13084 7500
rect 13136 7488 13142 7540
rect 13446 7528 13452 7540
rect 13407 7500 13452 7528
rect 13446 7488 13452 7500
rect 13504 7488 13510 7540
rect 13906 7528 13912 7540
rect 13867 7500 13912 7528
rect 13906 7488 13912 7500
rect 13964 7488 13970 7540
rect 13998 7488 14004 7540
rect 14056 7528 14062 7540
rect 14185 7531 14243 7537
rect 14185 7528 14197 7531
rect 14056 7500 14197 7528
rect 14056 7488 14062 7500
rect 14185 7497 14197 7500
rect 14231 7497 14243 7531
rect 16942 7528 16948 7540
rect 16903 7500 16948 7528
rect 14185 7491 14243 7497
rect 16942 7488 16948 7500
rect 17000 7488 17006 7540
rect 23934 7528 23940 7540
rect 23895 7500 23940 7528
rect 23934 7488 23940 7500
rect 23992 7488 23998 7540
rect 24026 7488 24032 7540
rect 24084 7528 24090 7540
rect 24397 7531 24455 7537
rect 24397 7528 24409 7531
rect 24084 7500 24409 7528
rect 24084 7488 24090 7500
rect 24397 7497 24409 7500
rect 24443 7497 24455 7531
rect 24397 7491 24455 7497
rect 24670 7488 24676 7540
rect 24728 7528 24734 7540
rect 24765 7531 24823 7537
rect 24765 7528 24777 7531
rect 24728 7500 24777 7528
rect 24728 7488 24734 7500
rect 24765 7497 24777 7500
rect 24811 7497 24823 7531
rect 24765 7491 24823 7497
rect 1578 7460 1584 7472
rect 1539 7432 1584 7460
rect 1578 7420 1584 7432
rect 1636 7420 1642 7472
rect 5629 7463 5687 7469
rect 5629 7429 5641 7463
rect 5675 7460 5687 7463
rect 6454 7460 6460 7472
rect 5675 7432 6460 7460
rect 5675 7429 5687 7432
rect 5629 7423 5687 7429
rect 6454 7420 6460 7432
rect 6512 7420 6518 7472
rect 9692 7460 9720 7488
rect 10689 7463 10747 7469
rect 10689 7460 10701 7463
rect 9692 7432 10701 7460
rect 10689 7429 10701 7432
rect 10735 7429 10747 7463
rect 10689 7423 10747 7429
rect 6365 7395 6423 7401
rect 6365 7361 6377 7395
rect 6411 7392 6423 7395
rect 6730 7392 6736 7404
rect 6411 7364 6736 7392
rect 6411 7361 6423 7364
rect 6365 7355 6423 7361
rect 6730 7352 6736 7364
rect 6788 7352 6794 7404
rect 8478 7352 8484 7404
rect 8536 7392 8542 7404
rect 8941 7395 8999 7401
rect 8941 7392 8953 7395
rect 8536 7364 8953 7392
rect 8536 7352 8542 7364
rect 8941 7361 8953 7364
rect 8987 7392 8999 7395
rect 9582 7392 9588 7404
rect 8987 7364 9588 7392
rect 8987 7361 8999 7364
rect 8941 7355 8999 7361
rect 9582 7352 9588 7364
rect 9640 7352 9646 7404
rect 9674 7352 9680 7404
rect 9732 7392 9738 7404
rect 10137 7395 10195 7401
rect 10137 7392 10149 7395
rect 9732 7364 10149 7392
rect 9732 7352 9738 7364
rect 10137 7361 10149 7364
rect 10183 7361 10195 7395
rect 10137 7355 10195 7361
rect 1394 7324 1400 7336
rect 1355 7296 1400 7324
rect 1394 7284 1400 7296
rect 1452 7284 1458 7336
rect 7561 7327 7619 7333
rect 7561 7293 7573 7327
rect 7607 7324 7619 7327
rect 8662 7324 8668 7336
rect 7607 7296 8668 7324
rect 7607 7293 7619 7296
rect 7561 7287 7619 7293
rect 8662 7284 8668 7296
rect 8720 7324 8726 7336
rect 9033 7327 9091 7333
rect 9033 7324 9045 7327
rect 8720 7296 9045 7324
rect 8720 7284 8726 7296
rect 9033 7293 9045 7296
rect 9079 7293 9091 7327
rect 9950 7324 9956 7336
rect 9911 7296 9956 7324
rect 9033 7287 9091 7293
rect 9950 7284 9956 7296
rect 10008 7284 10014 7336
rect 17218 7284 17224 7336
rect 17276 7324 17282 7336
rect 18049 7327 18107 7333
rect 18049 7324 18061 7327
rect 17276 7296 18061 7324
rect 17276 7284 17282 7296
rect 18049 7293 18061 7296
rect 18095 7324 18107 7327
rect 18601 7327 18659 7333
rect 18601 7324 18613 7327
rect 18095 7296 18613 7324
rect 18095 7293 18107 7296
rect 18049 7287 18107 7293
rect 18601 7293 18613 7296
rect 18647 7293 18659 7327
rect 18601 7287 18659 7293
rect 23842 7284 23848 7336
rect 23900 7324 23906 7336
rect 24581 7327 24639 7333
rect 24581 7324 24593 7327
rect 23900 7296 24593 7324
rect 23900 7284 23906 7296
rect 24581 7293 24593 7296
rect 24627 7324 24639 7327
rect 25133 7327 25191 7333
rect 25133 7324 25145 7327
rect 24627 7296 25145 7324
rect 24627 7293 24639 7296
rect 24581 7287 24639 7293
rect 25133 7293 25145 7296
rect 25179 7293 25191 7327
rect 25133 7287 25191 7293
rect 8386 7216 8392 7268
rect 8444 7256 8450 7268
rect 8941 7259 8999 7265
rect 8941 7256 8953 7259
rect 8444 7228 8953 7256
rect 8444 7216 8450 7228
rect 8941 7225 8953 7228
rect 8987 7225 8999 7259
rect 8941 7219 8999 7225
rect 18230 7188 18236 7200
rect 18191 7160 18236 7188
rect 18230 7148 18236 7160
rect 18288 7148 18294 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1394 6944 1400 6996
rect 1452 6984 1458 6996
rect 1581 6987 1639 6993
rect 1581 6984 1593 6987
rect 1452 6956 1593 6984
rect 1452 6944 1458 6956
rect 1581 6953 1593 6956
rect 1627 6953 1639 6987
rect 8478 6984 8484 6996
rect 8439 6956 8484 6984
rect 1581 6947 1639 6953
rect 8478 6944 8484 6956
rect 8536 6944 8542 6996
rect 8662 6944 8668 6996
rect 8720 6984 8726 6996
rect 8757 6987 8815 6993
rect 8757 6984 8769 6987
rect 8720 6956 8769 6984
rect 8720 6944 8726 6956
rect 8757 6953 8769 6956
rect 8803 6953 8815 6987
rect 9858 6984 9864 6996
rect 9819 6956 9864 6984
rect 8757 6947 8815 6953
rect 9858 6944 9864 6956
rect 9916 6944 9922 6996
rect 9950 6944 9956 6996
rect 10008 6984 10014 6996
rect 10229 6987 10287 6993
rect 10229 6984 10241 6987
rect 10008 6956 10241 6984
rect 10008 6944 10014 6956
rect 10229 6953 10241 6956
rect 10275 6953 10287 6987
rect 10229 6947 10287 6953
rect 11977 6987 12035 6993
rect 11977 6953 11989 6987
rect 12023 6984 12035 6987
rect 12250 6984 12256 6996
rect 12023 6956 12256 6984
rect 12023 6953 12035 6956
rect 11977 6947 12035 6953
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 24762 6984 24768 6996
rect 24723 6956 24768 6984
rect 24762 6944 24768 6956
rect 24820 6944 24826 6996
rect 4890 6916 4896 6928
rect 4632 6888 4896 6916
rect 4632 6857 4660 6888
rect 4890 6876 4896 6888
rect 4948 6876 4954 6928
rect 4617 6851 4675 6857
rect 4617 6817 4629 6851
rect 4663 6817 4675 6851
rect 4617 6811 4675 6817
rect 8113 6851 8171 6857
rect 8113 6817 8125 6851
rect 8159 6848 8171 6851
rect 8294 6848 8300 6860
rect 8159 6820 8300 6848
rect 8159 6817 8171 6820
rect 8113 6811 8171 6817
rect 8294 6808 8300 6820
rect 8352 6808 8358 6860
rect 24578 6848 24584 6860
rect 24539 6820 24584 6848
rect 24578 6808 24584 6820
rect 24636 6808 24642 6860
rect 4798 6780 4804 6792
rect 4759 6752 4804 6780
rect 4798 6740 4804 6752
rect 4856 6740 4862 6792
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 4709 6443 4767 6449
rect 4709 6409 4721 6443
rect 4755 6440 4767 6443
rect 4798 6440 4804 6452
rect 4755 6412 4804 6440
rect 4755 6409 4767 6412
rect 4709 6403 4767 6409
rect 4065 6239 4123 6245
rect 4065 6205 4077 6239
rect 4111 6236 4123 6239
rect 4724 6236 4752 6403
rect 4798 6400 4804 6412
rect 4856 6400 4862 6452
rect 4982 6440 4988 6452
rect 4943 6412 4988 6440
rect 4982 6400 4988 6412
rect 5040 6400 5046 6452
rect 9309 6443 9367 6449
rect 9309 6409 9321 6443
rect 9355 6440 9367 6443
rect 9582 6440 9588 6452
rect 9355 6412 9588 6440
rect 9355 6409 9367 6412
rect 9309 6403 9367 6409
rect 4111 6208 4752 6236
rect 8665 6239 8723 6245
rect 4111 6205 4123 6208
rect 4065 6199 4123 6205
rect 8665 6205 8677 6239
rect 8711 6236 8723 6239
rect 9324 6236 9352 6403
rect 9582 6400 9588 6412
rect 9640 6400 9646 6452
rect 24762 6440 24768 6452
rect 24723 6412 24768 6440
rect 24762 6400 24768 6412
rect 24820 6400 24826 6452
rect 24489 6375 24547 6381
rect 24489 6341 24501 6375
rect 24535 6372 24547 6375
rect 24670 6372 24676 6384
rect 24535 6344 24676 6372
rect 24535 6341 24547 6344
rect 24489 6335 24547 6341
rect 24670 6332 24676 6344
rect 24728 6332 24734 6384
rect 8711 6208 9352 6236
rect 8711 6205 8723 6208
rect 8665 6199 8723 6205
rect 24210 6196 24216 6248
rect 24268 6236 24274 6248
rect 24581 6239 24639 6245
rect 24581 6236 24593 6239
rect 24268 6208 24593 6236
rect 24268 6196 24274 6208
rect 24581 6205 24593 6208
rect 24627 6236 24639 6239
rect 25133 6239 25191 6245
rect 25133 6236 25145 6239
rect 24627 6208 25145 6236
rect 24627 6205 24639 6208
rect 24581 6199 24639 6205
rect 25133 6205 25145 6208
rect 25179 6205 25191 6239
rect 25133 6199 25191 6205
rect 4246 6100 4252 6112
rect 4207 6072 4252 6100
rect 4246 6060 4252 6072
rect 4304 6060 4310 6112
rect 8846 6100 8852 6112
rect 8807 6072 8852 6100
rect 8846 6060 8852 6072
rect 8904 6060 8910 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 24762 5896 24768 5908
rect 24723 5868 24768 5896
rect 24762 5856 24768 5868
rect 24820 5856 24826 5908
rect 20714 5720 20720 5772
rect 20772 5760 20778 5772
rect 20901 5763 20959 5769
rect 20901 5760 20913 5763
rect 20772 5732 20913 5760
rect 20772 5720 20778 5732
rect 20901 5729 20913 5732
rect 20947 5729 20959 5763
rect 24578 5760 24584 5772
rect 24539 5732 24584 5760
rect 20901 5723 20959 5729
rect 24578 5720 24584 5732
rect 24636 5720 24642 5772
rect 21082 5692 21088 5704
rect 21043 5664 21088 5692
rect 21082 5652 21088 5664
rect 21140 5652 21146 5704
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 20714 5312 20720 5364
rect 20772 5352 20778 5364
rect 20901 5355 20959 5361
rect 20901 5352 20913 5355
rect 20772 5324 20913 5352
rect 20772 5312 20778 5324
rect 20901 5321 20913 5324
rect 20947 5321 20959 5355
rect 24762 5352 24768 5364
rect 24723 5324 24768 5352
rect 20901 5315 20959 5321
rect 24762 5312 24768 5324
rect 24820 5312 24826 5364
rect 24489 5287 24547 5293
rect 24489 5253 24501 5287
rect 24535 5284 24547 5287
rect 24670 5284 24676 5296
rect 24535 5256 24676 5284
rect 24535 5253 24547 5256
rect 24489 5247 24547 5253
rect 24670 5244 24676 5256
rect 24728 5244 24734 5296
rect 24578 5148 24584 5160
rect 24539 5120 24584 5148
rect 24578 5108 24584 5120
rect 24636 5148 24642 5160
rect 25133 5151 25191 5157
rect 25133 5148 25145 5151
rect 24636 5120 25145 5148
rect 24636 5108 24642 5120
rect 25133 5117 25145 5120
rect 25179 5117 25191 5151
rect 25133 5111 25191 5117
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 21266 4808 21272 4820
rect 21227 4780 21272 4808
rect 21266 4768 21272 4780
rect 21324 4768 21330 4820
rect 21082 4672 21088 4684
rect 21043 4644 21088 4672
rect 21082 4632 21088 4644
rect 21140 4632 21146 4684
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 21082 4264 21088 4276
rect 21043 4236 21088 4264
rect 21082 4224 21088 4236
rect 21140 4224 21146 4276
rect 2406 4128 2412 4140
rect 1688 4100 2412 4128
rect 1688 4069 1716 4100
rect 2406 4088 2412 4100
rect 2464 4088 2470 4140
rect 1673 4063 1731 4069
rect 1673 4029 1685 4063
rect 1719 4029 1731 4063
rect 1673 4023 1731 4029
rect 1394 3952 1400 4004
rect 1452 3992 1458 4004
rect 1949 3995 2007 4001
rect 1949 3992 1961 3995
rect 1452 3964 1961 3992
rect 1452 3952 1458 3964
rect 1949 3961 1961 3964
rect 1995 3961 2007 3995
rect 1949 3955 2007 3961
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1394 3584 1400 3596
rect 1355 3556 1400 3584
rect 1394 3544 1400 3556
rect 1452 3544 1458 3596
rect 23569 3587 23627 3593
rect 23569 3553 23581 3587
rect 23615 3584 23627 3587
rect 23750 3584 23756 3596
rect 23615 3556 23756 3584
rect 23615 3553 23627 3556
rect 23569 3547 23627 3553
rect 23750 3544 23756 3556
rect 23808 3544 23814 3596
rect 24854 3584 24860 3596
rect 24815 3556 24860 3584
rect 24854 3544 24860 3556
rect 24912 3544 24918 3596
rect 23845 3519 23903 3525
rect 23845 3485 23857 3519
rect 23891 3516 23903 3519
rect 25130 3516 25136 3528
rect 23891 3488 25136 3516
rect 23891 3485 23903 3488
rect 23845 3479 23903 3485
rect 25130 3476 25136 3488
rect 25188 3476 25194 3528
rect 1578 3448 1584 3460
rect 1539 3420 1584 3448
rect 1578 3408 1584 3420
rect 1636 3408 1642 3460
rect 25038 3380 25044 3392
rect 24999 3352 25044 3380
rect 25038 3340 25044 3352
rect 25096 3340 25102 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1394 3136 1400 3188
rect 1452 3176 1458 3188
rect 1581 3179 1639 3185
rect 1581 3176 1593 3179
rect 1452 3148 1593 3176
rect 1452 3136 1458 3148
rect 1581 3145 1593 3148
rect 1627 3145 1639 3179
rect 1581 3139 1639 3145
rect 4525 3179 4583 3185
rect 4525 3145 4537 3179
rect 4571 3176 4583 3179
rect 4614 3176 4620 3188
rect 4571 3148 4620 3176
rect 4571 3145 4583 3148
rect 4525 3139 4583 3145
rect 3697 2975 3755 2981
rect 3697 2941 3709 2975
rect 3743 2972 3755 2975
rect 4540 2972 4568 3139
rect 4614 3136 4620 3148
rect 4672 3136 4678 3188
rect 23109 3179 23167 3185
rect 23109 3145 23121 3179
rect 23155 3176 23167 3179
rect 23750 3176 23756 3188
rect 23155 3148 23756 3176
rect 23155 3145 23167 3148
rect 23109 3139 23167 3145
rect 23750 3136 23756 3148
rect 23808 3136 23814 3188
rect 24854 3176 24860 3188
rect 24815 3148 24860 3176
rect 24854 3136 24860 3148
rect 24912 3136 24918 3188
rect 8110 2972 8116 2984
rect 3743 2944 4568 2972
rect 8071 2944 8116 2972
rect 3743 2941 3755 2944
rect 3697 2935 3755 2941
rect 8110 2932 8116 2944
rect 8168 2972 8174 2984
rect 8849 2975 8907 2981
rect 8849 2972 8861 2975
rect 8168 2944 8861 2972
rect 8168 2932 8174 2944
rect 8849 2941 8861 2944
rect 8895 2941 8907 2975
rect 8849 2935 8907 2941
rect 23477 2975 23535 2981
rect 23477 2941 23489 2975
rect 23523 2972 23535 2975
rect 23842 2972 23848 2984
rect 23523 2944 23848 2972
rect 23523 2941 23535 2944
rect 23477 2935 23535 2941
rect 23842 2932 23848 2944
rect 23900 2932 23906 2984
rect 24121 2975 24179 2981
rect 24121 2941 24133 2975
rect 24167 2972 24179 2975
rect 24854 2972 24860 2984
rect 24167 2944 24860 2972
rect 24167 2941 24179 2944
rect 24121 2935 24179 2941
rect 24854 2932 24860 2944
rect 24912 2932 24918 2984
rect 25130 2972 25136 2984
rect 25091 2944 25136 2972
rect 25130 2932 25136 2944
rect 25188 2972 25194 2984
rect 25685 2975 25743 2981
rect 25685 2972 25697 2975
rect 25188 2944 25697 2972
rect 25188 2932 25194 2944
rect 25685 2941 25697 2944
rect 25731 2941 25743 2975
rect 25685 2935 25743 2941
rect 2682 2864 2688 2916
rect 2740 2904 2746 2916
rect 3973 2907 4031 2913
rect 3973 2904 3985 2907
rect 2740 2876 3985 2904
rect 2740 2864 2746 2876
rect 3973 2873 3985 2876
rect 4019 2873 4031 2907
rect 3973 2867 4031 2873
rect 8202 2864 8208 2916
rect 8260 2904 8266 2916
rect 8389 2907 8447 2913
rect 8389 2904 8401 2907
rect 8260 2876 8401 2904
rect 8260 2864 8266 2876
rect 8389 2873 8401 2876
rect 8435 2873 8447 2907
rect 8389 2867 8447 2873
rect 25314 2836 25320 2848
rect 25275 2808 25320 2836
rect 25314 2796 25320 2808
rect 25372 2796 25378 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 2041 2635 2099 2641
rect 2041 2601 2053 2635
rect 2087 2632 2099 2635
rect 2682 2632 2688 2644
rect 2087 2604 2688 2632
rect 2087 2601 2099 2604
rect 2041 2595 2099 2601
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2496 1455 2499
rect 2056 2496 2084 2595
rect 2682 2592 2688 2604
rect 2740 2592 2746 2644
rect 8021 2635 8079 2641
rect 8021 2601 8033 2635
rect 8067 2632 8079 2635
rect 8202 2632 8208 2644
rect 8067 2604 8208 2632
rect 8067 2601 8079 2604
rect 8021 2595 8079 2601
rect 1443 2468 2084 2496
rect 7377 2499 7435 2505
rect 1443 2465 1455 2468
rect 1397 2459 1455 2465
rect 7377 2465 7389 2499
rect 7423 2496 7435 2499
rect 8036 2496 8064 2595
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 7423 2468 8064 2496
rect 22833 2499 22891 2505
rect 7423 2465 7435 2468
rect 7377 2459 7435 2465
rect 22833 2465 22845 2499
rect 22879 2496 22891 2499
rect 24029 2499 24087 2505
rect 22879 2468 23520 2496
rect 22879 2465 22891 2468
rect 22833 2459 22891 2465
rect 23492 2437 23520 2468
rect 24029 2465 24041 2499
rect 24075 2496 24087 2499
rect 24118 2496 24124 2508
rect 24075 2468 24124 2496
rect 24075 2465 24087 2468
rect 24029 2459 24087 2465
rect 24118 2456 24124 2468
rect 24176 2496 24182 2508
rect 24765 2499 24823 2505
rect 24765 2496 24777 2499
rect 24176 2468 24777 2496
rect 24176 2456 24182 2468
rect 24765 2465 24777 2468
rect 24811 2465 24823 2499
rect 24765 2459 24823 2465
rect 24854 2456 24860 2508
rect 24912 2496 24918 2508
rect 25317 2499 25375 2505
rect 25317 2496 25329 2499
rect 24912 2468 25329 2496
rect 24912 2456 24918 2468
rect 25317 2465 25329 2468
rect 25363 2496 25375 2499
rect 25869 2499 25927 2505
rect 25869 2496 25881 2499
rect 25363 2468 25881 2496
rect 25363 2465 25375 2468
rect 25317 2459 25375 2465
rect 25869 2465 25881 2468
rect 25915 2465 25927 2499
rect 25869 2459 25927 2465
rect 23477 2431 23535 2437
rect 23477 2397 23489 2431
rect 23523 2428 23535 2431
rect 24213 2431 24271 2437
rect 24213 2428 24225 2431
rect 23523 2400 24225 2428
rect 23523 2397 23535 2400
rect 23477 2391 23535 2397
rect 24213 2397 24225 2400
rect 24259 2397 24271 2431
rect 24213 2391 24271 2397
rect 1578 2292 1584 2304
rect 1539 2264 1584 2292
rect 1578 2252 1584 2264
rect 1636 2252 1642 2304
rect 7558 2292 7564 2304
rect 7519 2264 7564 2292
rect 7558 2252 7564 2264
rect 7616 2252 7622 2304
rect 23014 2292 23020 2304
rect 22975 2264 23020 2292
rect 23014 2252 23020 2264
rect 23072 2252 23078 2304
rect 25498 2292 25504 2304
rect 25459 2264 25504 2292
rect 25498 2252 25504 2264
rect 25556 2252 25562 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
<< via1 >>
rect 9772 26392 9824 26444
rect 24768 26392 24820 26444
rect 8208 26324 8260 26376
rect 23572 26324 23624 26376
rect 7380 26256 7432 26308
rect 24308 26256 24360 26308
rect 4068 25780 4120 25832
rect 13728 25780 13780 25832
rect 12900 25712 12952 25764
rect 21732 25712 21784 25764
rect 8576 25644 8628 25696
rect 25964 25644 26016 25696
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 12900 25440 12952 25492
rect 8392 25372 8444 25424
rect 15660 25440 15712 25492
rect 16856 25440 16908 25492
rect 20076 25440 20128 25492
rect 22192 25440 22244 25492
rect 25412 25440 25464 25492
rect 7104 25304 7156 25356
rect 10692 25304 10744 25356
rect 11336 25347 11388 25356
rect 11336 25313 11345 25347
rect 11345 25313 11379 25347
rect 11379 25313 11388 25347
rect 11336 25304 11388 25313
rect 1676 25279 1728 25288
rect 1676 25245 1685 25279
rect 1685 25245 1719 25279
rect 1719 25245 1728 25279
rect 1676 25236 1728 25245
rect 5080 25236 5132 25288
rect 8484 25279 8536 25288
rect 8484 25245 8493 25279
rect 8493 25245 8527 25279
rect 8527 25245 8536 25279
rect 8484 25236 8536 25245
rect 8760 25236 8812 25288
rect 14740 25304 14792 25356
rect 15292 25304 15344 25356
rect 23480 25372 23532 25424
rect 16304 25304 16356 25356
rect 16948 25347 17000 25356
rect 16948 25313 16957 25347
rect 16957 25313 16991 25347
rect 16991 25313 17000 25347
rect 16948 25304 17000 25313
rect 18236 25304 18288 25356
rect 19432 25347 19484 25356
rect 19432 25313 19441 25347
rect 19441 25313 19475 25347
rect 19475 25313 19484 25347
rect 19432 25304 19484 25313
rect 21088 25304 21140 25356
rect 15660 25236 15712 25288
rect 3976 25168 4028 25220
rect 10600 25168 10652 25220
rect 4712 25100 4764 25152
rect 7840 25100 7892 25152
rect 9404 25100 9456 25152
rect 11336 25100 11388 25152
rect 14096 25100 14148 25152
rect 17224 25236 17276 25288
rect 22652 25304 22704 25356
rect 24032 25347 24084 25356
rect 24032 25313 24041 25347
rect 24041 25313 24075 25347
rect 24075 25313 24084 25347
rect 24032 25304 24084 25313
rect 25688 25304 25740 25356
rect 17408 25168 17460 25220
rect 20628 25168 20680 25220
rect 20168 25100 20220 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 8392 24896 8444 24948
rect 13084 24896 13136 24948
rect 22652 24939 22704 24948
rect 1584 24803 1636 24812
rect 1584 24769 1593 24803
rect 1593 24769 1627 24803
rect 1627 24769 1636 24803
rect 1584 24760 1636 24769
rect 1768 24692 1820 24744
rect 3792 24760 3844 24812
rect 4712 24803 4764 24812
rect 4712 24769 4721 24803
rect 4721 24769 4755 24803
rect 4755 24769 4764 24803
rect 4712 24760 4764 24769
rect 8484 24828 8536 24880
rect 10600 24803 10652 24812
rect 10600 24769 10609 24803
rect 10609 24769 10643 24803
rect 10643 24769 10652 24803
rect 10600 24760 10652 24769
rect 10968 24760 11020 24812
rect 11336 24760 11388 24812
rect 11612 24760 11664 24812
rect 15568 24803 15620 24812
rect 15568 24769 15577 24803
rect 15577 24769 15611 24803
rect 15611 24769 15620 24803
rect 15568 24760 15620 24769
rect 21088 24828 21140 24880
rect 22652 24905 22661 24939
rect 22661 24905 22695 24939
rect 22695 24905 22704 24939
rect 22652 24896 22704 24905
rect 24768 24828 24820 24880
rect 23480 24803 23532 24812
rect 2412 24667 2464 24676
rect 2412 24633 2421 24667
rect 2421 24633 2455 24667
rect 2455 24633 2464 24667
rect 2412 24624 2464 24633
rect 3700 24624 3752 24676
rect 7012 24624 7064 24676
rect 7840 24624 7892 24676
rect 8300 24667 8352 24676
rect 8300 24633 8309 24667
rect 8309 24633 8343 24667
rect 8343 24633 8352 24667
rect 8300 24624 8352 24633
rect 1400 24556 1452 24608
rect 4344 24556 4396 24608
rect 5080 24599 5132 24608
rect 5080 24565 5089 24599
rect 5089 24565 5123 24599
rect 5123 24565 5132 24599
rect 5080 24556 5132 24565
rect 5540 24556 5592 24608
rect 7104 24599 7156 24608
rect 7104 24565 7113 24599
rect 7113 24565 7147 24599
rect 7147 24565 7156 24599
rect 7104 24556 7156 24565
rect 7748 24599 7800 24608
rect 7748 24565 7781 24599
rect 7781 24565 7800 24599
rect 7748 24556 7800 24565
rect 10692 24624 10744 24676
rect 10876 24624 10928 24676
rect 13452 24692 13504 24744
rect 14096 24692 14148 24744
rect 15384 24692 15436 24744
rect 18052 24735 18104 24744
rect 18052 24701 18061 24735
rect 18061 24701 18095 24735
rect 18095 24701 18104 24735
rect 18052 24692 18104 24701
rect 19340 24735 19392 24744
rect 19340 24701 19349 24735
rect 19349 24701 19383 24735
rect 19383 24701 19392 24735
rect 19340 24692 19392 24701
rect 20628 24735 20680 24744
rect 20628 24701 20637 24735
rect 20637 24701 20671 24735
rect 20671 24701 20680 24735
rect 23480 24769 23489 24803
rect 23489 24769 23523 24803
rect 23523 24769 23532 24803
rect 23480 24760 23532 24769
rect 20628 24692 20680 24701
rect 24768 24735 24820 24744
rect 24768 24701 24777 24735
rect 24777 24701 24811 24735
rect 24811 24701 24820 24735
rect 24768 24692 24820 24701
rect 11704 24624 11756 24676
rect 12532 24624 12584 24676
rect 12808 24667 12860 24676
rect 12808 24633 12817 24667
rect 12817 24633 12851 24667
rect 12851 24633 12860 24667
rect 12808 24624 12860 24633
rect 15476 24624 15528 24676
rect 18236 24624 18288 24676
rect 20536 24624 20588 24676
rect 9588 24556 9640 24608
rect 13360 24556 13412 24608
rect 14464 24556 14516 24608
rect 14832 24556 14884 24608
rect 15292 24599 15344 24608
rect 15292 24565 15301 24599
rect 15301 24565 15335 24599
rect 15335 24565 15344 24599
rect 15292 24556 15344 24565
rect 16396 24556 16448 24608
rect 16948 24599 17000 24608
rect 16948 24565 16957 24599
rect 16957 24565 16991 24599
rect 16991 24565 17000 24599
rect 16948 24556 17000 24565
rect 18328 24556 18380 24608
rect 20812 24599 20864 24608
rect 20812 24565 20821 24599
rect 20821 24565 20855 24599
rect 20855 24565 20864 24599
rect 20812 24556 20864 24565
rect 21916 24599 21968 24608
rect 21916 24565 21925 24599
rect 21925 24565 21959 24599
rect 21959 24565 21968 24599
rect 21916 24556 21968 24565
rect 23848 24599 23900 24608
rect 23848 24565 23857 24599
rect 23857 24565 23891 24599
rect 23891 24565 23900 24599
rect 23848 24556 23900 24565
rect 24032 24556 24084 24608
rect 24952 24599 25004 24608
rect 24952 24565 24961 24599
rect 24961 24565 24995 24599
rect 24995 24565 25004 24599
rect 24952 24556 25004 24565
rect 25688 24599 25740 24608
rect 25688 24565 25697 24599
rect 25697 24565 25731 24599
rect 25731 24565 25740 24599
rect 25688 24556 25740 24565
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 1676 24284 1728 24336
rect 8300 24352 8352 24404
rect 10876 24395 10928 24404
rect 10876 24361 10885 24395
rect 10885 24361 10919 24395
rect 10919 24361 10928 24395
rect 10876 24352 10928 24361
rect 11612 24352 11664 24404
rect 13360 24352 13412 24404
rect 14832 24352 14884 24404
rect 19432 24395 19484 24404
rect 2044 24327 2096 24336
rect 2044 24293 2053 24327
rect 2053 24293 2087 24327
rect 2087 24293 2096 24327
rect 2044 24284 2096 24293
rect 7932 24327 7984 24336
rect 7932 24293 7941 24327
rect 7941 24293 7975 24327
rect 7975 24293 7984 24327
rect 7932 24284 7984 24293
rect 8116 24284 8168 24336
rect 8576 24284 8628 24336
rect 11520 24284 11572 24336
rect 13820 24284 13872 24336
rect 17592 24284 17644 24336
rect 19432 24361 19441 24395
rect 19441 24361 19475 24395
rect 19475 24361 19484 24395
rect 19432 24352 19484 24361
rect 24860 24395 24912 24404
rect 24860 24361 24869 24395
rect 24869 24361 24903 24395
rect 24903 24361 24912 24395
rect 24860 24352 24912 24361
rect 19340 24284 19392 24336
rect 23112 24284 23164 24336
rect 664 24216 716 24268
rect 4988 24216 5040 24268
rect 5172 24259 5224 24268
rect 5172 24225 5206 24259
rect 5206 24225 5224 24259
rect 5172 24216 5224 24225
rect 7748 24259 7800 24268
rect 7748 24225 7757 24259
rect 7757 24225 7791 24259
rect 7791 24225 7800 24259
rect 7748 24216 7800 24225
rect 13176 24216 13228 24268
rect 13636 24216 13688 24268
rect 15568 24259 15620 24268
rect 15568 24225 15577 24259
rect 15577 24225 15611 24259
rect 15611 24225 15620 24259
rect 15568 24216 15620 24225
rect 3424 24148 3476 24200
rect 4160 24148 4212 24200
rect 11060 24191 11112 24200
rect 11060 24157 11069 24191
rect 11069 24157 11103 24191
rect 11103 24157 11112 24191
rect 11060 24148 11112 24157
rect 13912 24148 13964 24200
rect 14004 24148 14056 24200
rect 16028 24148 16080 24200
rect 17500 24191 17552 24200
rect 17500 24157 17509 24191
rect 17509 24157 17543 24191
rect 17543 24157 17552 24191
rect 17500 24148 17552 24157
rect 18328 24216 18380 24268
rect 1768 24080 1820 24132
rect 12808 24080 12860 24132
rect 13636 24080 13688 24132
rect 14188 24080 14240 24132
rect 14556 24080 14608 24132
rect 17132 24080 17184 24132
rect 4528 24012 4580 24064
rect 6276 24055 6328 24064
rect 6276 24021 6285 24055
rect 6285 24021 6319 24055
rect 6319 24021 6328 24055
rect 6276 24012 6328 24021
rect 7196 24012 7248 24064
rect 13728 24055 13780 24064
rect 13728 24021 13737 24055
rect 13737 24021 13771 24055
rect 13771 24021 13780 24055
rect 13728 24012 13780 24021
rect 14740 24055 14792 24064
rect 14740 24021 14749 24055
rect 14749 24021 14783 24055
rect 14783 24021 14792 24055
rect 14740 24012 14792 24021
rect 16948 24012 17000 24064
rect 21916 24216 21968 24268
rect 24216 24216 24268 24268
rect 24952 24216 25004 24268
rect 19432 24148 19484 24200
rect 19800 24191 19852 24200
rect 19800 24157 19809 24191
rect 19809 24157 19843 24191
rect 19843 24157 19852 24191
rect 19800 24148 19852 24157
rect 22100 24191 22152 24200
rect 22100 24157 22109 24191
rect 22109 24157 22143 24191
rect 22143 24157 22152 24191
rect 23572 24191 23624 24200
rect 22100 24148 22152 24157
rect 23572 24157 23581 24191
rect 23581 24157 23615 24191
rect 23615 24157 23624 24191
rect 23572 24148 23624 24157
rect 20444 24080 20496 24132
rect 18512 24012 18564 24064
rect 19340 24012 19392 24064
rect 20352 24055 20404 24064
rect 20352 24021 20361 24055
rect 20361 24021 20395 24055
rect 20395 24021 20404 24055
rect 20352 24012 20404 24021
rect 22928 24055 22980 24064
rect 22928 24021 22937 24055
rect 22937 24021 22971 24055
rect 22971 24021 22980 24055
rect 22928 24012 22980 24021
rect 23388 24012 23440 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 4160 23851 4212 23860
rect 4160 23817 4169 23851
rect 4169 23817 4203 23851
rect 4203 23817 4212 23851
rect 4160 23808 4212 23817
rect 8116 23808 8168 23860
rect 8392 23808 8444 23860
rect 9404 23851 9456 23860
rect 1400 23715 1452 23724
rect 1400 23681 1409 23715
rect 1409 23681 1443 23715
rect 1443 23681 1452 23715
rect 1400 23672 1452 23681
rect 9404 23817 9413 23851
rect 9413 23817 9447 23851
rect 9447 23817 9456 23851
rect 9404 23808 9456 23817
rect 10048 23851 10100 23860
rect 10048 23817 10057 23851
rect 10057 23817 10091 23851
rect 10091 23817 10100 23851
rect 10048 23808 10100 23817
rect 12716 23851 12768 23860
rect 12716 23817 12725 23851
rect 12725 23817 12759 23851
rect 12759 23817 12768 23851
rect 12716 23808 12768 23817
rect 16488 23851 16540 23860
rect 16488 23817 16497 23851
rect 16497 23817 16531 23851
rect 16531 23817 16540 23851
rect 16488 23808 16540 23817
rect 21456 23851 21508 23860
rect 21456 23817 21465 23851
rect 21465 23817 21499 23851
rect 21499 23817 21508 23851
rect 21456 23808 21508 23817
rect 23112 23851 23164 23860
rect 23112 23817 23121 23851
rect 23121 23817 23155 23851
rect 23155 23817 23164 23851
rect 23112 23808 23164 23817
rect 17500 23740 17552 23792
rect 4528 23647 4580 23656
rect 4528 23613 4562 23647
rect 4562 23613 4580 23647
rect 4528 23604 4580 23613
rect 7472 23647 7524 23656
rect 7472 23613 7481 23647
rect 7481 23613 7515 23647
rect 7515 23613 7524 23647
rect 7472 23604 7524 23613
rect 9404 23604 9456 23656
rect 1584 23536 1636 23588
rect 4344 23536 4396 23588
rect 5172 23536 5224 23588
rect 7104 23536 7156 23588
rect 7932 23536 7984 23588
rect 10048 23536 10100 23588
rect 10876 23604 10928 23656
rect 11060 23604 11112 23656
rect 11888 23604 11940 23656
rect 12164 23647 12216 23656
rect 12164 23613 12173 23647
rect 12173 23613 12207 23647
rect 12207 23613 12216 23647
rect 12164 23604 12216 23613
rect 2780 23511 2832 23520
rect 2780 23477 2789 23511
rect 2789 23477 2823 23511
rect 2823 23477 2832 23511
rect 3424 23511 3476 23520
rect 2780 23468 2832 23477
rect 3424 23477 3433 23511
rect 3433 23477 3467 23511
rect 3467 23477 3476 23511
rect 3424 23468 3476 23477
rect 4712 23468 4764 23520
rect 5632 23511 5684 23520
rect 5632 23477 5641 23511
rect 5641 23477 5675 23511
rect 5675 23477 5684 23511
rect 5632 23468 5684 23477
rect 5816 23468 5868 23520
rect 11520 23511 11572 23520
rect 11520 23477 11529 23511
rect 11529 23477 11563 23511
rect 11563 23477 11572 23511
rect 11520 23468 11572 23477
rect 11888 23468 11940 23520
rect 16304 23604 16356 23656
rect 13912 23579 13964 23588
rect 13912 23545 13946 23579
rect 13946 23545 13964 23579
rect 13912 23536 13964 23545
rect 13820 23468 13872 23520
rect 15476 23536 15528 23588
rect 16672 23536 16724 23588
rect 17500 23604 17552 23656
rect 18880 23740 18932 23792
rect 20536 23715 20588 23724
rect 20536 23681 20545 23715
rect 20545 23681 20579 23715
rect 20579 23681 20588 23715
rect 20536 23672 20588 23681
rect 23020 23740 23072 23792
rect 25412 23808 25464 23860
rect 27620 23808 27672 23860
rect 21824 23647 21876 23656
rect 21824 23613 21833 23647
rect 21833 23613 21867 23647
rect 21867 23613 21876 23647
rect 21824 23604 21876 23613
rect 17132 23536 17184 23588
rect 17776 23536 17828 23588
rect 18420 23579 18472 23588
rect 18420 23545 18429 23579
rect 18429 23545 18463 23579
rect 18463 23545 18472 23579
rect 18420 23536 18472 23545
rect 18512 23536 18564 23588
rect 20352 23536 20404 23588
rect 22008 23536 22060 23588
rect 22928 23536 22980 23588
rect 14280 23468 14332 23520
rect 17592 23468 17644 23520
rect 18144 23468 18196 23520
rect 19984 23468 20036 23520
rect 21824 23468 21876 23520
rect 25044 23468 25096 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 3424 23264 3476 23316
rect 4160 23264 4212 23316
rect 5816 23307 5868 23316
rect 1860 23196 1912 23248
rect 1400 23128 1452 23180
rect 3516 23171 3568 23180
rect 3516 23137 3525 23171
rect 3525 23137 3559 23171
rect 3559 23137 3568 23171
rect 3516 23128 3568 23137
rect 5816 23273 5825 23307
rect 5825 23273 5859 23307
rect 5859 23273 5868 23307
rect 5816 23264 5868 23273
rect 7748 23264 7800 23316
rect 12808 23264 12860 23316
rect 16212 23307 16264 23316
rect 16212 23273 16221 23307
rect 16221 23273 16255 23307
rect 16255 23273 16264 23307
rect 16212 23264 16264 23273
rect 16672 23307 16724 23316
rect 16672 23273 16681 23307
rect 16681 23273 16715 23307
rect 16715 23273 16724 23307
rect 16672 23264 16724 23273
rect 23572 23264 23624 23316
rect 24952 23264 25004 23316
rect 4712 23239 4764 23248
rect 4712 23205 4746 23239
rect 4746 23205 4764 23239
rect 4712 23196 4764 23205
rect 7012 23239 7064 23248
rect 7012 23205 7021 23239
rect 7021 23205 7055 23239
rect 7055 23205 7064 23239
rect 7012 23196 7064 23205
rect 7472 23239 7524 23248
rect 7472 23205 7481 23239
rect 7481 23205 7515 23239
rect 7515 23205 7524 23239
rect 7472 23196 7524 23205
rect 8116 23196 8168 23248
rect 8576 23239 8628 23248
rect 8576 23205 8585 23239
rect 8585 23205 8619 23239
rect 8619 23205 8628 23239
rect 8576 23196 8628 23205
rect 9496 23239 9548 23248
rect 9496 23205 9505 23239
rect 9505 23205 9539 23239
rect 9539 23205 9548 23239
rect 9496 23196 9548 23205
rect 11152 23239 11204 23248
rect 11152 23205 11186 23239
rect 11186 23205 11204 23239
rect 11152 23196 11204 23205
rect 11612 23196 11664 23248
rect 13820 23196 13872 23248
rect 14188 23239 14240 23248
rect 14188 23205 14197 23239
rect 14197 23205 14231 23239
rect 14231 23205 14240 23239
rect 14188 23196 14240 23205
rect 15752 23239 15804 23248
rect 15752 23205 15761 23239
rect 15761 23205 15795 23239
rect 15795 23205 15804 23239
rect 15752 23196 15804 23205
rect 17224 23196 17276 23248
rect 19800 23239 19852 23248
rect 19800 23205 19809 23239
rect 19809 23205 19843 23239
rect 19843 23205 19852 23239
rect 19800 23196 19852 23205
rect 20352 23196 20404 23248
rect 22284 23196 22336 23248
rect 23388 23196 23440 23248
rect 23480 23196 23532 23248
rect 7932 23171 7984 23180
rect 7932 23137 7941 23171
rect 7941 23137 7975 23171
rect 7975 23137 7984 23171
rect 7932 23128 7984 23137
rect 10600 23128 10652 23180
rect 10876 23171 10928 23180
rect 10876 23137 10885 23171
rect 10885 23137 10919 23171
rect 10919 23137 10928 23171
rect 10876 23128 10928 23137
rect 14280 23171 14332 23180
rect 14280 23137 14289 23171
rect 14289 23137 14323 23171
rect 14323 23137 14332 23171
rect 14280 23128 14332 23137
rect 8668 23103 8720 23112
rect 8668 23069 8677 23103
rect 8677 23069 8711 23103
rect 8711 23069 8720 23103
rect 8668 23060 8720 23069
rect 9588 23060 9640 23112
rect 13544 23103 13596 23112
rect 13544 23069 13553 23103
rect 13553 23069 13587 23103
rect 13587 23069 13596 23103
rect 13544 23060 13596 23069
rect 14004 23060 14056 23112
rect 10048 22992 10100 23044
rect 13728 23035 13780 23044
rect 13728 23001 13737 23035
rect 13737 23001 13771 23035
rect 13771 23001 13780 23035
rect 13728 22992 13780 23001
rect 3792 22967 3844 22976
rect 3792 22933 3801 22967
rect 3801 22933 3835 22967
rect 3835 22933 3844 22967
rect 3792 22924 3844 22933
rect 10876 22924 10928 22976
rect 12164 22924 12216 22976
rect 13268 22924 13320 22976
rect 14832 22924 14884 22976
rect 17684 23128 17736 23180
rect 21548 23128 21600 23180
rect 23020 23128 23072 23180
rect 25688 23196 25740 23248
rect 24952 23171 25004 23180
rect 24952 23137 24961 23171
rect 24961 23137 24995 23171
rect 24995 23137 25004 23171
rect 24952 23128 25004 23137
rect 17408 23103 17460 23112
rect 17408 23069 17417 23103
rect 17417 23069 17451 23103
rect 17451 23069 17460 23103
rect 17408 23060 17460 23069
rect 16672 22992 16724 23044
rect 20076 23060 20128 23112
rect 24032 23103 24084 23112
rect 24032 23069 24041 23103
rect 24041 23069 24075 23103
rect 24075 23069 24084 23103
rect 24032 23060 24084 23069
rect 19984 22992 20036 23044
rect 18144 22967 18196 22976
rect 18144 22933 18153 22967
rect 18153 22933 18187 22967
rect 18187 22933 18196 22967
rect 18144 22924 18196 22933
rect 18972 22924 19024 22976
rect 19156 22967 19208 22976
rect 19156 22933 19165 22967
rect 19165 22933 19199 22967
rect 19199 22933 19208 22967
rect 19156 22924 19208 22933
rect 19340 22967 19392 22976
rect 19340 22933 19349 22967
rect 19349 22933 19383 22967
rect 19383 22933 19392 22967
rect 19340 22924 19392 22933
rect 20536 22924 20588 22976
rect 23572 22924 23624 22976
rect 24216 22924 24268 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 2044 22720 2096 22772
rect 4160 22763 4212 22772
rect 4160 22729 4169 22763
rect 4169 22729 4203 22763
rect 4203 22729 4212 22763
rect 4160 22720 4212 22729
rect 5080 22720 5132 22772
rect 5448 22763 5500 22772
rect 5448 22729 5457 22763
rect 5457 22729 5491 22763
rect 5491 22729 5500 22763
rect 5448 22720 5500 22729
rect 5540 22720 5592 22772
rect 8576 22720 8628 22772
rect 8852 22720 8904 22772
rect 9956 22720 10008 22772
rect 10600 22763 10652 22772
rect 572 22652 624 22704
rect 1400 22584 1452 22636
rect 2872 22627 2924 22636
rect 2872 22593 2881 22627
rect 2881 22593 2915 22627
rect 2915 22593 2924 22627
rect 2872 22584 2924 22593
rect 3240 22627 3292 22636
rect 3240 22593 3249 22627
rect 3249 22593 3283 22627
rect 3283 22593 3292 22627
rect 3240 22584 3292 22593
rect 8116 22695 8168 22704
rect 8116 22661 8125 22695
rect 8125 22661 8159 22695
rect 8159 22661 8168 22695
rect 8116 22652 8168 22661
rect 7472 22584 7524 22636
rect 1768 22559 1820 22568
rect 1768 22525 1777 22559
rect 1777 22525 1811 22559
rect 1811 22525 1820 22559
rect 1768 22516 1820 22525
rect 2964 22559 3016 22568
rect 2964 22525 2973 22559
rect 2973 22525 3007 22559
rect 3007 22525 3016 22559
rect 2964 22516 3016 22525
rect 3792 22516 3844 22568
rect 5172 22516 5224 22568
rect 5448 22516 5500 22568
rect 6184 22516 6236 22568
rect 6828 22559 6880 22568
rect 6828 22525 6837 22559
rect 6837 22525 6871 22559
rect 6871 22525 6880 22559
rect 6828 22516 6880 22525
rect 1860 22448 1912 22500
rect 2136 22380 2188 22432
rect 3056 22380 3108 22432
rect 4344 22448 4396 22500
rect 7104 22491 7156 22500
rect 7104 22457 7113 22491
rect 7113 22457 7147 22491
rect 7147 22457 7156 22491
rect 7104 22448 7156 22457
rect 8392 22448 8444 22500
rect 10600 22729 10609 22763
rect 10609 22729 10643 22763
rect 10643 22729 10652 22763
rect 10600 22720 10652 22729
rect 10968 22720 11020 22772
rect 14188 22720 14240 22772
rect 16304 22763 16356 22772
rect 16304 22729 16313 22763
rect 16313 22729 16347 22763
rect 16347 22729 16356 22763
rect 16304 22720 16356 22729
rect 17684 22763 17736 22772
rect 17684 22729 17693 22763
rect 17693 22729 17727 22763
rect 17727 22729 17736 22763
rect 17684 22720 17736 22729
rect 18052 22720 18104 22772
rect 21640 22763 21692 22772
rect 11336 22652 11388 22704
rect 14740 22652 14792 22704
rect 14924 22652 14976 22704
rect 18788 22695 18840 22704
rect 18788 22661 18797 22695
rect 18797 22661 18831 22695
rect 18831 22661 18840 22695
rect 18788 22652 18840 22661
rect 21640 22729 21649 22763
rect 21649 22729 21683 22763
rect 21683 22729 21692 22763
rect 21640 22720 21692 22729
rect 23020 22763 23072 22772
rect 23020 22729 23029 22763
rect 23029 22729 23063 22763
rect 23063 22729 23072 22763
rect 23020 22720 23072 22729
rect 24952 22720 25004 22772
rect 25320 22720 25372 22772
rect 19800 22652 19852 22704
rect 23756 22652 23808 22704
rect 10968 22584 11020 22636
rect 12256 22584 12308 22636
rect 12624 22584 12676 22636
rect 13268 22584 13320 22636
rect 13728 22584 13780 22636
rect 13912 22584 13964 22636
rect 16764 22627 16816 22636
rect 16764 22593 16773 22627
rect 16773 22593 16807 22627
rect 16807 22593 16816 22627
rect 16764 22584 16816 22593
rect 16856 22627 16908 22636
rect 16856 22593 16865 22627
rect 16865 22593 16899 22627
rect 16899 22593 16908 22627
rect 16856 22584 16908 22593
rect 17408 22584 17460 22636
rect 18972 22584 19024 22636
rect 11060 22516 11112 22568
rect 12992 22516 13044 22568
rect 12164 22448 12216 22500
rect 12440 22448 12492 22500
rect 12900 22448 12952 22500
rect 14188 22448 14240 22500
rect 14740 22516 14792 22568
rect 15384 22516 15436 22568
rect 18880 22516 18932 22568
rect 24676 22584 24728 22636
rect 25596 22627 25648 22636
rect 25596 22593 25605 22627
rect 25605 22593 25639 22627
rect 25639 22593 25648 22627
rect 25596 22584 25648 22593
rect 20536 22559 20588 22568
rect 20536 22525 20570 22559
rect 20570 22525 20588 22559
rect 16212 22448 16264 22500
rect 18972 22448 19024 22500
rect 19156 22448 19208 22500
rect 20536 22516 20588 22525
rect 24032 22516 24084 22568
rect 21548 22448 21600 22500
rect 23664 22448 23716 22500
rect 24216 22448 24268 22500
rect 25044 22448 25096 22500
rect 3516 22380 3568 22432
rect 3792 22423 3844 22432
rect 3792 22389 3801 22423
rect 3801 22389 3835 22423
rect 3835 22389 3844 22423
rect 3792 22380 3844 22389
rect 6368 22380 6420 22432
rect 11336 22423 11388 22432
rect 11336 22389 11345 22423
rect 11345 22389 11379 22423
rect 11379 22389 11388 22423
rect 11336 22380 11388 22389
rect 11612 22380 11664 22432
rect 17224 22423 17276 22432
rect 17224 22389 17233 22423
rect 17233 22389 17267 22423
rect 17267 22389 17276 22423
rect 17224 22380 17276 22389
rect 19984 22380 20036 22432
rect 22284 22423 22336 22432
rect 22284 22389 22293 22423
rect 22293 22389 22327 22423
rect 22327 22389 22336 22423
rect 22284 22380 22336 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 3516 22176 3568 22228
rect 5172 22219 5224 22228
rect 5172 22185 5181 22219
rect 5181 22185 5215 22219
rect 5215 22185 5224 22219
rect 5172 22176 5224 22185
rect 5448 22219 5500 22228
rect 5448 22185 5457 22219
rect 5457 22185 5491 22219
rect 5491 22185 5500 22219
rect 5448 22176 5500 22185
rect 2872 22108 2924 22160
rect 4252 22108 4304 22160
rect 1400 22040 1452 22092
rect 3424 22040 3476 22092
rect 4344 22083 4396 22092
rect 4344 22049 4353 22083
rect 4353 22049 4387 22083
rect 4387 22049 4396 22083
rect 5632 22108 5684 22160
rect 6828 22108 6880 22160
rect 4344 22040 4396 22049
rect 4620 22015 4672 22024
rect 4620 21981 4629 22015
rect 4629 21981 4663 22015
rect 4663 21981 4672 22015
rect 4620 21972 4672 21981
rect 2780 21904 2832 21956
rect 2228 21836 2280 21888
rect 4896 21836 4948 21888
rect 7472 22176 7524 22228
rect 7932 22108 7984 22160
rect 8116 22151 8168 22160
rect 8116 22117 8125 22151
rect 8125 22117 8159 22151
rect 8159 22117 8168 22151
rect 8116 22108 8168 22117
rect 7748 22040 7800 22092
rect 8024 22040 8076 22092
rect 8392 22176 8444 22228
rect 9772 22176 9824 22228
rect 11152 22219 11204 22228
rect 11152 22185 11161 22219
rect 11161 22185 11195 22219
rect 11195 22185 11204 22219
rect 11152 22176 11204 22185
rect 13544 22176 13596 22228
rect 13728 22176 13780 22228
rect 13820 22176 13872 22228
rect 16672 22176 16724 22228
rect 16856 22176 16908 22228
rect 20076 22219 20128 22228
rect 20076 22185 20085 22219
rect 20085 22185 20119 22219
rect 20119 22185 20128 22219
rect 20076 22176 20128 22185
rect 23112 22176 23164 22228
rect 23480 22219 23532 22228
rect 23480 22185 23489 22219
rect 23489 22185 23523 22219
rect 23523 22185 23532 22219
rect 23480 22176 23532 22185
rect 10048 22108 10100 22160
rect 9496 22083 9548 22092
rect 9496 22049 9505 22083
rect 9505 22049 9539 22083
rect 9539 22049 9548 22083
rect 9496 22040 9548 22049
rect 10784 22040 10836 22092
rect 12900 22108 12952 22160
rect 13452 22108 13504 22160
rect 14280 22151 14332 22160
rect 14280 22117 14289 22151
rect 14289 22117 14323 22151
rect 14323 22117 14332 22151
rect 14280 22108 14332 22117
rect 15292 22108 15344 22160
rect 18788 22108 18840 22160
rect 11704 22040 11756 22092
rect 11980 22040 12032 22092
rect 13728 22040 13780 22092
rect 15568 22040 15620 22092
rect 17408 22040 17460 22092
rect 19524 22108 19576 22160
rect 19984 22108 20036 22160
rect 21548 22151 21600 22160
rect 21548 22117 21557 22151
rect 21557 22117 21591 22151
rect 21591 22117 21600 22151
rect 21548 22108 21600 22117
rect 6368 21972 6420 22024
rect 8116 22015 8168 22024
rect 8116 21981 8125 22015
rect 8125 21981 8159 22015
rect 8159 21981 8168 22015
rect 8116 21972 8168 21981
rect 8484 21972 8536 22024
rect 10048 21972 10100 22024
rect 10232 22015 10284 22024
rect 10232 21981 10241 22015
rect 10241 21981 10275 22015
rect 10275 21981 10284 22015
rect 10232 21972 10284 21981
rect 9680 21904 9732 21956
rect 9956 21904 10008 21956
rect 10968 21972 11020 22024
rect 11152 21972 11204 22024
rect 11888 21972 11940 22024
rect 15844 22015 15896 22024
rect 15844 21981 15853 22015
rect 15853 21981 15887 22015
rect 15887 21981 15896 22015
rect 15844 21972 15896 21981
rect 19432 22040 19484 22092
rect 20628 22040 20680 22092
rect 20904 22083 20956 22092
rect 20904 22049 20913 22083
rect 20913 22049 20947 22083
rect 20947 22049 20956 22083
rect 20904 22040 20956 22049
rect 21916 22040 21968 22092
rect 23296 22040 23348 22092
rect 23848 22108 23900 22160
rect 24032 22108 24084 22160
rect 24216 22108 24268 22160
rect 24584 22108 24636 22160
rect 24768 22108 24820 22160
rect 19892 21972 19944 22024
rect 20260 21972 20312 22024
rect 23020 21972 23072 22024
rect 25412 22040 25464 22092
rect 14280 21904 14332 21956
rect 14924 21904 14976 21956
rect 16856 21904 16908 21956
rect 23664 21904 23716 21956
rect 6092 21879 6144 21888
rect 6092 21845 6101 21879
rect 6101 21845 6135 21879
rect 6135 21845 6144 21879
rect 6092 21836 6144 21845
rect 7012 21879 7064 21888
rect 7012 21845 7021 21879
rect 7021 21845 7055 21879
rect 7055 21845 7064 21879
rect 7012 21836 7064 21845
rect 10784 21879 10836 21888
rect 10784 21845 10793 21879
rect 10793 21845 10827 21879
rect 10827 21845 10836 21879
rect 10784 21836 10836 21845
rect 11060 21836 11112 21888
rect 12900 21836 12952 21888
rect 13176 21836 13228 21888
rect 13912 21836 13964 21888
rect 14188 21836 14240 21888
rect 14648 21879 14700 21888
rect 14648 21845 14657 21879
rect 14657 21845 14691 21879
rect 14691 21845 14700 21879
rect 14648 21836 14700 21845
rect 15384 21879 15436 21888
rect 15384 21845 15393 21879
rect 15393 21845 15427 21879
rect 15427 21845 15436 21879
rect 15384 21836 15436 21845
rect 17776 21836 17828 21888
rect 19064 21836 19116 21888
rect 19432 21836 19484 21888
rect 20720 21836 20772 21888
rect 21088 21879 21140 21888
rect 21088 21845 21097 21879
rect 21097 21845 21131 21879
rect 21131 21845 21140 21879
rect 21088 21836 21140 21845
rect 22652 21836 22704 21888
rect 22928 21836 22980 21888
rect 23296 21836 23348 21888
rect 24032 21836 24084 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 2872 21675 2924 21684
rect 2872 21641 2881 21675
rect 2881 21641 2915 21675
rect 2915 21641 2924 21675
rect 2872 21632 2924 21641
rect 3424 21632 3476 21684
rect 8116 21632 8168 21684
rect 9588 21632 9640 21684
rect 10416 21675 10468 21684
rect 10416 21641 10425 21675
rect 10425 21641 10459 21675
rect 10459 21641 10468 21675
rect 10416 21632 10468 21641
rect 10692 21632 10744 21684
rect 11888 21675 11940 21684
rect 11888 21641 11897 21675
rect 11897 21641 11931 21675
rect 11931 21641 11940 21675
rect 11888 21632 11940 21641
rect 12532 21675 12584 21684
rect 12532 21641 12541 21675
rect 12541 21641 12575 21675
rect 12575 21641 12584 21675
rect 12532 21632 12584 21641
rect 14740 21632 14792 21684
rect 16396 21632 16448 21684
rect 17500 21632 17552 21684
rect 18972 21675 19024 21684
rect 18972 21641 18981 21675
rect 18981 21641 19015 21675
rect 19015 21641 19024 21675
rect 18972 21632 19024 21641
rect 19892 21675 19944 21684
rect 19892 21641 19901 21675
rect 19901 21641 19935 21675
rect 19935 21641 19944 21675
rect 19892 21632 19944 21641
rect 21916 21675 21968 21684
rect 21916 21641 21925 21675
rect 21925 21641 21959 21675
rect 21959 21641 21968 21675
rect 21916 21632 21968 21641
rect 23112 21675 23164 21684
rect 23112 21641 23121 21675
rect 23121 21641 23155 21675
rect 23155 21641 23164 21675
rect 23112 21632 23164 21641
rect 24216 21632 24268 21684
rect 24676 21675 24728 21684
rect 24676 21641 24685 21675
rect 24685 21641 24719 21675
rect 24719 21641 24728 21675
rect 24676 21632 24728 21641
rect 1492 21607 1544 21616
rect 1492 21573 1501 21607
rect 1501 21573 1535 21607
rect 1535 21573 1544 21607
rect 1492 21564 1544 21573
rect 3792 21564 3844 21616
rect 5540 21564 5592 21616
rect 8208 21607 8260 21616
rect 8208 21573 8217 21607
rect 8217 21573 8251 21607
rect 8251 21573 8260 21607
rect 8208 21564 8260 21573
rect 12348 21564 12400 21616
rect 3700 21496 3752 21548
rect 6092 21496 6144 21548
rect 10784 21496 10836 21548
rect 11980 21496 12032 21548
rect 2504 21428 2556 21480
rect 2780 21428 2832 21480
rect 6460 21428 6512 21480
rect 6644 21428 6696 21480
rect 7472 21428 7524 21480
rect 14556 21564 14608 21616
rect 19984 21564 20036 21616
rect 23296 21564 23348 21616
rect 23664 21564 23716 21616
rect 23940 21564 23992 21616
rect 14188 21496 14240 21548
rect 14648 21539 14700 21548
rect 14648 21505 14657 21539
rect 14657 21505 14691 21539
rect 14691 21505 14700 21539
rect 14648 21496 14700 21505
rect 16856 21539 16908 21548
rect 16856 21505 16865 21539
rect 16865 21505 16899 21539
rect 16899 21505 16908 21539
rect 16856 21496 16908 21505
rect 20076 21496 20128 21548
rect 20720 21496 20772 21548
rect 21364 21496 21416 21548
rect 22192 21496 22244 21548
rect 23756 21496 23808 21548
rect 15292 21471 15344 21480
rect 1768 21403 1820 21412
rect 1768 21369 1777 21403
rect 1777 21369 1811 21403
rect 1811 21369 1820 21403
rect 1768 21360 1820 21369
rect 2228 21360 2280 21412
rect 2964 21360 3016 21412
rect 5264 21360 5316 21412
rect 15292 21437 15301 21471
rect 15301 21437 15335 21471
rect 15335 21437 15344 21471
rect 15292 21428 15344 21437
rect 15936 21428 15988 21480
rect 7564 21360 7616 21412
rect 7748 21360 7800 21412
rect 10876 21403 10928 21412
rect 10876 21369 10885 21403
rect 10885 21369 10919 21403
rect 10919 21369 10928 21403
rect 10876 21360 10928 21369
rect 13084 21403 13136 21412
rect 13084 21369 13093 21403
rect 13093 21369 13127 21403
rect 13127 21369 13136 21403
rect 13084 21360 13136 21369
rect 13452 21360 13504 21412
rect 14556 21360 14608 21412
rect 2320 21292 2372 21344
rect 6644 21335 6696 21344
rect 6644 21301 6653 21335
rect 6653 21301 6687 21335
rect 6687 21301 6696 21335
rect 6644 21292 6696 21301
rect 8484 21292 8536 21344
rect 9680 21292 9732 21344
rect 9772 21292 9824 21344
rect 10692 21292 10744 21344
rect 11060 21335 11112 21344
rect 11060 21301 11069 21335
rect 11069 21301 11103 21335
rect 11103 21301 11112 21335
rect 11060 21292 11112 21301
rect 12624 21292 12676 21344
rect 14004 21335 14056 21344
rect 14004 21301 14013 21335
rect 14013 21301 14047 21335
rect 14047 21301 14056 21335
rect 15108 21360 15160 21412
rect 15844 21360 15896 21412
rect 16488 21360 16540 21412
rect 17500 21428 17552 21480
rect 19064 21428 19116 21480
rect 20352 21428 20404 21480
rect 22652 21471 22704 21480
rect 22652 21437 22661 21471
rect 22661 21437 22695 21471
rect 22695 21437 22704 21471
rect 22652 21428 22704 21437
rect 24124 21428 24176 21480
rect 24676 21428 24728 21480
rect 24860 21428 24912 21480
rect 14004 21292 14056 21301
rect 17960 21360 18012 21412
rect 19340 21360 19392 21412
rect 20444 21360 20496 21412
rect 22008 21360 22060 21412
rect 23020 21360 23072 21412
rect 23940 21360 23992 21412
rect 25044 21360 25096 21412
rect 17132 21292 17184 21344
rect 17408 21335 17460 21344
rect 17408 21301 17417 21335
rect 17417 21301 17451 21335
rect 17451 21301 17460 21335
rect 17408 21292 17460 21301
rect 20260 21335 20312 21344
rect 20260 21301 20269 21335
rect 20269 21301 20303 21335
rect 20303 21301 20312 21335
rect 20260 21292 20312 21301
rect 22560 21335 22612 21344
rect 22560 21301 22569 21335
rect 22569 21301 22603 21335
rect 22603 21301 22612 21335
rect 22560 21292 22612 21301
rect 23756 21335 23808 21344
rect 23756 21301 23765 21335
rect 23765 21301 23799 21335
rect 23799 21301 23808 21335
rect 23756 21292 23808 21301
rect 24124 21292 24176 21344
rect 25136 21335 25188 21344
rect 25136 21301 25145 21335
rect 25145 21301 25179 21335
rect 25179 21301 25188 21335
rect 25136 21292 25188 21301
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 2320 21088 2372 21140
rect 2964 21131 3016 21140
rect 2964 21097 2973 21131
rect 2973 21097 3007 21131
rect 3007 21097 3016 21131
rect 2964 21088 3016 21097
rect 3700 21088 3752 21140
rect 6460 21131 6512 21140
rect 6460 21097 6469 21131
rect 6469 21097 6503 21131
rect 6503 21097 6512 21131
rect 6460 21088 6512 21097
rect 7932 21088 7984 21140
rect 9956 21131 10008 21140
rect 9956 21097 9965 21131
rect 9965 21097 9999 21131
rect 9999 21097 10008 21131
rect 9956 21088 10008 21097
rect 11980 21131 12032 21140
rect 11980 21097 11989 21131
rect 11989 21097 12023 21131
rect 12023 21097 12032 21131
rect 11980 21088 12032 21097
rect 13360 21088 13412 21140
rect 13728 21088 13780 21140
rect 14556 21131 14608 21140
rect 14556 21097 14565 21131
rect 14565 21097 14599 21131
rect 14599 21097 14608 21131
rect 14556 21088 14608 21097
rect 16396 21131 16448 21140
rect 16396 21097 16405 21131
rect 16405 21097 16439 21131
rect 16439 21097 16448 21131
rect 16396 21088 16448 21097
rect 16580 21088 16632 21140
rect 16672 21088 16724 21140
rect 17868 21088 17920 21140
rect 18512 21131 18564 21140
rect 18512 21097 18521 21131
rect 18521 21097 18555 21131
rect 18555 21097 18564 21131
rect 18512 21088 18564 21097
rect 19524 21088 19576 21140
rect 20444 21131 20496 21140
rect 20444 21097 20453 21131
rect 20453 21097 20487 21131
rect 20487 21097 20496 21131
rect 20444 21088 20496 21097
rect 22284 21131 22336 21140
rect 22284 21097 22293 21131
rect 22293 21097 22327 21131
rect 22327 21097 22336 21131
rect 22284 21088 22336 21097
rect 22560 21088 22612 21140
rect 23388 21088 23440 21140
rect 24860 21088 24912 21140
rect 1492 21020 1544 21072
rect 2688 21020 2740 21072
rect 8116 21020 8168 21072
rect 8392 21063 8444 21072
rect 8392 21029 8401 21063
rect 8401 21029 8435 21063
rect 8435 21029 8444 21063
rect 8392 21020 8444 21029
rect 8484 21063 8536 21072
rect 8484 21029 8493 21063
rect 8493 21029 8527 21063
rect 8527 21029 8536 21063
rect 8484 21020 8536 21029
rect 10784 21020 10836 21072
rect 11704 21020 11756 21072
rect 12808 21020 12860 21072
rect 15752 21020 15804 21072
rect 20904 21020 20956 21072
rect 24216 21063 24268 21072
rect 24216 21029 24225 21063
rect 24225 21029 24259 21063
rect 24259 21029 24268 21063
rect 24216 21020 24268 21029
rect 2044 20952 2096 21004
rect 4896 20952 4948 21004
rect 7656 20952 7708 21004
rect 11152 20952 11204 21004
rect 12440 20952 12492 21004
rect 13728 20995 13780 21004
rect 13728 20961 13737 20995
rect 13737 20961 13771 20995
rect 13771 20961 13780 20995
rect 13728 20952 13780 20961
rect 15292 20952 15344 21004
rect 17040 20952 17092 21004
rect 17776 20952 17828 21004
rect 19340 20952 19392 21004
rect 20168 20952 20220 21004
rect 20996 20952 21048 21004
rect 24032 20952 24084 21004
rect 2688 20884 2740 20936
rect 5080 20927 5132 20936
rect 5080 20893 5089 20927
rect 5089 20893 5123 20927
rect 5123 20893 5132 20927
rect 5080 20884 5132 20893
rect 9312 20884 9364 20936
rect 12164 20884 12216 20936
rect 12992 20884 13044 20936
rect 14740 20884 14792 20936
rect 16948 20884 17000 20936
rect 17132 20927 17184 20936
rect 17132 20893 17141 20927
rect 17141 20893 17175 20927
rect 17175 20893 17184 20927
rect 17132 20884 17184 20893
rect 20904 20927 20956 20936
rect 20904 20893 20913 20927
rect 20913 20893 20947 20927
rect 20947 20893 20956 20927
rect 20904 20884 20956 20893
rect 1676 20859 1728 20868
rect 1676 20825 1685 20859
rect 1685 20825 1719 20859
rect 1719 20825 1728 20859
rect 1676 20816 1728 20825
rect 3700 20791 3752 20800
rect 3700 20757 3709 20791
rect 3709 20757 3743 20791
rect 3743 20757 3752 20791
rect 3700 20748 3752 20757
rect 4896 20791 4948 20800
rect 4896 20757 4905 20791
rect 4905 20757 4939 20791
rect 4939 20757 4948 20791
rect 4896 20748 4948 20757
rect 6828 20816 6880 20868
rect 12440 20816 12492 20868
rect 14648 20816 14700 20868
rect 24676 20884 24728 20936
rect 24952 21020 25004 21072
rect 25228 20995 25280 21004
rect 25228 20961 25237 20995
rect 25237 20961 25271 20995
rect 25271 20961 25280 20995
rect 25228 20952 25280 20961
rect 24860 20816 24912 20868
rect 5448 20748 5500 20800
rect 10324 20791 10376 20800
rect 10324 20757 10333 20791
rect 10333 20757 10367 20791
rect 10367 20757 10376 20791
rect 10324 20748 10376 20757
rect 12624 20791 12676 20800
rect 12624 20757 12633 20791
rect 12633 20757 12667 20791
rect 12667 20757 12676 20791
rect 12624 20748 12676 20757
rect 13084 20748 13136 20800
rect 13544 20748 13596 20800
rect 15568 20748 15620 20800
rect 18604 20748 18656 20800
rect 23480 20791 23532 20800
rect 23480 20757 23489 20791
rect 23489 20757 23523 20791
rect 23523 20757 23532 20791
rect 23480 20748 23532 20757
rect 25136 20791 25188 20800
rect 25136 20757 25145 20791
rect 25145 20757 25179 20791
rect 25179 20757 25188 20791
rect 25136 20748 25188 20757
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 2780 20544 2832 20596
rect 5264 20587 5316 20596
rect 5264 20553 5273 20587
rect 5273 20553 5307 20587
rect 5307 20553 5316 20587
rect 5264 20544 5316 20553
rect 7288 20587 7340 20596
rect 7288 20553 7297 20587
rect 7297 20553 7331 20587
rect 7331 20553 7340 20587
rect 7288 20544 7340 20553
rect 8116 20544 8168 20596
rect 9312 20587 9364 20596
rect 9312 20553 9321 20587
rect 9321 20553 9355 20587
rect 9355 20553 9364 20587
rect 9312 20544 9364 20553
rect 12348 20544 12400 20596
rect 13360 20544 13412 20596
rect 14096 20544 14148 20596
rect 14740 20544 14792 20596
rect 18328 20587 18380 20596
rect 18328 20553 18337 20587
rect 18337 20553 18371 20587
rect 18371 20553 18380 20587
rect 18328 20544 18380 20553
rect 20996 20544 21048 20596
rect 22192 20587 22244 20596
rect 22192 20553 22201 20587
rect 22201 20553 22235 20587
rect 22235 20553 22244 20587
rect 22192 20544 22244 20553
rect 22836 20544 22888 20596
rect 25228 20544 25280 20596
rect 2872 20476 2924 20528
rect 1400 20408 1452 20460
rect 5448 20408 5500 20460
rect 5816 20408 5868 20460
rect 2228 20340 2280 20392
rect 3700 20340 3752 20392
rect 6644 20340 6696 20392
rect 7656 20383 7708 20392
rect 7656 20349 7690 20383
rect 7690 20349 7708 20383
rect 7656 20340 7708 20349
rect 9864 20383 9916 20392
rect 9864 20349 9873 20383
rect 9873 20349 9907 20383
rect 9907 20349 9916 20383
rect 9864 20340 9916 20349
rect 12164 20383 12216 20392
rect 2964 20272 3016 20324
rect 4896 20272 4948 20324
rect 4252 20204 4304 20256
rect 5080 20204 5132 20256
rect 5724 20247 5776 20256
rect 5724 20213 5733 20247
rect 5733 20213 5767 20247
rect 5767 20213 5776 20247
rect 5724 20204 5776 20213
rect 6276 20204 6328 20256
rect 9588 20204 9640 20256
rect 12164 20349 12173 20383
rect 12173 20349 12207 20383
rect 12207 20349 12216 20383
rect 12164 20340 12216 20349
rect 13636 20383 13688 20392
rect 13636 20349 13645 20383
rect 13645 20349 13679 20383
rect 13679 20349 13688 20383
rect 13636 20340 13688 20349
rect 13820 20340 13872 20392
rect 14556 20340 14608 20392
rect 22652 20408 22704 20460
rect 16580 20383 16632 20392
rect 16580 20349 16589 20383
rect 16589 20349 16623 20383
rect 16623 20349 16632 20383
rect 16580 20340 16632 20349
rect 16948 20340 17000 20392
rect 10324 20272 10376 20324
rect 15016 20272 15068 20324
rect 16856 20315 16908 20324
rect 10784 20204 10836 20256
rect 11336 20204 11388 20256
rect 14648 20204 14700 20256
rect 15752 20247 15804 20256
rect 15752 20213 15761 20247
rect 15761 20213 15795 20247
rect 15795 20213 15804 20247
rect 15752 20204 15804 20213
rect 16856 20281 16865 20315
rect 16865 20281 16899 20315
rect 16899 20281 16908 20315
rect 16856 20272 16908 20281
rect 18052 20272 18104 20324
rect 18604 20315 18656 20324
rect 18604 20281 18613 20315
rect 18613 20281 18647 20315
rect 18647 20281 18656 20315
rect 18604 20272 18656 20281
rect 22100 20340 22152 20392
rect 23756 20340 23808 20392
rect 24032 20340 24084 20392
rect 20628 20272 20680 20324
rect 19064 20204 19116 20256
rect 20260 20204 20312 20256
rect 20904 20204 20956 20256
rect 22376 20204 22428 20256
rect 25504 20204 25556 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 1400 20000 1452 20052
rect 2044 20043 2096 20052
rect 2044 20009 2053 20043
rect 2053 20009 2087 20043
rect 2087 20009 2096 20043
rect 2044 20000 2096 20009
rect 3700 20000 3752 20052
rect 3792 20043 3844 20052
rect 3792 20009 3801 20043
rect 3801 20009 3835 20043
rect 3835 20009 3844 20043
rect 3792 20000 3844 20009
rect 5724 20000 5776 20052
rect 6828 20000 6880 20052
rect 9772 20000 9824 20052
rect 13820 20000 13872 20052
rect 14740 20043 14792 20052
rect 14740 20009 14749 20043
rect 14749 20009 14783 20043
rect 14783 20009 14792 20043
rect 14740 20000 14792 20009
rect 15108 20043 15160 20052
rect 15108 20009 15117 20043
rect 15117 20009 15151 20043
rect 15151 20009 15160 20043
rect 15108 20000 15160 20009
rect 15844 20000 15896 20052
rect 2780 19932 2832 19984
rect 8392 19975 8444 19984
rect 8392 19941 8401 19975
rect 8401 19941 8435 19975
rect 8435 19941 8444 19975
rect 8392 19932 8444 19941
rect 8484 19975 8536 19984
rect 8484 19941 8493 19975
rect 8493 19941 8527 19975
rect 8527 19941 8536 19975
rect 8484 19932 8536 19941
rect 9680 19932 9732 19984
rect 4160 19864 4212 19916
rect 4344 19907 4396 19916
rect 4344 19873 4378 19907
rect 4378 19873 4396 19907
rect 4344 19864 4396 19873
rect 5540 19864 5592 19916
rect 6184 19864 6236 19916
rect 2596 19796 2648 19848
rect 2964 19839 3016 19848
rect 2964 19805 2973 19839
rect 2973 19805 3007 19839
rect 3007 19805 3016 19839
rect 2964 19796 3016 19805
rect 3700 19796 3752 19848
rect 6736 19839 6788 19848
rect 2412 19728 2464 19780
rect 6736 19805 6745 19839
rect 6745 19805 6779 19839
rect 6779 19805 6788 19839
rect 6736 19796 6788 19805
rect 8576 19796 8628 19848
rect 13544 19932 13596 19984
rect 16856 20000 16908 20052
rect 17040 20043 17092 20052
rect 17040 20009 17049 20043
rect 17049 20009 17083 20043
rect 17083 20009 17092 20043
rect 17040 20000 17092 20009
rect 17960 20000 18012 20052
rect 20536 20000 20588 20052
rect 21180 20000 21232 20052
rect 22100 20000 22152 20052
rect 24216 20000 24268 20052
rect 25412 20043 25464 20052
rect 25412 20009 25421 20043
rect 25421 20009 25455 20043
rect 25455 20009 25464 20043
rect 25412 20000 25464 20009
rect 9864 19864 9916 19916
rect 11888 19864 11940 19916
rect 13636 19864 13688 19916
rect 17132 19932 17184 19984
rect 17868 19932 17920 19984
rect 19340 19932 19392 19984
rect 20996 19932 21048 19984
rect 23756 19932 23808 19984
rect 24032 19932 24084 19984
rect 24860 19932 24912 19984
rect 16764 19864 16816 19916
rect 21732 19864 21784 19916
rect 22376 19907 22428 19916
rect 22376 19873 22385 19907
rect 22385 19873 22419 19907
rect 22419 19873 22428 19907
rect 22376 19864 22428 19873
rect 23020 19864 23072 19916
rect 10140 19796 10192 19848
rect 5816 19728 5868 19780
rect 10876 19728 10928 19780
rect 16304 19796 16356 19848
rect 17040 19796 17092 19848
rect 20812 19796 20864 19848
rect 25504 19839 25556 19848
rect 25504 19805 25513 19839
rect 25513 19805 25547 19839
rect 25547 19805 25556 19839
rect 25504 19796 25556 19805
rect 7380 19660 7432 19712
rect 7564 19703 7616 19712
rect 7564 19669 7573 19703
rect 7573 19669 7607 19703
rect 7607 19669 7616 19703
rect 7564 19660 7616 19669
rect 9128 19703 9180 19712
rect 9128 19669 9137 19703
rect 9137 19669 9171 19703
rect 9171 19669 9180 19703
rect 9128 19660 9180 19669
rect 11336 19703 11388 19712
rect 11336 19669 11345 19703
rect 11345 19669 11379 19703
rect 11379 19669 11388 19703
rect 11336 19660 11388 19669
rect 12072 19660 12124 19712
rect 15568 19660 15620 19712
rect 19064 19703 19116 19712
rect 19064 19669 19073 19703
rect 19073 19669 19107 19703
rect 19107 19669 19116 19703
rect 19064 19660 19116 19669
rect 20168 19703 20220 19712
rect 20168 19669 20177 19703
rect 20177 19669 20211 19703
rect 20211 19669 20220 19703
rect 20168 19660 20220 19669
rect 23388 19660 23440 19712
rect 25872 19660 25924 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 1400 19456 1452 19508
rect 6184 19499 6236 19508
rect 6184 19465 6193 19499
rect 6193 19465 6227 19499
rect 6227 19465 6236 19499
rect 6184 19456 6236 19465
rect 8484 19456 8536 19508
rect 9772 19456 9824 19508
rect 10968 19456 11020 19508
rect 11888 19456 11940 19508
rect 14096 19456 14148 19508
rect 4252 19388 4304 19440
rect 3792 19320 3844 19372
rect 2688 19252 2740 19304
rect 7656 19320 7708 19372
rect 2596 19184 2648 19236
rect 2964 19116 3016 19168
rect 4344 19184 4396 19236
rect 4988 19227 5040 19236
rect 4160 19116 4212 19168
rect 4988 19193 4997 19227
rect 4997 19193 5031 19227
rect 5031 19193 5040 19227
rect 4988 19184 5040 19193
rect 6920 19252 6972 19304
rect 5356 19184 5408 19236
rect 7380 19227 7432 19236
rect 7380 19193 7389 19227
rect 7389 19193 7423 19227
rect 7423 19193 7432 19227
rect 8300 19252 8352 19304
rect 9128 19295 9180 19304
rect 9128 19261 9137 19295
rect 9137 19261 9171 19295
rect 9171 19261 9180 19295
rect 9128 19252 9180 19261
rect 9404 19295 9456 19304
rect 9404 19261 9413 19295
rect 9413 19261 9447 19295
rect 9447 19261 9456 19295
rect 9404 19252 9456 19261
rect 9496 19252 9548 19304
rect 11336 19320 11388 19372
rect 12532 19363 12584 19372
rect 12532 19329 12557 19363
rect 12557 19329 12584 19363
rect 12532 19320 12584 19329
rect 9680 19252 9732 19304
rect 10968 19252 11020 19304
rect 11612 19252 11664 19304
rect 7380 19184 7432 19193
rect 4528 19116 4580 19168
rect 7564 19116 7616 19168
rect 8116 19184 8168 19236
rect 10232 19184 10284 19236
rect 11152 19184 11204 19236
rect 8484 19159 8536 19168
rect 8484 19125 8493 19159
rect 8493 19125 8527 19159
rect 8527 19125 8536 19159
rect 8484 19116 8536 19125
rect 9864 19116 9916 19168
rect 12072 19184 12124 19236
rect 19432 19320 19484 19372
rect 20260 19456 20312 19508
rect 22376 19499 22428 19508
rect 22376 19465 22385 19499
rect 22385 19465 22419 19499
rect 22419 19465 22428 19499
rect 22376 19456 22428 19465
rect 23020 19499 23072 19508
rect 23020 19465 23029 19499
rect 23029 19465 23063 19499
rect 23063 19465 23072 19499
rect 23020 19456 23072 19465
rect 24216 19456 24268 19508
rect 24860 19456 24912 19508
rect 25504 19388 25556 19440
rect 25412 19320 25464 19372
rect 12808 19227 12860 19236
rect 12808 19193 12817 19227
rect 12817 19193 12851 19227
rect 12851 19193 12860 19227
rect 12808 19184 12860 19193
rect 13636 19184 13688 19236
rect 16488 19252 16540 19304
rect 18972 19252 19024 19304
rect 17040 19184 17092 19236
rect 18328 19227 18380 19236
rect 18328 19193 18337 19227
rect 18337 19193 18371 19227
rect 18371 19193 18380 19227
rect 19984 19252 20036 19304
rect 20168 19252 20220 19304
rect 24032 19252 24084 19304
rect 18328 19184 18380 19193
rect 19524 19184 19576 19236
rect 20076 19184 20128 19236
rect 24676 19184 24728 19236
rect 13268 19116 13320 19168
rect 13544 19159 13596 19168
rect 13544 19125 13553 19159
rect 13553 19125 13587 19159
rect 13587 19125 13596 19159
rect 13544 19116 13596 19125
rect 15384 19116 15436 19168
rect 16304 19159 16356 19168
rect 16304 19125 16313 19159
rect 16313 19125 16347 19159
rect 16347 19125 16356 19159
rect 16304 19116 16356 19125
rect 16764 19159 16816 19168
rect 16764 19125 16773 19159
rect 16773 19125 16807 19159
rect 16807 19125 16816 19159
rect 16764 19116 16816 19125
rect 19248 19116 19300 19168
rect 20720 19116 20772 19168
rect 22560 19159 22612 19168
rect 22560 19125 22569 19159
rect 22569 19125 22603 19159
rect 22603 19125 22612 19159
rect 22560 19116 22612 19125
rect 24032 19159 24084 19168
rect 24032 19125 24041 19159
rect 24041 19125 24075 19159
rect 24075 19125 24084 19159
rect 24032 19116 24084 19125
rect 24768 19159 24820 19168
rect 24768 19125 24777 19159
rect 24777 19125 24811 19159
rect 24811 19125 24820 19159
rect 24768 19116 24820 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 2688 18912 2740 18964
rect 3700 18955 3752 18964
rect 3700 18921 3709 18955
rect 3709 18921 3743 18955
rect 3743 18921 3752 18955
rect 3700 18912 3752 18921
rect 4344 18955 4396 18964
rect 4344 18921 4353 18955
rect 4353 18921 4387 18955
rect 4387 18921 4396 18955
rect 4344 18912 4396 18921
rect 7656 18955 7708 18964
rect 7656 18921 7665 18955
rect 7665 18921 7699 18955
rect 7699 18921 7708 18955
rect 7656 18912 7708 18921
rect 8392 18912 8444 18964
rect 9496 18955 9548 18964
rect 9496 18921 9505 18955
rect 9505 18921 9539 18955
rect 9539 18921 9548 18955
rect 9496 18912 9548 18921
rect 10140 18955 10192 18964
rect 10140 18921 10149 18955
rect 10149 18921 10183 18955
rect 10183 18921 10192 18955
rect 10140 18912 10192 18921
rect 10784 18912 10836 18964
rect 11336 18955 11388 18964
rect 2964 18887 3016 18896
rect 2964 18853 2973 18887
rect 2973 18853 3007 18887
rect 3007 18853 3016 18887
rect 5264 18887 5316 18896
rect 2964 18844 3016 18853
rect 5264 18853 5273 18887
rect 5273 18853 5307 18887
rect 5307 18853 5316 18887
rect 5264 18844 5316 18853
rect 11336 18921 11345 18955
rect 11345 18921 11379 18955
rect 11379 18921 11388 18955
rect 11336 18912 11388 18921
rect 12624 18912 12676 18964
rect 12808 18912 12860 18964
rect 12992 18912 13044 18964
rect 13912 18912 13964 18964
rect 15844 18912 15896 18964
rect 17132 18955 17184 18964
rect 17132 18921 17141 18955
rect 17141 18921 17175 18955
rect 17175 18921 17184 18955
rect 17132 18912 17184 18921
rect 18604 18955 18656 18964
rect 18604 18921 18613 18955
rect 18613 18921 18647 18955
rect 18647 18921 18656 18955
rect 18604 18912 18656 18921
rect 20812 18912 20864 18964
rect 21456 18955 21508 18964
rect 21456 18921 21465 18955
rect 21465 18921 21499 18955
rect 21499 18921 21508 18955
rect 21456 18912 21508 18921
rect 11704 18887 11756 18896
rect 11704 18853 11713 18887
rect 11713 18853 11747 18887
rect 11747 18853 11756 18887
rect 11704 18844 11756 18853
rect 12348 18844 12400 18896
rect 12532 18844 12584 18896
rect 14648 18844 14700 18896
rect 16212 18887 16264 18896
rect 16212 18853 16221 18887
rect 16221 18853 16255 18887
rect 16255 18853 16264 18887
rect 16212 18844 16264 18853
rect 17868 18844 17920 18896
rect 21364 18844 21416 18896
rect 23388 18844 23440 18896
rect 25044 18844 25096 18896
rect 3148 18776 3200 18828
rect 3608 18776 3660 18828
rect 4160 18776 4212 18828
rect 5448 18776 5500 18828
rect 7012 18776 7064 18828
rect 9864 18776 9916 18828
rect 12808 18776 12860 18828
rect 13728 18776 13780 18828
rect 16028 18819 16080 18828
rect 16028 18785 16037 18819
rect 16037 18785 16071 18819
rect 16071 18785 16080 18819
rect 16028 18776 16080 18785
rect 21180 18776 21232 18828
rect 22376 18819 22428 18828
rect 22376 18785 22385 18819
rect 22385 18785 22419 18819
rect 22419 18785 22428 18819
rect 22376 18776 22428 18785
rect 25228 18819 25280 18828
rect 25228 18785 25237 18819
rect 25237 18785 25271 18819
rect 25271 18785 25280 18819
rect 25228 18776 25280 18785
rect 25780 18776 25832 18828
rect 2780 18751 2832 18760
rect 2780 18717 2789 18751
rect 2789 18717 2823 18751
rect 2823 18717 2832 18751
rect 5264 18751 5316 18760
rect 2780 18708 2832 18717
rect 5264 18717 5273 18751
rect 5273 18717 5307 18751
rect 5307 18717 5316 18751
rect 5264 18708 5316 18717
rect 6184 18708 6236 18760
rect 10968 18751 11020 18760
rect 10968 18717 10977 18751
rect 10977 18717 11011 18751
rect 11011 18717 11020 18751
rect 10968 18708 11020 18717
rect 12072 18708 12124 18760
rect 12532 18751 12584 18760
rect 2688 18640 2740 18692
rect 4804 18683 4856 18692
rect 4804 18649 4813 18683
rect 4813 18649 4847 18683
rect 4847 18649 4856 18683
rect 4804 18640 4856 18649
rect 12256 18640 12308 18692
rect 12532 18717 12541 18751
rect 12541 18717 12575 18751
rect 12575 18717 12584 18751
rect 12532 18708 12584 18717
rect 14004 18751 14056 18760
rect 14004 18717 14013 18751
rect 14013 18717 14047 18751
rect 14047 18717 14056 18751
rect 14004 18708 14056 18717
rect 14464 18708 14516 18760
rect 16120 18708 16172 18760
rect 13084 18640 13136 18692
rect 14924 18640 14976 18692
rect 15752 18683 15804 18692
rect 15752 18649 15761 18683
rect 15761 18649 15795 18683
rect 15795 18649 15804 18683
rect 15752 18640 15804 18649
rect 1584 18615 1636 18624
rect 1584 18581 1593 18615
rect 1593 18581 1627 18615
rect 1627 18581 1636 18615
rect 1584 18572 1636 18581
rect 1860 18572 1912 18624
rect 2504 18572 2556 18624
rect 5540 18572 5592 18624
rect 6092 18615 6144 18624
rect 6092 18581 6101 18615
rect 6101 18581 6135 18615
rect 6135 18581 6144 18615
rect 6092 18572 6144 18581
rect 8668 18615 8720 18624
rect 8668 18581 8677 18615
rect 8677 18581 8711 18615
rect 8711 18581 8720 18615
rect 8668 18572 8720 18581
rect 9036 18615 9088 18624
rect 9036 18581 9045 18615
rect 9045 18581 9079 18615
rect 9079 18581 9088 18615
rect 9036 18572 9088 18581
rect 11980 18615 12032 18624
rect 11980 18581 11989 18615
rect 11989 18581 12023 18615
rect 12023 18581 12032 18615
rect 11980 18572 12032 18581
rect 13544 18615 13596 18624
rect 13544 18581 13553 18615
rect 13553 18581 13587 18615
rect 13587 18581 13596 18615
rect 13544 18572 13596 18581
rect 13728 18572 13780 18624
rect 15384 18572 15436 18624
rect 17132 18708 17184 18760
rect 19340 18708 19392 18760
rect 25136 18708 25188 18760
rect 25504 18751 25556 18760
rect 25504 18717 25513 18751
rect 25513 18717 25547 18751
rect 25547 18717 25556 18751
rect 25504 18708 25556 18717
rect 23388 18640 23440 18692
rect 23848 18640 23900 18692
rect 24768 18640 24820 18692
rect 17040 18572 17092 18624
rect 19524 18615 19576 18624
rect 19524 18581 19533 18615
rect 19533 18581 19567 18615
rect 19567 18581 19576 18615
rect 19524 18572 19576 18581
rect 22100 18615 22152 18624
rect 22100 18581 22109 18615
rect 22109 18581 22143 18615
rect 22143 18581 22152 18615
rect 22100 18572 22152 18581
rect 23572 18572 23624 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 2872 18368 2924 18420
rect 5356 18368 5408 18420
rect 6644 18368 6696 18420
rect 7012 18411 7064 18420
rect 7012 18377 7021 18411
rect 7021 18377 7055 18411
rect 7055 18377 7064 18411
rect 7012 18368 7064 18377
rect 8668 18368 8720 18420
rect 10784 18368 10836 18420
rect 9864 18300 9916 18352
rect 12164 18368 12216 18420
rect 12808 18411 12860 18420
rect 12808 18377 12817 18411
rect 12817 18377 12851 18411
rect 12851 18377 12860 18411
rect 12808 18368 12860 18377
rect 14004 18368 14056 18420
rect 14648 18368 14700 18420
rect 14832 18368 14884 18420
rect 15476 18368 15528 18420
rect 16396 18368 16448 18420
rect 17868 18411 17920 18420
rect 17868 18377 17877 18411
rect 17877 18377 17911 18411
rect 17911 18377 17920 18411
rect 17868 18368 17920 18377
rect 19432 18411 19484 18420
rect 19432 18377 19441 18411
rect 19441 18377 19475 18411
rect 19475 18377 19484 18411
rect 19432 18368 19484 18377
rect 20168 18368 20220 18420
rect 21364 18368 21416 18420
rect 23480 18368 23532 18420
rect 25044 18411 25096 18420
rect 11704 18300 11756 18352
rect 13636 18300 13688 18352
rect 14740 18300 14792 18352
rect 13912 18275 13964 18284
rect 13912 18241 13921 18275
rect 13921 18241 13955 18275
rect 13955 18241 13964 18275
rect 13912 18232 13964 18241
rect 16580 18232 16632 18284
rect 19340 18232 19392 18284
rect 22192 18300 22244 18352
rect 22376 18300 22428 18352
rect 22560 18275 22612 18284
rect 22560 18241 22569 18275
rect 22569 18241 22603 18275
rect 22603 18241 22612 18275
rect 22560 18232 22612 18241
rect 23848 18275 23900 18284
rect 23848 18241 23857 18275
rect 23857 18241 23891 18275
rect 23891 18241 23900 18275
rect 23848 18232 23900 18241
rect 1584 18207 1636 18216
rect 1584 18173 1593 18207
rect 1593 18173 1627 18207
rect 1627 18173 1636 18207
rect 1584 18164 1636 18173
rect 1860 18207 1912 18216
rect 1860 18173 1894 18207
rect 1894 18173 1912 18207
rect 1860 18164 1912 18173
rect 4252 18207 4304 18216
rect 4252 18173 4261 18207
rect 4261 18173 4295 18207
rect 4295 18173 4304 18207
rect 4252 18164 4304 18173
rect 6184 18164 6236 18216
rect 3700 18096 3752 18148
rect 4344 18096 4396 18148
rect 3608 18071 3660 18080
rect 3608 18037 3617 18071
rect 3617 18037 3651 18071
rect 3651 18037 3660 18071
rect 3608 18028 3660 18037
rect 5540 18028 5592 18080
rect 6184 18028 6236 18080
rect 12992 18164 13044 18216
rect 16396 18164 16448 18216
rect 17040 18207 17092 18216
rect 17040 18173 17049 18207
rect 17049 18173 17083 18207
rect 17083 18173 17092 18207
rect 17040 18164 17092 18173
rect 22100 18164 22152 18216
rect 7840 18096 7892 18148
rect 10692 18139 10744 18148
rect 10692 18105 10701 18139
rect 10701 18105 10735 18139
rect 10735 18105 10744 18139
rect 10692 18096 10744 18105
rect 10784 18139 10836 18148
rect 10784 18105 10793 18139
rect 10793 18105 10827 18139
rect 10827 18105 10836 18139
rect 10784 18096 10836 18105
rect 9312 18028 9364 18080
rect 9772 18028 9824 18080
rect 12164 18096 12216 18148
rect 13360 18096 13412 18148
rect 15384 18139 15436 18148
rect 15384 18105 15393 18139
rect 15393 18105 15427 18139
rect 15427 18105 15436 18139
rect 15384 18096 15436 18105
rect 16948 18139 17000 18148
rect 16948 18105 16957 18139
rect 16957 18105 16991 18139
rect 16991 18105 17000 18139
rect 16948 18096 17000 18105
rect 19432 18096 19484 18148
rect 12532 18028 12584 18080
rect 16028 18028 16080 18080
rect 16672 18028 16724 18080
rect 17132 18028 17184 18080
rect 18604 18071 18656 18080
rect 18604 18037 18613 18071
rect 18613 18037 18647 18071
rect 18647 18037 18656 18071
rect 18604 18028 18656 18037
rect 22100 18028 22152 18080
rect 24032 18096 24084 18148
rect 25044 18377 25053 18411
rect 25053 18377 25087 18411
rect 25087 18377 25096 18411
rect 25044 18368 25096 18377
rect 25780 18368 25832 18420
rect 23848 18028 23900 18080
rect 24584 18071 24636 18080
rect 24584 18037 24593 18071
rect 24593 18037 24627 18071
rect 24627 18037 24636 18071
rect 24584 18028 24636 18037
rect 25504 18028 25556 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 2780 17867 2832 17876
rect 2780 17833 2789 17867
rect 2789 17833 2823 17867
rect 2823 17833 2832 17867
rect 2780 17824 2832 17833
rect 2964 17824 3016 17876
rect 4160 17824 4212 17876
rect 4344 17867 4396 17876
rect 4344 17833 4353 17867
rect 4353 17833 4387 17867
rect 4387 17833 4396 17867
rect 4344 17824 4396 17833
rect 5264 17867 5316 17876
rect 5264 17833 5273 17867
rect 5273 17833 5307 17867
rect 5307 17833 5316 17867
rect 5264 17824 5316 17833
rect 5448 17824 5500 17876
rect 6920 17824 6972 17876
rect 8668 17824 8720 17876
rect 9312 17867 9364 17876
rect 9312 17833 9321 17867
rect 9321 17833 9355 17867
rect 9355 17833 9364 17867
rect 9312 17824 9364 17833
rect 10784 17824 10836 17876
rect 13360 17867 13412 17876
rect 13360 17833 13369 17867
rect 13369 17833 13403 17867
rect 13403 17833 13412 17867
rect 13360 17824 13412 17833
rect 14556 17824 14608 17876
rect 16120 17867 16172 17876
rect 16120 17833 16129 17867
rect 16129 17833 16163 17867
rect 16163 17833 16172 17867
rect 16120 17824 16172 17833
rect 16488 17867 16540 17876
rect 16488 17833 16497 17867
rect 16497 17833 16531 17867
rect 16531 17833 16540 17867
rect 16488 17824 16540 17833
rect 18972 17824 19024 17876
rect 19524 17824 19576 17876
rect 3240 17756 3292 17808
rect 4528 17756 4580 17808
rect 4804 17756 4856 17808
rect 7840 17756 7892 17808
rect 15660 17756 15712 17808
rect 19616 17756 19668 17808
rect 21180 17824 21232 17876
rect 22100 17867 22152 17876
rect 22100 17833 22109 17867
rect 22109 17833 22143 17867
rect 22143 17833 22152 17867
rect 22100 17824 22152 17833
rect 23480 17756 23532 17808
rect 24584 17756 24636 17808
rect 24952 17756 25004 17808
rect 25044 17756 25096 17808
rect 5540 17688 5592 17740
rect 11060 17731 11112 17740
rect 11060 17697 11094 17731
rect 11094 17697 11112 17731
rect 11060 17688 11112 17697
rect 13912 17688 13964 17740
rect 15292 17731 15344 17740
rect 15292 17697 15301 17731
rect 15301 17697 15335 17731
rect 15335 17697 15344 17731
rect 15292 17688 15344 17697
rect 16948 17731 17000 17740
rect 16948 17697 16982 17731
rect 16982 17697 17000 17731
rect 16948 17688 17000 17697
rect 21456 17688 21508 17740
rect 23572 17688 23624 17740
rect 2228 17663 2280 17672
rect 2228 17629 2237 17663
rect 2237 17629 2271 17663
rect 2271 17629 2280 17663
rect 2228 17620 2280 17629
rect 2688 17620 2740 17672
rect 8668 17663 8720 17672
rect 1768 17595 1820 17604
rect 1768 17561 1777 17595
rect 1777 17561 1811 17595
rect 1811 17561 1820 17595
rect 1768 17552 1820 17561
rect 8208 17552 8260 17604
rect 8668 17629 8677 17663
rect 8677 17629 8711 17663
rect 8711 17629 8720 17663
rect 8668 17620 8720 17629
rect 9680 17663 9732 17672
rect 9680 17629 9689 17663
rect 9689 17629 9723 17663
rect 9723 17629 9732 17663
rect 9680 17620 9732 17629
rect 10784 17663 10836 17672
rect 10784 17629 10793 17663
rect 10793 17629 10827 17663
rect 10827 17629 10836 17663
rect 10784 17620 10836 17629
rect 13636 17620 13688 17672
rect 14188 17663 14240 17672
rect 14188 17629 14197 17663
rect 14197 17629 14231 17663
rect 14231 17629 14240 17663
rect 14188 17620 14240 17629
rect 16672 17663 16724 17672
rect 16672 17629 16681 17663
rect 16681 17629 16715 17663
rect 16715 17629 16724 17663
rect 16672 17620 16724 17629
rect 19984 17620 20036 17672
rect 22192 17663 22244 17672
rect 22192 17629 22201 17663
rect 22201 17629 22235 17663
rect 22235 17629 22244 17663
rect 22192 17620 22244 17629
rect 25136 17663 25188 17672
rect 25136 17629 25145 17663
rect 25145 17629 25179 17663
rect 25179 17629 25188 17663
rect 25136 17620 25188 17629
rect 25504 17620 25556 17672
rect 9036 17552 9088 17604
rect 9588 17552 9640 17604
rect 13728 17595 13780 17604
rect 13728 17561 13737 17595
rect 13737 17561 13771 17595
rect 13771 17561 13780 17595
rect 13728 17552 13780 17561
rect 24032 17552 24084 17604
rect 24676 17552 24728 17604
rect 6184 17484 6236 17536
rect 10968 17484 11020 17536
rect 12164 17527 12216 17536
rect 12164 17493 12173 17527
rect 12173 17493 12207 17527
rect 12207 17493 12216 17527
rect 12164 17484 12216 17493
rect 12532 17484 12584 17536
rect 14832 17527 14884 17536
rect 14832 17493 14841 17527
rect 14841 17493 14875 17527
rect 14875 17493 14884 17527
rect 14832 17484 14884 17493
rect 18052 17527 18104 17536
rect 18052 17493 18061 17527
rect 18061 17493 18095 17527
rect 18095 17493 18104 17527
rect 18052 17484 18104 17493
rect 20168 17484 20220 17536
rect 23388 17484 23440 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 5172 17280 5224 17332
rect 7196 17280 7248 17332
rect 8024 17280 8076 17332
rect 8668 17280 8720 17332
rect 11060 17280 11112 17332
rect 15844 17280 15896 17332
rect 16580 17280 16632 17332
rect 18052 17280 18104 17332
rect 19524 17280 19576 17332
rect 21456 17323 21508 17332
rect 21456 17289 21465 17323
rect 21465 17289 21499 17323
rect 21499 17289 21508 17323
rect 21456 17280 21508 17289
rect 22192 17280 22244 17332
rect 23020 17323 23072 17332
rect 23020 17289 23029 17323
rect 23029 17289 23063 17323
rect 23063 17289 23072 17323
rect 23020 17280 23072 17289
rect 5540 17212 5592 17264
rect 4804 17144 4856 17196
rect 19616 17212 19668 17264
rect 20352 17212 20404 17264
rect 22836 17212 22888 17264
rect 23940 17212 23992 17264
rect 22560 17187 22612 17196
rect 2412 17119 2464 17128
rect 2412 17085 2421 17119
rect 2421 17085 2455 17119
rect 2455 17085 2464 17119
rect 2412 17076 2464 17085
rect 2688 17119 2740 17128
rect 1676 17008 1728 17060
rect 2688 17085 2722 17119
rect 2722 17085 2740 17119
rect 2688 17076 2740 17085
rect 1584 16940 1636 16992
rect 2412 16940 2464 16992
rect 3424 16940 3476 16992
rect 4160 16940 4212 16992
rect 5540 17051 5592 17060
rect 5540 17017 5549 17051
rect 5549 17017 5583 17051
rect 5583 17017 5592 17051
rect 5540 17008 5592 17017
rect 6184 17008 6236 17060
rect 6920 17076 6972 17128
rect 8208 16983 8260 16992
rect 8208 16949 8217 16983
rect 8217 16949 8251 16983
rect 8251 16949 8260 16983
rect 8208 16940 8260 16949
rect 9036 16940 9088 16992
rect 9404 17076 9456 17128
rect 10140 17076 10192 17128
rect 10784 16940 10836 16992
rect 15200 17076 15252 17128
rect 12532 17008 12584 17060
rect 13544 17008 13596 17060
rect 13360 16940 13412 16992
rect 15200 16940 15252 16992
rect 16672 16940 16724 16992
rect 22560 17153 22569 17187
rect 22569 17153 22603 17187
rect 22603 17153 22612 17187
rect 22560 17144 22612 17153
rect 25228 17187 25280 17196
rect 25228 17153 25237 17187
rect 25237 17153 25271 17187
rect 25271 17153 25280 17187
rect 25228 17144 25280 17153
rect 20996 17008 21048 17060
rect 22744 17008 22796 17060
rect 24032 17051 24084 17060
rect 24032 17017 24041 17051
rect 24041 17017 24075 17051
rect 24075 17017 24084 17051
rect 24032 17008 24084 17017
rect 24124 17008 24176 17060
rect 19432 16983 19484 16992
rect 19432 16949 19441 16983
rect 19441 16949 19475 16983
rect 19475 16949 19484 16983
rect 19432 16940 19484 16949
rect 21824 16983 21876 16992
rect 21824 16949 21833 16983
rect 21833 16949 21867 16983
rect 21867 16949 21876 16983
rect 21824 16940 21876 16949
rect 23388 16983 23440 16992
rect 23388 16949 23397 16983
rect 23397 16949 23431 16983
rect 23431 16949 23440 16983
rect 25136 17008 25188 17060
rect 25044 16983 25096 16992
rect 23388 16940 23440 16949
rect 25044 16949 25053 16983
rect 25053 16949 25087 16983
rect 25087 16949 25096 16983
rect 25044 16940 25096 16949
rect 25504 16940 25556 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1676 16779 1728 16788
rect 1676 16745 1685 16779
rect 1685 16745 1719 16779
rect 1719 16745 1728 16779
rect 1676 16736 1728 16745
rect 1768 16736 1820 16788
rect 2228 16736 2280 16788
rect 5448 16779 5500 16788
rect 5448 16745 5457 16779
rect 5457 16745 5491 16779
rect 5491 16745 5500 16779
rect 5448 16736 5500 16745
rect 5540 16736 5592 16788
rect 6920 16779 6972 16788
rect 6920 16745 6929 16779
rect 6929 16745 6963 16779
rect 6963 16745 6972 16779
rect 6920 16736 6972 16745
rect 8760 16736 8812 16788
rect 9128 16779 9180 16788
rect 9128 16745 9137 16779
rect 9137 16745 9171 16779
rect 9171 16745 9180 16779
rect 9128 16736 9180 16745
rect 9864 16736 9916 16788
rect 12348 16736 12400 16788
rect 3424 16668 3476 16720
rect 8208 16668 8260 16720
rect 1952 16600 2004 16652
rect 2136 16643 2188 16652
rect 2136 16609 2145 16643
rect 2145 16609 2179 16643
rect 2179 16609 2188 16643
rect 2136 16600 2188 16609
rect 2872 16643 2924 16652
rect 2872 16609 2881 16643
rect 2881 16609 2915 16643
rect 2915 16609 2924 16643
rect 2872 16600 2924 16609
rect 3240 16643 3292 16652
rect 3240 16609 3249 16643
rect 3249 16609 3283 16643
rect 3283 16609 3292 16643
rect 3240 16600 3292 16609
rect 4804 16600 4856 16652
rect 8392 16643 8444 16652
rect 8392 16609 8401 16643
rect 8401 16609 8435 16643
rect 8435 16609 8444 16643
rect 8392 16600 8444 16609
rect 9772 16668 9824 16720
rect 12256 16711 12308 16720
rect 12256 16677 12265 16711
rect 12265 16677 12299 16711
rect 12299 16677 12308 16711
rect 12256 16668 12308 16677
rect 13084 16711 13136 16720
rect 13084 16677 13093 16711
rect 13093 16677 13127 16711
rect 13127 16677 13136 16711
rect 13084 16668 13136 16677
rect 13728 16668 13780 16720
rect 13912 16711 13964 16720
rect 13912 16677 13921 16711
rect 13921 16677 13955 16711
rect 13955 16677 13964 16711
rect 13912 16668 13964 16677
rect 14188 16736 14240 16788
rect 19156 16736 19208 16788
rect 19524 16736 19576 16788
rect 21824 16736 21876 16788
rect 15292 16668 15344 16720
rect 9496 16600 9548 16652
rect 9220 16532 9272 16584
rect 10968 16600 11020 16652
rect 14556 16600 14608 16652
rect 15844 16668 15896 16720
rect 18144 16711 18196 16720
rect 18144 16677 18153 16711
rect 18153 16677 18187 16711
rect 18187 16677 18196 16711
rect 18144 16668 18196 16677
rect 18328 16711 18380 16720
rect 18328 16677 18337 16711
rect 18337 16677 18371 16711
rect 18371 16677 18380 16711
rect 18328 16668 18380 16677
rect 19984 16668 20036 16720
rect 10140 16532 10192 16584
rect 9588 16464 9640 16516
rect 11980 16464 12032 16516
rect 13084 16532 13136 16584
rect 13360 16532 13412 16584
rect 14648 16532 14700 16584
rect 15292 16575 15344 16584
rect 15292 16541 15301 16575
rect 15301 16541 15335 16575
rect 15335 16541 15344 16575
rect 15292 16532 15344 16541
rect 6736 16396 6788 16448
rect 7104 16396 7156 16448
rect 8116 16439 8168 16448
rect 8116 16405 8125 16439
rect 8125 16405 8159 16439
rect 8159 16405 8168 16439
rect 8116 16396 8168 16405
rect 11336 16396 11388 16448
rect 15476 16396 15528 16448
rect 16948 16600 17000 16652
rect 17500 16532 17552 16584
rect 18696 16600 18748 16652
rect 22376 16736 22428 16788
rect 23388 16736 23440 16788
rect 23664 16736 23716 16788
rect 22284 16711 22336 16720
rect 22284 16677 22293 16711
rect 22293 16677 22327 16711
rect 22327 16677 22336 16711
rect 22284 16668 22336 16677
rect 22560 16668 22612 16720
rect 23296 16668 23348 16720
rect 22744 16600 22796 16652
rect 24032 16600 24084 16652
rect 22468 16532 22520 16584
rect 23020 16532 23072 16584
rect 17868 16439 17920 16448
rect 17868 16405 17877 16439
rect 17877 16405 17911 16439
rect 17911 16405 17920 16439
rect 17868 16396 17920 16405
rect 21824 16439 21876 16448
rect 21824 16405 21833 16439
rect 21833 16405 21867 16439
rect 21867 16405 21876 16439
rect 21824 16396 21876 16405
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2228 16192 2280 16244
rect 3424 16235 3476 16244
rect 3424 16201 3433 16235
rect 3433 16201 3467 16235
rect 3467 16201 3476 16235
rect 3424 16192 3476 16201
rect 8944 16235 8996 16244
rect 8944 16201 8953 16235
rect 8953 16201 8987 16235
rect 8987 16201 8996 16235
rect 8944 16192 8996 16201
rect 9220 16235 9272 16244
rect 9220 16201 9229 16235
rect 9229 16201 9263 16235
rect 9263 16201 9272 16235
rect 9220 16192 9272 16201
rect 10140 16235 10192 16244
rect 10140 16201 10149 16235
rect 10149 16201 10183 16235
rect 10183 16201 10192 16235
rect 10140 16192 10192 16201
rect 13084 16192 13136 16244
rect 13820 16192 13872 16244
rect 14648 16235 14700 16244
rect 14648 16201 14657 16235
rect 14657 16201 14691 16235
rect 14691 16201 14700 16235
rect 14648 16192 14700 16201
rect 14740 16192 14792 16244
rect 15292 16192 15344 16244
rect 15844 16192 15896 16244
rect 16212 16192 16264 16244
rect 17500 16235 17552 16244
rect 17500 16201 17509 16235
rect 17509 16201 17543 16235
rect 17543 16201 17552 16235
rect 17500 16192 17552 16201
rect 18144 16192 18196 16244
rect 18328 16235 18380 16244
rect 18328 16201 18337 16235
rect 18337 16201 18371 16235
rect 18371 16201 18380 16235
rect 18328 16192 18380 16201
rect 23020 16192 23072 16244
rect 24032 16192 24084 16244
rect 4252 16124 4304 16176
rect 4620 16124 4672 16176
rect 7380 16167 7432 16176
rect 7380 16133 7389 16167
rect 7389 16133 7423 16167
rect 7423 16133 7432 16167
rect 7380 16124 7432 16133
rect 11980 16124 12032 16176
rect 18880 16167 18932 16176
rect 3056 16099 3108 16108
rect 3056 16065 3065 16099
rect 3065 16065 3099 16099
rect 3099 16065 3108 16099
rect 3056 16056 3108 16065
rect 6736 16056 6788 16108
rect 9404 16056 9456 16108
rect 9588 16099 9640 16108
rect 9588 16065 9597 16099
rect 9597 16065 9631 16099
rect 9631 16065 9640 16099
rect 9588 16056 9640 16065
rect 9864 16056 9916 16108
rect 12348 16056 12400 16108
rect 18880 16133 18889 16167
rect 18889 16133 18923 16167
rect 18923 16133 18932 16167
rect 18880 16124 18932 16133
rect 14832 16056 14884 16108
rect 16948 16099 17000 16108
rect 16948 16065 16957 16099
rect 16957 16065 16991 16099
rect 16991 16065 17000 16099
rect 16948 16056 17000 16065
rect 23572 16056 23624 16108
rect 24860 16056 24912 16108
rect 3332 15988 3384 16040
rect 6644 15988 6696 16040
rect 13176 16031 13228 16040
rect 13176 15997 13185 16031
rect 13185 15997 13219 16031
rect 13219 15997 13228 16031
rect 13176 15988 13228 15997
rect 14648 15988 14700 16040
rect 19156 16031 19208 16040
rect 19156 15997 19165 16031
rect 19165 15997 19199 16031
rect 19199 15997 19208 16031
rect 19156 15988 19208 15997
rect 20904 15988 20956 16040
rect 23020 15988 23072 16040
rect 8024 15920 8076 15972
rect 8944 15920 8996 15972
rect 10784 15920 10836 15972
rect 1400 15895 1452 15904
rect 1400 15861 1409 15895
rect 1409 15861 1443 15895
rect 1443 15861 1452 15895
rect 1400 15852 1452 15861
rect 3332 15852 3384 15904
rect 4804 15852 4856 15904
rect 6828 15852 6880 15904
rect 7012 15852 7064 15904
rect 8208 15852 8260 15904
rect 8392 15895 8444 15904
rect 8392 15861 8401 15895
rect 8401 15861 8435 15895
rect 8435 15861 8444 15895
rect 8392 15852 8444 15861
rect 11336 15895 11388 15904
rect 11336 15861 11345 15895
rect 11345 15861 11379 15895
rect 11379 15861 11388 15895
rect 11336 15852 11388 15861
rect 13636 15963 13688 15972
rect 13636 15929 13645 15963
rect 13645 15929 13679 15963
rect 13679 15929 13688 15963
rect 13636 15920 13688 15929
rect 13820 15963 13872 15972
rect 13820 15929 13829 15963
rect 13829 15929 13863 15963
rect 13863 15929 13872 15963
rect 13820 15920 13872 15929
rect 15476 15963 15528 15972
rect 15476 15929 15485 15963
rect 15485 15929 15519 15963
rect 15519 15929 15528 15963
rect 15476 15920 15528 15929
rect 15660 15920 15712 15972
rect 17040 15963 17092 15972
rect 17040 15929 17049 15963
rect 17049 15929 17083 15963
rect 17083 15929 17092 15963
rect 17040 15920 17092 15929
rect 18144 15920 18196 15972
rect 19984 15920 20036 15972
rect 21088 15963 21140 15972
rect 21088 15929 21122 15963
rect 21122 15929 21140 15963
rect 21088 15920 21140 15929
rect 22284 15920 22336 15972
rect 24216 15988 24268 16040
rect 24676 15988 24728 16040
rect 12348 15852 12400 15904
rect 15568 15852 15620 15904
rect 15844 15895 15896 15904
rect 15844 15861 15853 15895
rect 15853 15861 15887 15895
rect 15887 15861 15896 15895
rect 15844 15852 15896 15861
rect 16396 15852 16448 15904
rect 18604 15895 18656 15904
rect 18604 15861 18613 15895
rect 18613 15861 18647 15895
rect 18647 15861 18656 15895
rect 18604 15852 18656 15861
rect 20904 15852 20956 15904
rect 21916 15852 21968 15904
rect 23480 15852 23532 15904
rect 25688 15852 25740 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 2780 15648 2832 15700
rect 6644 15691 6696 15700
rect 6644 15657 6653 15691
rect 6653 15657 6687 15691
rect 6687 15657 6696 15691
rect 6644 15648 6696 15657
rect 7012 15648 7064 15700
rect 8300 15691 8352 15700
rect 8300 15657 8309 15691
rect 8309 15657 8343 15691
rect 8343 15657 8352 15691
rect 8300 15648 8352 15657
rect 8760 15691 8812 15700
rect 8760 15657 8769 15691
rect 8769 15657 8803 15691
rect 8803 15657 8812 15691
rect 8760 15648 8812 15657
rect 9588 15648 9640 15700
rect 10968 15648 11020 15700
rect 11980 15691 12032 15700
rect 11980 15657 11989 15691
rect 11989 15657 12023 15691
rect 12023 15657 12032 15691
rect 11980 15648 12032 15657
rect 13544 15648 13596 15700
rect 15568 15648 15620 15700
rect 15752 15691 15804 15700
rect 15752 15657 15761 15691
rect 15761 15657 15795 15691
rect 15795 15657 15804 15691
rect 15752 15648 15804 15657
rect 16856 15648 16908 15700
rect 17408 15648 17460 15700
rect 21272 15648 21324 15700
rect 22284 15648 22336 15700
rect 22468 15648 22520 15700
rect 23480 15648 23532 15700
rect 4804 15580 4856 15632
rect 1584 15512 1636 15564
rect 2872 15512 2924 15564
rect 4068 15555 4120 15564
rect 4068 15521 4077 15555
rect 4077 15521 4111 15555
rect 4111 15521 4120 15555
rect 4068 15512 4120 15521
rect 6092 15580 6144 15632
rect 9956 15580 10008 15632
rect 13912 15580 13964 15632
rect 15476 15580 15528 15632
rect 15660 15623 15712 15632
rect 15660 15589 15669 15623
rect 15669 15589 15703 15623
rect 15703 15589 15712 15623
rect 15660 15580 15712 15589
rect 18880 15623 18932 15632
rect 18880 15589 18889 15623
rect 18889 15589 18923 15623
rect 18923 15589 18932 15623
rect 18880 15580 18932 15589
rect 5540 15555 5592 15564
rect 5540 15521 5574 15555
rect 5574 15521 5592 15555
rect 5540 15512 5592 15521
rect 7104 15512 7156 15564
rect 8024 15512 8076 15564
rect 9680 15512 9732 15564
rect 12164 15512 12216 15564
rect 12992 15512 13044 15564
rect 15384 15512 15436 15564
rect 16396 15555 16448 15564
rect 16396 15521 16405 15555
rect 16405 15521 16439 15555
rect 16439 15521 16448 15555
rect 16396 15512 16448 15521
rect 8208 15487 8260 15496
rect 8208 15453 8217 15487
rect 8217 15453 8251 15487
rect 8251 15453 8260 15487
rect 8208 15444 8260 15453
rect 9404 15444 9456 15496
rect 9864 15444 9916 15496
rect 11704 15444 11756 15496
rect 12440 15487 12492 15496
rect 12440 15453 12449 15487
rect 12449 15453 12483 15487
rect 12483 15453 12492 15487
rect 12440 15444 12492 15453
rect 14556 15444 14608 15496
rect 16672 15512 16724 15564
rect 16580 15444 16632 15496
rect 18144 15444 18196 15496
rect 2504 15376 2556 15428
rect 9772 15419 9824 15428
rect 9772 15385 9781 15419
rect 9781 15385 9815 15419
rect 9815 15385 9824 15419
rect 9772 15376 9824 15385
rect 18880 15376 18932 15428
rect 22652 15580 22704 15632
rect 23020 15623 23072 15632
rect 23020 15589 23029 15623
rect 23029 15589 23063 15623
rect 23063 15589 23072 15623
rect 23020 15580 23072 15589
rect 23204 15580 23256 15632
rect 24400 15623 24452 15632
rect 24400 15589 24409 15623
rect 24409 15589 24443 15623
rect 24443 15589 24452 15623
rect 24400 15580 24452 15589
rect 20812 15512 20864 15564
rect 22008 15512 22060 15564
rect 19156 15487 19208 15496
rect 19156 15453 19165 15487
rect 19165 15453 19199 15487
rect 19199 15453 19208 15487
rect 19156 15444 19208 15453
rect 19984 15444 20036 15496
rect 21916 15444 21968 15496
rect 23480 15512 23532 15564
rect 25136 15580 25188 15632
rect 24860 15512 24912 15564
rect 20996 15419 21048 15428
rect 20996 15385 21005 15419
rect 21005 15385 21039 15419
rect 21039 15385 21048 15419
rect 20996 15376 21048 15385
rect 2596 15308 2648 15360
rect 3792 15308 3844 15360
rect 5080 15351 5132 15360
rect 5080 15317 5089 15351
rect 5089 15317 5123 15351
rect 5123 15317 5132 15351
rect 5080 15308 5132 15317
rect 7840 15351 7892 15360
rect 7840 15317 7849 15351
rect 7849 15317 7883 15351
rect 7883 15317 7892 15351
rect 7840 15308 7892 15317
rect 10692 15351 10744 15360
rect 10692 15317 10701 15351
rect 10701 15317 10735 15351
rect 10735 15317 10744 15351
rect 10692 15308 10744 15317
rect 19248 15308 19300 15360
rect 20720 15308 20772 15360
rect 24768 15308 24820 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 2136 15104 2188 15156
rect 2872 15147 2924 15156
rect 2872 15113 2881 15147
rect 2881 15113 2915 15147
rect 2915 15113 2924 15147
rect 2872 15104 2924 15113
rect 3608 15147 3660 15156
rect 3608 15113 3617 15147
rect 3617 15113 3651 15147
rect 3651 15113 3660 15147
rect 3608 15104 3660 15113
rect 4160 15147 4212 15156
rect 4160 15113 4169 15147
rect 4169 15113 4203 15147
rect 4203 15113 4212 15147
rect 4160 15104 4212 15113
rect 5540 15104 5592 15156
rect 6184 15147 6236 15156
rect 6184 15113 6193 15147
rect 6193 15113 6227 15147
rect 6227 15113 6236 15147
rect 6184 15104 6236 15113
rect 6920 15147 6972 15156
rect 6920 15113 6929 15147
rect 6929 15113 6963 15147
rect 6963 15113 6972 15147
rect 6920 15104 6972 15113
rect 7012 15104 7064 15156
rect 8300 15104 8352 15156
rect 10140 15104 10192 15156
rect 1768 14968 1820 15020
rect 2504 15036 2556 15088
rect 11428 15104 11480 15156
rect 2688 14968 2740 15020
rect 3056 14900 3108 14952
rect 3608 14900 3660 14952
rect 4068 14900 4120 14952
rect 4804 14900 4856 14952
rect 6736 14900 6788 14952
rect 9036 14943 9088 14952
rect 9036 14909 9045 14943
rect 9045 14909 9079 14943
rect 9079 14909 9088 14943
rect 9036 14900 9088 14909
rect 11704 14900 11756 14952
rect 12440 15104 12492 15156
rect 16488 15147 16540 15156
rect 16488 15113 16497 15147
rect 16497 15113 16531 15147
rect 16531 15113 16540 15147
rect 16488 15104 16540 15113
rect 16672 15104 16724 15156
rect 17408 15147 17460 15156
rect 17408 15113 17417 15147
rect 17417 15113 17451 15147
rect 17451 15113 17460 15147
rect 17408 15104 17460 15113
rect 19984 15147 20036 15156
rect 19984 15113 19993 15147
rect 19993 15113 20027 15147
rect 20027 15113 20036 15147
rect 19984 15104 20036 15113
rect 20812 15104 20864 15156
rect 21272 15104 21324 15156
rect 21640 15104 21692 15156
rect 21916 15147 21968 15156
rect 21916 15113 21925 15147
rect 21925 15113 21959 15147
rect 21959 15113 21968 15147
rect 21916 15104 21968 15113
rect 22652 15147 22704 15156
rect 22652 15113 22661 15147
rect 22661 15113 22695 15147
rect 22695 15113 22704 15147
rect 22652 15104 22704 15113
rect 23480 15147 23532 15156
rect 23480 15113 23489 15147
rect 23489 15113 23523 15147
rect 23523 15113 23532 15147
rect 23480 15104 23532 15113
rect 24676 15147 24728 15156
rect 24676 15113 24685 15147
rect 24685 15113 24719 15147
rect 24719 15113 24728 15147
rect 24676 15104 24728 15113
rect 13268 15036 13320 15088
rect 15108 15079 15160 15088
rect 15108 15045 15117 15079
rect 15117 15045 15151 15079
rect 15151 15045 15160 15079
rect 15108 15036 15160 15045
rect 20628 15079 20680 15088
rect 20628 15045 20637 15079
rect 20637 15045 20671 15079
rect 20671 15045 20680 15079
rect 20628 15036 20680 15045
rect 23756 15079 23808 15088
rect 23756 15045 23765 15079
rect 23765 15045 23799 15079
rect 23799 15045 23808 15079
rect 23756 15036 23808 15045
rect 13084 15011 13136 15020
rect 13084 14977 13093 15011
rect 13093 14977 13127 15011
rect 13127 14977 13136 15011
rect 13912 15011 13964 15020
rect 13084 14968 13136 14977
rect 13912 14977 13921 15011
rect 13921 14977 13955 15011
rect 13955 14977 13964 15011
rect 13912 14968 13964 14977
rect 15384 14968 15436 15020
rect 20996 15011 21048 15020
rect 20996 14977 21005 15011
rect 21005 14977 21039 15011
rect 21039 14977 21048 15011
rect 20996 14968 21048 14977
rect 22100 15011 22152 15020
rect 22100 14977 22109 15011
rect 22109 14977 22143 15011
rect 22143 14977 22152 15011
rect 22100 14968 22152 14977
rect 1952 14875 2004 14884
rect 1952 14841 1961 14875
rect 1961 14841 1995 14875
rect 1995 14841 2004 14875
rect 1952 14832 2004 14841
rect 2596 14832 2648 14884
rect 4344 14832 4396 14884
rect 5080 14832 5132 14884
rect 7104 14832 7156 14884
rect 7380 14875 7432 14884
rect 7380 14841 7389 14875
rect 7389 14841 7423 14875
rect 7423 14841 7432 14875
rect 7380 14832 7432 14841
rect 7472 14875 7524 14884
rect 7472 14841 7481 14875
rect 7481 14841 7515 14875
rect 7515 14841 7524 14875
rect 8300 14875 8352 14884
rect 7472 14832 7524 14841
rect 8300 14841 8309 14875
rect 8309 14841 8343 14875
rect 8343 14841 8352 14875
rect 8300 14832 8352 14841
rect 9496 14832 9548 14884
rect 10692 14832 10744 14884
rect 13820 14900 13872 14952
rect 16396 14900 16448 14952
rect 15844 14832 15896 14884
rect 18144 14900 18196 14952
rect 19524 14832 19576 14884
rect 1584 14764 1636 14816
rect 2136 14764 2188 14816
rect 3148 14807 3200 14816
rect 3148 14773 3157 14807
rect 3157 14773 3191 14807
rect 3191 14773 3200 14807
rect 3148 14764 3200 14773
rect 8484 14807 8536 14816
rect 8484 14773 8493 14807
rect 8493 14773 8527 14807
rect 8527 14773 8536 14807
rect 8484 14764 8536 14773
rect 9588 14764 9640 14816
rect 9772 14807 9824 14816
rect 9772 14773 9781 14807
rect 9781 14773 9815 14807
rect 9815 14773 9824 14807
rect 9772 14764 9824 14773
rect 9956 14764 10008 14816
rect 11244 14807 11296 14816
rect 11244 14773 11253 14807
rect 11253 14773 11287 14807
rect 11287 14773 11296 14807
rect 11244 14764 11296 14773
rect 14464 14807 14516 14816
rect 14464 14773 14473 14807
rect 14473 14773 14507 14807
rect 14507 14773 14516 14807
rect 14464 14764 14516 14773
rect 16948 14807 17000 14816
rect 16948 14773 16957 14807
rect 16957 14773 16991 14807
rect 16991 14773 17000 14807
rect 16948 14764 17000 14773
rect 19156 14764 19208 14816
rect 19984 14900 20036 14952
rect 24032 14943 24084 14952
rect 24032 14909 24041 14943
rect 24041 14909 24075 14943
rect 24075 14909 24084 14943
rect 24032 14900 24084 14909
rect 24952 14900 25004 14952
rect 20720 14832 20772 14884
rect 21180 14875 21232 14884
rect 21180 14841 21189 14875
rect 21189 14841 21223 14875
rect 21223 14841 21232 14875
rect 21180 14832 21232 14841
rect 22836 14832 22888 14884
rect 25044 14875 25096 14884
rect 25044 14841 25053 14875
rect 25053 14841 25087 14875
rect 25087 14841 25096 14875
rect 25044 14832 25096 14841
rect 22100 14764 22152 14816
rect 23020 14764 23072 14816
rect 25596 14764 25648 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1400 14492 1452 14544
rect 2044 14535 2096 14544
rect 2044 14501 2053 14535
rect 2053 14501 2087 14535
rect 2087 14501 2096 14535
rect 2044 14492 2096 14501
rect 2228 14535 2280 14544
rect 2228 14501 2237 14535
rect 2237 14501 2271 14535
rect 2271 14501 2280 14535
rect 2228 14492 2280 14501
rect 2320 14535 2372 14544
rect 2320 14501 2329 14535
rect 2329 14501 2363 14535
rect 2363 14501 2372 14535
rect 2872 14560 2924 14612
rect 4344 14560 4396 14612
rect 5080 14560 5132 14612
rect 5540 14560 5592 14612
rect 7472 14560 7524 14612
rect 8392 14603 8444 14612
rect 8392 14569 8401 14603
rect 8401 14569 8435 14603
rect 8435 14569 8444 14603
rect 8392 14560 8444 14569
rect 8944 14560 8996 14612
rect 9404 14603 9456 14612
rect 9404 14569 9413 14603
rect 9413 14569 9447 14603
rect 9447 14569 9456 14603
rect 9404 14560 9456 14569
rect 9864 14560 9916 14612
rect 13084 14560 13136 14612
rect 14280 14560 14332 14612
rect 16948 14560 17000 14612
rect 18420 14560 18472 14612
rect 18880 14603 18932 14612
rect 18880 14569 18889 14603
rect 18889 14569 18923 14603
rect 18923 14569 18932 14603
rect 18880 14560 18932 14569
rect 19340 14560 19392 14612
rect 21180 14560 21232 14612
rect 22836 14603 22888 14612
rect 22836 14569 22845 14603
rect 22845 14569 22879 14603
rect 22879 14569 22888 14603
rect 22836 14560 22888 14569
rect 24032 14560 24084 14612
rect 2320 14492 2372 14501
rect 8116 14492 8168 14544
rect 2504 14424 2556 14476
rect 3332 14424 3384 14476
rect 7104 14424 7156 14476
rect 10232 14467 10284 14476
rect 10232 14433 10241 14467
rect 10241 14433 10275 14467
rect 10275 14433 10284 14467
rect 17316 14492 17368 14544
rect 17868 14492 17920 14544
rect 19156 14492 19208 14544
rect 23388 14492 23440 14544
rect 10232 14424 10284 14433
rect 12164 14424 12216 14476
rect 13452 14467 13504 14476
rect 13452 14433 13461 14467
rect 13461 14433 13495 14467
rect 13495 14433 13504 14467
rect 13452 14424 13504 14433
rect 15568 14424 15620 14476
rect 16396 14424 16448 14476
rect 19340 14424 19392 14476
rect 20628 14424 20680 14476
rect 20996 14424 21048 14476
rect 4068 14399 4120 14408
rect 4068 14365 4077 14399
rect 4077 14365 4111 14399
rect 4111 14365 4120 14399
rect 4068 14356 4120 14365
rect 10508 14399 10560 14408
rect 1768 14331 1820 14340
rect 1768 14297 1777 14331
rect 1777 14297 1811 14331
rect 1811 14297 1820 14331
rect 1768 14288 1820 14297
rect 6644 14288 6696 14340
rect 10508 14365 10517 14399
rect 10517 14365 10551 14399
rect 10551 14365 10560 14399
rect 10508 14356 10560 14365
rect 11244 14356 11296 14408
rect 8208 14288 8260 14340
rect 10968 14288 11020 14340
rect 3608 14220 3660 14272
rect 4068 14220 4120 14272
rect 7288 14263 7340 14272
rect 7288 14229 7297 14263
rect 7297 14229 7331 14263
rect 7331 14229 7340 14263
rect 7288 14220 7340 14229
rect 9036 14220 9088 14272
rect 11152 14220 11204 14272
rect 16028 14356 16080 14408
rect 17408 14399 17460 14408
rect 17408 14365 17417 14399
rect 17417 14365 17451 14399
rect 17451 14365 17460 14399
rect 17408 14356 17460 14365
rect 19892 14399 19944 14408
rect 19892 14365 19901 14399
rect 19901 14365 19935 14399
rect 19935 14365 19944 14399
rect 19892 14356 19944 14365
rect 20904 14399 20956 14408
rect 20904 14365 20913 14399
rect 20913 14365 20947 14399
rect 20947 14365 20956 14399
rect 20904 14356 20956 14365
rect 23388 14399 23440 14408
rect 23388 14365 23397 14399
rect 23397 14365 23431 14399
rect 23431 14365 23440 14399
rect 23388 14356 23440 14365
rect 15384 14331 15436 14340
rect 15384 14297 15393 14331
rect 15393 14297 15427 14331
rect 15427 14297 15436 14331
rect 15384 14288 15436 14297
rect 11704 14220 11756 14272
rect 16948 14263 17000 14272
rect 16948 14229 16957 14263
rect 16957 14229 16991 14263
rect 16991 14229 17000 14263
rect 16948 14220 17000 14229
rect 20536 14220 20588 14272
rect 22284 14263 22336 14272
rect 22284 14229 22293 14263
rect 22293 14229 22327 14263
rect 22327 14229 22336 14263
rect 22284 14220 22336 14229
rect 22836 14220 22888 14272
rect 24952 14220 25004 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1952 14016 2004 14068
rect 2044 14016 2096 14068
rect 3332 14059 3384 14068
rect 3332 14025 3341 14059
rect 3341 14025 3375 14059
rect 3375 14025 3384 14059
rect 3332 14016 3384 14025
rect 4160 14016 4212 14068
rect 6644 14059 6696 14068
rect 6644 14025 6653 14059
rect 6653 14025 6687 14059
rect 6687 14025 6696 14059
rect 6644 14016 6696 14025
rect 6920 14059 6972 14068
rect 6920 14025 6929 14059
rect 6929 14025 6963 14059
rect 6963 14025 6972 14059
rect 6920 14016 6972 14025
rect 10508 14016 10560 14068
rect 12164 14059 12216 14068
rect 12164 14025 12173 14059
rect 12173 14025 12207 14059
rect 12207 14025 12216 14059
rect 12164 14016 12216 14025
rect 2504 13991 2556 14000
rect 2504 13957 2513 13991
rect 2513 13957 2547 13991
rect 2547 13957 2556 13991
rect 2504 13948 2556 13957
rect 3608 13948 3660 14000
rect 8392 13948 8444 14000
rect 10140 13948 10192 14000
rect 10968 13948 11020 14000
rect 11060 13948 11112 14000
rect 14464 14016 14516 14068
rect 16396 14059 16448 14068
rect 16396 14025 16405 14059
rect 16405 14025 16439 14059
rect 16439 14025 16448 14059
rect 16396 14016 16448 14025
rect 17316 14059 17368 14068
rect 17316 14025 17325 14059
rect 17325 14025 17359 14059
rect 17359 14025 17368 14059
rect 17316 14016 17368 14025
rect 17408 14016 17460 14068
rect 19892 14016 19944 14068
rect 20996 14059 21048 14068
rect 20996 14025 21005 14059
rect 21005 14025 21039 14059
rect 21039 14025 21048 14059
rect 20996 14016 21048 14025
rect 25044 14059 25096 14068
rect 25044 14025 25053 14059
rect 25053 14025 25087 14059
rect 25087 14025 25096 14059
rect 25044 14016 25096 14025
rect 2320 13880 2372 13932
rect 2780 13880 2832 13932
rect 4068 13880 4120 13932
rect 5632 13923 5684 13932
rect 5632 13889 5641 13923
rect 5641 13889 5675 13923
rect 5675 13889 5684 13923
rect 5632 13880 5684 13889
rect 7288 13880 7340 13932
rect 11152 13880 11204 13932
rect 14280 13948 14332 14000
rect 17776 13991 17828 14000
rect 17776 13957 17785 13991
rect 17785 13957 17819 13991
rect 17819 13957 17828 13991
rect 19524 13991 19576 14000
rect 17776 13948 17828 13957
rect 1768 13855 1820 13864
rect 1768 13821 1777 13855
rect 1777 13821 1811 13855
rect 1811 13821 1820 13855
rect 1768 13812 1820 13821
rect 5540 13812 5592 13864
rect 6828 13812 6880 13864
rect 7472 13855 7524 13864
rect 7472 13821 7481 13855
rect 7481 13821 7515 13855
rect 7515 13821 7524 13855
rect 7472 13812 7524 13821
rect 8116 13812 8168 13864
rect 8760 13855 8812 13864
rect 8760 13821 8769 13855
rect 8769 13821 8803 13855
rect 8803 13821 8812 13855
rect 8760 13812 8812 13821
rect 9036 13855 9088 13864
rect 9036 13821 9045 13855
rect 9045 13821 9079 13855
rect 9079 13821 9088 13855
rect 9036 13812 9088 13821
rect 4068 13787 4120 13796
rect 4068 13753 4077 13787
rect 4077 13753 4111 13787
rect 4111 13753 4120 13787
rect 4068 13744 4120 13753
rect 4528 13744 4580 13796
rect 6736 13744 6788 13796
rect 8944 13787 8996 13796
rect 8944 13753 8953 13787
rect 8953 13753 8987 13787
rect 8987 13753 8996 13787
rect 8944 13744 8996 13753
rect 11336 13812 11388 13864
rect 13452 13812 13504 13864
rect 15016 13855 15068 13864
rect 15016 13821 15025 13855
rect 15025 13821 15059 13855
rect 15059 13821 15068 13855
rect 15016 13812 15068 13821
rect 16028 13812 16080 13864
rect 19524 13957 19533 13991
rect 19533 13957 19567 13991
rect 19567 13957 19576 13991
rect 19524 13948 19576 13957
rect 18696 13923 18748 13932
rect 18696 13889 18705 13923
rect 18705 13889 18739 13923
rect 18739 13889 18748 13923
rect 18696 13880 18748 13889
rect 18420 13855 18472 13864
rect 18420 13821 18429 13855
rect 18429 13821 18463 13855
rect 18463 13821 18472 13855
rect 18420 13812 18472 13821
rect 20904 13812 20956 13864
rect 23388 13855 23440 13864
rect 23388 13821 23397 13855
rect 23397 13821 23431 13855
rect 23431 13821 23440 13855
rect 23388 13812 23440 13821
rect 24952 13812 25004 13864
rect 18880 13744 18932 13796
rect 19984 13744 20036 13796
rect 1952 13719 2004 13728
rect 1952 13685 1961 13719
rect 1961 13685 1995 13719
rect 1995 13685 2004 13719
rect 1952 13676 2004 13685
rect 3608 13676 3660 13728
rect 5632 13719 5684 13728
rect 5632 13685 5641 13719
rect 5641 13685 5675 13719
rect 5675 13685 5684 13719
rect 5632 13676 5684 13685
rect 7840 13676 7892 13728
rect 10140 13676 10192 13728
rect 11704 13676 11756 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 1768 13472 1820 13524
rect 2044 13404 2096 13456
rect 3056 13472 3108 13524
rect 3884 13472 3936 13524
rect 4068 13472 4120 13524
rect 5448 13515 5500 13524
rect 5448 13481 5457 13515
rect 5457 13481 5491 13515
rect 5491 13481 5500 13515
rect 5448 13472 5500 13481
rect 6828 13472 6880 13524
rect 7104 13472 7156 13524
rect 7840 13515 7892 13524
rect 7840 13481 7849 13515
rect 7849 13481 7883 13515
rect 7883 13481 7892 13515
rect 7840 13472 7892 13481
rect 8024 13472 8076 13524
rect 9864 13472 9916 13524
rect 11152 13472 11204 13524
rect 12348 13472 12400 13524
rect 18696 13472 18748 13524
rect 19248 13472 19300 13524
rect 19984 13472 20036 13524
rect 20996 13472 21048 13524
rect 23296 13472 23348 13524
rect 23572 13472 23624 13524
rect 2964 13447 3016 13456
rect 2964 13413 2973 13447
rect 2973 13413 3007 13447
rect 3007 13413 3016 13447
rect 2964 13404 3016 13413
rect 3976 13404 4028 13456
rect 4436 13404 4488 13456
rect 5540 13404 5592 13456
rect 5816 13447 5868 13456
rect 5816 13413 5850 13447
rect 5850 13413 5868 13447
rect 5816 13404 5868 13413
rect 8484 13404 8536 13456
rect 10692 13404 10744 13456
rect 12808 13404 12860 13456
rect 15568 13447 15620 13456
rect 15568 13413 15577 13447
rect 15577 13413 15611 13447
rect 15611 13413 15620 13447
rect 15568 13404 15620 13413
rect 16396 13404 16448 13456
rect 19340 13404 19392 13456
rect 19708 13404 19760 13456
rect 22560 13447 22612 13456
rect 22560 13413 22569 13447
rect 22569 13413 22603 13447
rect 22603 13413 22612 13447
rect 22560 13404 22612 13413
rect 22836 13404 22888 13456
rect 24124 13447 24176 13456
rect 24124 13413 24133 13447
rect 24133 13413 24167 13447
rect 24167 13413 24176 13447
rect 24124 13404 24176 13413
rect 24860 13404 24912 13456
rect 25044 13404 25096 13456
rect 4068 13379 4120 13388
rect 4068 13345 4077 13379
rect 4077 13345 4111 13379
rect 4111 13345 4120 13379
rect 4068 13336 4120 13345
rect 3240 13268 3292 13320
rect 5356 13268 5408 13320
rect 8760 13268 8812 13320
rect 9496 13268 9548 13320
rect 9864 13268 9916 13320
rect 10600 13268 10652 13320
rect 11704 13336 11756 13388
rect 12992 13336 13044 13388
rect 13728 13311 13780 13320
rect 13728 13277 13737 13311
rect 13737 13277 13771 13311
rect 13771 13277 13780 13311
rect 13728 13268 13780 13277
rect 19432 13336 19484 13388
rect 22468 13336 22520 13388
rect 13912 13268 13964 13320
rect 14280 13268 14332 13320
rect 15016 13311 15068 13320
rect 15016 13277 15025 13311
rect 15025 13277 15059 13311
rect 15059 13277 15068 13311
rect 15016 13268 15068 13277
rect 15844 13268 15896 13320
rect 16028 13268 16080 13320
rect 19064 13268 19116 13320
rect 4528 13200 4580 13252
rect 4712 13243 4764 13252
rect 4712 13209 4721 13243
rect 4721 13209 4755 13243
rect 4755 13209 4764 13243
rect 4712 13200 4764 13209
rect 8208 13200 8260 13252
rect 12532 13200 12584 13252
rect 25044 13268 25096 13320
rect 23664 13243 23716 13252
rect 23664 13209 23673 13243
rect 23673 13209 23707 13243
rect 23707 13209 23716 13243
rect 23664 13200 23716 13209
rect 1952 13175 2004 13184
rect 1952 13141 1961 13175
rect 1961 13141 1995 13175
rect 1995 13141 2004 13175
rect 1952 13132 2004 13141
rect 3976 13132 4028 13184
rect 9588 13132 9640 13184
rect 10140 13175 10192 13184
rect 10140 13141 10149 13175
rect 10149 13141 10183 13175
rect 10183 13141 10192 13175
rect 10140 13132 10192 13141
rect 17592 13175 17644 13184
rect 17592 13141 17601 13175
rect 17601 13141 17635 13175
rect 17635 13141 17644 13175
rect 17592 13132 17644 13141
rect 19800 13132 19852 13184
rect 21456 13175 21508 13184
rect 21456 13141 21465 13175
rect 21465 13141 21499 13175
rect 21499 13141 21508 13175
rect 21456 13132 21508 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 2872 12928 2924 12980
rect 3332 12928 3384 12980
rect 4160 12928 4212 12980
rect 6000 12971 6052 12980
rect 6000 12937 6009 12971
rect 6009 12937 6043 12971
rect 6043 12937 6052 12971
rect 6000 12928 6052 12937
rect 12808 12928 12860 12980
rect 13360 12971 13412 12980
rect 13360 12937 13369 12971
rect 13369 12937 13403 12971
rect 13403 12937 13412 12971
rect 13360 12928 13412 12937
rect 2044 12903 2096 12912
rect 2044 12869 2053 12903
rect 2053 12869 2087 12903
rect 2087 12869 2096 12903
rect 2044 12860 2096 12869
rect 6828 12860 6880 12912
rect 8024 12903 8076 12912
rect 8024 12869 8033 12903
rect 8033 12869 8067 12903
rect 8067 12869 8076 12903
rect 8024 12860 8076 12869
rect 14556 12928 14608 12980
rect 16396 12928 16448 12980
rect 16948 12928 17000 12980
rect 19064 12928 19116 12980
rect 19340 12971 19392 12980
rect 19340 12937 19349 12971
rect 19349 12937 19383 12971
rect 19383 12937 19392 12971
rect 19340 12928 19392 12937
rect 19708 12928 19760 12980
rect 22192 12928 22244 12980
rect 22560 12928 22612 12980
rect 22836 12971 22888 12980
rect 22836 12937 22845 12971
rect 22845 12937 22879 12971
rect 22879 12937 22888 12971
rect 22836 12928 22888 12937
rect 24124 12928 24176 12980
rect 25044 12971 25096 12980
rect 25044 12937 25053 12971
rect 25053 12937 25087 12971
rect 25087 12937 25096 12971
rect 25044 12928 25096 12937
rect 16028 12903 16080 12912
rect 4068 12792 4120 12844
rect 5172 12835 5224 12844
rect 5172 12801 5181 12835
rect 5181 12801 5215 12835
rect 5215 12801 5224 12835
rect 5172 12792 5224 12801
rect 5448 12792 5500 12844
rect 7472 12835 7524 12844
rect 7472 12801 7481 12835
rect 7481 12801 7515 12835
rect 7515 12801 7524 12835
rect 7472 12792 7524 12801
rect 8300 12792 8352 12844
rect 16028 12869 16037 12903
rect 16037 12869 16071 12903
rect 16071 12869 16080 12903
rect 16028 12860 16080 12869
rect 16488 12860 16540 12912
rect 13912 12835 13964 12844
rect 13912 12801 13921 12835
rect 13921 12801 13955 12835
rect 13955 12801 13964 12835
rect 13912 12792 13964 12801
rect 19524 12903 19576 12912
rect 19524 12869 19533 12903
rect 19533 12869 19567 12903
rect 19567 12869 19576 12903
rect 19524 12860 19576 12869
rect 21088 12903 21140 12912
rect 21088 12869 21097 12903
rect 21097 12869 21131 12903
rect 21131 12869 21140 12903
rect 21088 12860 21140 12869
rect 22468 12903 22520 12912
rect 22468 12869 22477 12903
rect 22477 12869 22511 12903
rect 22511 12869 22520 12903
rect 22468 12860 22520 12869
rect 2136 12767 2188 12776
rect 2136 12733 2145 12767
rect 2145 12733 2179 12767
rect 2179 12733 2188 12767
rect 2136 12724 2188 12733
rect 3884 12656 3936 12708
rect 4068 12656 4120 12708
rect 4712 12656 4764 12708
rect 10600 12724 10652 12776
rect 10784 12724 10836 12776
rect 8300 12656 8352 12708
rect 10876 12656 10928 12708
rect 17592 12724 17644 12776
rect 19800 12767 19852 12776
rect 19800 12733 19809 12767
rect 19809 12733 19843 12767
rect 19843 12733 19852 12767
rect 19800 12724 19852 12733
rect 21456 12792 21508 12844
rect 22008 12792 22060 12844
rect 14004 12656 14056 12708
rect 16764 12699 16816 12708
rect 16764 12665 16773 12699
rect 16773 12665 16807 12699
rect 16807 12665 16816 12699
rect 16764 12656 16816 12665
rect 18604 12699 18656 12708
rect 18604 12665 18613 12699
rect 18613 12665 18647 12699
rect 18647 12665 18656 12699
rect 18604 12656 18656 12665
rect 20076 12699 20128 12708
rect 20076 12665 20085 12699
rect 20085 12665 20119 12699
rect 20119 12665 20128 12699
rect 22100 12724 22152 12776
rect 22652 12724 22704 12776
rect 23112 12724 23164 12776
rect 20076 12656 20128 12665
rect 21548 12699 21600 12708
rect 21548 12665 21557 12699
rect 21557 12665 21591 12699
rect 21591 12665 21600 12699
rect 21548 12656 21600 12665
rect 5356 12588 5408 12640
rect 6092 12588 6144 12640
rect 7012 12588 7064 12640
rect 7748 12588 7800 12640
rect 8668 12588 8720 12640
rect 10692 12588 10744 12640
rect 11704 12588 11756 12640
rect 20812 12588 20864 12640
rect 23664 12724 23716 12776
rect 24216 12724 24268 12776
rect 24676 12724 24728 12776
rect 23388 12588 23440 12640
rect 23756 12588 23808 12640
rect 25412 12631 25464 12640
rect 25412 12597 25421 12631
rect 25421 12597 25455 12631
rect 25455 12597 25464 12631
rect 25412 12588 25464 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 2780 12384 2832 12436
rect 3240 12384 3292 12436
rect 8484 12427 8536 12436
rect 8484 12393 8493 12427
rect 8493 12393 8527 12427
rect 8527 12393 8536 12427
rect 8484 12384 8536 12393
rect 8760 12427 8812 12436
rect 8760 12393 8769 12427
rect 8769 12393 8803 12427
rect 8803 12393 8812 12427
rect 8760 12384 8812 12393
rect 11244 12384 11296 12436
rect 13820 12427 13872 12436
rect 13820 12393 13829 12427
rect 13829 12393 13863 12427
rect 13863 12393 13872 12427
rect 13820 12384 13872 12393
rect 16764 12427 16816 12436
rect 16764 12393 16773 12427
rect 16773 12393 16807 12427
rect 16807 12393 16816 12427
rect 16764 12384 16816 12393
rect 19984 12427 20036 12436
rect 19984 12393 19993 12427
rect 19993 12393 20027 12427
rect 20027 12393 20036 12427
rect 19984 12384 20036 12393
rect 22100 12384 22152 12436
rect 23756 12384 23808 12436
rect 23940 12384 23992 12436
rect 24676 12384 24728 12436
rect 3056 12359 3108 12368
rect 3056 12325 3065 12359
rect 3065 12325 3099 12359
rect 3099 12325 3108 12359
rect 3056 12316 3108 12325
rect 3332 12316 3384 12368
rect 7288 12316 7340 12368
rect 8944 12316 8996 12368
rect 14372 12316 14424 12368
rect 16212 12359 16264 12368
rect 16212 12325 16221 12359
rect 16221 12325 16255 12359
rect 16255 12325 16264 12359
rect 16212 12316 16264 12325
rect 17592 12316 17644 12368
rect 23112 12316 23164 12368
rect 24860 12316 24912 12368
rect 2136 12248 2188 12300
rect 5448 12248 5500 12300
rect 7380 12248 7432 12300
rect 7748 12291 7800 12300
rect 7748 12257 7757 12291
rect 7757 12257 7791 12291
rect 7791 12257 7800 12291
rect 7748 12248 7800 12257
rect 10048 12291 10100 12300
rect 10048 12257 10057 12291
rect 10057 12257 10091 12291
rect 10091 12257 10100 12291
rect 10048 12248 10100 12257
rect 12164 12291 12216 12300
rect 12164 12257 12198 12291
rect 12198 12257 12216 12291
rect 12164 12248 12216 12257
rect 15660 12248 15712 12300
rect 19432 12248 19484 12300
rect 21180 12291 21232 12300
rect 21180 12257 21214 12291
rect 21214 12257 21232 12291
rect 21180 12248 21232 12257
rect 1400 12223 1452 12232
rect 1400 12189 1409 12223
rect 1409 12189 1443 12223
rect 1443 12189 1452 12223
rect 1400 12180 1452 12189
rect 6000 12223 6052 12232
rect 6000 12189 6009 12223
rect 6009 12189 6043 12223
rect 6043 12189 6052 12223
rect 6000 12180 6052 12189
rect 7472 12180 7524 12232
rect 8024 12223 8076 12232
rect 8024 12189 8033 12223
rect 8033 12189 8067 12223
rect 8067 12189 8076 12223
rect 8024 12180 8076 12189
rect 9680 12180 9732 12232
rect 9864 12180 9916 12232
rect 10324 12223 10376 12232
rect 10324 12189 10333 12223
rect 10333 12189 10367 12223
rect 10367 12189 10376 12223
rect 10324 12180 10376 12189
rect 3332 12112 3384 12164
rect 7656 12112 7708 12164
rect 16120 12223 16172 12232
rect 16120 12189 16129 12223
rect 16129 12189 16163 12223
rect 16163 12189 16172 12223
rect 16120 12180 16172 12189
rect 16304 12223 16356 12232
rect 16304 12189 16313 12223
rect 16313 12189 16347 12223
rect 16347 12189 16356 12223
rect 16304 12180 16356 12189
rect 17224 12223 17276 12232
rect 17224 12189 17233 12223
rect 17233 12189 17267 12223
rect 17267 12189 17276 12223
rect 17224 12180 17276 12189
rect 20904 12223 20956 12232
rect 20904 12189 20913 12223
rect 20913 12189 20947 12223
rect 20947 12189 20956 12223
rect 20904 12180 20956 12189
rect 23848 12223 23900 12232
rect 23848 12189 23857 12223
rect 23857 12189 23891 12223
rect 23891 12189 23900 12223
rect 23848 12180 23900 12189
rect 13268 12155 13320 12164
rect 13268 12121 13277 12155
rect 13277 12121 13311 12155
rect 13311 12121 13320 12155
rect 13268 12112 13320 12121
rect 2412 12044 2464 12096
rect 3884 12087 3936 12096
rect 3884 12053 3893 12087
rect 3893 12053 3927 12087
rect 3927 12053 3936 12087
rect 3884 12044 3936 12053
rect 7012 12087 7064 12096
rect 7012 12053 7021 12087
rect 7021 12053 7055 12087
rect 7055 12053 7064 12087
rect 7012 12044 7064 12053
rect 7472 12087 7524 12096
rect 7472 12053 7481 12087
rect 7481 12053 7515 12087
rect 7515 12053 7524 12087
rect 7472 12044 7524 12053
rect 8300 12044 8352 12096
rect 9128 12087 9180 12096
rect 9128 12053 9137 12087
rect 9137 12053 9171 12087
rect 9171 12053 9180 12087
rect 9128 12044 9180 12053
rect 9680 12044 9732 12096
rect 10692 12087 10744 12096
rect 10692 12053 10701 12087
rect 10701 12053 10735 12087
rect 10735 12053 10744 12087
rect 10692 12044 10744 12053
rect 11704 12087 11756 12096
rect 11704 12053 11713 12087
rect 11713 12053 11747 12087
rect 11747 12053 11756 12087
rect 11704 12044 11756 12053
rect 15752 12087 15804 12096
rect 15752 12053 15761 12087
rect 15761 12053 15795 12087
rect 15795 12053 15804 12087
rect 15752 12044 15804 12053
rect 17960 12044 18012 12096
rect 20076 12044 20128 12096
rect 21824 12044 21876 12096
rect 25228 12087 25280 12096
rect 25228 12053 25237 12087
rect 25237 12053 25271 12087
rect 25271 12053 25280 12087
rect 25228 12044 25280 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 3056 11840 3108 11892
rect 3332 11883 3384 11892
rect 3332 11849 3341 11883
rect 3341 11849 3375 11883
rect 3375 11849 3384 11883
rect 3332 11840 3384 11849
rect 6092 11840 6144 11892
rect 6460 11840 6512 11892
rect 6828 11840 6880 11892
rect 7288 11840 7340 11892
rect 7656 11883 7708 11892
rect 7656 11849 7665 11883
rect 7665 11849 7699 11883
rect 7699 11849 7708 11883
rect 7656 11840 7708 11849
rect 11796 11883 11848 11892
rect 11796 11849 11805 11883
rect 11805 11849 11839 11883
rect 11839 11849 11848 11883
rect 11796 11840 11848 11849
rect 15660 11883 15712 11892
rect 15660 11849 15669 11883
rect 15669 11849 15703 11883
rect 15703 11849 15712 11883
rect 15660 11840 15712 11849
rect 16212 11883 16264 11892
rect 16212 11849 16221 11883
rect 16221 11849 16255 11883
rect 16255 11849 16264 11883
rect 16212 11840 16264 11849
rect 17592 11883 17644 11892
rect 17592 11849 17601 11883
rect 17601 11849 17635 11883
rect 17635 11849 17644 11883
rect 17592 11840 17644 11849
rect 18604 11840 18656 11892
rect 21180 11840 21232 11892
rect 23112 11883 23164 11892
rect 23112 11849 23121 11883
rect 23121 11849 23155 11883
rect 23155 11849 23164 11883
rect 23112 11840 23164 11849
rect 24860 11840 24912 11892
rect 1860 11772 1912 11824
rect 9220 11815 9272 11824
rect 9220 11781 9229 11815
rect 9229 11781 9263 11815
rect 9263 11781 9272 11815
rect 9220 11772 9272 11781
rect 10876 11815 10928 11824
rect 10876 11781 10885 11815
rect 10885 11781 10919 11815
rect 10919 11781 10928 11815
rect 10876 11772 10928 11781
rect 4068 11704 4120 11756
rect 5448 11747 5500 11756
rect 5448 11713 5457 11747
rect 5457 11713 5491 11747
rect 5491 11713 5500 11747
rect 5448 11704 5500 11713
rect 7932 11704 7984 11756
rect 8300 11704 8352 11756
rect 11152 11704 11204 11756
rect 13912 11772 13964 11824
rect 20812 11815 20864 11824
rect 20812 11781 20821 11815
rect 20821 11781 20855 11815
rect 20855 11781 20864 11815
rect 20812 11772 20864 11781
rect 21824 11772 21876 11824
rect 23848 11772 23900 11824
rect 13176 11747 13228 11756
rect 13176 11713 13185 11747
rect 13185 11713 13219 11747
rect 13219 11713 13228 11747
rect 13176 11704 13228 11713
rect 19432 11747 19484 11756
rect 19432 11713 19441 11747
rect 19441 11713 19475 11747
rect 19475 11713 19484 11747
rect 19432 11704 19484 11713
rect 21088 11704 21140 11756
rect 3884 11679 3936 11688
rect 3884 11645 3893 11679
rect 3893 11645 3927 11679
rect 3927 11645 3936 11679
rect 3884 11636 3936 11645
rect 4988 11636 5040 11688
rect 7472 11636 7524 11688
rect 8852 11636 8904 11688
rect 11704 11636 11756 11688
rect 14280 11679 14332 11688
rect 14280 11645 14289 11679
rect 14289 11645 14323 11679
rect 14323 11645 14332 11679
rect 14280 11636 14332 11645
rect 24216 11636 24268 11688
rect 25228 11636 25280 11688
rect 2136 11568 2188 11620
rect 2320 11611 2372 11620
rect 2320 11577 2329 11611
rect 2329 11577 2363 11611
rect 2363 11577 2372 11611
rect 2320 11568 2372 11577
rect 2872 11568 2924 11620
rect 2228 11543 2280 11552
rect 2228 11509 2237 11543
rect 2237 11509 2271 11543
rect 2271 11509 2280 11543
rect 2228 11500 2280 11509
rect 3332 11500 3384 11552
rect 7748 11568 7800 11620
rect 8024 11568 8076 11620
rect 5356 11543 5408 11552
rect 5356 11509 5365 11543
rect 5365 11509 5399 11543
rect 5399 11509 5408 11543
rect 5356 11500 5408 11509
rect 6644 11543 6696 11552
rect 6644 11509 6653 11543
rect 6653 11509 6687 11543
rect 6687 11509 6696 11543
rect 6644 11500 6696 11509
rect 7656 11500 7708 11552
rect 8116 11543 8168 11552
rect 8116 11509 8125 11543
rect 8125 11509 8159 11543
rect 8159 11509 8168 11543
rect 8116 11500 8168 11509
rect 9128 11568 9180 11620
rect 10324 11568 10376 11620
rect 9036 11543 9088 11552
rect 9036 11509 9045 11543
rect 9045 11509 9079 11543
rect 9079 11509 9088 11543
rect 9036 11500 9088 11509
rect 9680 11543 9732 11552
rect 9680 11509 9689 11543
rect 9689 11509 9723 11543
rect 9723 11509 9732 11543
rect 9680 11500 9732 11509
rect 9864 11500 9916 11552
rect 11244 11568 11296 11620
rect 11612 11568 11664 11620
rect 12072 11500 12124 11552
rect 14464 11568 14516 11620
rect 18788 11568 18840 11620
rect 21364 11611 21416 11620
rect 21364 11577 21373 11611
rect 21373 11577 21407 11611
rect 21407 11577 21416 11611
rect 21364 11568 21416 11577
rect 13268 11543 13320 11552
rect 13268 11509 13277 11543
rect 13277 11509 13311 11543
rect 13311 11509 13320 11543
rect 13268 11500 13320 11509
rect 16672 11500 16724 11552
rect 17224 11543 17276 11552
rect 17224 11509 17233 11543
rect 17233 11509 17267 11543
rect 17267 11509 17276 11543
rect 17224 11500 17276 11509
rect 18604 11543 18656 11552
rect 18604 11509 18613 11543
rect 18613 11509 18647 11543
rect 18647 11509 18656 11543
rect 18604 11500 18656 11509
rect 19524 11500 19576 11552
rect 21088 11500 21140 11552
rect 21824 11543 21876 11552
rect 21824 11509 21833 11543
rect 21833 11509 21867 11543
rect 21867 11509 21876 11543
rect 21824 11500 21876 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 2320 11296 2372 11348
rect 2964 11296 3016 11348
rect 4344 11296 4396 11348
rect 5448 11339 5500 11348
rect 4436 11271 4488 11280
rect 4436 11237 4445 11271
rect 4445 11237 4479 11271
rect 4479 11237 4488 11271
rect 4436 11228 4488 11237
rect 4528 11228 4580 11280
rect 5448 11305 5457 11339
rect 5457 11305 5491 11339
rect 5491 11305 5500 11339
rect 5448 11296 5500 11305
rect 6460 11339 6512 11348
rect 6460 11305 6469 11339
rect 6469 11305 6503 11339
rect 6503 11305 6512 11339
rect 6460 11296 6512 11305
rect 8392 11296 8444 11348
rect 8944 11339 8996 11348
rect 8944 11305 8953 11339
rect 8953 11305 8987 11339
rect 8987 11305 8996 11339
rect 8944 11296 8996 11305
rect 4988 11228 5040 11280
rect 8208 11228 8260 11280
rect 10784 11296 10836 11348
rect 10876 11296 10928 11348
rect 11336 11296 11388 11348
rect 11796 11296 11848 11348
rect 12164 11296 12216 11348
rect 14464 11296 14516 11348
rect 16120 11296 16172 11348
rect 18788 11339 18840 11348
rect 18788 11305 18797 11339
rect 18797 11305 18831 11339
rect 18831 11305 18840 11339
rect 18788 11296 18840 11305
rect 21088 11339 21140 11348
rect 21088 11305 21097 11339
rect 21097 11305 21131 11339
rect 21131 11305 21140 11339
rect 21088 11296 21140 11305
rect 22100 11296 22152 11348
rect 23756 11339 23808 11348
rect 23756 11305 23765 11339
rect 23765 11305 23799 11339
rect 23799 11305 23808 11339
rect 23756 11296 23808 11305
rect 24216 11339 24268 11348
rect 24216 11305 24225 11339
rect 24225 11305 24259 11339
rect 24259 11305 24268 11339
rect 24216 11296 24268 11305
rect 25136 11296 25188 11348
rect 10232 11271 10284 11280
rect 10232 11237 10241 11271
rect 10241 11237 10275 11271
rect 10275 11237 10284 11271
rect 10232 11228 10284 11237
rect 12348 11228 12400 11280
rect 19340 11228 19392 11280
rect 24676 11271 24728 11280
rect 24676 11237 24685 11271
rect 24685 11237 24719 11271
rect 24719 11237 24728 11271
rect 24676 11228 24728 11237
rect 24860 11271 24912 11280
rect 24860 11237 24869 11271
rect 24869 11237 24903 11271
rect 24903 11237 24912 11271
rect 24860 11228 24912 11237
rect 24952 11271 25004 11280
rect 24952 11237 24961 11271
rect 24961 11237 24995 11271
rect 24995 11237 25004 11271
rect 24952 11228 25004 11237
rect 1400 11203 1452 11212
rect 1400 11169 1409 11203
rect 1409 11169 1443 11203
rect 1443 11169 1452 11203
rect 1400 11160 1452 11169
rect 2780 11160 2832 11212
rect 6276 11203 6328 11212
rect 6276 11169 6285 11203
rect 6285 11169 6319 11203
rect 6319 11169 6328 11203
rect 6276 11160 6328 11169
rect 6644 11160 6696 11212
rect 9036 11160 9088 11212
rect 16304 11160 16356 11212
rect 16948 11203 17000 11212
rect 16948 11169 16982 11203
rect 16982 11169 17000 11203
rect 16948 11160 17000 11169
rect 19524 11160 19576 11212
rect 21364 11160 21416 11212
rect 22100 11203 22152 11212
rect 22100 11169 22134 11203
rect 22134 11169 22152 11203
rect 22100 11160 22152 11169
rect 23388 11160 23440 11212
rect 24216 11160 24268 11212
rect 2872 11092 2924 11144
rect 4160 11092 4212 11144
rect 6552 11135 6604 11144
rect 6552 11101 6561 11135
rect 6561 11101 6595 11135
rect 6595 11101 6604 11135
rect 6552 11092 6604 11101
rect 7656 11135 7708 11144
rect 7656 11101 7665 11135
rect 7665 11101 7699 11135
rect 7699 11101 7708 11135
rect 7656 11092 7708 11101
rect 10324 11135 10376 11144
rect 10324 11101 10333 11135
rect 10333 11101 10367 11135
rect 10367 11101 10376 11135
rect 10324 11092 10376 11101
rect 11704 11135 11756 11144
rect 11704 11101 11713 11135
rect 11713 11101 11747 11135
rect 11747 11101 11756 11135
rect 11704 11092 11756 11101
rect 16672 11135 16724 11144
rect 16672 11101 16681 11135
rect 16681 11101 16715 11135
rect 16715 11101 16724 11135
rect 16672 11092 16724 11101
rect 19432 11092 19484 11144
rect 21824 11135 21876 11144
rect 21824 11101 21833 11135
rect 21833 11101 21867 11135
rect 21867 11101 21876 11135
rect 21824 11092 21876 11101
rect 24124 11092 24176 11144
rect 2320 11024 2372 11076
rect 4068 11024 4120 11076
rect 5540 11024 5592 11076
rect 7012 11024 7064 11076
rect 10048 11024 10100 11076
rect 11152 11024 11204 11076
rect 18880 11024 18932 11076
rect 5172 10999 5224 11008
rect 5172 10965 5181 10999
rect 5181 10965 5215 10999
rect 5215 10965 5224 10999
rect 5172 10956 5224 10965
rect 7196 10956 7248 11008
rect 8576 10956 8628 11008
rect 13084 10999 13136 11008
rect 13084 10965 13093 10999
rect 13093 10965 13127 10999
rect 13127 10965 13136 10999
rect 13084 10956 13136 10965
rect 19524 10956 19576 11008
rect 21456 10999 21508 11008
rect 21456 10965 21465 10999
rect 21465 10965 21499 10999
rect 21499 10965 21508 10999
rect 21456 10956 21508 10965
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 3792 10795 3844 10804
rect 3792 10761 3801 10795
rect 3801 10761 3835 10795
rect 3835 10761 3844 10795
rect 3792 10752 3844 10761
rect 4436 10752 4488 10804
rect 6552 10752 6604 10804
rect 6828 10752 6880 10804
rect 7012 10795 7064 10804
rect 7012 10761 7021 10795
rect 7021 10761 7055 10795
rect 7055 10761 7064 10795
rect 7012 10752 7064 10761
rect 8392 10752 8444 10804
rect 8944 10752 8996 10804
rect 10784 10752 10836 10804
rect 11060 10752 11112 10804
rect 14280 10752 14332 10804
rect 16672 10795 16724 10804
rect 2688 10727 2740 10736
rect 2688 10693 2697 10727
rect 2697 10693 2731 10727
rect 2731 10693 2740 10727
rect 2688 10684 2740 10693
rect 2780 10684 2832 10736
rect 3976 10684 4028 10736
rect 4620 10684 4672 10736
rect 8208 10684 8260 10736
rect 8484 10684 8536 10736
rect 10876 10727 10928 10736
rect 10876 10693 10885 10727
rect 10885 10693 10919 10727
rect 10919 10693 10928 10727
rect 10876 10684 10928 10693
rect 12532 10727 12584 10736
rect 12532 10693 12541 10727
rect 12541 10693 12575 10727
rect 12575 10693 12584 10727
rect 12532 10684 12584 10693
rect 5172 10616 5224 10668
rect 7104 10616 7156 10668
rect 7564 10616 7616 10668
rect 9956 10616 10008 10668
rect 1952 10548 2004 10600
rect 2872 10548 2924 10600
rect 3608 10591 3660 10600
rect 3608 10557 3617 10591
rect 3617 10557 3651 10591
rect 3651 10557 3660 10591
rect 3608 10548 3660 10557
rect 4160 10548 4212 10600
rect 5448 10548 5500 10600
rect 13176 10616 13228 10668
rect 16672 10761 16681 10795
rect 16681 10761 16715 10795
rect 16715 10761 16724 10795
rect 16672 10752 16724 10761
rect 19616 10795 19668 10804
rect 19616 10761 19625 10795
rect 19625 10761 19659 10795
rect 19659 10761 19668 10795
rect 19616 10752 19668 10761
rect 20812 10795 20864 10804
rect 20812 10761 20821 10795
rect 20821 10761 20855 10795
rect 20855 10761 20864 10795
rect 20812 10752 20864 10761
rect 18052 10684 18104 10736
rect 20628 10684 20680 10736
rect 20720 10684 20772 10736
rect 21824 10752 21876 10804
rect 21916 10684 21968 10736
rect 22008 10659 22060 10668
rect 22008 10625 22017 10659
rect 22017 10625 22051 10659
rect 22051 10625 22060 10659
rect 22008 10616 22060 10625
rect 25504 10752 25556 10804
rect 24952 10684 25004 10736
rect 11888 10591 11940 10600
rect 7472 10523 7524 10532
rect 7472 10489 7481 10523
rect 7481 10489 7515 10523
rect 7515 10489 7524 10523
rect 7472 10480 7524 10489
rect 8392 10480 8444 10532
rect 10048 10480 10100 10532
rect 10324 10480 10376 10532
rect 11336 10523 11388 10532
rect 11336 10489 11345 10523
rect 11345 10489 11379 10523
rect 11379 10489 11388 10523
rect 11336 10480 11388 10489
rect 11888 10557 11897 10591
rect 11897 10557 11931 10591
rect 11931 10557 11940 10591
rect 11888 10548 11940 10557
rect 13728 10548 13780 10600
rect 17684 10548 17736 10600
rect 1768 10412 1820 10464
rect 2044 10455 2096 10464
rect 2044 10421 2053 10455
rect 2053 10421 2087 10455
rect 2087 10421 2096 10455
rect 2044 10412 2096 10421
rect 2228 10412 2280 10464
rect 3516 10412 3568 10464
rect 4528 10412 4580 10464
rect 5448 10412 5500 10464
rect 9956 10412 10008 10464
rect 10784 10412 10836 10464
rect 12716 10480 12768 10532
rect 13084 10523 13136 10532
rect 13084 10489 13093 10523
rect 13093 10489 13127 10523
rect 13127 10489 13136 10523
rect 13084 10480 13136 10489
rect 14648 10480 14700 10532
rect 16948 10480 17000 10532
rect 17868 10480 17920 10532
rect 20076 10548 20128 10600
rect 23756 10548 23808 10600
rect 13452 10455 13504 10464
rect 13452 10421 13461 10455
rect 13461 10421 13495 10455
rect 13495 10421 13504 10455
rect 13452 10412 13504 10421
rect 14464 10412 14516 10464
rect 15568 10412 15620 10464
rect 17776 10455 17828 10464
rect 17776 10421 17785 10455
rect 17785 10421 17819 10455
rect 17819 10421 17828 10455
rect 19524 10480 19576 10532
rect 19616 10480 19668 10532
rect 19984 10480 20036 10532
rect 20444 10523 20496 10532
rect 20444 10489 20453 10523
rect 20453 10489 20487 10523
rect 20487 10489 20496 10523
rect 20444 10480 20496 10489
rect 20904 10480 20956 10532
rect 21456 10480 21508 10532
rect 18604 10455 18656 10464
rect 17776 10412 17828 10421
rect 18604 10421 18613 10455
rect 18613 10421 18647 10455
rect 18647 10421 18656 10455
rect 18604 10412 18656 10421
rect 20260 10412 20312 10464
rect 20812 10412 20864 10464
rect 22100 10412 22152 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1400 10208 1452 10260
rect 2596 10208 2648 10260
rect 3332 10251 3384 10260
rect 3332 10217 3341 10251
rect 3341 10217 3375 10251
rect 3375 10217 3384 10251
rect 3332 10208 3384 10217
rect 3608 10251 3660 10260
rect 3608 10217 3617 10251
rect 3617 10217 3651 10251
rect 3651 10217 3660 10251
rect 3608 10208 3660 10217
rect 4344 10251 4396 10260
rect 4344 10217 4353 10251
rect 4353 10217 4387 10251
rect 4387 10217 4396 10251
rect 4344 10208 4396 10217
rect 6184 10251 6236 10260
rect 6184 10217 6193 10251
rect 6193 10217 6227 10251
rect 6227 10217 6236 10251
rect 6184 10208 6236 10217
rect 7564 10208 7616 10260
rect 8852 10251 8904 10260
rect 8852 10217 8861 10251
rect 8861 10217 8895 10251
rect 8895 10217 8904 10251
rect 8852 10208 8904 10217
rect 10140 10208 10192 10260
rect 12440 10251 12492 10260
rect 12440 10217 12449 10251
rect 12449 10217 12483 10251
rect 12483 10217 12492 10251
rect 13084 10251 13136 10260
rect 12440 10208 12492 10217
rect 13084 10217 13093 10251
rect 13093 10217 13127 10251
rect 13127 10217 13136 10251
rect 13084 10208 13136 10217
rect 14648 10251 14700 10260
rect 14648 10217 14657 10251
rect 14657 10217 14691 10251
rect 14691 10217 14700 10251
rect 14648 10208 14700 10217
rect 15844 10251 15896 10260
rect 15844 10217 15853 10251
rect 15853 10217 15887 10251
rect 15887 10217 15896 10251
rect 15844 10208 15896 10217
rect 18604 10208 18656 10260
rect 18788 10208 18840 10260
rect 19524 10251 19576 10260
rect 19524 10217 19533 10251
rect 19533 10217 19567 10251
rect 19567 10217 19576 10251
rect 19524 10208 19576 10217
rect 23296 10251 23348 10260
rect 23296 10217 23305 10251
rect 23305 10217 23339 10251
rect 23339 10217 23348 10251
rect 23296 10208 23348 10217
rect 23572 10208 23624 10260
rect 23848 10208 23900 10260
rect 24676 10208 24728 10260
rect 25136 10251 25188 10260
rect 25136 10217 25145 10251
rect 25145 10217 25179 10251
rect 25179 10217 25188 10251
rect 25136 10208 25188 10217
rect 5172 10140 5224 10192
rect 8208 10140 8260 10192
rect 8392 10183 8444 10192
rect 8392 10149 8401 10183
rect 8401 10149 8435 10183
rect 8435 10149 8444 10183
rect 8392 10140 8444 10149
rect 12532 10140 12584 10192
rect 12716 10140 12768 10192
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 2688 10072 2740 10124
rect 7656 10072 7708 10124
rect 8668 10072 8720 10124
rect 9956 10072 10008 10124
rect 10692 10072 10744 10124
rect 11336 10115 11388 10124
rect 11336 10081 11345 10115
rect 11345 10081 11379 10115
rect 11379 10081 11388 10115
rect 11336 10072 11388 10081
rect 11888 10072 11940 10124
rect 14464 10140 14516 10192
rect 15660 10183 15712 10192
rect 15660 10149 15669 10183
rect 15669 10149 15703 10183
rect 15703 10149 15712 10183
rect 15660 10140 15712 10149
rect 15292 10072 15344 10124
rect 16948 10140 17000 10192
rect 17684 10140 17736 10192
rect 23020 10140 23072 10192
rect 21732 10072 21784 10124
rect 23664 10072 23716 10124
rect 24124 10072 24176 10124
rect 24952 10115 25004 10124
rect 24952 10081 24961 10115
rect 24961 10081 24995 10115
rect 24995 10081 25004 10115
rect 24952 10072 25004 10081
rect 4804 10047 4856 10056
rect 4804 10013 4813 10047
rect 4813 10013 4847 10047
rect 4847 10013 4856 10047
rect 4804 10004 4856 10013
rect 10784 10004 10836 10056
rect 11612 10047 11664 10056
rect 11612 10013 11621 10047
rect 11621 10013 11655 10047
rect 11655 10013 11664 10047
rect 11612 10004 11664 10013
rect 13084 10004 13136 10056
rect 13452 10004 13504 10056
rect 17500 10047 17552 10056
rect 17500 10013 17509 10047
rect 17509 10013 17543 10047
rect 17543 10013 17552 10047
rect 17500 10004 17552 10013
rect 20720 10004 20772 10056
rect 2688 9979 2740 9988
rect 2688 9945 2697 9979
rect 2697 9945 2731 9979
rect 2731 9945 2740 9979
rect 2688 9936 2740 9945
rect 10968 9936 11020 9988
rect 11704 9936 11756 9988
rect 23480 9979 23532 9988
rect 23480 9945 23489 9979
rect 23489 9945 23523 9979
rect 23523 9945 23532 9979
rect 23480 9936 23532 9945
rect 23848 9936 23900 9988
rect 24032 9936 24084 9988
rect 1676 9868 1728 9920
rect 5448 9868 5500 9920
rect 7840 9911 7892 9920
rect 7840 9877 7849 9911
rect 7849 9877 7883 9911
rect 7883 9877 7892 9911
rect 7840 9868 7892 9877
rect 10048 9868 10100 9920
rect 10784 9911 10836 9920
rect 10784 9877 10793 9911
rect 10793 9877 10827 9911
rect 10827 9877 10836 9911
rect 10784 9868 10836 9877
rect 11060 9911 11112 9920
rect 11060 9877 11069 9911
rect 11069 9877 11103 9911
rect 11103 9877 11112 9911
rect 11060 9868 11112 9877
rect 11336 9868 11388 9920
rect 15384 9911 15436 9920
rect 15384 9877 15393 9911
rect 15393 9877 15427 9911
rect 15427 9877 15436 9911
rect 15384 9868 15436 9877
rect 19892 9911 19944 9920
rect 19892 9877 19901 9911
rect 19901 9877 19935 9911
rect 19935 9877 19944 9911
rect 19892 9868 19944 9877
rect 22100 9868 22152 9920
rect 22928 9911 22980 9920
rect 22928 9877 22937 9911
rect 22937 9877 22971 9911
rect 22971 9877 22980 9911
rect 22928 9868 22980 9877
rect 24860 9911 24912 9920
rect 24860 9877 24869 9911
rect 24869 9877 24903 9911
rect 24903 9877 24912 9911
rect 24860 9868 24912 9877
rect 25228 9868 25280 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 5172 9664 5224 9716
rect 2504 9596 2556 9648
rect 4068 9596 4120 9648
rect 2872 9528 2924 9580
rect 6828 9664 6880 9716
rect 7656 9707 7708 9716
rect 7656 9673 7665 9707
rect 7665 9673 7699 9707
rect 7699 9673 7708 9707
rect 7656 9664 7708 9673
rect 11888 9707 11940 9716
rect 11888 9673 11897 9707
rect 11897 9673 11931 9707
rect 11931 9673 11940 9707
rect 11888 9664 11940 9673
rect 9956 9596 10008 9648
rect 13820 9639 13872 9648
rect 13820 9605 13829 9639
rect 13829 9605 13863 9639
rect 13863 9605 13872 9639
rect 13820 9596 13872 9605
rect 14004 9596 14056 9648
rect 4252 9503 4304 9512
rect 4252 9469 4261 9503
rect 4261 9469 4295 9503
rect 4295 9469 4304 9503
rect 4252 9460 4304 9469
rect 4344 9460 4396 9512
rect 10968 9528 11020 9580
rect 11152 9528 11204 9580
rect 6092 9460 6144 9512
rect 7932 9460 7984 9512
rect 8392 9460 8444 9512
rect 2872 9392 2924 9444
rect 8208 9392 8260 9444
rect 9496 9392 9548 9444
rect 11060 9460 11112 9512
rect 12164 9503 12216 9512
rect 12164 9469 12173 9503
rect 12173 9469 12207 9503
rect 12207 9469 12216 9503
rect 12164 9460 12216 9469
rect 15292 9664 15344 9716
rect 15660 9664 15712 9716
rect 16672 9664 16724 9716
rect 17500 9707 17552 9716
rect 17500 9673 17509 9707
rect 17509 9673 17543 9707
rect 17543 9673 17552 9707
rect 17500 9664 17552 9673
rect 20720 9707 20772 9716
rect 20720 9673 20729 9707
rect 20729 9673 20763 9707
rect 20763 9673 20772 9707
rect 20720 9664 20772 9673
rect 20904 9707 20956 9716
rect 20904 9673 20913 9707
rect 20913 9673 20947 9707
rect 20947 9673 20956 9707
rect 20904 9664 20956 9673
rect 23296 9664 23348 9716
rect 15752 9596 15804 9648
rect 18144 9639 18196 9648
rect 18144 9605 18153 9639
rect 18153 9605 18187 9639
rect 18187 9605 18196 9639
rect 18144 9596 18196 9605
rect 19156 9639 19208 9648
rect 19156 9605 19165 9639
rect 19165 9605 19199 9639
rect 19199 9605 19208 9639
rect 19156 9596 19208 9605
rect 19432 9596 19484 9648
rect 20444 9596 20496 9648
rect 21732 9596 21784 9648
rect 23020 9639 23072 9648
rect 23020 9605 23029 9639
rect 23029 9605 23063 9639
rect 23063 9605 23072 9639
rect 23020 9596 23072 9605
rect 23572 9664 23624 9716
rect 24952 9707 25004 9716
rect 24952 9673 24961 9707
rect 24961 9673 24995 9707
rect 24995 9673 25004 9707
rect 24952 9664 25004 9673
rect 23756 9639 23808 9648
rect 15568 9571 15620 9580
rect 10876 9435 10928 9444
rect 10876 9401 10885 9435
rect 10885 9401 10919 9435
rect 10919 9401 10928 9435
rect 10876 9392 10928 9401
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 2780 9324 2832 9376
rect 3240 9324 3292 9376
rect 6276 9367 6328 9376
rect 6276 9333 6285 9367
rect 6285 9333 6319 9367
rect 6319 9333 6328 9367
rect 6276 9324 6328 9333
rect 7196 9324 7248 9376
rect 9220 9367 9272 9376
rect 9220 9333 9229 9367
rect 9229 9333 9263 9367
rect 9263 9333 9272 9367
rect 9220 9324 9272 9333
rect 10140 9367 10192 9376
rect 10140 9333 10149 9367
rect 10149 9333 10183 9367
rect 10183 9333 10192 9367
rect 11704 9392 11756 9444
rect 12348 9392 12400 9444
rect 15568 9537 15577 9571
rect 15577 9537 15611 9571
rect 15611 9537 15620 9571
rect 15568 9528 15620 9537
rect 17776 9528 17828 9580
rect 18788 9528 18840 9580
rect 22008 9528 22060 9580
rect 22376 9571 22428 9580
rect 22376 9537 22385 9571
rect 22385 9537 22419 9571
rect 22419 9537 22428 9571
rect 22376 9528 22428 9537
rect 23756 9605 23765 9639
rect 23765 9605 23799 9639
rect 23799 9605 23808 9639
rect 23756 9596 23808 9605
rect 25504 9596 25556 9648
rect 13084 9392 13136 9444
rect 15476 9435 15528 9444
rect 15476 9401 15485 9435
rect 15485 9401 15519 9435
rect 15519 9401 15528 9435
rect 15476 9392 15528 9401
rect 17224 9392 17276 9444
rect 18052 9392 18104 9444
rect 10140 9324 10192 9333
rect 11980 9324 12032 9376
rect 20720 9460 20772 9512
rect 25044 9460 25096 9512
rect 22928 9392 22980 9444
rect 18880 9324 18932 9376
rect 21088 9324 21140 9376
rect 23112 9324 23164 9376
rect 24768 9392 24820 9444
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 1400 9120 1452 9172
rect 4344 9163 4396 9172
rect 4344 9129 4353 9163
rect 4353 9129 4387 9163
rect 4387 9129 4396 9163
rect 4344 9120 4396 9129
rect 5172 9163 5224 9172
rect 5172 9129 5181 9163
rect 5181 9129 5215 9163
rect 5215 9129 5224 9163
rect 5172 9120 5224 9129
rect 6920 9120 6972 9172
rect 7932 9120 7984 9172
rect 9496 9163 9548 9172
rect 9496 9129 9505 9163
rect 9505 9129 9539 9163
rect 9539 9129 9548 9163
rect 9496 9120 9548 9129
rect 10876 9120 10928 9172
rect 11980 9163 12032 9172
rect 11980 9129 11989 9163
rect 11989 9129 12023 9163
rect 12023 9129 12032 9163
rect 11980 9120 12032 9129
rect 13636 9163 13688 9172
rect 13636 9129 13645 9163
rect 13645 9129 13679 9163
rect 13679 9129 13688 9163
rect 13636 9120 13688 9129
rect 14188 9163 14240 9172
rect 14188 9129 14197 9163
rect 14197 9129 14231 9163
rect 14231 9129 14240 9163
rect 14188 9120 14240 9129
rect 15476 9120 15528 9172
rect 15844 9120 15896 9172
rect 17224 9163 17276 9172
rect 17224 9129 17233 9163
rect 17233 9129 17267 9163
rect 17267 9129 17276 9163
rect 17224 9120 17276 9129
rect 17684 9120 17736 9172
rect 18696 9120 18748 9172
rect 23112 9163 23164 9172
rect 23112 9129 23121 9163
rect 23121 9129 23155 9163
rect 23155 9129 23164 9163
rect 23112 9120 23164 9129
rect 24124 9120 24176 9172
rect 24952 9163 25004 9172
rect 24952 9129 24961 9163
rect 24961 9129 24995 9163
rect 24995 9129 25004 9163
rect 24952 9120 25004 9129
rect 4252 9052 4304 9104
rect 4804 9095 4856 9104
rect 4804 9061 4813 9095
rect 4813 9061 4847 9095
rect 4847 9061 4856 9095
rect 4804 9052 4856 9061
rect 10048 9052 10100 9104
rect 10692 9052 10744 9104
rect 13544 9052 13596 9104
rect 18788 9095 18840 9104
rect 18788 9061 18797 9095
rect 18797 9061 18831 9095
rect 18831 9061 18840 9095
rect 18788 9052 18840 9061
rect 21548 9095 21600 9104
rect 21548 9061 21557 9095
rect 21557 9061 21591 9095
rect 21591 9061 21600 9095
rect 21548 9052 21600 9061
rect 23572 9095 23624 9104
rect 23572 9061 23581 9095
rect 23581 9061 23615 9095
rect 23615 9061 23624 9095
rect 23572 9052 23624 9061
rect 2044 8984 2096 9036
rect 6184 8984 6236 9036
rect 10876 9027 10928 9036
rect 10876 8993 10910 9027
rect 10910 8993 10928 9027
rect 10876 8984 10928 8993
rect 12348 8984 12400 9036
rect 17960 8984 18012 9036
rect 21364 9027 21416 9036
rect 21364 8993 21373 9027
rect 21373 8993 21407 9027
rect 21407 8993 21416 9027
rect 21364 8984 21416 8993
rect 23020 8984 23072 9036
rect 24676 9052 24728 9104
rect 24768 9027 24820 9036
rect 24768 8993 24777 9027
rect 24777 8993 24811 9027
rect 24811 8993 24820 9027
rect 24768 8984 24820 8993
rect 6092 8916 6144 8968
rect 1492 8780 1544 8832
rect 9312 8780 9364 8832
rect 13176 8891 13228 8900
rect 13176 8857 13185 8891
rect 13185 8857 13219 8891
rect 13219 8857 13228 8891
rect 13176 8848 13228 8857
rect 11704 8780 11756 8832
rect 13084 8780 13136 8832
rect 17316 8916 17368 8968
rect 18880 8959 18932 8968
rect 18604 8848 18656 8900
rect 18880 8925 18889 8959
rect 18889 8925 18923 8959
rect 18923 8925 18932 8959
rect 18880 8916 18932 8925
rect 21732 8916 21784 8968
rect 23848 8959 23900 8968
rect 23848 8925 23857 8959
rect 23857 8925 23891 8959
rect 23891 8925 23900 8959
rect 23848 8916 23900 8925
rect 19156 8848 19208 8900
rect 21088 8891 21140 8900
rect 21088 8857 21097 8891
rect 21097 8857 21131 8891
rect 21131 8857 21140 8891
rect 21088 8848 21140 8857
rect 22928 8848 22980 8900
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 2044 8619 2096 8628
rect 2044 8585 2053 8619
rect 2053 8585 2087 8619
rect 2087 8585 2096 8619
rect 2044 8576 2096 8585
rect 6184 8576 6236 8628
rect 6276 8576 6328 8628
rect 7932 8576 7984 8628
rect 9312 8576 9364 8628
rect 10048 8576 10100 8628
rect 11796 8619 11848 8628
rect 11796 8585 11805 8619
rect 11805 8585 11839 8619
rect 11839 8585 11848 8619
rect 11796 8576 11848 8585
rect 13636 8576 13688 8628
rect 18788 8576 18840 8628
rect 21548 8576 21600 8628
rect 21732 8619 21784 8628
rect 21732 8585 21741 8619
rect 21741 8585 21775 8619
rect 21775 8585 21784 8619
rect 21732 8576 21784 8585
rect 22468 8576 22520 8628
rect 23848 8576 23900 8628
rect 24860 8619 24912 8628
rect 24860 8585 24869 8619
rect 24869 8585 24903 8619
rect 24903 8585 24912 8619
rect 24860 8576 24912 8585
rect 25136 8619 25188 8628
rect 25136 8585 25145 8619
rect 25145 8585 25179 8619
rect 25179 8585 25188 8619
rect 25136 8576 25188 8585
rect 9220 8440 9272 8492
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 6092 8372 6144 8424
rect 7196 8415 7248 8424
rect 7196 8381 7205 8415
rect 7205 8381 7239 8415
rect 7239 8381 7248 8415
rect 7196 8372 7248 8381
rect 11704 8508 11756 8560
rect 12440 8508 12492 8560
rect 13452 8440 13504 8492
rect 12256 8415 12308 8424
rect 12256 8381 12265 8415
rect 12265 8381 12299 8415
rect 12299 8381 12308 8415
rect 12256 8372 12308 8381
rect 23020 8508 23072 8560
rect 14464 8440 14516 8492
rect 21364 8440 21416 8492
rect 7656 8304 7708 8356
rect 8392 8304 8444 8356
rect 9496 8304 9548 8356
rect 10140 8304 10192 8356
rect 12716 8304 12768 8356
rect 14188 8372 14240 8424
rect 18144 8372 18196 8424
rect 23664 8415 23716 8424
rect 23664 8381 23673 8415
rect 23673 8381 23707 8415
rect 23707 8381 23716 8415
rect 23664 8372 23716 8381
rect 24952 8415 25004 8424
rect 24952 8381 24961 8415
rect 24961 8381 24995 8415
rect 24995 8381 25004 8415
rect 24952 8372 25004 8381
rect 14096 8304 14148 8356
rect 14556 8347 14608 8356
rect 14556 8313 14565 8347
rect 14565 8313 14599 8347
rect 14599 8313 14608 8347
rect 14556 8304 14608 8313
rect 18512 8347 18564 8356
rect 18512 8313 18521 8347
rect 18521 8313 18555 8347
rect 18555 8313 18564 8347
rect 18512 8304 18564 8313
rect 19156 8304 19208 8356
rect 23940 8347 23992 8356
rect 23940 8313 23949 8347
rect 23949 8313 23983 8347
rect 23983 8313 23992 8347
rect 23940 8304 23992 8313
rect 7380 8279 7432 8288
rect 7380 8245 7389 8279
rect 7389 8245 7423 8279
rect 7423 8245 7432 8279
rect 7380 8236 7432 8245
rect 7840 8236 7892 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1584 8075 1636 8084
rect 1584 8041 1593 8075
rect 1593 8041 1627 8075
rect 1627 8041 1636 8075
rect 1584 8032 1636 8041
rect 6736 8032 6788 8084
rect 7196 8032 7248 8084
rect 7380 8075 7432 8084
rect 7380 8041 7389 8075
rect 7389 8041 7423 8075
rect 7423 8041 7432 8075
rect 7380 8032 7432 8041
rect 9864 8032 9916 8084
rect 10876 8032 10928 8084
rect 13912 8032 13964 8084
rect 14464 8075 14516 8084
rect 14464 8041 14473 8075
rect 14473 8041 14507 8075
rect 14507 8041 14516 8075
rect 14464 8032 14516 8041
rect 18880 8032 18932 8084
rect 23388 8032 23440 8084
rect 24768 8075 24820 8084
rect 24768 8041 24777 8075
rect 24777 8041 24811 8075
rect 24811 8041 24820 8075
rect 24768 8032 24820 8041
rect 6828 7964 6880 8016
rect 7932 7964 7984 8016
rect 8484 7964 8536 8016
rect 9496 8007 9548 8016
rect 9496 7973 9505 8007
rect 9505 7973 9539 8007
rect 9539 7973 9548 8007
rect 9496 7964 9548 7973
rect 11612 7964 11664 8016
rect 2044 7896 2096 7948
rect 8300 7896 8352 7948
rect 9680 7896 9732 7948
rect 12256 7939 12308 7948
rect 12256 7905 12265 7939
rect 12265 7905 12299 7939
rect 12299 7905 12308 7939
rect 12256 7896 12308 7905
rect 16580 7896 16632 7948
rect 16948 7939 17000 7948
rect 16948 7905 16957 7939
rect 16957 7905 16991 7939
rect 16991 7905 17000 7939
rect 16948 7896 17000 7905
rect 23940 7896 23992 7948
rect 24032 7896 24084 7948
rect 6460 7871 6512 7880
rect 6460 7837 6469 7871
rect 6469 7837 6503 7871
rect 6503 7837 6512 7871
rect 6460 7828 6512 7837
rect 8668 7871 8720 7880
rect 8668 7837 8677 7871
rect 8677 7837 8711 7871
rect 8711 7837 8720 7871
rect 8668 7828 8720 7837
rect 10324 7871 10376 7880
rect 10324 7837 10333 7871
rect 10333 7837 10367 7871
rect 10367 7837 10376 7871
rect 10324 7828 10376 7837
rect 12072 7828 12124 7880
rect 12624 7828 12676 7880
rect 13544 7828 13596 7880
rect 14004 7871 14056 7880
rect 14004 7837 14013 7871
rect 14013 7837 14047 7871
rect 14047 7837 14056 7871
rect 14004 7828 14056 7837
rect 17224 7871 17276 7880
rect 5448 7760 5500 7812
rect 9772 7803 9824 7812
rect 9772 7769 9781 7803
rect 9781 7769 9815 7803
rect 9815 7769 9824 7803
rect 9772 7760 9824 7769
rect 13452 7760 13504 7812
rect 17224 7837 17233 7871
rect 17233 7837 17267 7871
rect 17267 7837 17276 7871
rect 17224 7828 17276 7837
rect 11980 7735 12032 7744
rect 11980 7701 11989 7735
rect 11989 7701 12023 7735
rect 12023 7701 12032 7735
rect 11980 7692 12032 7701
rect 23664 7735 23716 7744
rect 23664 7701 23673 7735
rect 23673 7701 23707 7735
rect 23707 7701 23716 7735
rect 23664 7692 23716 7701
rect 23848 7692 23900 7744
rect 24124 7692 24176 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 2044 7531 2096 7540
rect 2044 7497 2053 7531
rect 2053 7497 2087 7531
rect 2087 7497 2096 7531
rect 2044 7488 2096 7497
rect 6828 7488 6880 7540
rect 7932 7531 7984 7540
rect 7932 7497 7941 7531
rect 7941 7497 7975 7531
rect 7975 7497 7984 7531
rect 7932 7488 7984 7497
rect 8392 7488 8444 7540
rect 9680 7488 9732 7540
rect 10324 7488 10376 7540
rect 11612 7531 11664 7540
rect 11612 7497 11621 7531
rect 11621 7497 11655 7531
rect 11655 7497 11664 7531
rect 11612 7488 11664 7497
rect 12072 7488 12124 7540
rect 12716 7531 12768 7540
rect 12716 7497 12725 7531
rect 12725 7497 12759 7531
rect 12759 7497 12768 7531
rect 12716 7488 12768 7497
rect 13084 7531 13136 7540
rect 13084 7497 13093 7531
rect 13093 7497 13127 7531
rect 13127 7497 13136 7531
rect 13084 7488 13136 7497
rect 13452 7531 13504 7540
rect 13452 7497 13461 7531
rect 13461 7497 13495 7531
rect 13495 7497 13504 7531
rect 13452 7488 13504 7497
rect 13912 7531 13964 7540
rect 13912 7497 13921 7531
rect 13921 7497 13955 7531
rect 13955 7497 13964 7531
rect 13912 7488 13964 7497
rect 14004 7488 14056 7540
rect 16948 7531 17000 7540
rect 16948 7497 16957 7531
rect 16957 7497 16991 7531
rect 16991 7497 17000 7531
rect 16948 7488 17000 7497
rect 23940 7531 23992 7540
rect 23940 7497 23949 7531
rect 23949 7497 23983 7531
rect 23983 7497 23992 7531
rect 23940 7488 23992 7497
rect 24032 7488 24084 7540
rect 24676 7488 24728 7540
rect 1584 7463 1636 7472
rect 1584 7429 1593 7463
rect 1593 7429 1627 7463
rect 1627 7429 1636 7463
rect 1584 7420 1636 7429
rect 6460 7420 6512 7472
rect 6736 7352 6788 7404
rect 8484 7352 8536 7404
rect 9588 7352 9640 7404
rect 9680 7352 9732 7404
rect 1400 7327 1452 7336
rect 1400 7293 1409 7327
rect 1409 7293 1443 7327
rect 1443 7293 1452 7327
rect 1400 7284 1452 7293
rect 8668 7284 8720 7336
rect 9956 7327 10008 7336
rect 9956 7293 9965 7327
rect 9965 7293 9999 7327
rect 9999 7293 10008 7327
rect 9956 7284 10008 7293
rect 17224 7284 17276 7336
rect 23848 7284 23900 7336
rect 8392 7216 8444 7268
rect 18236 7191 18288 7200
rect 18236 7157 18245 7191
rect 18245 7157 18279 7191
rect 18279 7157 18288 7191
rect 18236 7148 18288 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 1400 6944 1452 6996
rect 8484 6987 8536 6996
rect 8484 6953 8493 6987
rect 8493 6953 8527 6987
rect 8527 6953 8536 6987
rect 8484 6944 8536 6953
rect 8668 6944 8720 6996
rect 9864 6987 9916 6996
rect 9864 6953 9873 6987
rect 9873 6953 9907 6987
rect 9907 6953 9916 6987
rect 9864 6944 9916 6953
rect 9956 6944 10008 6996
rect 12256 6944 12308 6996
rect 24768 6987 24820 6996
rect 24768 6953 24777 6987
rect 24777 6953 24811 6987
rect 24811 6953 24820 6987
rect 24768 6944 24820 6953
rect 4896 6876 4948 6928
rect 8300 6808 8352 6860
rect 24584 6851 24636 6860
rect 24584 6817 24593 6851
rect 24593 6817 24627 6851
rect 24627 6817 24636 6851
rect 24584 6808 24636 6817
rect 4804 6783 4856 6792
rect 4804 6749 4813 6783
rect 4813 6749 4847 6783
rect 4847 6749 4856 6783
rect 4804 6740 4856 6749
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 4804 6400 4856 6452
rect 4988 6443 5040 6452
rect 4988 6409 4997 6443
rect 4997 6409 5031 6443
rect 5031 6409 5040 6443
rect 4988 6400 5040 6409
rect 9588 6400 9640 6452
rect 24768 6443 24820 6452
rect 24768 6409 24777 6443
rect 24777 6409 24811 6443
rect 24811 6409 24820 6443
rect 24768 6400 24820 6409
rect 24676 6332 24728 6384
rect 24216 6196 24268 6248
rect 4252 6103 4304 6112
rect 4252 6069 4261 6103
rect 4261 6069 4295 6103
rect 4295 6069 4304 6103
rect 4252 6060 4304 6069
rect 8852 6103 8904 6112
rect 8852 6069 8861 6103
rect 8861 6069 8895 6103
rect 8895 6069 8904 6103
rect 8852 6060 8904 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 24768 5899 24820 5908
rect 24768 5865 24777 5899
rect 24777 5865 24811 5899
rect 24811 5865 24820 5899
rect 24768 5856 24820 5865
rect 20720 5720 20772 5772
rect 24584 5763 24636 5772
rect 24584 5729 24593 5763
rect 24593 5729 24627 5763
rect 24627 5729 24636 5763
rect 24584 5720 24636 5729
rect 21088 5695 21140 5704
rect 21088 5661 21097 5695
rect 21097 5661 21131 5695
rect 21131 5661 21140 5695
rect 21088 5652 21140 5661
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 20720 5312 20772 5364
rect 24768 5355 24820 5364
rect 24768 5321 24777 5355
rect 24777 5321 24811 5355
rect 24811 5321 24820 5355
rect 24768 5312 24820 5321
rect 24676 5244 24728 5296
rect 24584 5151 24636 5160
rect 24584 5117 24593 5151
rect 24593 5117 24627 5151
rect 24627 5117 24636 5151
rect 24584 5108 24636 5117
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 21272 4811 21324 4820
rect 21272 4777 21281 4811
rect 21281 4777 21315 4811
rect 21315 4777 21324 4811
rect 21272 4768 21324 4777
rect 21088 4675 21140 4684
rect 21088 4641 21097 4675
rect 21097 4641 21131 4675
rect 21131 4641 21140 4675
rect 21088 4632 21140 4641
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 21088 4267 21140 4276
rect 21088 4233 21097 4267
rect 21097 4233 21131 4267
rect 21131 4233 21140 4267
rect 21088 4224 21140 4233
rect 2412 4131 2464 4140
rect 2412 4097 2421 4131
rect 2421 4097 2455 4131
rect 2455 4097 2464 4131
rect 2412 4088 2464 4097
rect 1400 3952 1452 4004
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 1400 3587 1452 3596
rect 1400 3553 1409 3587
rect 1409 3553 1443 3587
rect 1443 3553 1452 3587
rect 1400 3544 1452 3553
rect 23756 3544 23808 3596
rect 24860 3587 24912 3596
rect 24860 3553 24869 3587
rect 24869 3553 24903 3587
rect 24903 3553 24912 3587
rect 24860 3544 24912 3553
rect 25136 3476 25188 3528
rect 1584 3451 1636 3460
rect 1584 3417 1593 3451
rect 1593 3417 1627 3451
rect 1627 3417 1636 3451
rect 1584 3408 1636 3417
rect 25044 3383 25096 3392
rect 25044 3349 25053 3383
rect 25053 3349 25087 3383
rect 25087 3349 25096 3383
rect 25044 3340 25096 3349
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1400 3136 1452 3188
rect 4620 3136 4672 3188
rect 23756 3136 23808 3188
rect 24860 3179 24912 3188
rect 24860 3145 24869 3179
rect 24869 3145 24903 3179
rect 24903 3145 24912 3179
rect 24860 3136 24912 3145
rect 8116 2975 8168 2984
rect 8116 2941 8125 2975
rect 8125 2941 8159 2975
rect 8159 2941 8168 2975
rect 8116 2932 8168 2941
rect 23848 2975 23900 2984
rect 23848 2941 23857 2975
rect 23857 2941 23891 2975
rect 23891 2941 23900 2975
rect 23848 2932 23900 2941
rect 24860 2932 24912 2984
rect 25136 2975 25188 2984
rect 25136 2941 25145 2975
rect 25145 2941 25179 2975
rect 25179 2941 25188 2975
rect 25136 2932 25188 2941
rect 2688 2864 2740 2916
rect 8208 2864 8260 2916
rect 25320 2839 25372 2848
rect 25320 2805 25329 2839
rect 25329 2805 25363 2839
rect 25363 2805 25372 2839
rect 25320 2796 25372 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 2688 2592 2740 2644
rect 8208 2592 8260 2644
rect 24124 2456 24176 2508
rect 24860 2456 24912 2508
rect 1584 2295 1636 2304
rect 1584 2261 1593 2295
rect 1593 2261 1627 2295
rect 1627 2261 1636 2295
rect 1584 2252 1636 2261
rect 7564 2295 7616 2304
rect 7564 2261 7573 2295
rect 7573 2261 7607 2295
rect 7607 2261 7616 2295
rect 7564 2252 7616 2261
rect 23020 2295 23072 2304
rect 23020 2261 23029 2295
rect 23029 2261 23063 2295
rect 23063 2261 23072 2295
rect 23020 2252 23072 2261
rect 25504 2295 25556 2304
rect 25504 2261 25513 2295
rect 25513 2261 25547 2295
rect 25547 2261 25556 2295
rect 25504 2252 25556 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
<< metal2 >>
rect 202 27520 258 28000
rect 662 27520 718 28000
rect 1214 27520 1270 28000
rect 1306 27704 1362 27713
rect 1306 27639 1362 27648
rect 216 22137 244 27520
rect 676 24274 704 27520
rect 1228 24857 1256 27520
rect 1214 24848 1270 24857
rect 1214 24783 1270 24792
rect 664 24268 716 24274
rect 664 24210 716 24216
rect 572 22704 624 22710
rect 572 22646 624 22652
rect 584 22409 612 22646
rect 570 22400 626 22409
rect 570 22335 626 22344
rect 202 22128 258 22137
rect 202 22063 258 22072
rect 1320 18873 1348 27639
rect 1766 27520 1822 28000
rect 2318 27520 2374 28000
rect 2870 27520 2926 28000
rect 3422 27520 3478 28000
rect 3882 27520 3938 28000
rect 4434 27520 4490 28000
rect 4986 27520 5042 28000
rect 5538 27520 5594 28000
rect 6090 27520 6146 28000
rect 6642 27520 6698 28000
rect 7194 27520 7250 28000
rect 7654 27520 7710 28000
rect 8206 27520 8262 28000
rect 8758 27520 8814 28000
rect 9310 27520 9366 28000
rect 9862 27520 9918 28000
rect 10414 27520 10470 28000
rect 10874 27520 10930 28000
rect 11426 27520 11482 28000
rect 11978 27520 12034 28000
rect 12530 27520 12586 28000
rect 13082 27520 13138 28000
rect 13634 27520 13690 28000
rect 14186 27520 14242 28000
rect 14646 27520 14702 28000
rect 15198 27520 15254 28000
rect 15750 27520 15806 28000
rect 16302 27520 16358 28000
rect 16854 27520 16910 28000
rect 17406 27520 17462 28000
rect 17866 27520 17922 28000
rect 18418 27520 18474 28000
rect 18970 27520 19026 28000
rect 19522 27520 19578 28000
rect 20074 27520 20130 28000
rect 20626 27520 20682 28000
rect 21178 27520 21234 28000
rect 21638 27520 21694 28000
rect 22190 27520 22246 28000
rect 22742 27520 22798 28000
rect 23294 27520 23350 28000
rect 23570 27704 23626 27713
rect 23570 27639 23626 27648
rect 1582 27024 1638 27033
rect 1582 26959 1638 26968
rect 1596 24818 1624 26959
rect 1676 25288 1728 25294
rect 1676 25230 1728 25236
rect 1584 24812 1636 24818
rect 1584 24754 1636 24760
rect 1400 24608 1452 24614
rect 1400 24550 1452 24556
rect 1412 23730 1440 24550
rect 1400 23724 1452 23730
rect 1400 23666 1452 23672
rect 1412 23186 1440 23666
rect 1596 23594 1624 24754
rect 1688 24342 1716 25230
rect 1780 25208 1808 27520
rect 1780 25180 2176 25208
rect 1768 24744 1820 24750
rect 1768 24686 1820 24692
rect 1676 24336 1728 24342
rect 1676 24278 1728 24284
rect 1780 24138 1808 24686
rect 2044 24336 2096 24342
rect 2044 24278 2096 24284
rect 1768 24132 1820 24138
rect 1768 24074 1820 24080
rect 1766 23760 1822 23769
rect 1766 23695 1822 23704
rect 1584 23588 1636 23594
rect 1584 23530 1636 23536
rect 1400 23180 1452 23186
rect 1400 23122 1452 23128
rect 1412 22642 1440 23122
rect 1400 22636 1452 22642
rect 1400 22578 1452 22584
rect 1412 22098 1440 22578
rect 1780 22574 1808 23695
rect 1860 23248 1912 23254
rect 1860 23190 1912 23196
rect 1768 22568 1820 22574
rect 1768 22510 1820 22516
rect 1872 22506 1900 23190
rect 2056 22778 2084 24278
rect 2044 22772 2096 22778
rect 2044 22714 2096 22720
rect 1950 22536 2006 22545
rect 1860 22500 1912 22506
rect 1950 22471 2006 22480
rect 1860 22442 1912 22448
rect 1400 22092 1452 22098
rect 1400 22034 1452 22040
rect 1412 20466 1440 22034
rect 1492 21616 1544 21622
rect 1492 21558 1544 21564
rect 1504 21078 1532 21558
rect 1674 21448 1730 21457
rect 1674 21383 1730 21392
rect 1768 21412 1820 21418
rect 1492 21072 1544 21078
rect 1492 21014 1544 21020
rect 1688 20874 1716 21383
rect 1768 21354 1820 21360
rect 1780 21185 1808 21354
rect 1766 21176 1822 21185
rect 1766 21111 1822 21120
rect 1676 20868 1728 20874
rect 1676 20810 1728 20816
rect 1400 20460 1452 20466
rect 1400 20402 1452 20408
rect 1412 20058 1440 20402
rect 1400 20052 1452 20058
rect 1400 19994 1452 20000
rect 1412 19514 1440 19994
rect 1400 19508 1452 19514
rect 1400 19450 1452 19456
rect 1306 18864 1362 18873
rect 1306 18799 1362 18808
rect 1412 18612 1440 19450
rect 1584 18624 1636 18630
rect 1412 18584 1584 18612
rect 1584 18566 1636 18572
rect 1860 18624 1912 18630
rect 1860 18566 1912 18572
rect 1490 18320 1546 18329
rect 1490 18255 1546 18264
rect 1400 15904 1452 15910
rect 1400 15846 1452 15852
rect 1412 14550 1440 15846
rect 1400 14544 1452 14550
rect 1400 14486 1452 14492
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1412 11529 1440 12174
rect 1398 11520 1454 11529
rect 1398 11455 1454 11464
rect 1398 11248 1454 11257
rect 1398 11183 1400 11192
rect 1452 11183 1454 11192
rect 1400 11154 1452 11160
rect 1412 10266 1440 11154
rect 1400 10260 1452 10266
rect 1400 10202 1452 10208
rect 1398 10160 1454 10169
rect 1398 10095 1400 10104
rect 1452 10095 1454 10104
rect 1400 10066 1452 10072
rect 1412 9178 1440 10066
rect 1400 9172 1452 9178
rect 1400 9114 1452 9120
rect 1504 9058 1532 18255
rect 1596 18222 1624 18566
rect 1872 18222 1900 18566
rect 1584 18216 1636 18222
rect 1860 18216 1912 18222
rect 1584 18158 1636 18164
rect 1766 18184 1822 18193
rect 1596 16998 1624 18158
rect 1860 18158 1912 18164
rect 1766 18119 1822 18128
rect 1780 17610 1808 18119
rect 1768 17604 1820 17610
rect 1768 17546 1820 17552
rect 1676 17060 1728 17066
rect 1676 17002 1728 17008
rect 1584 16992 1636 16998
rect 1584 16934 1636 16940
rect 1596 15570 1624 16934
rect 1688 16794 1716 17002
rect 1780 16794 1808 17546
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1768 16788 1820 16794
rect 1768 16730 1820 16736
rect 1964 16658 1992 22471
rect 2148 22438 2176 25180
rect 2136 22432 2188 22438
rect 2136 22374 2188 22380
rect 2228 21888 2280 21894
rect 2228 21830 2280 21836
rect 2240 21418 2268 21830
rect 2228 21412 2280 21418
rect 2228 21354 2280 21360
rect 2044 21004 2096 21010
rect 2044 20946 2096 20952
rect 2056 20058 2084 20946
rect 2240 20398 2268 21354
rect 2332 21350 2360 27520
rect 2412 24676 2464 24682
rect 2412 24618 2464 24624
rect 2424 24585 2452 24618
rect 2410 24576 2466 24585
rect 2884 24562 2912 27520
rect 3436 24562 3464 27520
rect 3790 26344 3846 26353
rect 3790 26279 3846 26288
rect 3698 24848 3754 24857
rect 3804 24818 3832 26279
rect 3698 24783 3754 24792
rect 3792 24812 3844 24818
rect 3712 24682 3740 24783
rect 3792 24754 3844 24760
rect 3700 24676 3752 24682
rect 3700 24618 3752 24624
rect 2884 24534 3188 24562
rect 2410 24511 2466 24520
rect 2780 23520 2832 23526
rect 2780 23462 2832 23468
rect 2410 21992 2466 22001
rect 2792 21962 2820 23462
rect 2872 22636 2924 22642
rect 2872 22578 2924 22584
rect 2884 22166 2912 22578
rect 2964 22568 3016 22574
rect 2962 22536 2964 22545
rect 3016 22536 3018 22545
rect 2962 22471 3018 22480
rect 3056 22432 3108 22438
rect 3056 22374 3108 22380
rect 3068 22273 3096 22374
rect 3054 22264 3110 22273
rect 3054 22199 3110 22208
rect 2872 22160 2924 22166
rect 2872 22102 2924 22108
rect 2962 22128 3018 22137
rect 2410 21927 2466 21936
rect 2780 21956 2832 21962
rect 2320 21344 2372 21350
rect 2320 21286 2372 21292
rect 2332 21146 2360 21286
rect 2320 21140 2372 21146
rect 2320 21082 2372 21088
rect 2228 20392 2280 20398
rect 2228 20334 2280 20340
rect 2044 20052 2096 20058
rect 2044 19994 2096 20000
rect 2332 19281 2360 21082
rect 2424 19786 2452 21927
rect 2780 21898 2832 21904
rect 2792 21486 2820 21898
rect 2884 21690 2912 22102
rect 2962 22063 3018 22072
rect 2872 21684 2924 21690
rect 2872 21626 2924 21632
rect 2504 21480 2556 21486
rect 2504 21422 2556 21428
rect 2780 21480 2832 21486
rect 2780 21422 2832 21428
rect 2412 19780 2464 19786
rect 2412 19722 2464 19728
rect 2318 19272 2374 19281
rect 2318 19207 2374 19216
rect 2516 18630 2544 21422
rect 2976 21418 3004 22063
rect 2964 21412 3016 21418
rect 2964 21354 3016 21360
rect 2976 21146 3004 21354
rect 2964 21140 3016 21146
rect 2964 21082 3016 21088
rect 2688 21072 2740 21078
rect 2740 21020 2912 21026
rect 2688 21014 2912 21020
rect 2700 20998 2912 21014
rect 2688 20936 2740 20942
rect 2688 20878 2740 20884
rect 2700 20618 2728 20878
rect 2700 20602 2820 20618
rect 2700 20596 2832 20602
rect 2700 20590 2780 20596
rect 2596 19848 2648 19854
rect 2596 19790 2648 19796
rect 2608 19242 2636 19790
rect 2700 19310 2728 20590
rect 2780 20538 2832 20544
rect 2884 20534 2912 20998
rect 2872 20528 2924 20534
rect 2872 20470 2924 20476
rect 2964 20324 3016 20330
rect 2964 20266 3016 20272
rect 2780 19984 2832 19990
rect 2780 19926 2832 19932
rect 2688 19304 2740 19310
rect 2688 19246 2740 19252
rect 2596 19236 2648 19242
rect 2596 19178 2648 19184
rect 2700 18970 2728 19246
rect 2688 18964 2740 18970
rect 2688 18906 2740 18912
rect 2792 18850 2820 19926
rect 2976 19854 3004 20266
rect 2964 19848 3016 19854
rect 2964 19790 3016 19796
rect 2964 19168 3016 19174
rect 2964 19110 3016 19116
rect 2976 18902 3004 19110
rect 2700 18822 2820 18850
rect 2964 18896 3016 18902
rect 2964 18838 3016 18844
rect 2700 18698 2728 18822
rect 2780 18760 2832 18766
rect 2780 18702 2832 18708
rect 2688 18692 2740 18698
rect 2688 18634 2740 18640
rect 2504 18624 2556 18630
rect 2792 18601 2820 18702
rect 2504 18566 2556 18572
rect 2778 18592 2834 18601
rect 2778 18527 2834 18536
rect 2792 17882 2820 18527
rect 2872 18420 2924 18426
rect 2872 18362 2924 18368
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 2228 17672 2280 17678
rect 2228 17614 2280 17620
rect 2688 17672 2740 17678
rect 2688 17614 2740 17620
rect 2240 16794 2268 17614
rect 2700 17134 2728 17614
rect 2412 17128 2464 17134
rect 2412 17070 2464 17076
rect 2688 17128 2740 17134
rect 2688 17070 2740 17076
rect 2424 16998 2452 17070
rect 2412 16992 2464 16998
rect 2412 16934 2464 16940
rect 2228 16788 2280 16794
rect 2228 16730 2280 16736
rect 2134 16688 2190 16697
rect 1952 16652 2004 16658
rect 2134 16623 2136 16632
rect 1952 16594 2004 16600
rect 2188 16623 2190 16632
rect 2136 16594 2188 16600
rect 1584 15564 1636 15570
rect 1584 15506 1636 15512
rect 1596 14822 1624 15506
rect 2148 15162 2176 16594
rect 2240 16250 2268 16730
rect 2228 16244 2280 16250
rect 2228 16186 2280 16192
rect 2700 15688 2728 17070
rect 2884 16658 2912 18362
rect 2976 17882 3004 18838
rect 3160 18834 3188 24534
rect 3344 24534 3464 24562
rect 3238 23624 3294 23633
rect 3238 23559 3294 23568
rect 3252 22642 3280 23559
rect 3240 22636 3292 22642
rect 3240 22578 3292 22584
rect 3148 18828 3200 18834
rect 3148 18770 3200 18776
rect 3344 18465 3372 24534
rect 3424 24200 3476 24206
rect 3424 24142 3476 24148
rect 3436 23526 3464 24142
rect 3424 23520 3476 23526
rect 3424 23462 3476 23468
rect 3436 23322 3464 23462
rect 3424 23316 3476 23322
rect 3424 23258 3476 23264
rect 3436 22098 3464 23258
rect 3514 23216 3570 23225
rect 3514 23151 3516 23160
rect 3568 23151 3570 23160
rect 3516 23122 3568 23128
rect 3528 22438 3556 23122
rect 3712 22545 3740 24618
rect 3792 22976 3844 22982
rect 3792 22918 3844 22924
rect 3804 22574 3832 22918
rect 3792 22568 3844 22574
rect 3698 22536 3754 22545
rect 3792 22510 3844 22516
rect 3698 22471 3754 22480
rect 3516 22432 3568 22438
rect 3516 22374 3568 22380
rect 3528 22234 3556 22374
rect 3516 22228 3568 22234
rect 3516 22170 3568 22176
rect 3424 22092 3476 22098
rect 3424 22034 3476 22040
rect 3436 21690 3464 22034
rect 3424 21684 3476 21690
rect 3424 21626 3476 21632
rect 3712 21554 3740 22471
rect 3792 22432 3844 22438
rect 3792 22374 3844 22380
rect 3804 22273 3832 22374
rect 3790 22264 3846 22273
rect 3790 22199 3846 22208
rect 3792 21616 3844 21622
rect 3792 21558 3844 21564
rect 3700 21548 3752 21554
rect 3700 21490 3752 21496
rect 3712 21146 3740 21490
rect 3700 21140 3752 21146
rect 3700 21082 3752 21088
rect 3700 20800 3752 20806
rect 3700 20742 3752 20748
rect 3712 20398 3740 20742
rect 3700 20392 3752 20398
rect 3700 20334 3752 20340
rect 3712 20058 3740 20334
rect 3804 20058 3832 21558
rect 3896 20233 3924 27520
rect 4068 25832 4120 25838
rect 4068 25774 4120 25780
rect 3974 25664 4030 25673
rect 3974 25599 4030 25608
rect 3988 25226 4016 25599
rect 3976 25220 4028 25226
rect 3976 25162 4028 25168
rect 4080 25129 4108 25774
rect 4066 25120 4122 25129
rect 4066 25055 4122 25064
rect 4344 24608 4396 24614
rect 4344 24550 4396 24556
rect 4160 24200 4212 24206
rect 4160 24142 4212 24148
rect 4172 23866 4200 24142
rect 4160 23860 4212 23866
rect 4160 23802 4212 23808
rect 4172 23322 4200 23802
rect 4356 23594 4384 24550
rect 4344 23588 4396 23594
rect 4344 23530 4396 23536
rect 4160 23316 4212 23322
rect 4160 23258 4212 23264
rect 4172 22778 4200 23258
rect 4160 22772 4212 22778
rect 4160 22714 4212 22720
rect 3974 22672 4030 22681
rect 4172 22658 4200 22714
rect 4172 22630 4292 22658
rect 3974 22607 4030 22616
rect 3988 22137 4016 22607
rect 4264 22166 4292 22630
rect 4356 22506 4384 23530
rect 4344 22500 4396 22506
rect 4344 22442 4396 22448
rect 4252 22160 4304 22166
rect 3974 22128 4030 22137
rect 4252 22102 4304 22108
rect 3974 22063 4030 22072
rect 4264 20262 4292 22102
rect 4344 22092 4396 22098
rect 4344 22034 4396 22040
rect 4356 22001 4384 22034
rect 4342 21992 4398 22001
rect 4342 21927 4398 21936
rect 4252 20256 4304 20262
rect 3882 20224 3938 20233
rect 4252 20198 4304 20204
rect 3882 20159 3938 20168
rect 3700 20052 3752 20058
rect 3700 19994 3752 20000
rect 3792 20052 3844 20058
rect 3792 19994 3844 20000
rect 3700 19848 3752 19854
rect 3700 19790 3752 19796
rect 3712 18970 3740 19790
rect 3804 19378 3832 19994
rect 4264 19938 4292 20198
rect 4172 19922 4292 19938
rect 4160 19916 4292 19922
rect 4212 19910 4292 19916
rect 4344 19916 4396 19922
rect 4160 19858 4212 19864
rect 4344 19858 4396 19864
rect 4172 19428 4200 19858
rect 4252 19440 4304 19446
rect 4172 19400 4252 19428
rect 4252 19382 4304 19388
rect 3792 19372 3844 19378
rect 3792 19314 3844 19320
rect 3790 19272 3846 19281
rect 3846 19230 4200 19258
rect 3790 19207 3846 19216
rect 4172 19174 4200 19230
rect 4160 19168 4212 19174
rect 4160 19110 4212 19116
rect 3700 18964 3752 18970
rect 3700 18906 3752 18912
rect 3608 18828 3660 18834
rect 3608 18770 3660 18776
rect 3330 18456 3386 18465
rect 3330 18391 3386 18400
rect 2964 17876 3016 17882
rect 2964 17818 3016 17824
rect 3240 17808 3292 17814
rect 3240 17750 3292 17756
rect 3252 16658 3280 17750
rect 2872 16652 2924 16658
rect 2872 16594 2924 16600
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 2884 16096 2912 16594
rect 3056 16108 3108 16114
rect 2884 16068 3056 16096
rect 2780 15700 2832 15706
rect 2700 15660 2780 15688
rect 2504 15428 2556 15434
rect 2504 15370 2556 15376
rect 2226 15328 2282 15337
rect 2226 15263 2282 15272
rect 2136 15156 2188 15162
rect 2136 15098 2188 15104
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1584 14816 1636 14822
rect 1584 14758 1636 14764
rect 1780 14346 1808 14962
rect 1952 14884 2004 14890
rect 1952 14826 2004 14832
rect 1768 14340 1820 14346
rect 1768 14282 1820 14288
rect 1964 14074 1992 14826
rect 2136 14816 2188 14822
rect 2136 14758 2188 14764
rect 2044 14544 2096 14550
rect 2044 14486 2096 14492
rect 2056 14074 2084 14486
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 2044 14068 2096 14074
rect 2044 14010 2096 14016
rect 1766 13968 1822 13977
rect 1766 13903 1822 13912
rect 1780 13870 1808 13903
rect 1768 13864 1820 13870
rect 1768 13806 1820 13812
rect 1780 13530 1808 13806
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1768 13524 1820 13530
rect 1768 13466 1820 13472
rect 1964 13190 1992 13670
rect 2044 13456 2096 13462
rect 2044 13398 2096 13404
rect 1952 13184 2004 13190
rect 1952 13126 2004 13132
rect 1860 11824 1912 11830
rect 1860 11766 1912 11772
rect 1768 10464 1820 10470
rect 1768 10406 1820 10412
rect 1676 9920 1728 9926
rect 1676 9862 1728 9868
rect 1582 9480 1638 9489
rect 1582 9415 1638 9424
rect 1596 9382 1624 9415
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1412 9030 1532 9058
rect 1412 8430 1440 9030
rect 1492 8832 1544 8838
rect 1492 8774 1544 8780
rect 1582 8800 1638 8809
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1398 7848 1454 7857
rect 1398 7783 1454 7792
rect 1412 7342 1440 7783
rect 1400 7336 1452 7342
rect 1400 7278 1452 7284
rect 1412 7002 1440 7278
rect 1400 6996 1452 7002
rect 1400 6938 1452 6944
rect 1504 4185 1532 8774
rect 1582 8735 1638 8744
rect 1596 8634 1624 8735
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1582 8120 1638 8129
rect 1582 8055 1584 8064
rect 1636 8055 1638 8064
rect 1584 8026 1636 8032
rect 1584 7472 1636 7478
rect 1582 7440 1584 7449
rect 1636 7440 1638 7449
rect 1582 7375 1638 7384
rect 1688 4865 1716 9862
rect 1674 4856 1730 4865
rect 1674 4791 1730 4800
rect 1490 4176 1546 4185
rect 1490 4111 1546 4120
rect 1400 4004 1452 4010
rect 1400 3946 1452 3952
rect 1412 3602 1440 3946
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 1412 3194 1440 3538
rect 1582 3496 1638 3505
rect 1582 3431 1584 3440
rect 1636 3431 1638 3440
rect 1584 3402 1636 3408
rect 1400 3188 1452 3194
rect 1400 3130 1452 3136
rect 1780 2961 1808 10406
rect 1872 3097 1900 11766
rect 1964 10606 1992 13126
rect 2056 12918 2084 13398
rect 2044 12912 2096 12918
rect 2044 12854 2096 12860
rect 2148 12782 2176 14758
rect 2240 14550 2268 15263
rect 2516 15094 2544 15370
rect 2596 15360 2648 15366
rect 2596 15302 2648 15308
rect 2504 15088 2556 15094
rect 2504 15030 2556 15036
rect 2608 14890 2636 15302
rect 2700 15026 2728 15660
rect 2780 15642 2832 15648
rect 2884 15570 2912 16068
rect 3056 16050 3108 16056
rect 3344 16046 3372 18391
rect 3620 18086 3648 18770
rect 3712 18154 3740 18906
rect 4160 18828 4212 18834
rect 4160 18770 4212 18776
rect 3700 18148 3752 18154
rect 3700 18090 3752 18096
rect 3608 18080 3660 18086
rect 3606 18048 3608 18057
rect 3660 18048 3662 18057
rect 3606 17983 3662 17992
rect 3974 17912 4030 17921
rect 4172 17882 4200 18770
rect 4264 18222 4292 19382
rect 4356 19242 4384 19858
rect 4344 19236 4396 19242
rect 4344 19178 4396 19184
rect 4356 18970 4384 19178
rect 4344 18964 4396 18970
rect 4344 18906 4396 18912
rect 4252 18216 4304 18222
rect 4252 18158 4304 18164
rect 4344 18148 4396 18154
rect 4344 18090 4396 18096
rect 4356 17882 4384 18090
rect 3974 17847 4030 17856
rect 4160 17876 4212 17882
rect 3424 16992 3476 16998
rect 3424 16934 3476 16940
rect 3436 16726 3464 16934
rect 3424 16720 3476 16726
rect 3424 16662 3476 16668
rect 3436 16250 3464 16662
rect 3424 16244 3476 16250
rect 3424 16186 3476 16192
rect 3332 16040 3384 16046
rect 3988 16017 4016 17847
rect 4160 17818 4212 17824
rect 4344 17876 4396 17882
rect 4344 17818 4396 17824
rect 4160 16992 4212 16998
rect 4080 16940 4160 16946
rect 4080 16934 4212 16940
rect 4080 16918 4200 16934
rect 3332 15982 3384 15988
rect 3974 16008 4030 16017
rect 3344 15910 3372 15982
rect 3974 15943 4030 15952
rect 3332 15904 3384 15910
rect 4080 15881 4108 16918
rect 4252 16176 4304 16182
rect 4158 16144 4214 16153
rect 4252 16118 4304 16124
rect 4158 16079 4214 16088
rect 3332 15846 3384 15852
rect 4066 15872 4122 15881
rect 4066 15807 4122 15816
rect 4172 15688 4200 16079
rect 4080 15660 4200 15688
rect 4080 15570 4108 15660
rect 2872 15564 2924 15570
rect 2872 15506 2924 15512
rect 4068 15564 4120 15570
rect 4068 15506 4120 15512
rect 2884 15162 2912 15506
rect 3606 15464 3662 15473
rect 3606 15399 3662 15408
rect 3620 15162 3648 15399
rect 3792 15360 3844 15366
rect 3792 15302 3844 15308
rect 2872 15156 2924 15162
rect 2872 15098 2924 15104
rect 3608 15156 3660 15162
rect 3608 15098 3660 15104
rect 2688 15020 2740 15026
rect 2688 14962 2740 14968
rect 2596 14884 2648 14890
rect 2596 14826 2648 14832
rect 2884 14618 2912 15098
rect 3514 15056 3570 15065
rect 3514 14991 3570 15000
rect 3056 14952 3108 14958
rect 3056 14894 3108 14900
rect 2872 14612 2924 14618
rect 2872 14554 2924 14560
rect 2228 14544 2280 14550
rect 2228 14486 2280 14492
rect 2320 14544 2372 14550
rect 2320 14486 2372 14492
rect 2332 13938 2360 14486
rect 2504 14476 2556 14482
rect 2504 14418 2556 14424
rect 2516 14385 2544 14418
rect 2502 14376 2558 14385
rect 2502 14311 2558 14320
rect 2516 14006 2544 14311
rect 2504 14000 2556 14006
rect 2504 13942 2556 13948
rect 2320 13932 2372 13938
rect 2320 13874 2372 13880
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2136 12776 2188 12782
rect 2136 12718 2188 12724
rect 2502 12744 2558 12753
rect 2148 12306 2176 12718
rect 2502 12679 2558 12688
rect 2136 12300 2188 12306
rect 2136 12242 2188 12248
rect 2412 12096 2464 12102
rect 2412 12038 2464 12044
rect 2136 11620 2188 11626
rect 2136 11562 2188 11568
rect 2320 11620 2372 11626
rect 2320 11562 2372 11568
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 2148 10554 2176 11562
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 2240 11064 2268 11494
rect 2332 11354 2360 11562
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 2320 11076 2372 11082
rect 2240 11036 2320 11064
rect 2320 11018 2372 11024
rect 2148 10526 2268 10554
rect 2240 10470 2268 10526
rect 2044 10464 2096 10470
rect 2044 10406 2096 10412
rect 2228 10464 2280 10470
rect 2228 10406 2280 10412
rect 2056 10305 2084 10406
rect 2042 10296 2098 10305
rect 2042 10231 2098 10240
rect 2044 9036 2096 9042
rect 2044 8978 2096 8984
rect 2056 8945 2084 8978
rect 2042 8936 2098 8945
rect 2042 8871 2098 8880
rect 2056 8634 2084 8871
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 2042 8120 2098 8129
rect 2042 8055 2098 8064
rect 2056 7954 2084 8055
rect 2240 7993 2268 10406
rect 2226 7984 2282 7993
rect 2044 7948 2096 7954
rect 2226 7919 2282 7928
rect 2044 7890 2096 7896
rect 2056 7546 2084 7890
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 2332 7449 2360 11018
rect 2318 7440 2374 7449
rect 2318 7375 2374 7384
rect 2424 4146 2452 12038
rect 2516 9654 2544 12679
rect 2792 12442 2820 13874
rect 3068 13530 3096 14894
rect 3148 14816 3200 14822
rect 3148 14758 3200 14764
rect 3238 14784 3294 14793
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 2964 13456 3016 13462
rect 2962 13424 2964 13433
rect 3016 13424 3018 13433
rect 2884 13382 2962 13410
rect 2884 12986 2912 13382
rect 2962 13359 3018 13368
rect 2872 12980 2924 12986
rect 2872 12922 2924 12928
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2792 12322 2820 12378
rect 2608 12294 2820 12322
rect 3056 12368 3108 12374
rect 3056 12310 3108 12316
rect 2608 10266 2636 12294
rect 3068 11898 3096 12310
rect 3056 11892 3108 11898
rect 3056 11834 3108 11840
rect 2870 11656 2926 11665
rect 2870 11591 2872 11600
rect 2924 11591 2926 11600
rect 2872 11562 2924 11568
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 2792 10742 2820 11154
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2688 10736 2740 10742
rect 2686 10704 2688 10713
rect 2780 10736 2832 10742
rect 2740 10704 2742 10713
rect 2780 10678 2832 10684
rect 2686 10639 2742 10648
rect 2884 10606 2912 11086
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 2700 10130 2820 10146
rect 2688 10124 2820 10130
rect 2740 10118 2820 10124
rect 2688 10066 2740 10072
rect 2686 10024 2742 10033
rect 2686 9959 2688 9968
rect 2740 9959 2742 9968
rect 2688 9930 2740 9936
rect 2504 9648 2556 9654
rect 2504 9590 2556 9596
rect 2792 9382 2820 10118
rect 2870 10024 2926 10033
rect 2870 9959 2926 9968
rect 2884 9586 2912 9959
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 2870 9480 2926 9489
rect 2870 9415 2872 9424
rect 2924 9415 2926 9424
rect 2872 9386 2924 9392
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2976 5545 3004 11290
rect 3160 6769 3188 14758
rect 3238 14719 3294 14728
rect 3252 13326 3280 14719
rect 3332 14476 3384 14482
rect 3332 14418 3384 14424
rect 3344 14074 3372 14418
rect 3332 14068 3384 14074
rect 3332 14010 3384 14016
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 3252 12442 3280 13262
rect 3344 12986 3372 14010
rect 3332 12980 3384 12986
rect 3332 12922 3384 12928
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 3344 12374 3372 12922
rect 3332 12368 3384 12374
rect 3332 12310 3384 12316
rect 3330 12200 3386 12209
rect 3330 12135 3332 12144
rect 3384 12135 3386 12144
rect 3332 12106 3384 12112
rect 3344 11898 3372 12106
rect 3332 11892 3384 11898
rect 3332 11834 3384 11840
rect 3332 11552 3384 11558
rect 3332 11494 3384 11500
rect 3344 10266 3372 11494
rect 3528 11257 3556 14991
rect 3620 14958 3648 15098
rect 3608 14952 3660 14958
rect 3608 14894 3660 14900
rect 3698 14648 3754 14657
rect 3698 14583 3754 14592
rect 3608 14272 3660 14278
rect 3608 14214 3660 14220
rect 3620 14006 3648 14214
rect 3608 14000 3660 14006
rect 3608 13942 3660 13948
rect 3620 13734 3648 13942
rect 3608 13728 3660 13734
rect 3608 13670 3660 13676
rect 3712 12889 3740 14583
rect 3804 13297 3832 15302
rect 4172 15162 4200 15660
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 4080 14414 4108 14894
rect 4068 14408 4120 14414
rect 4120 14368 4200 14396
rect 4068 14350 4120 14356
rect 4068 14272 4120 14278
rect 4068 14214 4120 14220
rect 4080 13938 4108 14214
rect 4172 14074 4200 14368
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4068 13932 4120 13938
rect 4120 13892 4200 13920
rect 4068 13874 4120 13880
rect 4068 13796 4120 13802
rect 4068 13738 4120 13744
rect 3974 13696 4030 13705
rect 3974 13631 4030 13640
rect 3884 13524 3936 13530
rect 3884 13466 3936 13472
rect 3790 13288 3846 13297
rect 3790 13223 3846 13232
rect 3698 12880 3754 12889
rect 3698 12815 3754 12824
rect 3896 12714 3924 13466
rect 3988 13462 4016 13631
rect 4080 13530 4108 13738
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 3976 13456 4028 13462
rect 3976 13398 4028 13404
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 3884 12708 3936 12714
rect 3884 12650 3936 12656
rect 3896 12102 3924 12650
rect 3884 12096 3936 12102
rect 3988 12073 4016 13126
rect 4080 12850 4108 13330
rect 4172 12986 4200 13892
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 4068 12708 4120 12714
rect 4068 12650 4120 12656
rect 3884 12038 3936 12044
rect 3974 12064 4030 12073
rect 3896 11694 3924 12038
rect 3974 11999 4030 12008
rect 4080 11914 4108 12650
rect 3988 11886 4108 11914
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 3790 11384 3846 11393
rect 3790 11319 3846 11328
rect 3514 11248 3570 11257
rect 3514 11183 3570 11192
rect 3804 10810 3832 11319
rect 3792 10804 3844 10810
rect 3792 10746 3844 10752
rect 3988 10742 4016 11886
rect 4264 11801 4292 16118
rect 4344 14884 4396 14890
rect 4344 14826 4396 14832
rect 4356 14793 4384 14826
rect 4342 14784 4398 14793
rect 4342 14719 4398 14728
rect 4356 14618 4384 14719
rect 4344 14612 4396 14618
rect 4344 14554 4396 14560
rect 4448 13462 4476 27520
rect 4712 25152 4764 25158
rect 4712 25094 4764 25100
rect 4724 24818 4752 25094
rect 5000 24857 5028 27520
rect 5080 25288 5132 25294
rect 5080 25230 5132 25236
rect 4986 24848 5042 24857
rect 4712 24812 4764 24818
rect 4986 24783 5042 24792
rect 4712 24754 4764 24760
rect 4528 24064 4580 24070
rect 4528 24006 4580 24012
rect 4540 23662 4568 24006
rect 4528 23656 4580 23662
rect 4528 23598 4580 23604
rect 4540 23497 4568 23598
rect 4724 23526 4752 24754
rect 5092 24614 5120 25230
rect 5552 24732 5580 27520
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5552 24704 6040 24732
rect 5080 24608 5132 24614
rect 5080 24550 5132 24556
rect 5540 24608 5592 24614
rect 5540 24550 5592 24556
rect 4802 24440 4858 24449
rect 4802 24375 4858 24384
rect 4712 23520 4764 23526
rect 4526 23488 4582 23497
rect 4712 23462 4764 23468
rect 4526 23423 4582 23432
rect 4724 23254 4752 23462
rect 4712 23248 4764 23254
rect 4712 23190 4764 23196
rect 4526 22536 4582 22545
rect 4526 22471 4582 22480
rect 4540 22137 4568 22471
rect 4526 22128 4582 22137
rect 4526 22063 4582 22072
rect 4620 22024 4672 22030
rect 4618 21992 4620 22001
rect 4672 21992 4674 22001
rect 4618 21927 4674 21936
rect 4816 20097 4844 24375
rect 4988 24268 5040 24274
rect 4988 24210 5040 24216
rect 4896 21888 4948 21894
rect 4896 21830 4948 21836
rect 4908 21010 4936 21830
rect 4896 21004 4948 21010
rect 4896 20946 4948 20952
rect 4908 20806 4936 20946
rect 4896 20800 4948 20806
rect 4896 20742 4948 20748
rect 4908 20330 4936 20742
rect 5000 20369 5028 24210
rect 5092 22778 5120 24550
rect 5172 24268 5224 24274
rect 5172 24210 5224 24216
rect 5184 23594 5212 24210
rect 5172 23588 5224 23594
rect 5172 23530 5224 23536
rect 5080 22772 5132 22778
rect 5080 22714 5132 22720
rect 5184 22574 5212 23530
rect 5552 23202 5580 24550
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5632 23520 5684 23526
rect 5632 23462 5684 23468
rect 5816 23520 5868 23526
rect 5816 23462 5868 23468
rect 5460 23174 5580 23202
rect 5460 22778 5488 23174
rect 5644 23066 5672 23462
rect 5828 23322 5856 23462
rect 6012 23361 6040 24704
rect 5998 23352 6054 23361
rect 5816 23316 5868 23322
rect 5998 23287 6054 23296
rect 5816 23258 5868 23264
rect 6104 23236 6132 27520
rect 6276 24064 6328 24070
rect 6276 24006 6328 24012
rect 5552 23038 5672 23066
rect 6012 23208 6132 23236
rect 6288 23225 6316 24006
rect 6274 23216 6330 23225
rect 5552 22778 5580 23038
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5448 22772 5500 22778
rect 5448 22714 5500 22720
rect 5540 22772 5592 22778
rect 5540 22714 5592 22720
rect 5172 22568 5224 22574
rect 5448 22568 5500 22574
rect 5172 22510 5224 22516
rect 5446 22536 5448 22545
rect 5500 22536 5502 22545
rect 5184 22234 5212 22510
rect 5446 22471 5502 22480
rect 5460 22234 5672 22250
rect 5172 22228 5224 22234
rect 5172 22170 5224 22176
rect 5448 22228 5672 22234
rect 5500 22222 5672 22228
rect 5448 22170 5500 22176
rect 5644 22166 5672 22222
rect 5632 22160 5684 22166
rect 5632 22102 5684 22108
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5540 21616 5592 21622
rect 5540 21558 5592 21564
rect 5264 21412 5316 21418
rect 5264 21354 5316 21360
rect 5080 20936 5132 20942
rect 5080 20878 5132 20884
rect 4986 20360 5042 20369
rect 4896 20324 4948 20330
rect 4986 20295 5042 20304
rect 4896 20266 4948 20272
rect 5092 20262 5120 20878
rect 5276 20602 5304 21354
rect 5448 20800 5500 20806
rect 5448 20742 5500 20748
rect 5264 20596 5316 20602
rect 5264 20538 5316 20544
rect 5460 20466 5488 20742
rect 5448 20460 5500 20466
rect 5448 20402 5500 20408
rect 5080 20256 5132 20262
rect 5080 20198 5132 20204
rect 4802 20088 4858 20097
rect 4802 20023 4858 20032
rect 5552 19922 5580 21558
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5816 20460 5868 20466
rect 5816 20402 5868 20408
rect 5724 20256 5776 20262
rect 5724 20198 5776 20204
rect 5736 20058 5764 20198
rect 5724 20052 5776 20058
rect 5724 19994 5776 20000
rect 5540 19916 5592 19922
rect 5540 19858 5592 19864
rect 5828 19786 5856 20402
rect 5816 19780 5868 19786
rect 5816 19722 5868 19728
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 4986 19272 5042 19281
rect 4986 19207 4988 19216
rect 5040 19207 5042 19216
rect 5356 19236 5408 19242
rect 4988 19178 5040 19184
rect 5356 19178 5408 19184
rect 4528 19168 4580 19174
rect 4528 19110 4580 19116
rect 4540 17814 4568 19110
rect 4710 19000 4766 19009
rect 4710 18935 4766 18944
rect 4724 18578 4752 18935
rect 5264 18896 5316 18902
rect 4986 18864 5042 18873
rect 5262 18864 5264 18873
rect 5316 18864 5318 18873
rect 4986 18799 5042 18808
rect 5184 18822 5262 18850
rect 4802 18728 4858 18737
rect 4802 18663 4804 18672
rect 4856 18663 4858 18672
rect 4804 18634 4856 18640
rect 4724 18550 4844 18578
rect 4816 18465 4844 18550
rect 4802 18456 4858 18465
rect 4802 18391 4858 18400
rect 4816 17814 4844 18391
rect 4528 17808 4580 17814
rect 4528 17750 4580 17756
rect 4804 17808 4856 17814
rect 4804 17750 4856 17756
rect 4816 17202 4844 17750
rect 4804 17196 4856 17202
rect 4804 17138 4856 17144
rect 4804 16652 4856 16658
rect 4804 16594 4856 16600
rect 4620 16176 4672 16182
rect 4620 16118 4672 16124
rect 4528 13796 4580 13802
rect 4528 13738 4580 13744
rect 4436 13456 4488 13462
rect 4436 13398 4488 13404
rect 4540 13258 4568 13738
rect 4528 13252 4580 13258
rect 4528 13194 4580 13200
rect 4632 12356 4660 16118
rect 4816 15910 4844 16594
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 4816 15638 4844 15846
rect 4804 15632 4856 15638
rect 4804 15574 4856 15580
rect 4816 14958 4844 15574
rect 4804 14952 4856 14958
rect 4804 14894 4856 14900
rect 4710 13288 4766 13297
rect 4710 13223 4712 13232
rect 4764 13223 4766 13232
rect 4712 13194 4764 13200
rect 4724 12714 4752 13194
rect 4712 12708 4764 12714
rect 4712 12650 4764 12656
rect 4632 12328 4752 12356
rect 4250 11792 4306 11801
rect 4068 11756 4120 11762
rect 4250 11727 4306 11736
rect 4068 11698 4120 11704
rect 4080 11082 4108 11698
rect 4434 11520 4490 11529
rect 4434 11455 4490 11464
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 4068 11076 4120 11082
rect 4068 11018 4120 11024
rect 3976 10736 4028 10742
rect 3976 10678 4028 10684
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3252 8537 3280 9318
rect 3238 8528 3294 8537
rect 3238 8463 3294 8472
rect 3146 6760 3202 6769
rect 3146 6695 3202 6704
rect 2962 5536 3018 5545
rect 2962 5471 3018 5480
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 1858 3088 1914 3097
rect 1858 3023 1914 3032
rect 1766 2952 1822 2961
rect 1766 2887 1822 2896
rect 2688 2916 2740 2922
rect 2688 2858 2740 2864
rect 2700 2650 2728 2858
rect 2688 2644 2740 2650
rect 2688 2586 2740 2592
rect 1584 2304 1636 2310
rect 1582 2272 1584 2281
rect 1636 2272 1638 2281
rect 1582 2207 1638 2216
rect 3528 377 3556 10406
rect 3620 10266 3648 10542
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 4080 9654 4108 11018
rect 4172 10606 4200 11086
rect 4160 10600 4212 10606
rect 4160 10542 4212 10548
rect 4356 10266 4384 11290
rect 4448 11286 4476 11455
rect 4436 11280 4488 11286
rect 4436 11222 4488 11228
rect 4528 11280 4580 11286
rect 4528 11222 4580 11228
rect 4448 10810 4476 11222
rect 4436 10804 4488 10810
rect 4436 10746 4488 10752
rect 4540 10470 4568 11222
rect 4620 10736 4672 10742
rect 4620 10678 4672 10684
rect 4528 10464 4580 10470
rect 4526 10432 4528 10441
rect 4580 10432 4582 10441
rect 4526 10367 4582 10376
rect 4344 10260 4396 10266
rect 4344 10202 4396 10208
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4344 9512 4396 9518
rect 4344 9454 4396 9460
rect 4264 9110 4292 9454
rect 4356 9178 4384 9454
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4252 9104 4304 9110
rect 4252 9046 4304 9052
rect 4250 6216 4306 6225
rect 4250 6151 4306 6160
rect 4264 6118 4292 6151
rect 4252 6112 4304 6118
rect 4252 6054 4304 6060
rect 4632 3194 4660 10678
rect 4724 9659 4752 12328
rect 5000 11694 5028 18799
rect 5184 17338 5212 18822
rect 5262 18799 5318 18808
rect 5264 18760 5316 18766
rect 5264 18702 5316 18708
rect 5276 17882 5304 18702
rect 5368 18426 5396 19178
rect 5448 18828 5500 18834
rect 5448 18770 5500 18776
rect 5356 18420 5408 18426
rect 5356 18362 5408 18368
rect 5460 17882 5488 18770
rect 5540 18624 5592 18630
rect 5540 18566 5592 18572
rect 5552 18193 5580 18566
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5538 18184 5594 18193
rect 5538 18119 5594 18128
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 5264 17876 5316 17882
rect 5264 17818 5316 17824
rect 5448 17876 5500 17882
rect 5448 17818 5500 17824
rect 5446 17776 5502 17785
rect 5552 17746 5580 18022
rect 5446 17711 5502 17720
rect 5540 17740 5592 17746
rect 5172 17332 5224 17338
rect 5172 17274 5224 17280
rect 5460 16794 5488 17711
rect 5540 17682 5592 17688
rect 5552 17270 5580 17682
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5540 17264 5592 17270
rect 5540 17206 5592 17212
rect 5552 17066 5580 17206
rect 5540 17060 5592 17066
rect 5540 17002 5592 17008
rect 5552 16794 5580 17002
rect 5448 16788 5500 16794
rect 5448 16730 5500 16736
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6012 15881 6040 23208
rect 6274 23151 6330 23160
rect 6656 22964 6684 27520
rect 7208 26466 7236 27520
rect 7208 26438 7604 26466
rect 7380 26308 7432 26314
rect 7380 26250 7432 26256
rect 7104 25356 7156 25362
rect 7104 25298 7156 25304
rect 7012 24676 7064 24682
rect 7012 24618 7064 24624
rect 7024 23254 7052 24618
rect 7116 24614 7144 25298
rect 7104 24608 7156 24614
rect 7104 24550 7156 24556
rect 7116 23594 7144 24550
rect 7196 24064 7248 24070
rect 7196 24006 7248 24012
rect 7104 23588 7156 23594
rect 7104 23530 7156 23536
rect 7012 23248 7064 23254
rect 7012 23190 7064 23196
rect 6656 22936 6776 22964
rect 6184 22568 6236 22574
rect 6184 22510 6236 22516
rect 6196 21978 6224 22510
rect 6368 22432 6420 22438
rect 6368 22374 6420 22380
rect 6380 22030 6408 22374
rect 6748 22080 6776 22936
rect 6828 22568 6880 22574
rect 6828 22510 6880 22516
rect 6840 22250 6868 22510
rect 7104 22500 7156 22506
rect 7104 22442 7156 22448
rect 6840 22222 7052 22250
rect 6828 22160 6880 22166
rect 6880 22108 6960 22114
rect 6828 22102 6960 22108
rect 6840 22086 6960 22102
rect 6564 22052 6776 22080
rect 6104 21950 6224 21978
rect 6368 22024 6420 22030
rect 6368 21966 6420 21972
rect 6104 21894 6132 21950
rect 6092 21888 6144 21894
rect 6092 21830 6144 21836
rect 6104 21554 6132 21830
rect 6092 21548 6144 21554
rect 6092 21490 6144 21496
rect 6460 21480 6512 21486
rect 6460 21422 6512 21428
rect 6472 21146 6500 21422
rect 6460 21140 6512 21146
rect 6460 21082 6512 21088
rect 6276 20256 6328 20262
rect 6276 20198 6328 20204
rect 6184 19916 6236 19922
rect 6184 19858 6236 19864
rect 6196 19514 6224 19858
rect 6184 19508 6236 19514
rect 6184 19450 6236 19456
rect 6184 18760 6236 18766
rect 6288 18748 6316 20198
rect 6236 18720 6316 18748
rect 6184 18702 6236 18708
rect 6092 18624 6144 18630
rect 6092 18566 6144 18572
rect 6104 16697 6132 18566
rect 6196 18222 6224 18702
rect 6184 18216 6236 18222
rect 6184 18158 6236 18164
rect 6196 18086 6224 18158
rect 6184 18080 6236 18086
rect 6184 18022 6236 18028
rect 6196 17542 6224 18022
rect 6184 17536 6236 17542
rect 6184 17478 6236 17484
rect 6196 17066 6224 17478
rect 6184 17060 6236 17066
rect 6184 17002 6236 17008
rect 6090 16688 6146 16697
rect 6090 16623 6146 16632
rect 5998 15872 6054 15881
rect 5998 15807 6054 15816
rect 6092 15632 6144 15638
rect 6196 15620 6224 17002
rect 6144 15592 6224 15620
rect 6092 15574 6144 15580
rect 5540 15564 5592 15570
rect 5540 15506 5592 15512
rect 5080 15360 5132 15366
rect 5080 15302 5132 15308
rect 5092 14890 5120 15302
rect 5552 15162 5580 15506
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 6196 15162 6224 15592
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 6184 15156 6236 15162
rect 6184 15098 6236 15104
rect 5080 14884 5132 14890
rect 5080 14826 5132 14832
rect 5092 14618 5120 14826
rect 5552 14618 5580 15098
rect 6564 14657 6592 22052
rect 6644 21480 6696 21486
rect 6644 21422 6696 21428
rect 6656 21350 6684 21422
rect 6644 21344 6696 21350
rect 6644 21286 6696 21292
rect 6656 20398 6684 21286
rect 6828 20868 6880 20874
rect 6828 20810 6880 20816
rect 6644 20392 6696 20398
rect 6644 20334 6696 20340
rect 6840 20058 6868 20810
rect 6828 20052 6880 20058
rect 6828 19994 6880 20000
rect 6736 19848 6788 19854
rect 6736 19790 6788 19796
rect 6644 18420 6696 18426
rect 6644 18362 6696 18368
rect 6656 16046 6684 18362
rect 6748 18329 6776 19790
rect 6932 19310 6960 22086
rect 7024 21894 7052 22222
rect 7012 21888 7064 21894
rect 7012 21830 7064 21836
rect 7024 21457 7052 21830
rect 7010 21448 7066 21457
rect 7010 21383 7066 21392
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 7012 18828 7064 18834
rect 7012 18770 7064 18776
rect 7024 18426 7052 18770
rect 7116 18737 7144 22442
rect 7102 18728 7158 18737
rect 7102 18663 7158 18672
rect 7012 18420 7064 18426
rect 7012 18362 7064 18368
rect 6734 18320 6790 18329
rect 6734 18255 6790 18264
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6932 17134 6960 17818
rect 7208 17490 7236 24006
rect 7286 23352 7342 23361
rect 7286 23287 7342 23296
rect 7300 20602 7328 23287
rect 7288 20596 7340 20602
rect 7288 20538 7340 20544
rect 7392 19718 7420 26250
rect 7472 23656 7524 23662
rect 7472 23598 7524 23604
rect 7484 23254 7512 23598
rect 7472 23248 7524 23254
rect 7472 23190 7524 23196
rect 7484 22642 7512 23190
rect 7472 22636 7524 22642
rect 7472 22578 7524 22584
rect 7484 22234 7512 22578
rect 7472 22228 7524 22234
rect 7472 22170 7524 22176
rect 7484 21486 7512 22170
rect 7472 21480 7524 21486
rect 7472 21422 7524 21428
rect 7576 21418 7604 26438
rect 7564 21412 7616 21418
rect 7564 21354 7616 21360
rect 7668 21128 7696 27520
rect 8220 26466 8248 27520
rect 8036 26438 8248 26466
rect 7840 25152 7892 25158
rect 7840 25094 7892 25100
rect 7852 24682 7880 25094
rect 7840 24676 7892 24682
rect 7840 24618 7892 24624
rect 7748 24608 7800 24614
rect 7748 24550 7800 24556
rect 7760 24274 7788 24550
rect 7932 24336 7984 24342
rect 7930 24304 7932 24313
rect 7984 24304 7986 24313
rect 7748 24268 7800 24274
rect 7930 24239 7986 24248
rect 7748 24210 7800 24216
rect 7760 23322 7788 24210
rect 7932 23588 7984 23594
rect 7932 23530 7984 23536
rect 7748 23316 7800 23322
rect 7748 23258 7800 23264
rect 7944 23186 7972 23530
rect 7932 23180 7984 23186
rect 7932 23122 7984 23128
rect 8036 22386 8064 26438
rect 8208 26376 8260 26382
rect 8208 26318 8260 26324
rect 8116 24336 8168 24342
rect 8116 24278 8168 24284
rect 8128 23866 8156 24278
rect 8116 23860 8168 23866
rect 8116 23802 8168 23808
rect 8116 23248 8168 23254
rect 8116 23190 8168 23196
rect 8128 22710 8156 23190
rect 8116 22704 8168 22710
rect 8114 22672 8116 22681
rect 8168 22672 8170 22681
rect 8114 22607 8170 22616
rect 7760 22358 8064 22386
rect 7760 22098 7788 22358
rect 7838 22264 7894 22273
rect 7838 22199 7894 22208
rect 7748 22092 7800 22098
rect 7748 22034 7800 22040
rect 7748 21412 7800 21418
rect 7748 21354 7800 21360
rect 7484 21100 7696 21128
rect 7380 19712 7432 19718
rect 7380 19654 7432 19660
rect 7380 19236 7432 19242
rect 7380 19178 7432 19184
rect 7208 17462 7328 17490
rect 7196 17332 7248 17338
rect 7196 17274 7248 17280
rect 6920 17128 6972 17134
rect 6920 17070 6972 17076
rect 6932 16794 6960 17070
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 6736 16448 6788 16454
rect 6736 16390 6788 16396
rect 7104 16448 7156 16454
rect 7104 16390 7156 16396
rect 6748 16114 6776 16390
rect 6736 16108 6788 16114
rect 6736 16050 6788 16056
rect 6644 16040 6696 16046
rect 6644 15982 6696 15988
rect 6656 15706 6684 15982
rect 6748 15722 6776 16050
rect 7024 15910 7052 15941
rect 6828 15904 6880 15910
rect 7012 15904 7064 15910
rect 6880 15864 6960 15892
rect 6828 15846 6880 15852
rect 6644 15700 6696 15706
rect 6748 15694 6868 15722
rect 6644 15642 6696 15648
rect 6840 15042 6868 15694
rect 6932 15162 6960 15864
rect 7010 15872 7012 15881
rect 7064 15872 7066 15881
rect 7010 15807 7066 15816
rect 7024 15706 7052 15807
rect 7012 15700 7064 15706
rect 7012 15642 7064 15648
rect 7116 15570 7144 16390
rect 7104 15564 7156 15570
rect 7104 15506 7156 15512
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 6840 15014 6960 15042
rect 6736 14952 6788 14958
rect 6736 14894 6788 14900
rect 6550 14648 6606 14657
rect 5080 14612 5132 14618
rect 5080 14554 5132 14560
rect 5540 14612 5592 14618
rect 6550 14583 6606 14592
rect 5540 14554 5592 14560
rect 6644 14340 6696 14346
rect 6644 14282 6696 14288
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 6656 14074 6684 14282
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 5632 13932 5684 13938
rect 5632 13874 5684 13880
rect 5540 13864 5592 13870
rect 5644 13841 5672 13874
rect 5540 13806 5592 13812
rect 5630 13832 5686 13841
rect 5552 13546 5580 13806
rect 6748 13802 6776 14894
rect 6932 14074 6960 15014
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 7024 13954 7052 15098
rect 7116 14890 7144 15506
rect 7104 14884 7156 14890
rect 7104 14826 7156 14832
rect 7116 14482 7144 14826
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 6932 13926 7052 13954
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 5630 13767 5686 13776
rect 6736 13796 6788 13802
rect 6736 13738 6788 13744
rect 5632 13728 5684 13734
rect 5630 13696 5632 13705
rect 5684 13696 5686 13705
rect 5630 13631 5686 13640
rect 5460 13530 5580 13546
rect 5448 13524 5580 13530
rect 5500 13518 5580 13524
rect 5814 13560 5870 13569
rect 6840 13530 6868 13806
rect 5814 13495 5870 13504
rect 6828 13524 6880 13530
rect 5448 13466 5500 13472
rect 5356 13320 5408 13326
rect 5356 13262 5408 13268
rect 5172 12844 5224 12850
rect 5172 12786 5224 12792
rect 5184 12753 5212 12786
rect 5170 12744 5226 12753
rect 5170 12679 5226 12688
rect 5368 12646 5396 13262
rect 5460 12850 5488 13466
rect 5828 13462 5856 13495
rect 6828 13466 6880 13472
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5816 13456 5868 13462
rect 5816 13398 5868 13404
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 5356 12640 5408 12646
rect 5356 12582 5408 12588
rect 5460 12306 5488 12786
rect 5552 12345 5580 13398
rect 5828 13274 5856 13398
rect 5828 13246 6040 13274
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6012 12986 6040 13246
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 6012 12866 6040 12922
rect 6828 12912 6880 12918
rect 6012 12838 6224 12866
rect 6828 12854 6880 12860
rect 6092 12640 6144 12646
rect 6092 12582 6144 12588
rect 5538 12336 5594 12345
rect 5448 12300 5500 12306
rect 5538 12271 5594 12280
rect 5448 12242 5500 12248
rect 5460 11762 5488 12242
rect 6000 12232 6052 12238
rect 5998 12200 6000 12209
rect 6052 12200 6054 12209
rect 5998 12135 6054 12144
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 6104 11898 6132 12582
rect 6092 11892 6144 11898
rect 6092 11834 6144 11840
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 4988 11688 5040 11694
rect 4988 11630 5040 11636
rect 5000 11286 5028 11630
rect 5356 11552 5408 11558
rect 5354 11520 5356 11529
rect 5408 11520 5410 11529
rect 5354 11455 5410 11464
rect 5460 11354 5488 11698
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 4988 11280 5040 11286
rect 4988 11222 5040 11228
rect 5540 11076 5592 11082
rect 5460 11036 5540 11064
rect 5172 11008 5224 11014
rect 5172 10950 5224 10956
rect 5184 10674 5212 10950
rect 5172 10668 5224 10674
rect 5172 10610 5224 10616
rect 5184 10198 5212 10610
rect 5460 10606 5488 11036
rect 5540 11018 5592 11024
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 5172 10192 5224 10198
rect 5172 10134 5224 10140
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 4710 9650 4766 9659
rect 4710 9585 4766 9594
rect 4816 9110 4844 9998
rect 5184 9722 5212 10134
rect 5460 9926 5488 10406
rect 6196 10266 6224 12838
rect 6734 12064 6790 12073
rect 6734 11999 6790 12008
rect 6460 11892 6512 11898
rect 6460 11834 6512 11840
rect 6472 11354 6500 11834
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6656 11218 6684 11494
rect 6276 11212 6328 11218
rect 6276 11154 6328 11160
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6184 10260 6236 10266
rect 6184 10202 6236 10208
rect 5448 9920 5500 9926
rect 5448 9862 5500 9868
rect 5172 9716 5224 9722
rect 5172 9658 5224 9664
rect 4894 9616 4950 9625
rect 4894 9551 4950 9560
rect 4804 9104 4856 9110
rect 4804 9046 4856 9052
rect 4908 6934 4936 9551
rect 5184 9178 5212 9658
rect 5172 9172 5224 9178
rect 5172 9114 5224 9120
rect 5460 7818 5488 9862
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 6092 9512 6144 9518
rect 6092 9454 6144 9460
rect 6104 8974 6132 9454
rect 6288 9382 6316 11154
rect 6552 11144 6604 11150
rect 6552 11086 6604 11092
rect 6564 10810 6592 11086
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6458 9752 6514 9761
rect 6458 9687 6514 9696
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 6104 8430 6132 8910
rect 6196 8634 6224 8978
rect 6288 8634 6316 9318
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6092 8424 6144 8430
rect 6092 8366 6144 8372
rect 6472 7886 6500 9687
rect 6748 8090 6776 11999
rect 6840 11898 6868 12854
rect 6828 11892 6880 11898
rect 6828 11834 6880 11840
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 6840 9722 6868 10746
rect 6932 10033 6960 13926
rect 7116 13530 7144 14418
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 7012 12640 7064 12646
rect 7012 12582 7064 12588
rect 7024 12102 7052 12582
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 7024 11082 7052 12038
rect 7208 11937 7236 17274
rect 7300 15065 7328 17462
rect 7392 16289 7420 19178
rect 7378 16280 7434 16289
rect 7378 16215 7434 16224
rect 7380 16176 7432 16182
rect 7380 16118 7432 16124
rect 7286 15056 7342 15065
rect 7286 14991 7342 15000
rect 7392 14890 7420 16118
rect 7484 15201 7512 21100
rect 7656 21004 7708 21010
rect 7656 20946 7708 20952
rect 7562 20496 7618 20505
rect 7562 20431 7618 20440
rect 7576 19961 7604 20431
rect 7668 20398 7696 20946
rect 7656 20392 7708 20398
rect 7656 20334 7708 20340
rect 7562 19952 7618 19961
rect 7562 19887 7618 19896
rect 7564 19712 7616 19718
rect 7564 19654 7616 19660
rect 7576 19174 7604 19654
rect 7656 19372 7708 19378
rect 7656 19314 7708 19320
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 7470 15192 7526 15201
rect 7470 15127 7526 15136
rect 7380 14884 7432 14890
rect 7380 14826 7432 14832
rect 7472 14884 7524 14890
rect 7472 14826 7524 14832
rect 7378 14784 7434 14793
rect 7378 14719 7434 14728
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7300 13938 7328 14214
rect 7288 13932 7340 13938
rect 7288 13874 7340 13880
rect 7392 13818 7420 14719
rect 7484 14618 7512 14826
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 7484 13870 7512 14554
rect 7300 13790 7420 13818
rect 7472 13864 7524 13870
rect 7472 13806 7524 13812
rect 7300 12374 7328 13790
rect 7576 13682 7604 19110
rect 7668 18970 7696 19314
rect 7656 18964 7708 18970
rect 7656 18906 7708 18912
rect 7654 17096 7710 17105
rect 7654 17031 7710 17040
rect 7392 13654 7604 13682
rect 7288 12368 7340 12374
rect 7288 12310 7340 12316
rect 7194 11928 7250 11937
rect 7300 11898 7328 12310
rect 7392 12306 7420 13654
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7484 12238 7512 12786
rect 7668 12288 7696 17031
rect 7760 12646 7788 21354
rect 7852 20913 7880 22199
rect 7932 22160 7984 22166
rect 7932 22102 7984 22108
rect 8116 22160 8168 22166
rect 8220 22148 8248 26318
rect 8576 25696 8628 25702
rect 8576 25638 8628 25644
rect 8392 25424 8444 25430
rect 8392 25366 8444 25372
rect 8404 24954 8432 25366
rect 8484 25288 8536 25294
rect 8484 25230 8536 25236
rect 8392 24948 8444 24954
rect 8392 24890 8444 24896
rect 8404 24857 8432 24890
rect 8496 24886 8524 25230
rect 8484 24880 8536 24886
rect 8390 24848 8446 24857
rect 8484 24822 8536 24828
rect 8390 24783 8446 24792
rect 8300 24676 8352 24682
rect 8300 24618 8352 24624
rect 8312 24410 8340 24618
rect 8300 24404 8352 24410
rect 8300 24346 8352 24352
rect 8312 23848 8340 24346
rect 8404 24041 8432 24783
rect 8390 24032 8446 24041
rect 8390 23967 8446 23976
rect 8392 23860 8444 23866
rect 8312 23820 8392 23848
rect 8392 23802 8444 23808
rect 8404 22506 8432 23802
rect 8496 23769 8524 24822
rect 8588 24342 8616 25638
rect 8772 25294 8800 27520
rect 8760 25288 8812 25294
rect 8760 25230 8812 25236
rect 8576 24336 8628 24342
rect 8576 24278 8628 24284
rect 8482 23760 8538 23769
rect 8482 23695 8538 23704
rect 8588 23338 8616 24278
rect 8588 23310 8892 23338
rect 8576 23248 8628 23254
rect 8576 23190 8628 23196
rect 8588 22953 8616 23190
rect 8668 23112 8720 23118
rect 8668 23054 8720 23060
rect 8574 22944 8630 22953
rect 8574 22879 8630 22888
rect 8588 22778 8616 22879
rect 8576 22772 8628 22778
rect 8576 22714 8628 22720
rect 8392 22500 8444 22506
rect 8392 22442 8444 22448
rect 8404 22234 8432 22442
rect 8392 22228 8444 22234
rect 8392 22170 8444 22176
rect 8168 22120 8248 22148
rect 8116 22102 8168 22108
rect 7944 21146 7972 22102
rect 8024 22092 8076 22098
rect 8024 22034 8076 22040
rect 7932 21140 7984 21146
rect 7932 21082 7984 21088
rect 7838 20904 7894 20913
rect 7838 20839 7894 20848
rect 7840 18148 7892 18154
rect 7840 18090 7892 18096
rect 7852 17814 7880 18090
rect 7840 17808 7892 17814
rect 7838 17776 7840 17785
rect 7892 17776 7894 17785
rect 7838 17711 7894 17720
rect 7840 15360 7892 15366
rect 7840 15302 7892 15308
rect 7852 13734 7880 15302
rect 7840 13728 7892 13734
rect 7840 13670 7892 13676
rect 7852 13530 7880 13670
rect 7840 13524 7892 13530
rect 7840 13466 7892 13472
rect 7748 12640 7800 12646
rect 7748 12582 7800 12588
rect 7576 12260 7696 12288
rect 7748 12300 7800 12306
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7194 11863 7250 11872
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7484 11694 7512 12038
rect 7472 11688 7524 11694
rect 7472 11630 7524 11636
rect 7102 11520 7158 11529
rect 7102 11455 7158 11464
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 7010 10976 7066 10985
rect 7010 10911 7066 10920
rect 7024 10810 7052 10911
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 7116 10674 7144 11455
rect 7576 11132 7604 12260
rect 7748 12242 7800 12248
rect 7656 12164 7708 12170
rect 7656 12106 7708 12112
rect 7668 11898 7696 12106
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7760 11626 7788 12242
rect 7944 11762 7972 21082
rect 8036 17338 8064 22034
rect 8116 22024 8168 22030
rect 8116 21966 8168 21972
rect 8484 22024 8536 22030
rect 8484 21966 8536 21972
rect 8128 21690 8156 21966
rect 8206 21856 8262 21865
rect 8206 21791 8262 21800
rect 8116 21684 8168 21690
rect 8116 21626 8168 21632
rect 8220 21622 8248 21791
rect 8208 21616 8260 21622
rect 8208 21558 8260 21564
rect 8496 21350 8524 21966
rect 8680 21865 8708 23054
rect 8864 22778 8892 23310
rect 8852 22772 8904 22778
rect 8852 22714 8904 22720
rect 8666 21856 8722 21865
rect 8666 21791 8722 21800
rect 9324 21706 9352 27520
rect 9772 26444 9824 26450
rect 9772 26386 9824 26392
rect 9404 25152 9456 25158
rect 9404 25094 9456 25100
rect 9416 23866 9444 25094
rect 9588 24608 9640 24614
rect 9640 24556 9720 24562
rect 9588 24550 9720 24556
rect 9600 24534 9720 24550
rect 9404 23860 9456 23866
rect 9404 23802 9456 23808
rect 9416 23662 9444 23802
rect 9404 23656 9456 23662
rect 9404 23598 9456 23604
rect 9496 23248 9548 23254
rect 9494 23216 9496 23225
rect 9548 23216 9550 23225
rect 9494 23151 9550 23160
rect 9588 23112 9640 23118
rect 9588 23054 9640 23060
rect 9494 22128 9550 22137
rect 9494 22063 9496 22072
rect 9548 22063 9550 22072
rect 9496 22034 9548 22040
rect 9494 21720 9550 21729
rect 9324 21678 9494 21706
rect 8484 21344 8536 21350
rect 8484 21286 8536 21292
rect 8496 21078 8524 21286
rect 8116 21072 8168 21078
rect 8392 21072 8444 21078
rect 8116 21014 8168 21020
rect 8390 21040 8392 21049
rect 8484 21072 8536 21078
rect 8444 21040 8446 21049
rect 8128 20602 8156 21014
rect 8484 21014 8536 21020
rect 8390 20975 8446 20984
rect 8206 20904 8262 20913
rect 8206 20839 8262 20848
rect 8116 20596 8168 20602
rect 8116 20538 8168 20544
rect 8220 19394 8248 20839
rect 8496 19990 8524 21014
rect 9324 20942 9352 21678
rect 9600 21690 9628 23054
rect 9692 21962 9720 24534
rect 9784 22234 9812 26386
rect 9772 22228 9824 22234
rect 9772 22170 9824 22176
rect 9680 21956 9732 21962
rect 9680 21898 9732 21904
rect 9494 21655 9550 21664
rect 9588 21684 9640 21690
rect 9588 21626 9640 21632
rect 9784 21350 9812 22170
rect 9680 21344 9732 21350
rect 9680 21286 9732 21292
rect 9772 21344 9824 21350
rect 9772 21286 9824 21292
rect 9312 20936 9364 20942
rect 9312 20878 9364 20884
rect 9324 20602 9352 20878
rect 9312 20596 9364 20602
rect 9312 20538 9364 20544
rect 9402 20496 9458 20505
rect 9402 20431 9458 20440
rect 8758 20224 8814 20233
rect 8758 20159 8814 20168
rect 8392 19984 8444 19990
rect 8392 19926 8444 19932
rect 8484 19984 8536 19990
rect 8484 19926 8536 19932
rect 8404 19553 8432 19926
rect 8390 19544 8446 19553
rect 8496 19514 8524 19926
rect 8576 19848 8628 19854
rect 8576 19790 8628 19796
rect 8390 19479 8446 19488
rect 8484 19508 8536 19514
rect 8128 19366 8248 19394
rect 8128 19242 8156 19366
rect 8300 19304 8352 19310
rect 8220 19264 8300 19292
rect 8116 19236 8168 19242
rect 8116 19178 8168 19184
rect 8220 17610 8248 19264
rect 8300 19246 8352 19252
rect 8404 18970 8432 19479
rect 8484 19450 8536 19456
rect 8588 19394 8616 19790
rect 8496 19366 8616 19394
rect 8496 19174 8524 19366
rect 8484 19168 8536 19174
rect 8484 19110 8536 19116
rect 8392 18964 8444 18970
rect 8392 18906 8444 18912
rect 8496 18465 8524 19110
rect 8668 18624 8720 18630
rect 8668 18566 8720 18572
rect 8482 18456 8538 18465
rect 8680 18426 8708 18566
rect 8482 18391 8538 18400
rect 8668 18420 8720 18426
rect 8208 17604 8260 17610
rect 8208 17546 8260 17552
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 8208 16992 8260 16998
rect 8208 16934 8260 16940
rect 8220 16726 8248 16934
rect 8208 16720 8260 16726
rect 8208 16662 8260 16668
rect 8496 16674 8524 18391
rect 8668 18362 8720 18368
rect 8680 17882 8708 18362
rect 8668 17876 8720 17882
rect 8668 17818 8720 17824
rect 8668 17672 8720 17678
rect 8668 17614 8720 17620
rect 8680 17338 8708 17614
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 8772 16794 8800 20159
rect 9128 19712 9180 19718
rect 9128 19654 9180 19660
rect 9140 19310 9168 19654
rect 9416 19310 9444 20431
rect 9588 20256 9640 20262
rect 9586 20224 9588 20233
rect 9640 20224 9642 20233
rect 9586 20159 9642 20168
rect 9692 19990 9720 21286
rect 9876 20482 9904 27520
rect 10428 25752 10456 27520
rect 10152 25724 10456 25752
rect 9954 24576 10010 24585
rect 9954 24511 10010 24520
rect 9968 24177 9996 24511
rect 10046 24304 10102 24313
rect 10046 24239 10102 24248
rect 9954 24168 10010 24177
rect 9954 24103 10010 24112
rect 10060 23866 10088 24239
rect 10048 23860 10100 23866
rect 10048 23802 10100 23808
rect 10048 23588 10100 23594
rect 10048 23530 10100 23536
rect 9954 23488 10010 23497
rect 9954 23423 10010 23432
rect 9968 22778 9996 23423
rect 10060 23050 10088 23530
rect 10048 23044 10100 23050
rect 10048 22986 10100 22992
rect 9956 22772 10008 22778
rect 9956 22714 10008 22720
rect 10046 22264 10102 22273
rect 10046 22199 10102 22208
rect 10060 22166 10088 22199
rect 10048 22160 10100 22166
rect 10048 22102 10100 22108
rect 10048 22024 10100 22030
rect 10048 21966 10100 21972
rect 9956 21956 10008 21962
rect 9956 21898 10008 21904
rect 9968 21865 9996 21898
rect 9954 21856 10010 21865
rect 9954 21791 10010 21800
rect 9968 21146 9996 21791
rect 9956 21140 10008 21146
rect 9956 21082 10008 21088
rect 9876 20454 9996 20482
rect 9864 20392 9916 20398
rect 9864 20334 9916 20340
rect 9770 20088 9826 20097
rect 9770 20023 9772 20032
rect 9824 20023 9826 20032
rect 9772 19994 9824 20000
rect 9680 19984 9732 19990
rect 9680 19926 9732 19932
rect 9784 19514 9812 19994
rect 9876 19922 9904 20334
rect 9864 19916 9916 19922
rect 9864 19858 9916 19864
rect 9772 19508 9824 19514
rect 9772 19450 9824 19456
rect 9128 19304 9180 19310
rect 9128 19246 9180 19252
rect 9404 19304 9456 19310
rect 9404 19246 9456 19252
rect 9496 19304 9548 19310
rect 9496 19246 9548 19252
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9508 18970 9536 19246
rect 9496 18964 9548 18970
rect 9496 18906 9548 18912
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 9048 17610 9076 18566
rect 9312 18080 9364 18086
rect 9312 18022 9364 18028
rect 9324 17882 9352 18022
rect 9312 17876 9364 17882
rect 9312 17818 9364 17824
rect 9126 17776 9182 17785
rect 9126 17711 9182 17720
rect 9036 17604 9088 17610
rect 9036 17546 9088 17552
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 8760 16788 8812 16794
rect 8760 16730 8812 16736
rect 8392 16652 8444 16658
rect 8496 16646 8708 16674
rect 8392 16594 8444 16600
rect 8116 16448 8168 16454
rect 8116 16390 8168 16396
rect 8298 16416 8354 16425
rect 8024 15972 8076 15978
rect 8024 15914 8076 15920
rect 8036 15570 8064 15914
rect 8024 15564 8076 15570
rect 8024 15506 8076 15512
rect 8128 15337 8156 16390
rect 8298 16351 8354 16360
rect 8206 16280 8262 16289
rect 8206 16215 8262 16224
rect 8220 15910 8248 16215
rect 8208 15904 8260 15910
rect 8208 15846 8260 15852
rect 8312 15706 8340 16351
rect 8404 15910 8432 16594
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 8114 15328 8170 15337
rect 8114 15263 8170 15272
rect 8220 14906 8248 15438
rect 8312 15162 8340 15642
rect 8404 15609 8432 15846
rect 8390 15600 8446 15609
rect 8390 15535 8446 15544
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8298 14920 8354 14929
rect 8220 14878 8298 14906
rect 8298 14855 8300 14864
rect 8352 14855 8354 14864
rect 8300 14826 8352 14832
rect 8484 14816 8536 14822
rect 8484 14758 8536 14764
rect 8390 14648 8446 14657
rect 8390 14583 8392 14592
rect 8444 14583 8446 14592
rect 8392 14554 8444 14560
rect 8116 14544 8168 14550
rect 8116 14486 8168 14492
rect 8128 13870 8156 14486
rect 8208 14340 8260 14346
rect 8208 14282 8260 14288
rect 8220 14226 8248 14282
rect 8220 14198 8340 14226
rect 8206 14104 8262 14113
rect 8206 14039 8262 14048
rect 8116 13864 8168 13870
rect 8116 13806 8168 13812
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 8036 12918 8064 13466
rect 8024 12912 8076 12918
rect 8022 12880 8024 12889
rect 8076 12880 8078 12889
rect 8022 12815 8078 12824
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 8036 11626 8064 12174
rect 7748 11620 7800 11626
rect 7748 11562 7800 11568
rect 8024 11620 8076 11626
rect 8024 11562 8076 11568
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7668 11150 7696 11494
rect 7484 11104 7604 11132
rect 7656 11144 7708 11150
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 6918 10024 6974 10033
rect 6918 9959 6974 9968
rect 6828 9716 6880 9722
rect 6828 9658 6880 9664
rect 6840 9194 6868 9658
rect 7208 9466 7236 10950
rect 7484 10538 7512 11104
rect 7656 11086 7708 11092
rect 7668 10849 7696 11086
rect 7654 10840 7710 10849
rect 7654 10775 7710 10784
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7472 10532 7524 10538
rect 7472 10474 7524 10480
rect 7576 10266 7604 10610
rect 7654 10432 7710 10441
rect 7654 10367 7710 10376
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7576 10033 7604 10202
rect 7668 10130 7696 10367
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7562 10024 7618 10033
rect 7562 9959 7618 9968
rect 7668 9722 7696 10066
rect 7656 9716 7708 9722
rect 7656 9658 7708 9664
rect 7116 9438 7236 9466
rect 6840 9178 6960 9194
rect 6840 9172 6972 9178
rect 6840 9166 6920 9172
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 6472 7478 6500 7822
rect 6460 7472 6512 7478
rect 6460 7414 6512 7420
rect 6748 7410 6776 8026
rect 6840 8022 6868 9166
rect 6920 9114 6972 9120
rect 6828 8016 6880 8022
rect 6828 7958 6880 7964
rect 6840 7546 6868 7958
rect 7116 7857 7144 9438
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7208 8430 7236 9318
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 7208 8090 7236 8366
rect 7668 8362 7696 9658
rect 7760 8945 7788 11562
rect 8128 11558 8156 13806
rect 8220 13258 8248 14039
rect 8208 13252 8260 13258
rect 8208 13194 8260 13200
rect 8312 12850 8340 14198
rect 8392 14000 8444 14006
rect 8392 13942 8444 13948
rect 8404 13705 8432 13942
rect 8390 13696 8446 13705
rect 8390 13631 8446 13640
rect 8496 13462 8524 14758
rect 8574 14376 8630 14385
rect 8574 14311 8630 14320
rect 8484 13456 8536 13462
rect 8484 13398 8536 13404
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 8300 12708 8352 12714
rect 8300 12650 8352 12656
rect 8312 12102 8340 12650
rect 8496 12442 8524 13398
rect 8588 13297 8616 14311
rect 8574 13288 8630 13297
rect 8574 13223 8630 13232
rect 8680 13172 8708 16646
rect 8772 15706 8800 16730
rect 8942 16552 8998 16561
rect 8942 16487 8998 16496
rect 8956 16250 8984 16487
rect 8944 16244 8996 16250
rect 8944 16186 8996 16192
rect 8956 15978 8984 16186
rect 8944 15972 8996 15978
rect 8944 15914 8996 15920
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 8758 15056 8814 15065
rect 8758 14991 8814 15000
rect 8772 13870 8800 14991
rect 9048 14958 9076 16934
rect 9140 16794 9168 17711
rect 9324 17116 9352 17818
rect 9692 17762 9720 19246
rect 9784 18086 9812 19450
rect 9864 19168 9916 19174
rect 9864 19110 9916 19116
rect 9876 19009 9904 19110
rect 9862 19000 9918 19009
rect 9862 18935 9918 18944
rect 9876 18834 9904 18935
rect 9864 18828 9916 18834
rect 9864 18770 9916 18776
rect 9876 18358 9904 18770
rect 9864 18352 9916 18358
rect 9864 18294 9916 18300
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9508 17734 9720 17762
rect 9404 17128 9456 17134
rect 9324 17088 9404 17116
rect 9404 17070 9456 17076
rect 9508 16946 9536 17734
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 9588 17604 9640 17610
rect 9588 17546 9640 17552
rect 9324 16918 9536 16946
rect 9128 16788 9180 16794
rect 9128 16730 9180 16736
rect 9220 16584 9272 16590
rect 9126 16552 9182 16561
rect 9220 16526 9272 16532
rect 9126 16487 9182 16496
rect 9140 16289 9168 16487
rect 9126 16280 9182 16289
rect 9232 16250 9260 16526
rect 9126 16215 9182 16224
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 9036 14952 9088 14958
rect 9036 14894 9088 14900
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 8956 14521 8984 14554
rect 8942 14512 8998 14521
rect 8942 14447 8998 14456
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8956 13802 8984 14447
rect 9036 14272 9088 14278
rect 9036 14214 9088 14220
rect 9048 13870 9076 14214
rect 9036 13864 9088 13870
rect 9036 13806 9088 13812
rect 8944 13796 8996 13802
rect 8944 13738 8996 13744
rect 9048 13569 9076 13806
rect 9034 13560 9090 13569
rect 9034 13495 9090 13504
rect 8760 13320 8812 13326
rect 8760 13262 8812 13268
rect 8588 13144 8708 13172
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 8390 12200 8446 12209
rect 8390 12135 8446 12144
rect 8300 12096 8352 12102
rect 8300 12038 8352 12044
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 8208 11280 8260 11286
rect 8208 11222 8260 11228
rect 8220 10742 8248 11222
rect 8208 10736 8260 10742
rect 8208 10678 8260 10684
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7746 8936 7802 8945
rect 7746 8871 7802 8880
rect 7656 8356 7708 8362
rect 7656 8298 7708 8304
rect 7852 8294 7880 9862
rect 8220 9625 8248 10134
rect 8206 9616 8262 9625
rect 8206 9551 8262 9560
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7944 9178 7972 9454
rect 8220 9450 8248 9551
rect 8208 9444 8260 9450
rect 8208 9386 8260 9392
rect 7932 9172 7984 9178
rect 7932 9114 7984 9120
rect 7944 8634 7972 9114
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7840 8288 7892 8294
rect 7840 8230 7892 8236
rect 7392 8090 7420 8230
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7932 8016 7984 8022
rect 7932 7958 7984 7964
rect 7102 7848 7158 7857
rect 7102 7783 7158 7792
rect 7944 7546 7972 7958
rect 8312 7954 8340 11698
rect 8404 11354 8432 12135
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8404 10810 8432 11290
rect 8588 11014 8616 13144
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 8484 10736 8536 10742
rect 8484 10678 8536 10684
rect 8392 10532 8444 10538
rect 8392 10474 8444 10480
rect 8404 10198 8432 10474
rect 8392 10192 8444 10198
rect 8392 10134 8444 10140
rect 8404 9518 8432 10134
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 4896 6928 4948 6934
rect 4948 6876 5028 6882
rect 4896 6870 5028 6876
rect 4908 6854 5028 6870
rect 8312 6866 8340 7890
rect 8404 7546 8432 8298
rect 8496 8022 8524 10678
rect 8680 10130 8708 12582
rect 8772 12442 8800 13262
rect 9324 12753 9352 16918
rect 9496 16652 9548 16658
rect 9496 16594 9548 16600
rect 9402 16280 9458 16289
rect 9402 16215 9458 16224
rect 9416 16114 9444 16215
rect 9404 16108 9456 16114
rect 9404 16050 9456 16056
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 9416 14618 9444 15438
rect 9508 14890 9536 16594
rect 9600 16522 9628 17546
rect 9588 16516 9640 16522
rect 9588 16458 9640 16464
rect 9692 16266 9720 17614
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 9772 16720 9824 16726
rect 9772 16662 9824 16668
rect 9600 16238 9720 16266
rect 9600 16114 9628 16238
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9600 15706 9628 16050
rect 9588 15700 9640 15706
rect 9588 15642 9640 15648
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9496 14884 9548 14890
rect 9496 14826 9548 14832
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 9508 13326 9536 14826
rect 9588 14816 9640 14822
rect 9692 14770 9720 15506
rect 9784 15434 9812 16662
rect 9876 16114 9904 16730
rect 9968 16289 9996 20454
rect 9954 16280 10010 16289
rect 9954 16215 10010 16224
rect 9864 16108 9916 16114
rect 9864 16050 9916 16056
rect 9876 15502 9904 16050
rect 9956 15632 10008 15638
rect 9956 15574 10008 15580
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9772 15428 9824 15434
rect 9772 15370 9824 15376
rect 9862 15328 9918 15337
rect 9862 15263 9918 15272
rect 9640 14764 9720 14770
rect 9588 14758 9720 14764
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 9600 14742 9720 14758
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9310 12744 9366 12753
rect 9310 12679 9366 12688
rect 8760 12436 8812 12442
rect 8760 12378 8812 12384
rect 8944 12368 8996 12374
rect 8944 12310 8996 12316
rect 8852 11688 8904 11694
rect 8852 11630 8904 11636
rect 8864 10266 8892 11630
rect 8956 11354 8984 12310
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 9140 11626 9168 12038
rect 9220 11824 9272 11830
rect 9220 11766 9272 11772
rect 9128 11620 9180 11626
rect 9128 11562 9180 11568
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 8956 10810 8984 11290
rect 9048 11218 9076 11494
rect 9036 11212 9088 11218
rect 9036 11154 9088 11160
rect 8944 10804 8996 10810
rect 8944 10746 8996 10752
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 8668 10124 8720 10130
rect 8668 10066 8720 10072
rect 9140 9636 9168 11562
rect 9232 9761 9260 11766
rect 9600 11642 9628 13126
rect 9692 12238 9720 14742
rect 9784 12753 9812 14758
rect 9876 14618 9904 15263
rect 9968 14822 9996 15574
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9876 13530 9904 14554
rect 9864 13524 9916 13530
rect 9864 13466 9916 13472
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 9770 12744 9826 12753
rect 9770 12679 9826 12688
rect 9876 12594 9904 13262
rect 9784 12566 9904 12594
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9680 12096 9732 12102
rect 9678 12064 9680 12073
rect 9732 12064 9734 12073
rect 9678 11999 9734 12008
rect 9600 11614 9720 11642
rect 9692 11558 9720 11614
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9692 10985 9720 11494
rect 9678 10976 9734 10985
rect 9678 10911 9734 10920
rect 9784 9874 9812 12566
rect 10060 12424 10088 21966
rect 10152 19972 10180 25724
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10692 25356 10744 25362
rect 10692 25298 10744 25304
rect 10600 25220 10652 25226
rect 10600 25162 10652 25168
rect 10612 24818 10640 25162
rect 10600 24812 10652 24818
rect 10600 24754 10652 24760
rect 10704 24682 10732 25298
rect 10888 24834 10916 27520
rect 11336 25356 11388 25362
rect 11336 25298 11388 25304
rect 11348 25265 11376 25298
rect 11334 25256 11390 25265
rect 11334 25191 11390 25200
rect 11336 25152 11388 25158
rect 11336 25094 11388 25100
rect 10796 24806 10916 24834
rect 11348 24818 11376 25094
rect 10968 24812 11020 24818
rect 10692 24676 10744 24682
rect 10692 24618 10744 24624
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10600 23180 10652 23186
rect 10600 23122 10652 23128
rect 10612 22778 10640 23122
rect 10600 22772 10652 22778
rect 10600 22714 10652 22720
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10232 22024 10284 22030
rect 10232 21966 10284 21972
rect 10244 21842 10272 21966
rect 10414 21856 10470 21865
rect 10244 21814 10414 21842
rect 10414 21791 10470 21800
rect 10428 21690 10456 21791
rect 10704 21690 10732 24618
rect 10796 22098 10824 24806
rect 10968 24754 11020 24760
rect 11336 24812 11388 24818
rect 11336 24754 11388 24760
rect 10876 24676 10928 24682
rect 10876 24618 10928 24624
rect 10888 24410 10916 24618
rect 10876 24404 10928 24410
rect 10876 24346 10928 24352
rect 10876 23656 10928 23662
rect 10876 23598 10928 23604
rect 10888 23186 10916 23598
rect 10980 23474 11008 24754
rect 11060 24200 11112 24206
rect 11060 24142 11112 24148
rect 11072 23662 11100 24142
rect 11060 23656 11112 23662
rect 11060 23598 11112 23604
rect 10980 23446 11100 23474
rect 10966 23352 11022 23361
rect 10966 23287 11022 23296
rect 10876 23180 10928 23186
rect 10876 23122 10928 23128
rect 10876 22976 10928 22982
rect 10876 22918 10928 22924
rect 10784 22092 10836 22098
rect 10784 22034 10836 22040
rect 10784 21888 10836 21894
rect 10784 21830 10836 21836
rect 10416 21684 10468 21690
rect 10416 21626 10468 21632
rect 10692 21684 10744 21690
rect 10692 21626 10744 21632
rect 10796 21554 10824 21830
rect 10784 21548 10836 21554
rect 10784 21490 10836 21496
rect 10888 21418 10916 22918
rect 10980 22778 11008 23287
rect 11072 23225 11100 23446
rect 11152 23248 11204 23254
rect 11058 23216 11114 23225
rect 11152 23190 11204 23196
rect 11058 23151 11114 23160
rect 10968 22772 11020 22778
rect 10968 22714 11020 22720
rect 10968 22636 11020 22642
rect 10968 22578 11020 22584
rect 10980 22030 11008 22578
rect 11072 22574 11100 23151
rect 11060 22568 11112 22574
rect 11060 22510 11112 22516
rect 11164 22234 11192 23190
rect 11242 23080 11298 23089
rect 11242 23015 11298 23024
rect 11256 22409 11284 23015
rect 11336 22704 11388 22710
rect 11336 22646 11388 22652
rect 11348 22438 11376 22646
rect 11336 22432 11388 22438
rect 11242 22400 11298 22409
rect 11336 22374 11388 22380
rect 11242 22335 11298 22344
rect 11152 22228 11204 22234
rect 11152 22170 11204 22176
rect 11348 22137 11376 22374
rect 11334 22128 11390 22137
rect 11334 22063 11390 22072
rect 10968 22024 11020 22030
rect 10968 21966 11020 21972
rect 11152 22024 11204 22030
rect 11152 21966 11204 21972
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 10876 21412 10928 21418
rect 10876 21354 10928 21360
rect 10692 21344 10744 21350
rect 10692 21286 10744 21292
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10324 20800 10376 20806
rect 10324 20742 10376 20748
rect 10336 20641 10364 20742
rect 10322 20632 10378 20641
rect 10322 20567 10378 20576
rect 10336 20330 10364 20567
rect 10324 20324 10376 20330
rect 10324 20266 10376 20272
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10152 19944 10272 19972
rect 10140 19848 10192 19854
rect 10140 19790 10192 19796
rect 10152 18970 10180 19790
rect 10244 19242 10272 19944
rect 10704 19666 10732 21286
rect 10784 21072 10836 21078
rect 10784 21014 10836 21020
rect 10796 20262 10824 21014
rect 10784 20256 10836 20262
rect 10784 20198 10836 20204
rect 10888 19786 10916 21354
rect 11072 21350 11100 21830
rect 11060 21344 11112 21350
rect 10980 21304 11060 21332
rect 10876 19780 10928 19786
rect 10876 19722 10928 19728
rect 10704 19638 10916 19666
rect 10782 19272 10838 19281
rect 10232 19236 10284 19242
rect 10782 19207 10838 19216
rect 10232 19178 10284 19184
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10796 18970 10824 19207
rect 10140 18964 10192 18970
rect 10140 18906 10192 18912
rect 10784 18964 10836 18970
rect 10784 18906 10836 18912
rect 10796 18426 10824 18906
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 10690 18184 10746 18193
rect 10690 18119 10692 18128
rect 10744 18119 10746 18128
rect 10784 18148 10836 18154
rect 10692 18090 10744 18096
rect 10784 18090 10836 18096
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10796 17882 10824 18090
rect 10784 17876 10836 17882
rect 10784 17818 10836 17824
rect 10784 17672 10836 17678
rect 10784 17614 10836 17620
rect 10140 17128 10192 17134
rect 10140 17070 10192 17076
rect 10152 16590 10180 17070
rect 10796 16998 10824 17614
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10152 16250 10180 16526
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10784 15972 10836 15978
rect 10784 15914 10836 15920
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10692 15360 10744 15366
rect 10796 15337 10824 15914
rect 10692 15302 10744 15308
rect 10782 15328 10838 15337
rect 10138 15192 10194 15201
rect 10138 15127 10140 15136
rect 10192 15127 10194 15136
rect 10140 15098 10192 15104
rect 10152 14006 10180 15098
rect 10704 14890 10732 15302
rect 10782 15263 10838 15272
rect 10692 14884 10744 14890
rect 10692 14826 10744 14832
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 10244 14113 10272 14418
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 10230 14104 10286 14113
rect 10520 14074 10548 14350
rect 10230 14039 10286 14048
rect 10508 14068 10560 14074
rect 10508 14010 10560 14016
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 10152 13734 10180 13942
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 10782 13696 10838 13705
rect 10289 13628 10585 13648
rect 10782 13631 10838 13640
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10692 13456 10744 13462
rect 10692 13398 10744 13404
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 10140 13184 10192 13190
rect 10140 13126 10192 13132
rect 9968 12396 10088 12424
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 9876 11558 9904 12174
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9692 9846 9812 9874
rect 9218 9752 9274 9761
rect 9692 9738 9720 9846
rect 9218 9687 9274 9696
rect 9600 9710 9720 9738
rect 9140 9608 9260 9636
rect 9232 9382 9260 9608
rect 9496 9444 9548 9450
rect 9496 9386 9548 9392
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 9232 8498 9260 9318
rect 9508 9178 9536 9386
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 9324 8634 9352 8774
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9496 8356 9548 8362
rect 9496 8298 9548 8304
rect 9508 8022 9536 8298
rect 8484 8016 8536 8022
rect 8484 7958 8536 7964
rect 9496 8016 9548 8022
rect 9496 7958 9548 7964
rect 8668 7880 8720 7886
rect 8666 7848 8668 7857
rect 8720 7848 8722 7857
rect 8666 7783 8722 7792
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8404 7274 8432 7482
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 8392 7268 8444 7274
rect 8392 7210 8444 7216
rect 8496 7002 8524 7346
rect 8680 7342 8708 7783
rect 9600 7410 9628 9710
rect 9876 9081 9904 11494
rect 9968 10674 9996 12396
rect 10152 12322 10180 13126
rect 10612 12782 10640 13262
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 10704 12646 10732 13398
rect 10796 13161 10824 13631
rect 10782 13152 10838 13161
rect 10782 13087 10838 13096
rect 10888 12866 10916 19638
rect 10980 19514 11008 21304
rect 11060 21286 11112 21292
rect 11164 21010 11192 21966
rect 11242 21448 11298 21457
rect 11242 21383 11298 21392
rect 11152 21004 11204 21010
rect 11152 20946 11204 20952
rect 11256 20913 11284 21383
rect 11242 20904 11298 20913
rect 11242 20839 11298 20848
rect 11058 20360 11114 20369
rect 11058 20295 11114 20304
rect 11072 19825 11100 20295
rect 11336 20256 11388 20262
rect 11336 20198 11388 20204
rect 11150 20088 11206 20097
rect 11150 20023 11206 20032
rect 11058 19816 11114 19825
rect 11058 19751 11114 19760
rect 11164 19689 11192 20023
rect 11348 19718 11376 20198
rect 11336 19712 11388 19718
rect 11150 19680 11206 19689
rect 11336 19654 11388 19660
rect 11150 19615 11206 19624
rect 10968 19508 11020 19514
rect 10968 19450 11020 19456
rect 10966 19408 11022 19417
rect 11348 19378 11376 19654
rect 10966 19343 11022 19352
rect 11336 19372 11388 19378
rect 10980 19310 11008 19343
rect 11336 19314 11388 19320
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 11058 19272 11114 19281
rect 11058 19207 11114 19216
rect 11152 19236 11204 19242
rect 10968 18760 11020 18766
rect 10968 18702 11020 18708
rect 10980 17542 11008 18702
rect 11072 18329 11100 19207
rect 11152 19178 11204 19184
rect 11058 18320 11114 18329
rect 11058 18255 11114 18264
rect 11060 17740 11112 17746
rect 11060 17682 11112 17688
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 11072 17338 11100 17682
rect 11060 17332 11112 17338
rect 11060 17274 11112 17280
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 10980 15706 11008 16594
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 11164 15065 11192 19178
rect 11348 18970 11376 19314
rect 11336 18964 11388 18970
rect 11336 18906 11388 18912
rect 11336 16448 11388 16454
rect 11336 16390 11388 16396
rect 11348 15910 11376 16390
rect 11336 15904 11388 15910
rect 11336 15846 11388 15852
rect 11348 15065 11376 15846
rect 11440 15162 11468 27520
rect 11992 24834 12020 27520
rect 11612 24812 11664 24818
rect 11612 24754 11664 24760
rect 11808 24806 12020 24834
rect 12544 24834 12572 27520
rect 12900 25764 12952 25770
rect 12900 25706 12952 25712
rect 12912 25498 12940 25706
rect 12900 25492 12952 25498
rect 12900 25434 12952 25440
rect 13096 25106 13124 27520
rect 12912 25078 13124 25106
rect 12714 24848 12770 24857
rect 12544 24806 12664 24834
rect 11624 24410 11652 24754
rect 11704 24676 11756 24682
rect 11704 24618 11756 24624
rect 11612 24404 11664 24410
rect 11612 24346 11664 24352
rect 11520 24336 11572 24342
rect 11520 24278 11572 24284
rect 11532 23526 11560 24278
rect 11520 23520 11572 23526
rect 11518 23488 11520 23497
rect 11572 23488 11574 23497
rect 11518 23423 11574 23432
rect 11624 23254 11652 24346
rect 11612 23248 11664 23254
rect 11612 23190 11664 23196
rect 11716 23066 11744 24618
rect 11532 23038 11744 23066
rect 11532 17921 11560 23038
rect 11610 22808 11666 22817
rect 11610 22743 11666 22752
rect 11624 22438 11652 22743
rect 11612 22432 11664 22438
rect 11612 22374 11664 22380
rect 11624 19310 11652 22374
rect 11704 22092 11756 22098
rect 11704 22034 11756 22040
rect 11716 21078 11744 22034
rect 11704 21072 11756 21078
rect 11704 21014 11756 21020
rect 11612 19304 11664 19310
rect 11612 19246 11664 19252
rect 11704 18896 11756 18902
rect 11702 18864 11704 18873
rect 11756 18864 11758 18873
rect 11702 18799 11758 18808
rect 11704 18352 11756 18358
rect 11704 18294 11756 18300
rect 11518 17912 11574 17921
rect 11518 17847 11574 17856
rect 11716 17785 11744 18294
rect 11702 17776 11758 17785
rect 11702 17711 11758 17720
rect 11518 15600 11574 15609
rect 11518 15535 11574 15544
rect 11428 15156 11480 15162
rect 11428 15098 11480 15104
rect 11150 15056 11206 15065
rect 11072 15014 11150 15042
rect 10966 14784 11022 14793
rect 10966 14719 11022 14728
rect 10980 14346 11008 14719
rect 10968 14340 11020 14346
rect 10968 14282 11020 14288
rect 11072 14006 11100 15014
rect 11150 14991 11206 15000
rect 11334 15056 11390 15065
rect 11334 14991 11390 15000
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 11256 14414 11284 14758
rect 11440 14532 11468 15098
rect 11348 14504 11468 14532
rect 11244 14408 11296 14414
rect 11244 14350 11296 14356
rect 11152 14272 11204 14278
rect 11152 14214 11204 14220
rect 10968 14000 11020 14006
rect 10968 13942 11020 13948
rect 11060 14000 11112 14006
rect 11060 13942 11112 13948
rect 10980 13002 11008 13942
rect 11164 13938 11192 14214
rect 11152 13932 11204 13938
rect 11152 13874 11204 13880
rect 11164 13530 11192 13874
rect 11348 13870 11376 14504
rect 11336 13864 11388 13870
rect 11336 13806 11388 13812
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 10980 12974 11284 13002
rect 10888 12838 11008 12866
rect 10784 12776 10836 12782
rect 10784 12718 10836 12724
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10060 12306 10180 12322
rect 10048 12300 10180 12306
rect 10100 12294 10180 12300
rect 10048 12242 10100 12248
rect 10060 11082 10088 12242
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10336 11626 10364 12174
rect 10704 12102 10732 12582
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10704 11665 10732 12038
rect 10690 11656 10746 11665
rect 10324 11620 10376 11626
rect 10690 11591 10746 11600
rect 10324 11562 10376 11568
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10796 11354 10824 12718
rect 10876 12708 10928 12714
rect 10876 12650 10928 12656
rect 10888 12481 10916 12650
rect 10874 12472 10930 12481
rect 10874 12407 10930 12416
rect 10980 12209 11008 12838
rect 11256 12442 11284 12974
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 10966 12200 11022 12209
rect 10966 12135 11022 12144
rect 10876 11824 10928 11830
rect 10876 11766 10928 11772
rect 10888 11354 10916 11766
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 10232 11280 10284 11286
rect 10232 11222 10284 11228
rect 10244 11121 10272 11222
rect 10324 11144 10376 11150
rect 10230 11112 10286 11121
rect 10048 11076 10100 11082
rect 10048 11018 10100 11024
rect 10152 11070 10230 11098
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 9954 10568 10010 10577
rect 9954 10503 10010 10512
rect 10048 10532 10100 10538
rect 9968 10470 9996 10503
rect 10048 10474 10100 10480
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9968 10130 9996 10406
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 10060 9926 10088 10474
rect 10152 10266 10180 11070
rect 10324 11086 10376 11092
rect 10230 11047 10286 11056
rect 10336 10538 10364 11086
rect 10796 10810 10824 11290
rect 10980 10826 11008 12135
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 11164 11082 11192 11698
rect 11256 11626 11284 12378
rect 11244 11620 11296 11626
rect 11244 11562 11296 11568
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 11152 11076 11204 11082
rect 11152 11018 11204 11024
rect 10980 10810 11100 10826
rect 10784 10804 10836 10810
rect 10704 10764 10784 10792
rect 10324 10532 10376 10538
rect 10324 10474 10376 10480
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10140 10260 10192 10266
rect 10704 10248 10732 10764
rect 10980 10804 11112 10810
rect 10980 10798 11060 10804
rect 10784 10746 10836 10752
rect 11060 10746 11112 10752
rect 10876 10736 10928 10742
rect 10876 10678 10928 10684
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10140 10202 10192 10208
rect 10612 10220 10732 10248
rect 10048 9920 10100 9926
rect 10612 9897 10640 10220
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10048 9862 10100 9868
rect 10598 9888 10654 9897
rect 9956 9648 10008 9654
rect 9956 9590 10008 9596
rect 9862 9072 9918 9081
rect 9862 9007 9918 9016
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9770 7984 9826 7993
rect 9680 7948 9732 7954
rect 9770 7919 9826 7928
rect 9680 7890 9732 7896
rect 9692 7546 9720 7890
rect 9784 7818 9812 7919
rect 9772 7812 9824 7818
rect 9772 7754 9824 7760
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8680 7002 8708 7278
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 8668 6996 8720 7002
rect 8668 6938 8720 6944
rect 4804 6792 4856 6798
rect 4804 6734 4856 6740
rect 4816 6458 4844 6734
rect 5000 6458 5028 6854
rect 8300 6860 8352 6866
rect 8300 6802 8352 6808
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 9692 6474 9720 7346
rect 9876 7002 9904 8026
rect 9968 7342 9996 9590
rect 10060 9110 10088 9862
rect 10598 9823 10654 9832
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10048 9104 10100 9110
rect 10048 9046 10100 9052
rect 10060 8634 10088 9046
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 10152 8362 10180 9318
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10704 9110 10732 10066
rect 10796 10062 10824 10406
rect 10784 10056 10836 10062
rect 10784 9998 10836 10004
rect 10796 9926 10824 9998
rect 10784 9920 10836 9926
rect 10784 9862 10836 9868
rect 10692 9104 10744 9110
rect 10692 9046 10744 9052
rect 10796 9058 10824 9862
rect 10888 9450 10916 10678
rect 10968 9988 11020 9994
rect 10968 9930 11020 9936
rect 10980 9586 11008 9930
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 11072 9518 11100 9862
rect 11164 9586 11192 11018
rect 11348 10538 11376 11290
rect 11532 11257 11560 15535
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11716 14958 11744 15438
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11716 14278 11744 14894
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11716 13734 11744 14214
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11716 13394 11744 13670
rect 11808 13569 11836 24806
rect 12532 24676 12584 24682
rect 12532 24618 12584 24624
rect 12346 24032 12402 24041
rect 12346 23967 12402 23976
rect 11888 23656 11940 23662
rect 12164 23656 12216 23662
rect 11888 23598 11940 23604
rect 12162 23624 12164 23633
rect 12360 23633 12388 23967
rect 12216 23624 12218 23633
rect 11900 23526 11928 23598
rect 12162 23559 12218 23568
rect 12346 23624 12402 23633
rect 12346 23559 12402 23568
rect 11888 23520 11940 23526
rect 11888 23462 11940 23468
rect 12164 22976 12216 22982
rect 12164 22918 12216 22924
rect 12176 22506 12204 22918
rect 12254 22672 12310 22681
rect 12254 22607 12256 22616
rect 12308 22607 12310 22616
rect 12256 22578 12308 22584
rect 12346 22536 12402 22545
rect 12164 22500 12216 22506
rect 12346 22471 12402 22480
rect 12440 22500 12492 22506
rect 12164 22442 12216 22448
rect 11980 22092 12032 22098
rect 11980 22034 12032 22040
rect 11888 22024 11940 22030
rect 11888 21966 11940 21972
rect 11900 21690 11928 21966
rect 11888 21684 11940 21690
rect 11888 21626 11940 21632
rect 11900 19922 11928 21626
rect 11992 21554 12020 22034
rect 12070 21856 12126 21865
rect 12070 21791 12126 21800
rect 11980 21548 12032 21554
rect 11980 21490 12032 21496
rect 11992 21146 12020 21490
rect 11980 21140 12032 21146
rect 11980 21082 12032 21088
rect 12084 21026 12112 21791
rect 12360 21622 12388 22471
rect 12440 22442 12492 22448
rect 12348 21616 12400 21622
rect 12348 21558 12400 21564
rect 12452 21457 12480 22442
rect 12544 21690 12572 24618
rect 12636 24177 12664 24806
rect 12714 24783 12770 24792
rect 12622 24168 12678 24177
rect 12622 24103 12678 24112
rect 12728 23866 12756 24783
rect 12808 24676 12860 24682
rect 12808 24618 12860 24624
rect 12820 24138 12848 24618
rect 12808 24132 12860 24138
rect 12808 24074 12860 24080
rect 12716 23860 12768 23866
rect 12716 23802 12768 23808
rect 12912 23746 12940 25078
rect 13084 24948 13136 24954
rect 13084 24890 13136 24896
rect 12990 24168 13046 24177
rect 12990 24103 13046 24112
rect 12728 23718 12940 23746
rect 12624 22636 12676 22642
rect 12624 22578 12676 22584
rect 12636 22545 12664 22578
rect 12622 22536 12678 22545
rect 12622 22471 12678 22480
rect 12532 21684 12584 21690
rect 12532 21626 12584 21632
rect 12438 21448 12494 21457
rect 12438 21383 12494 21392
rect 12624 21344 12676 21350
rect 12624 21286 12676 21292
rect 11992 20998 12112 21026
rect 12440 21004 12492 21010
rect 11888 19916 11940 19922
rect 11888 19858 11940 19864
rect 11900 19514 11928 19858
rect 11888 19508 11940 19514
rect 11888 19450 11940 19456
rect 11992 19394 12020 20998
rect 12360 20964 12440 20992
rect 12164 20936 12216 20942
rect 12164 20878 12216 20884
rect 12176 20398 12204 20878
rect 12360 20602 12388 20964
rect 12440 20946 12492 20952
rect 12440 20868 12492 20874
rect 12440 20810 12492 20816
rect 12348 20596 12400 20602
rect 12348 20538 12400 20544
rect 12164 20392 12216 20398
rect 12164 20334 12216 20340
rect 12072 19712 12124 19718
rect 12072 19654 12124 19660
rect 11900 19366 12020 19394
rect 11794 13560 11850 13569
rect 11794 13495 11850 13504
rect 11900 13410 11928 19366
rect 12084 19242 12112 19654
rect 12452 19394 12480 20810
rect 12636 20806 12664 21286
rect 12624 20800 12676 20806
rect 12624 20742 12676 20748
rect 12176 19366 12480 19394
rect 12532 19372 12584 19378
rect 12072 19236 12124 19242
rect 12072 19178 12124 19184
rect 12084 18766 12112 19178
rect 12072 18760 12124 18766
rect 12072 18702 12124 18708
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11992 16833 12020 18566
rect 12176 18426 12204 19366
rect 12532 19314 12584 19320
rect 12544 18902 12572 19314
rect 12636 18970 12664 20742
rect 12728 19825 12756 23718
rect 12808 23316 12860 23322
rect 12808 23258 12860 23264
rect 12820 21078 12848 23258
rect 13004 22953 13032 24103
rect 12990 22944 13046 22953
rect 12990 22879 13046 22888
rect 12992 22568 13044 22574
rect 12992 22510 13044 22516
rect 12900 22500 12952 22506
rect 12900 22442 12952 22448
rect 12912 22166 12940 22442
rect 12900 22160 12952 22166
rect 12900 22102 12952 22108
rect 12900 21888 12952 21894
rect 12900 21830 12952 21836
rect 12808 21072 12860 21078
rect 12808 21014 12860 21020
rect 12714 19816 12770 19825
rect 12714 19751 12770 19760
rect 12728 19553 12756 19751
rect 12714 19544 12770 19553
rect 12714 19479 12770 19488
rect 12820 19242 12848 21014
rect 12808 19236 12860 19242
rect 12808 19178 12860 19184
rect 12820 18970 12848 19178
rect 12624 18964 12676 18970
rect 12624 18906 12676 18912
rect 12808 18964 12860 18970
rect 12808 18906 12860 18912
rect 12348 18896 12400 18902
rect 12348 18838 12400 18844
rect 12532 18896 12584 18902
rect 12532 18838 12584 18844
rect 12256 18692 12308 18698
rect 12256 18634 12308 18640
rect 12164 18420 12216 18426
rect 12164 18362 12216 18368
rect 12164 18148 12216 18154
rect 12164 18090 12216 18096
rect 12176 17785 12204 18090
rect 12162 17776 12218 17785
rect 12162 17711 12218 17720
rect 12164 17536 12216 17542
rect 12164 17478 12216 17484
rect 11978 16824 12034 16833
rect 11978 16759 12034 16768
rect 11980 16516 12032 16522
rect 11980 16458 12032 16464
rect 11992 16182 12020 16458
rect 11980 16176 12032 16182
rect 11980 16118 12032 16124
rect 11992 15706 12020 16118
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 12176 15570 12204 17478
rect 12268 16726 12296 18634
rect 12360 16794 12388 18838
rect 12808 18828 12860 18834
rect 12808 18770 12860 18776
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12544 18086 12572 18702
rect 12820 18426 12848 18770
rect 12808 18420 12860 18426
rect 12808 18362 12860 18368
rect 12532 18080 12584 18086
rect 12532 18022 12584 18028
rect 12544 17542 12572 18022
rect 12912 17762 12940 21830
rect 13004 20942 13032 22510
rect 13096 21706 13124 24890
rect 13452 24744 13504 24750
rect 13452 24686 13504 24692
rect 13360 24608 13412 24614
rect 13360 24550 13412 24556
rect 13372 24410 13400 24550
rect 13360 24404 13412 24410
rect 13360 24346 13412 24352
rect 13176 24268 13228 24274
rect 13176 24210 13228 24216
rect 13188 21894 13216 24210
rect 13268 22976 13320 22982
rect 13268 22918 13320 22924
rect 13280 22642 13308 22918
rect 13268 22636 13320 22642
rect 13268 22578 13320 22584
rect 13176 21888 13228 21894
rect 13176 21830 13228 21836
rect 13096 21678 13216 21706
rect 13084 21412 13136 21418
rect 13084 21354 13136 21360
rect 12992 20936 13044 20942
rect 12992 20878 13044 20884
rect 13004 18970 13032 20878
rect 13096 20806 13124 21354
rect 13084 20800 13136 20806
rect 13084 20742 13136 20748
rect 12992 18964 13044 18970
rect 12992 18906 13044 18912
rect 13004 18222 13032 18906
rect 13084 18692 13136 18698
rect 13084 18634 13136 18640
rect 12992 18216 13044 18222
rect 12992 18158 13044 18164
rect 12728 17734 12940 17762
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12544 17066 12572 17478
rect 12532 17060 12584 17066
rect 12532 17002 12584 17008
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12256 16720 12308 16726
rect 12256 16662 12308 16668
rect 12544 16130 12572 17002
rect 12360 16114 12572 16130
rect 12348 16108 12572 16114
rect 12400 16102 12572 16108
rect 12348 16050 12400 16056
rect 12348 15904 12400 15910
rect 12400 15864 12572 15892
rect 12728 15881 12756 17734
rect 12806 17640 12862 17649
rect 12806 17575 12862 17584
rect 12348 15846 12400 15852
rect 12164 15564 12216 15570
rect 12164 15506 12216 15512
rect 12440 15496 12492 15502
rect 12440 15438 12492 15444
rect 12254 15328 12310 15337
rect 12254 15263 12310 15272
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 12176 14074 12204 14418
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11808 13382 11928 13410
rect 11716 12646 11744 13330
rect 11704 12640 11756 12646
rect 11704 12582 11756 12588
rect 11610 12336 11666 12345
rect 11610 12271 11666 12280
rect 11624 11626 11652 12271
rect 11716 12102 11744 12582
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11808 12050 11836 13382
rect 12070 12336 12126 12345
rect 12070 12271 12126 12280
rect 12164 12300 12216 12306
rect 11716 11694 11744 12038
rect 11808 12022 12020 12050
rect 11794 11928 11850 11937
rect 11794 11863 11796 11872
rect 11848 11863 11850 11872
rect 11796 11834 11848 11840
rect 11704 11688 11756 11694
rect 11704 11630 11756 11636
rect 11612 11620 11664 11626
rect 11612 11562 11664 11568
rect 11518 11248 11574 11257
rect 11518 11183 11574 11192
rect 11716 11150 11744 11630
rect 11796 11348 11848 11354
rect 11796 11290 11848 11296
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11336 10532 11388 10538
rect 11336 10474 11388 10480
rect 11242 10296 11298 10305
rect 11242 10231 11298 10240
rect 11256 10033 11284 10231
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 11242 10024 11298 10033
rect 11242 9959 11298 9968
rect 11348 9926 11376 10066
rect 11612 10056 11664 10062
rect 11612 9998 11664 10004
rect 11336 9920 11388 9926
rect 11336 9862 11388 9868
rect 11624 9625 11652 9998
rect 11716 9994 11744 11086
rect 11704 9988 11756 9994
rect 11704 9930 11756 9936
rect 11610 9616 11666 9625
rect 11152 9580 11204 9586
rect 11610 9551 11666 9560
rect 11152 9522 11204 9528
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 11716 9450 11744 9930
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 11704 9444 11756 9450
rect 11704 9386 11756 9392
rect 10888 9178 10916 9386
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 10796 9042 10916 9058
rect 10796 9036 10928 9042
rect 10796 9030 10876 9036
rect 10876 8978 10928 8984
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10888 8090 10916 8978
rect 11716 8838 11744 9386
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11716 8566 11744 8774
rect 11808 8634 11836 11290
rect 11886 10840 11942 10849
rect 11886 10775 11942 10784
rect 11900 10606 11928 10775
rect 11888 10600 11940 10606
rect 11888 10542 11940 10548
rect 11992 10418 12020 12022
rect 12084 11558 12112 12271
rect 12164 12242 12216 12248
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 12176 11354 12204 12242
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 12162 10432 12218 10441
rect 11992 10390 12162 10418
rect 12162 10367 12218 10376
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 11900 9722 11928 10066
rect 12176 9761 12204 10367
rect 12162 9752 12218 9761
rect 11888 9716 11940 9722
rect 12162 9687 12218 9696
rect 11888 9658 11940 9664
rect 12176 9518 12204 9687
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 11992 9178 12020 9318
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 12268 9081 12296 15263
rect 12452 15162 12480 15438
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 12348 13524 12400 13530
rect 12348 13466 12400 13472
rect 12360 11286 12388 13466
rect 12544 13258 12572 15864
rect 12714 15872 12770 15881
rect 12714 15807 12770 15816
rect 12728 13433 12756 15807
rect 12820 13462 12848 17575
rect 13096 17105 13124 18634
rect 13082 17096 13138 17105
rect 13082 17031 13138 17040
rect 13082 16824 13138 16833
rect 13082 16759 13138 16768
rect 13096 16726 13124 16759
rect 13084 16720 13136 16726
rect 13084 16662 13136 16668
rect 13084 16584 13136 16590
rect 13084 16526 13136 16532
rect 13096 16250 13124 16526
rect 13084 16244 13136 16250
rect 13084 16186 13136 16192
rect 13188 16130 13216 21678
rect 13266 21448 13322 21457
rect 13266 21383 13322 21392
rect 13280 20913 13308 21383
rect 13372 21146 13400 24346
rect 13464 22166 13492 24686
rect 13648 24274 13676 27520
rect 13728 25832 13780 25838
rect 13728 25774 13780 25780
rect 13740 24834 13768 25774
rect 14096 25152 14148 25158
rect 14096 25094 14148 25100
rect 13740 24806 13860 24834
rect 13832 24342 13860 24806
rect 14108 24750 14136 25094
rect 14096 24744 14148 24750
rect 14096 24686 14148 24692
rect 13820 24336 13872 24342
rect 13820 24278 13872 24284
rect 13636 24268 13688 24274
rect 13636 24210 13688 24216
rect 13636 24132 13688 24138
rect 13636 24074 13688 24080
rect 13544 23112 13596 23118
rect 13544 23054 13596 23060
rect 13556 22234 13584 23054
rect 13544 22228 13596 22234
rect 13544 22170 13596 22176
rect 13452 22160 13504 22166
rect 13452 22102 13504 22108
rect 13648 21593 13676 24074
rect 13728 24064 13780 24070
rect 13728 24006 13780 24012
rect 13740 23338 13768 24006
rect 13832 23526 13860 24278
rect 13912 24200 13964 24206
rect 13912 24142 13964 24148
rect 14004 24200 14056 24206
rect 14004 24142 14056 24148
rect 13924 23594 13952 24142
rect 13912 23588 13964 23594
rect 13912 23530 13964 23536
rect 13820 23520 13872 23526
rect 13820 23462 13872 23468
rect 13740 23310 13860 23338
rect 13832 23254 13860 23310
rect 13820 23248 13872 23254
rect 13726 23216 13782 23225
rect 13820 23190 13872 23196
rect 13726 23151 13782 23160
rect 13740 23050 13768 23151
rect 13728 23044 13780 23050
rect 13728 22986 13780 22992
rect 13728 22636 13780 22642
rect 13728 22578 13780 22584
rect 13740 22234 13768 22578
rect 13832 22234 13860 23190
rect 13924 22642 13952 23530
rect 14016 23118 14044 24142
rect 14004 23112 14056 23118
rect 14004 23054 14056 23060
rect 14002 22944 14058 22953
rect 14002 22879 14058 22888
rect 13912 22636 13964 22642
rect 13912 22578 13964 22584
rect 13728 22228 13780 22234
rect 13728 22170 13780 22176
rect 13820 22228 13872 22234
rect 13820 22170 13872 22176
rect 13728 22092 13780 22098
rect 14016 22080 14044 22879
rect 13728 22034 13780 22040
rect 13832 22052 14044 22080
rect 13634 21584 13690 21593
rect 13634 21519 13690 21528
rect 13452 21412 13504 21418
rect 13452 21354 13504 21360
rect 13360 21140 13412 21146
rect 13360 21082 13412 21088
rect 13266 20904 13322 20913
rect 13266 20839 13322 20848
rect 13372 20602 13400 21082
rect 13360 20596 13412 20602
rect 13360 20538 13412 20544
rect 13372 19281 13400 20538
rect 13358 19272 13414 19281
rect 13358 19207 13414 19216
rect 13268 19168 13320 19174
rect 13268 19110 13320 19116
rect 13280 18057 13308 19110
rect 13372 18154 13400 19207
rect 13464 18329 13492 21354
rect 13740 21146 13768 22034
rect 13832 21865 13860 22052
rect 13912 21888 13964 21894
rect 13818 21856 13874 21865
rect 13912 21830 13964 21836
rect 13818 21791 13874 21800
rect 13728 21140 13780 21146
rect 13780 21100 13860 21128
rect 13728 21082 13780 21088
rect 13728 21004 13780 21010
rect 13728 20946 13780 20952
rect 13544 20800 13596 20806
rect 13544 20742 13596 20748
rect 13556 19990 13584 20742
rect 13636 20392 13688 20398
rect 13636 20334 13688 20340
rect 13544 19984 13596 19990
rect 13544 19926 13596 19932
rect 13556 19174 13584 19926
rect 13648 19922 13676 20334
rect 13636 19916 13688 19922
rect 13636 19858 13688 19864
rect 13648 19242 13676 19858
rect 13636 19236 13688 19242
rect 13636 19178 13688 19184
rect 13544 19168 13596 19174
rect 13542 19136 13544 19145
rect 13596 19136 13598 19145
rect 13542 19071 13598 19080
rect 13740 18834 13768 20946
rect 13832 20398 13860 21100
rect 13820 20392 13872 20398
rect 13924 20369 13952 21830
rect 14004 21344 14056 21350
rect 14004 21286 14056 21292
rect 14016 20641 14044 21286
rect 14002 20632 14058 20641
rect 14108 20602 14136 24686
rect 14200 24138 14228 27520
rect 14660 24698 14688 27520
rect 15212 25480 15240 27520
rect 15660 25492 15712 25498
rect 15212 25452 15424 25480
rect 14740 25356 14792 25362
rect 14740 25298 14792 25304
rect 15292 25356 15344 25362
rect 15292 25298 15344 25304
rect 14384 24670 14688 24698
rect 14188 24132 14240 24138
rect 14188 24074 14240 24080
rect 14292 23526 14320 23557
rect 14280 23520 14332 23526
rect 14278 23488 14280 23497
rect 14332 23488 14334 23497
rect 14278 23423 14334 23432
rect 14188 23248 14240 23254
rect 14188 23190 14240 23196
rect 14200 22778 14228 23190
rect 14292 23186 14320 23423
rect 14280 23180 14332 23186
rect 14280 23122 14332 23128
rect 14188 22772 14240 22778
rect 14188 22714 14240 22720
rect 14188 22500 14240 22506
rect 14188 22442 14240 22448
rect 14200 21894 14228 22442
rect 14292 22166 14320 23122
rect 14280 22160 14332 22166
rect 14280 22102 14332 22108
rect 14280 21956 14332 21962
rect 14280 21898 14332 21904
rect 14188 21888 14240 21894
rect 14188 21830 14240 21836
rect 14188 21548 14240 21554
rect 14188 21490 14240 21496
rect 14002 20567 14058 20576
rect 14096 20596 14148 20602
rect 14096 20538 14148 20544
rect 13820 20334 13872 20340
rect 13910 20360 13966 20369
rect 13832 20058 13860 20334
rect 13910 20295 13966 20304
rect 13820 20052 13872 20058
rect 13820 19994 13872 20000
rect 13924 19938 13952 20295
rect 13832 19910 13952 19938
rect 13728 18828 13780 18834
rect 13728 18770 13780 18776
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 13728 18624 13780 18630
rect 13728 18566 13780 18572
rect 13450 18320 13506 18329
rect 13450 18255 13506 18264
rect 13360 18148 13412 18154
rect 13360 18090 13412 18096
rect 13266 18048 13322 18057
rect 13266 17983 13322 17992
rect 13372 17882 13400 18090
rect 13464 18034 13492 18255
rect 13556 18193 13584 18566
rect 13636 18352 13688 18358
rect 13636 18294 13688 18300
rect 13542 18184 13598 18193
rect 13542 18119 13598 18128
rect 13464 18006 13584 18034
rect 13450 17912 13506 17921
rect 13360 17876 13412 17882
rect 13450 17847 13506 17856
rect 13360 17818 13412 17824
rect 13266 17096 13322 17105
rect 13266 17031 13322 17040
rect 12912 16102 13216 16130
rect 12912 14929 12940 16102
rect 13176 16040 13228 16046
rect 13174 16008 13176 16017
rect 13228 16008 13230 16017
rect 13174 15943 13230 15952
rect 12992 15564 13044 15570
rect 12992 15506 13044 15512
rect 12898 14920 12954 14929
rect 12898 14855 12954 14864
rect 12808 13456 12860 13462
rect 12714 13424 12770 13433
rect 12808 13398 12860 13404
rect 12714 13359 12770 13368
rect 12532 13252 12584 13258
rect 12532 13194 12584 13200
rect 12820 12986 12848 13398
rect 13004 13394 13032 15506
rect 13280 15094 13308 17031
rect 13360 16992 13412 16998
rect 13360 16934 13412 16940
rect 13372 16590 13400 16934
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 13268 15088 13320 15094
rect 13268 15030 13320 15036
rect 13358 15056 13414 15065
rect 13084 15020 13136 15026
rect 13358 14991 13414 15000
rect 13084 14962 13136 14968
rect 13096 14618 13124 14962
rect 13084 14612 13136 14618
rect 13084 14554 13136 14560
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 13372 12986 13400 14991
rect 13464 14657 13492 17847
rect 13556 17524 13584 18006
rect 13648 17678 13676 18294
rect 13636 17672 13688 17678
rect 13636 17614 13688 17620
rect 13740 17610 13768 18566
rect 13832 18170 13860 19910
rect 14108 19514 14136 20538
rect 14096 19508 14148 19514
rect 14096 19450 14148 19456
rect 13912 18964 13964 18970
rect 13912 18906 13964 18912
rect 13924 18290 13952 18906
rect 14004 18760 14056 18766
rect 14004 18702 14056 18708
rect 14016 18426 14044 18702
rect 14004 18420 14056 18426
rect 14004 18362 14056 18368
rect 13912 18284 13964 18290
rect 13912 18226 13964 18232
rect 13832 18142 14044 18170
rect 13912 17740 13964 17746
rect 13912 17682 13964 17688
rect 13728 17604 13780 17610
rect 13728 17546 13780 17552
rect 13556 17496 13676 17524
rect 13544 17060 13596 17066
rect 13544 17002 13596 17008
rect 13556 15706 13584 17002
rect 13648 16572 13676 17496
rect 13924 16726 13952 17682
rect 14016 17354 14044 18142
rect 14200 17762 14228 21490
rect 14292 20505 14320 21898
rect 14278 20496 14334 20505
rect 14278 20431 14334 20440
rect 14200 17734 14320 17762
rect 14188 17672 14240 17678
rect 14188 17614 14240 17620
rect 14016 17326 14136 17354
rect 13728 16720 13780 16726
rect 13912 16720 13964 16726
rect 13780 16680 13860 16708
rect 13728 16662 13780 16668
rect 13648 16544 13768 16572
rect 13636 15972 13688 15978
rect 13636 15914 13688 15920
rect 13648 15745 13676 15914
rect 13634 15736 13690 15745
rect 13544 15700 13596 15706
rect 13634 15671 13690 15680
rect 13544 15642 13596 15648
rect 13740 15620 13768 16544
rect 13832 16250 13860 16680
rect 13912 16662 13964 16668
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13818 16144 13874 16153
rect 13818 16079 13874 16088
rect 13832 15978 13860 16079
rect 13820 15972 13872 15978
rect 13820 15914 13872 15920
rect 13924 15638 13952 16662
rect 14108 16425 14136 17326
rect 14200 16794 14228 17614
rect 14188 16788 14240 16794
rect 14188 16730 14240 16736
rect 14094 16416 14150 16425
rect 14094 16351 14150 16360
rect 13648 15592 13768 15620
rect 13912 15632 13964 15638
rect 13542 14920 13598 14929
rect 13542 14855 13598 14864
rect 13450 14648 13506 14657
rect 13450 14583 13506 14592
rect 13450 14512 13506 14521
rect 13450 14447 13452 14456
rect 13504 14447 13506 14456
rect 13452 14418 13504 14424
rect 13464 13870 13492 14418
rect 13452 13864 13504 13870
rect 13452 13806 13504 13812
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 13360 12980 13412 12986
rect 13360 12922 13412 12928
rect 12622 12472 12678 12481
rect 12622 12407 12678 12416
rect 13266 12472 13322 12481
rect 13266 12407 13322 12416
rect 12348 11280 12400 11286
rect 12348 11222 12400 11228
rect 12360 11132 12388 11222
rect 12360 11104 12480 11132
rect 12452 10266 12480 11104
rect 12532 10736 12584 10742
rect 12532 10678 12584 10684
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12544 10198 12572 10678
rect 12532 10192 12584 10198
rect 12532 10134 12584 10140
rect 12348 9444 12400 9450
rect 12348 9386 12400 9392
rect 12254 9072 12310 9081
rect 12360 9042 12388 9386
rect 12254 9007 12310 9016
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 12254 8936 12310 8945
rect 12254 8871 12310 8880
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11704 8560 11756 8566
rect 11704 8502 11756 8508
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 11612 8016 11664 8022
rect 11612 7958 11664 7964
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10336 7546 10364 7822
rect 11624 7546 11652 7958
rect 11808 7857 11836 8570
rect 12268 8430 12296 8871
rect 12440 8560 12492 8566
rect 12440 8502 12492 8508
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 12256 7948 12308 7954
rect 12452 7936 12480 8502
rect 12308 7908 12480 7936
rect 12256 7890 12308 7896
rect 12072 7880 12124 7886
rect 11794 7848 11850 7857
rect 12072 7822 12124 7828
rect 11794 7783 11850 7792
rect 11980 7744 12032 7750
rect 11980 7686 12032 7692
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 11612 7540 11664 7546
rect 11612 7482 11664 7488
rect 11992 7449 12020 7686
rect 12084 7546 12112 7822
rect 12072 7540 12124 7546
rect 12072 7482 12124 7488
rect 11978 7440 12034 7449
rect 11978 7375 12034 7384
rect 9956 7336 10008 7342
rect 9956 7278 10008 7284
rect 9968 7002 9996 7278
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 12268 7002 12296 7890
rect 12636 7886 12664 12407
rect 13280 12170 13308 12407
rect 13268 12164 13320 12170
rect 13268 12106 13320 12112
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 13188 11393 13216 11698
rect 13268 11552 13320 11558
rect 13266 11520 13268 11529
rect 13320 11520 13322 11529
rect 13266 11455 13322 11464
rect 13174 11384 13230 11393
rect 13174 11319 13230 11328
rect 13084 11008 13136 11014
rect 13084 10950 13136 10956
rect 13096 10538 13124 10950
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 12716 10532 12768 10538
rect 12716 10474 12768 10480
rect 13084 10532 13136 10538
rect 13084 10474 13136 10480
rect 12728 10198 12756 10474
rect 13082 10432 13138 10441
rect 13082 10367 13138 10376
rect 13096 10266 13124 10367
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 12716 10192 12768 10198
rect 12716 10134 12768 10140
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 13096 9450 13124 9998
rect 13084 9444 13136 9450
rect 13084 9386 13136 9392
rect 13096 8838 13124 9386
rect 13188 8906 13216 10610
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 13464 10062 13492 10406
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13556 9110 13584 14855
rect 13648 9178 13676 15592
rect 13912 15574 13964 15580
rect 13910 15056 13966 15065
rect 13910 14991 13912 15000
rect 13964 14991 13966 15000
rect 13912 14962 13964 14968
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13832 13410 13860 14894
rect 14292 14618 14320 17734
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 14292 14006 14320 14554
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 14292 13841 14320 13942
rect 14278 13832 14334 13841
rect 14278 13767 14334 13776
rect 13740 13382 13860 13410
rect 13740 13326 13768 13382
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13832 12442 13860 13382
rect 13912 13320 13964 13326
rect 13912 13262 13964 13268
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 13924 12850 13952 13262
rect 14002 12880 14058 12889
rect 13912 12844 13964 12850
rect 14002 12815 14058 12824
rect 13912 12786 13964 12792
rect 14016 12714 14044 12815
rect 14004 12708 14056 12714
rect 14004 12650 14056 12656
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13912 11824 13964 11830
rect 13912 11766 13964 11772
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13740 9466 13768 10542
rect 13820 9648 13872 9654
rect 13818 9616 13820 9625
rect 13872 9616 13874 9625
rect 13818 9551 13874 9560
rect 13740 9438 13860 9466
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13544 9104 13596 9110
rect 13544 9046 13596 9052
rect 13176 8900 13228 8906
rect 13176 8842 13228 8848
rect 13084 8832 13136 8838
rect 13084 8774 13136 8780
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 12728 7546 12756 8298
rect 13096 7546 13124 8774
rect 13452 8492 13504 8498
rect 13452 8434 13504 8440
rect 13464 7818 13492 8434
rect 13556 7886 13584 9046
rect 13648 8634 13676 9114
rect 13636 8628 13688 8634
rect 13636 8570 13688 8576
rect 13648 8537 13676 8570
rect 13634 8528 13690 8537
rect 13634 8463 13690 8472
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13452 7812 13504 7818
rect 13452 7754 13504 7760
rect 13464 7546 13492 7754
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 13084 7540 13136 7546
rect 13084 7482 13136 7488
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13832 7426 13860 9438
rect 13924 8090 13952 11766
rect 14292 11694 14320 13262
rect 14384 12374 14412 24670
rect 14464 24608 14516 24614
rect 14464 24550 14516 24556
rect 14476 21434 14504 24550
rect 14556 24132 14608 24138
rect 14556 24074 14608 24080
rect 14568 21622 14596 24074
rect 14752 24070 14780 25298
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15304 24614 15332 25298
rect 15396 24857 15424 25452
rect 15764 25480 15792 27520
rect 15712 25452 15792 25480
rect 15660 25434 15712 25440
rect 16316 25362 16344 27520
rect 16868 25498 16896 27520
rect 16856 25492 16908 25498
rect 16856 25434 16908 25440
rect 16304 25356 16356 25362
rect 16304 25298 16356 25304
rect 16948 25356 17000 25362
rect 16948 25298 17000 25304
rect 15660 25288 15712 25294
rect 15660 25230 15712 25236
rect 15382 24848 15438 24857
rect 15382 24783 15438 24792
rect 15568 24812 15620 24818
rect 15568 24754 15620 24760
rect 15384 24744 15436 24750
rect 15384 24686 15436 24692
rect 14832 24608 14884 24614
rect 14832 24550 14884 24556
rect 15292 24608 15344 24614
rect 15292 24550 15344 24556
rect 14844 24410 14872 24550
rect 14832 24404 14884 24410
rect 14832 24346 14884 24352
rect 14740 24064 14792 24070
rect 14740 24006 14792 24012
rect 14752 22710 14780 24006
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15304 23225 15332 24550
rect 15290 23216 15346 23225
rect 15290 23151 15346 23160
rect 14832 22976 14884 22982
rect 14832 22918 14884 22924
rect 14740 22704 14792 22710
rect 14740 22646 14792 22652
rect 14740 22568 14792 22574
rect 14740 22510 14792 22516
rect 14648 21888 14700 21894
rect 14648 21830 14700 21836
rect 14556 21616 14608 21622
rect 14556 21558 14608 21564
rect 14660 21554 14688 21830
rect 14752 21690 14780 22510
rect 14740 21684 14792 21690
rect 14740 21626 14792 21632
rect 14648 21548 14700 21554
rect 14648 21490 14700 21496
rect 14476 21418 14596 21434
rect 14476 21412 14608 21418
rect 14476 21406 14556 21412
rect 14556 21354 14608 21360
rect 14462 21312 14518 21321
rect 14462 21247 14518 21256
rect 14476 20777 14504 21247
rect 14568 21146 14596 21354
rect 14556 21140 14608 21146
rect 14556 21082 14608 21088
rect 14660 20874 14688 21490
rect 14740 20936 14792 20942
rect 14740 20878 14792 20884
rect 14648 20868 14700 20874
rect 14648 20810 14700 20816
rect 14462 20768 14518 20777
rect 14462 20703 14518 20712
rect 14476 18766 14504 20703
rect 14752 20602 14780 20878
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 14556 20392 14608 20398
rect 14556 20334 14608 20340
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 14568 17882 14596 20334
rect 14648 20256 14700 20262
rect 14646 20224 14648 20233
rect 14700 20224 14702 20233
rect 14646 20159 14702 20168
rect 14660 18902 14688 20159
rect 14752 20058 14780 20538
rect 14740 20052 14792 20058
rect 14740 19994 14792 20000
rect 14648 18896 14700 18902
rect 14648 18838 14700 18844
rect 14660 18426 14688 18838
rect 14844 18426 14872 22918
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14924 22704 14976 22710
rect 14924 22646 14976 22652
rect 14936 21962 14964 22646
rect 15396 22574 15424 24686
rect 15476 24676 15528 24682
rect 15476 24618 15528 24624
rect 15488 24154 15516 24618
rect 15580 24274 15608 24754
rect 15568 24268 15620 24274
rect 15568 24210 15620 24216
rect 15488 24126 15608 24154
rect 15476 23588 15528 23594
rect 15476 23530 15528 23536
rect 15488 22817 15516 23530
rect 15474 22808 15530 22817
rect 15474 22743 15530 22752
rect 15580 22692 15608 24126
rect 15488 22664 15608 22692
rect 15384 22568 15436 22574
rect 15384 22510 15436 22516
rect 15292 22160 15344 22166
rect 15292 22102 15344 22108
rect 14924 21956 14976 21962
rect 14924 21898 14976 21904
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15304 21486 15332 22102
rect 15384 21888 15436 21894
rect 15384 21830 15436 21836
rect 15396 21593 15424 21830
rect 15382 21584 15438 21593
rect 15382 21519 15438 21528
rect 15292 21480 15344 21486
rect 15292 21422 15344 21428
rect 15108 21412 15160 21418
rect 15108 21354 15160 21360
rect 15120 21128 15148 21354
rect 15120 21100 15424 21128
rect 15292 21004 15344 21010
rect 15292 20946 15344 20952
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15016 20324 15068 20330
rect 15304 20312 15332 20946
rect 15068 20284 15332 20312
rect 15016 20266 15068 20272
rect 15120 20058 15148 20284
rect 15290 20224 15346 20233
rect 15290 20159 15346 20168
rect 15108 20052 15160 20058
rect 15108 19994 15160 20000
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15304 19428 15332 20159
rect 14936 19400 15332 19428
rect 14936 19281 14964 19400
rect 14922 19272 14978 19281
rect 14922 19207 14978 19216
rect 14936 18698 14964 19207
rect 15396 19174 15424 21100
rect 15488 20233 15516 22664
rect 15568 22092 15620 22098
rect 15568 22034 15620 22040
rect 15580 20806 15608 22034
rect 15568 20800 15620 20806
rect 15568 20742 15620 20748
rect 15474 20224 15530 20233
rect 15474 20159 15530 20168
rect 15474 20088 15530 20097
rect 15474 20023 15530 20032
rect 15384 19168 15436 19174
rect 15384 19110 15436 19116
rect 14924 18692 14976 18698
rect 14924 18634 14976 18640
rect 15384 18624 15436 18630
rect 15384 18566 15436 18572
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14648 18420 14700 18426
rect 14648 18362 14700 18368
rect 14832 18420 14884 18426
rect 14832 18362 14884 18368
rect 14740 18352 14792 18358
rect 14740 18294 14792 18300
rect 14556 17876 14608 17882
rect 14556 17818 14608 17824
rect 14568 16658 14596 17818
rect 14556 16652 14608 16658
rect 14556 16594 14608 16600
rect 14648 16584 14700 16590
rect 14648 16526 14700 16532
rect 14554 16280 14610 16289
rect 14660 16250 14688 16526
rect 14752 16250 14780 18294
rect 15396 18154 15424 18566
rect 15488 18426 15516 20023
rect 15568 19712 15620 19718
rect 15568 19654 15620 19660
rect 15476 18420 15528 18426
rect 15476 18362 15528 18368
rect 15384 18148 15436 18154
rect 15384 18090 15436 18096
rect 15382 18048 15438 18057
rect 15382 17983 15438 17992
rect 15292 17740 15344 17746
rect 15292 17682 15344 17688
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 14554 16215 14610 16224
rect 14648 16244 14700 16250
rect 14568 15502 14596 16215
rect 14648 16186 14700 16192
rect 14740 16244 14792 16250
rect 14740 16186 14792 16192
rect 14660 16046 14688 16186
rect 14844 16114 14872 17478
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15200 17128 15252 17134
rect 15200 17070 15252 17076
rect 15212 16998 15240 17070
rect 15200 16992 15252 16998
rect 15200 16934 15252 16940
rect 15212 16572 15240 16934
rect 15304 16726 15332 17682
rect 15292 16720 15344 16726
rect 15292 16662 15344 16668
rect 15292 16584 15344 16590
rect 15212 16544 15292 16572
rect 15292 16526 15344 16532
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15304 16250 15332 16526
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 14648 16040 14700 16046
rect 14648 15982 14700 15988
rect 15396 15570 15424 17983
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15488 15978 15516 16390
rect 15476 15972 15528 15978
rect 15476 15914 15528 15920
rect 15488 15638 15516 15914
rect 15580 15910 15608 19654
rect 15672 17814 15700 25230
rect 16486 24712 16542 24721
rect 16486 24647 16542 24656
rect 16396 24608 16448 24614
rect 16396 24550 16448 24556
rect 16028 24200 16080 24206
rect 16028 24142 16080 24148
rect 15750 23352 15806 23361
rect 15750 23287 15806 23296
rect 15764 23254 15792 23287
rect 15752 23248 15804 23254
rect 15752 23190 15804 23196
rect 15750 22400 15806 22409
rect 15750 22335 15806 22344
rect 15764 21078 15792 22335
rect 15844 22024 15896 22030
rect 15844 21966 15896 21972
rect 15856 21418 15884 21966
rect 15936 21480 15988 21486
rect 15936 21422 15988 21428
rect 15844 21412 15896 21418
rect 15844 21354 15896 21360
rect 15842 21176 15898 21185
rect 15842 21111 15898 21120
rect 15752 21072 15804 21078
rect 15752 21014 15804 21020
rect 15764 20262 15792 21014
rect 15856 20777 15884 21111
rect 15842 20768 15898 20777
rect 15842 20703 15898 20712
rect 15752 20256 15804 20262
rect 15750 20224 15752 20233
rect 15804 20224 15806 20233
rect 15750 20159 15806 20168
rect 15844 20052 15896 20058
rect 15844 19994 15896 20000
rect 15750 19680 15806 19689
rect 15750 19615 15806 19624
rect 15764 18698 15792 19615
rect 15856 18970 15884 19994
rect 15844 18964 15896 18970
rect 15844 18906 15896 18912
rect 15752 18692 15804 18698
rect 15752 18634 15804 18640
rect 15660 17808 15712 17814
rect 15660 17750 15712 17756
rect 15856 17338 15884 18906
rect 15844 17332 15896 17338
rect 15844 17274 15896 17280
rect 15856 16726 15884 17274
rect 15844 16720 15896 16726
rect 15844 16662 15896 16668
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 15660 15972 15712 15978
rect 15660 15914 15712 15920
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15580 15706 15608 15846
rect 15568 15700 15620 15706
rect 15568 15642 15620 15648
rect 15672 15638 15700 15914
rect 15856 15910 15884 16186
rect 15844 15904 15896 15910
rect 15844 15846 15896 15852
rect 15750 15736 15806 15745
rect 15750 15671 15752 15680
rect 15804 15671 15806 15680
rect 15752 15642 15804 15648
rect 15476 15632 15528 15638
rect 15476 15574 15528 15580
rect 15660 15632 15712 15638
rect 15660 15574 15712 15580
rect 15384 15564 15436 15570
rect 15384 15506 15436 15512
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15108 15088 15160 15094
rect 15108 15030 15160 15036
rect 14554 14920 14610 14929
rect 14554 14855 14610 14864
rect 14464 14816 14516 14822
rect 14464 14758 14516 14764
rect 14476 14074 14504 14758
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14568 12986 14596 14855
rect 15120 14385 15148 15030
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 15106 14376 15162 14385
rect 15396 14346 15424 14962
rect 15856 14890 15884 15846
rect 15844 14884 15896 14890
rect 15844 14826 15896 14832
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 15106 14311 15162 14320
rect 15384 14340 15436 14346
rect 15384 14282 15436 14288
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 15028 13326 15056 13806
rect 15474 13560 15530 13569
rect 15474 13495 15530 13504
rect 15016 13320 15068 13326
rect 15016 13262 15068 13268
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15488 13025 15516 13495
rect 15580 13462 15608 14418
rect 15568 13456 15620 13462
rect 15566 13424 15568 13433
rect 15620 13424 15622 13433
rect 15566 13359 15622 13368
rect 15856 13326 15884 14826
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 15474 13016 15530 13025
rect 14556 12980 14608 12986
rect 15474 12951 15530 12960
rect 14556 12922 14608 12928
rect 14372 12368 14424 12374
rect 14372 12310 14424 12316
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14292 10810 14320 11630
rect 14384 11121 14412 12310
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14464 11620 14516 11626
rect 14464 11562 14516 11568
rect 14476 11354 14504 11562
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14370 11112 14426 11121
rect 14370 11047 14426 11056
rect 14280 10804 14332 10810
rect 14280 10746 14332 10752
rect 14476 10470 14504 11290
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14648 10532 14700 10538
rect 14648 10474 14700 10480
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14186 10296 14242 10305
rect 14186 10231 14242 10240
rect 14200 10033 14228 10231
rect 14476 10198 14504 10406
rect 14660 10305 14688 10474
rect 14646 10296 14702 10305
rect 14646 10231 14648 10240
rect 14700 10231 14702 10240
rect 14648 10202 14700 10208
rect 14464 10192 14516 10198
rect 14660 10171 14688 10202
rect 14464 10134 14516 10140
rect 14186 10024 14242 10033
rect 14186 9959 14242 9968
rect 14004 9648 14056 9654
rect 14004 9590 14056 9596
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 13924 7546 13952 8026
rect 14016 7886 14044 9590
rect 14094 9480 14150 9489
rect 14094 9415 14150 9424
rect 14108 8362 14136 9415
rect 14200 9178 14228 9959
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 14200 8430 14228 9114
rect 14476 8498 14504 10134
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15304 9722 15332 10066
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15396 9761 15424 9862
rect 15382 9752 15438 9761
rect 15292 9716 15344 9722
rect 15382 9687 15438 9696
rect 15292 9658 15344 9664
rect 15488 9450 15516 12951
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15672 11898 15700 12242
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 15764 11665 15792 12038
rect 15750 11656 15806 11665
rect 15750 11591 15806 11600
rect 15750 10976 15806 10985
rect 15750 10911 15806 10920
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15580 9586 15608 10406
rect 15660 10192 15712 10198
rect 15764 10169 15792 10911
rect 15948 10849 15976 21422
rect 16040 21185 16068 24142
rect 16304 23656 16356 23662
rect 16304 23598 16356 23604
rect 16212 23316 16264 23322
rect 16212 23258 16264 23264
rect 16224 22506 16252 23258
rect 16316 22778 16344 23598
rect 16304 22772 16356 22778
rect 16304 22714 16356 22720
rect 16212 22500 16264 22506
rect 16212 22442 16264 22448
rect 16408 21690 16436 24550
rect 16500 23866 16528 24647
rect 16960 24614 16988 25298
rect 17224 25288 17276 25294
rect 17222 25256 17224 25265
rect 17276 25256 17278 25265
rect 17420 25226 17448 27520
rect 17222 25191 17278 25200
rect 17408 25220 17460 25226
rect 17408 25162 17460 25168
rect 17880 24857 17908 27520
rect 18236 25356 18288 25362
rect 18236 25298 18288 25304
rect 17866 24848 17922 24857
rect 17866 24783 17922 24792
rect 18052 24744 18104 24750
rect 18050 24712 18052 24721
rect 18104 24712 18106 24721
rect 18248 24682 18276 25298
rect 18432 24721 18460 27520
rect 18418 24712 18474 24721
rect 18050 24647 18106 24656
rect 18236 24676 18288 24682
rect 18418 24647 18474 24656
rect 18236 24618 18288 24624
rect 16948 24608 17000 24614
rect 16948 24550 17000 24556
rect 17592 24336 17644 24342
rect 17592 24278 17644 24284
rect 17500 24200 17552 24206
rect 17498 24168 17500 24177
rect 17552 24168 17554 24177
rect 17132 24132 17184 24138
rect 17498 24103 17554 24112
rect 17132 24074 17184 24080
rect 16948 24064 17000 24070
rect 16948 24006 17000 24012
rect 16488 23860 16540 23866
rect 16488 23802 16540 23808
rect 16672 23588 16724 23594
rect 16672 23530 16724 23536
rect 16684 23322 16712 23530
rect 16672 23316 16724 23322
rect 16672 23258 16724 23264
rect 16684 23050 16712 23258
rect 16672 23044 16724 23050
rect 16672 22986 16724 22992
rect 16764 22636 16816 22642
rect 16764 22578 16816 22584
rect 16856 22636 16908 22642
rect 16856 22578 16908 22584
rect 16776 22545 16804 22578
rect 16762 22536 16818 22545
rect 16762 22471 16818 22480
rect 16868 22234 16896 22578
rect 16672 22228 16724 22234
rect 16672 22170 16724 22176
rect 16856 22228 16908 22234
rect 16856 22170 16908 22176
rect 16396 21684 16448 21690
rect 16396 21626 16448 21632
rect 16488 21412 16540 21418
rect 16488 21354 16540 21360
rect 16394 21312 16450 21321
rect 16394 21247 16450 21256
rect 16026 21176 16082 21185
rect 16408 21146 16436 21247
rect 16026 21111 16082 21120
rect 16396 21140 16448 21146
rect 16396 21082 16448 21088
rect 16394 20224 16450 20233
rect 16394 20159 16450 20168
rect 16304 19848 16356 19854
rect 16304 19790 16356 19796
rect 16316 19174 16344 19790
rect 16304 19168 16356 19174
rect 16304 19110 16356 19116
rect 16212 18896 16264 18902
rect 16212 18838 16264 18844
rect 16028 18828 16080 18834
rect 16028 18770 16080 18776
rect 16040 18086 16068 18770
rect 16120 18760 16172 18766
rect 16120 18702 16172 18708
rect 16028 18080 16080 18086
rect 16028 18022 16080 18028
rect 16040 17377 16068 18022
rect 16132 17882 16160 18702
rect 16224 18057 16252 18838
rect 16210 18048 16266 18057
rect 16210 17983 16266 17992
rect 16120 17876 16172 17882
rect 16120 17818 16172 17824
rect 16026 17368 16082 17377
rect 16026 17303 16082 17312
rect 16224 16250 16252 17983
rect 16316 16697 16344 19110
rect 16408 18426 16436 20159
rect 16500 19310 16528 21354
rect 16684 21146 16712 22170
rect 16960 22114 16988 24006
rect 17144 23594 17172 24074
rect 17512 23798 17540 24103
rect 17500 23792 17552 23798
rect 17500 23734 17552 23740
rect 17500 23656 17552 23662
rect 17500 23598 17552 23604
rect 17132 23588 17184 23594
rect 17132 23530 17184 23536
rect 17224 23248 17276 23254
rect 17224 23190 17276 23196
rect 17236 22438 17264 23190
rect 17408 23112 17460 23118
rect 17408 23054 17460 23060
rect 17420 22953 17448 23054
rect 17406 22944 17462 22953
rect 17406 22879 17462 22888
rect 17420 22642 17448 22879
rect 17408 22636 17460 22642
rect 17408 22578 17460 22584
rect 17224 22432 17276 22438
rect 17224 22374 17276 22380
rect 16868 22086 16988 22114
rect 16868 21962 16896 22086
rect 16856 21956 16908 21962
rect 16856 21898 16908 21904
rect 16868 21554 16896 21898
rect 16856 21548 16908 21554
rect 16856 21490 16908 21496
rect 17132 21344 17184 21350
rect 17132 21286 17184 21292
rect 16580 21140 16632 21146
rect 16580 21082 16632 21088
rect 16672 21140 16724 21146
rect 16672 21082 16724 21088
rect 16592 20398 16620 21082
rect 17040 21004 17092 21010
rect 17040 20946 17092 20952
rect 16948 20936 17000 20942
rect 16948 20878 17000 20884
rect 16960 20398 16988 20878
rect 16580 20392 16632 20398
rect 16580 20334 16632 20340
rect 16948 20392 17000 20398
rect 16948 20334 17000 20340
rect 16856 20324 16908 20330
rect 16856 20266 16908 20272
rect 16868 20058 16896 20266
rect 16856 20052 16908 20058
rect 16856 19994 16908 20000
rect 16960 19938 16988 20334
rect 17052 20058 17080 20946
rect 17144 20942 17172 21286
rect 17132 20936 17184 20942
rect 17132 20878 17184 20884
rect 17040 20052 17092 20058
rect 17040 19994 17092 20000
rect 17132 19984 17184 19990
rect 16764 19916 16816 19922
rect 16960 19910 17080 19938
rect 17236 19961 17264 22374
rect 17408 22092 17460 22098
rect 17408 22034 17460 22040
rect 17420 21350 17448 22034
rect 17512 21690 17540 23598
rect 17604 23526 17632 24278
rect 17682 23760 17738 23769
rect 17682 23695 17738 23704
rect 17592 23520 17644 23526
rect 17592 23462 17644 23468
rect 17500 21684 17552 21690
rect 17500 21626 17552 21632
rect 17512 21486 17540 21626
rect 17500 21480 17552 21486
rect 17500 21422 17552 21428
rect 17408 21344 17460 21350
rect 17408 21286 17460 21292
rect 17498 20768 17554 20777
rect 17604 20754 17632 23462
rect 17696 23186 17724 23695
rect 17776 23588 17828 23594
rect 17776 23530 17828 23536
rect 17684 23180 17736 23186
rect 17684 23122 17736 23128
rect 17696 22778 17724 23122
rect 17684 22772 17736 22778
rect 17684 22714 17736 22720
rect 17788 21894 17816 23530
rect 18144 23520 18196 23526
rect 18144 23462 18196 23468
rect 18156 22982 18184 23462
rect 18248 23361 18276 24618
rect 18328 24608 18380 24614
rect 18328 24550 18380 24556
rect 18340 24274 18368 24550
rect 18328 24268 18380 24274
rect 18328 24210 18380 24216
rect 18234 23352 18290 23361
rect 18234 23287 18290 23296
rect 18144 22976 18196 22982
rect 18144 22918 18196 22924
rect 18052 22772 18104 22778
rect 18052 22714 18104 22720
rect 17776 21888 17828 21894
rect 17776 21830 17828 21836
rect 17788 21010 17816 21830
rect 17960 21412 18012 21418
rect 17960 21354 18012 21360
rect 17868 21140 17920 21146
rect 17868 21082 17920 21088
rect 17776 21004 17828 21010
rect 17776 20946 17828 20952
rect 17554 20726 17632 20754
rect 17498 20703 17554 20712
rect 17132 19926 17184 19932
rect 17222 19952 17278 19961
rect 16764 19858 16816 19864
rect 16488 19304 16540 19310
rect 16488 19246 16540 19252
rect 16776 19174 16804 19858
rect 17052 19854 17080 19910
rect 17040 19848 17092 19854
rect 17040 19790 17092 19796
rect 17052 19242 17080 19790
rect 17040 19236 17092 19242
rect 17040 19178 17092 19184
rect 16764 19168 16816 19174
rect 16764 19110 16816 19116
rect 16396 18420 16448 18426
rect 16396 18362 16448 18368
rect 16580 18284 16632 18290
rect 16580 18226 16632 18232
rect 16396 18216 16448 18222
rect 16396 18158 16448 18164
rect 16408 17320 16436 18158
rect 16592 17898 16620 18226
rect 16672 18080 16724 18086
rect 16672 18022 16724 18028
rect 16500 17882 16620 17898
rect 16488 17876 16620 17882
rect 16540 17870 16620 17876
rect 16488 17818 16540 17824
rect 16684 17678 16712 18022
rect 16672 17672 16724 17678
rect 16672 17614 16724 17620
rect 16580 17332 16632 17338
rect 16408 17292 16580 17320
rect 16580 17274 16632 17280
rect 16684 16998 16712 17614
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16302 16688 16358 16697
rect 16302 16623 16358 16632
rect 16212 16244 16264 16250
rect 16212 16186 16264 16192
rect 16396 15904 16448 15910
rect 16396 15846 16448 15852
rect 16408 15570 16436 15846
rect 16776 15586 16804 19110
rect 17052 18748 17080 19178
rect 17144 18970 17172 19926
rect 17222 19887 17278 19896
rect 17132 18964 17184 18970
rect 17132 18906 17184 18912
rect 17132 18760 17184 18766
rect 17052 18720 17132 18748
rect 17132 18702 17184 18708
rect 17040 18624 17092 18630
rect 16946 18592 17002 18601
rect 17040 18566 17092 18572
rect 16946 18527 17002 18536
rect 16960 18154 16988 18527
rect 17052 18329 17080 18566
rect 17038 18320 17094 18329
rect 17038 18255 17094 18264
rect 17052 18222 17080 18255
rect 17040 18216 17092 18222
rect 17040 18158 17092 18164
rect 16948 18148 17000 18154
rect 16948 18090 17000 18096
rect 17144 18086 17172 18702
rect 17132 18080 17184 18086
rect 17132 18022 17184 18028
rect 16948 17740 17000 17746
rect 16948 17682 17000 17688
rect 16960 16658 16988 17682
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 16854 16552 16910 16561
rect 16854 16487 16910 16496
rect 17038 16552 17094 16561
rect 17038 16487 17094 16496
rect 16868 15706 16896 16487
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 16856 15700 16908 15706
rect 16856 15642 16908 15648
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16672 15564 16724 15570
rect 16776 15558 16896 15586
rect 16672 15506 16724 15512
rect 16580 15496 16632 15502
rect 16500 15444 16580 15450
rect 16500 15438 16632 15444
rect 16500 15422 16620 15438
rect 16500 15162 16528 15422
rect 16684 15162 16712 15506
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 16672 15156 16724 15162
rect 16672 15098 16724 15104
rect 16396 14952 16448 14958
rect 16396 14894 16448 14900
rect 16408 14482 16436 14894
rect 16396 14476 16448 14482
rect 16396 14418 16448 14424
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 16040 13977 16068 14350
rect 16408 14074 16436 14418
rect 16762 14376 16818 14385
rect 16868 14362 16896 15558
rect 16960 15473 16988 16050
rect 17052 15978 17080 16487
rect 17040 15972 17092 15978
rect 17040 15914 17092 15920
rect 16946 15464 17002 15473
rect 16946 15399 17002 15408
rect 16948 14816 17000 14822
rect 16948 14758 17000 14764
rect 16960 14618 16988 14758
rect 16948 14612 17000 14618
rect 16948 14554 17000 14560
rect 17038 14376 17094 14385
rect 16868 14334 17038 14362
rect 16762 14311 16818 14320
rect 17038 14311 17094 14320
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16026 13968 16082 13977
rect 16026 13903 16082 13912
rect 16040 13870 16068 13903
rect 16028 13864 16080 13870
rect 16028 13806 16080 13812
rect 16408 13462 16436 14010
rect 16396 13456 16448 13462
rect 16396 13398 16448 13404
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 16040 12918 16068 13262
rect 16408 12986 16436 13398
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16028 12912 16080 12918
rect 16028 12854 16080 12860
rect 16488 12912 16540 12918
rect 16488 12854 16540 12860
rect 16212 12368 16264 12374
rect 16118 12336 16174 12345
rect 16212 12310 16264 12316
rect 16118 12271 16174 12280
rect 16132 12238 16160 12271
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 16132 11354 16160 12174
rect 16224 11898 16252 12310
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16316 11218 16344 12174
rect 16304 11212 16356 11218
rect 16304 11154 16356 11160
rect 15934 10840 15990 10849
rect 15934 10775 15990 10784
rect 15842 10568 15898 10577
rect 15842 10503 15898 10512
rect 15856 10266 15884 10503
rect 15844 10260 15896 10266
rect 15844 10202 15896 10208
rect 15660 10134 15712 10140
rect 15750 10160 15806 10169
rect 15672 9722 15700 10134
rect 15750 10095 15806 10104
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 15764 9654 15792 10095
rect 15752 9648 15804 9654
rect 15752 9590 15804 9596
rect 15568 9580 15620 9586
rect 15568 9522 15620 9528
rect 15476 9444 15528 9450
rect 15476 9386 15528 9392
rect 15488 9178 15516 9386
rect 15856 9178 15884 10202
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 15844 9172 15896 9178
rect 15844 9114 15896 9120
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 14096 8356 14148 8362
rect 14096 8298 14148 8304
rect 14476 8090 14504 8434
rect 14554 8392 14610 8401
rect 16500 8378 16528 12854
rect 16776 12714 16804 14311
rect 16948 14272 17000 14278
rect 16948 14214 17000 14220
rect 16960 12986 16988 14214
rect 17052 13705 17080 14311
rect 17038 13696 17094 13705
rect 17038 13631 17094 13640
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 16764 12708 16816 12714
rect 16764 12650 16816 12656
rect 16776 12442 16804 12650
rect 16764 12436 16816 12442
rect 17236 12424 17264 19887
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17512 16250 17540 16526
rect 17500 16244 17552 16250
rect 17500 16186 17552 16192
rect 17408 15700 17460 15706
rect 17408 15642 17460 15648
rect 17420 15162 17448 15642
rect 17408 15156 17460 15162
rect 17408 15098 17460 15104
rect 17316 14544 17368 14550
rect 17316 14486 17368 14492
rect 17328 14074 17356 14486
rect 17408 14408 17460 14414
rect 17408 14350 17460 14356
rect 17420 14074 17448 14350
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17604 13569 17632 20726
rect 17880 19990 17908 21082
rect 17972 20058 18000 21354
rect 18064 20330 18092 22714
rect 18156 21321 18184 22918
rect 18142 21312 18198 21321
rect 18142 21247 18198 21256
rect 18142 20632 18198 20641
rect 18340 20602 18368 24210
rect 18512 24064 18564 24070
rect 18512 24006 18564 24012
rect 18524 23594 18552 24006
rect 18880 23792 18932 23798
rect 18880 23734 18932 23740
rect 18420 23588 18472 23594
rect 18420 23530 18472 23536
rect 18512 23588 18564 23594
rect 18512 23530 18564 23536
rect 18142 20567 18198 20576
rect 18328 20596 18380 20602
rect 18052 20324 18104 20330
rect 18052 20266 18104 20272
rect 17960 20052 18012 20058
rect 17960 19994 18012 20000
rect 17868 19984 17920 19990
rect 17868 19926 17920 19932
rect 17972 19360 18000 19994
rect 17880 19332 18000 19360
rect 17880 18902 17908 19332
rect 17868 18896 17920 18902
rect 17868 18838 17920 18844
rect 17880 18426 17908 18838
rect 17868 18420 17920 18426
rect 17868 18362 17920 18368
rect 18052 17536 18104 17542
rect 18052 17478 18104 17484
rect 18064 17338 18092 17478
rect 18052 17332 18104 17338
rect 18052 17274 18104 17280
rect 18156 16726 18184 20567
rect 18328 20538 18380 20544
rect 18234 20496 18290 20505
rect 18234 20431 18290 20440
rect 18144 16720 18196 16726
rect 18144 16662 18196 16668
rect 17868 16448 17920 16454
rect 17868 16390 17920 16396
rect 17774 14648 17830 14657
rect 17774 14583 17830 14592
rect 17788 14006 17816 14583
rect 17880 14550 17908 16390
rect 18156 16289 18184 16662
rect 18142 16280 18198 16289
rect 18142 16215 18144 16224
rect 18196 16215 18198 16224
rect 18144 16186 18196 16192
rect 18156 16155 18184 16186
rect 18144 15972 18196 15978
rect 18144 15914 18196 15920
rect 18156 15502 18184 15914
rect 18144 15496 18196 15502
rect 18144 15438 18196 15444
rect 18156 14958 18184 15438
rect 18144 14952 18196 14958
rect 18144 14894 18196 14900
rect 18248 14793 18276 20431
rect 18326 19816 18382 19825
rect 18326 19751 18382 19760
rect 18340 19242 18368 19751
rect 18328 19236 18380 19242
rect 18328 19178 18380 19184
rect 18432 17241 18460 23530
rect 18524 21146 18552 23530
rect 18788 22704 18840 22710
rect 18788 22646 18840 22652
rect 18800 22166 18828 22646
rect 18892 22574 18920 23734
rect 18984 23066 19012 27520
rect 19432 25356 19484 25362
rect 19432 25298 19484 25304
rect 19340 24744 19392 24750
rect 19340 24686 19392 24692
rect 19352 24342 19380 24686
rect 19444 24410 19472 25298
rect 19432 24404 19484 24410
rect 19432 24346 19484 24352
rect 19340 24336 19392 24342
rect 19340 24278 19392 24284
rect 19432 24200 19484 24206
rect 19352 24177 19432 24188
rect 19338 24168 19432 24177
rect 19394 24160 19432 24168
rect 19432 24142 19484 24148
rect 19338 24103 19394 24112
rect 19340 24064 19392 24070
rect 19340 24006 19392 24012
rect 19352 23225 19380 24006
rect 19338 23216 19394 23225
rect 19338 23151 19394 23160
rect 18984 23038 19288 23066
rect 18972 22976 19024 22982
rect 18972 22918 19024 22924
rect 19156 22976 19208 22982
rect 19156 22918 19208 22924
rect 18984 22642 19012 22918
rect 18972 22636 19024 22642
rect 18972 22578 19024 22584
rect 18880 22568 18932 22574
rect 18880 22510 18932 22516
rect 19168 22506 19196 22918
rect 18972 22500 19024 22506
rect 18972 22442 19024 22448
rect 19156 22500 19208 22506
rect 19156 22442 19208 22448
rect 18788 22160 18840 22166
rect 18788 22102 18840 22108
rect 18984 21690 19012 22442
rect 19260 22250 19288 23038
rect 19340 22976 19392 22982
rect 19340 22918 19392 22924
rect 19168 22222 19288 22250
rect 19064 21888 19116 21894
rect 19168 21865 19196 22222
rect 19246 22128 19302 22137
rect 19246 22063 19302 22072
rect 19064 21830 19116 21836
rect 19154 21856 19210 21865
rect 18972 21684 19024 21690
rect 18972 21626 19024 21632
rect 19076 21486 19104 21830
rect 19154 21791 19210 21800
rect 19064 21480 19116 21486
rect 19064 21422 19116 21428
rect 18512 21140 18564 21146
rect 18512 21082 18564 21088
rect 18604 20800 18656 20806
rect 18604 20742 18656 20748
rect 18616 20330 18644 20742
rect 18604 20324 18656 20330
rect 18604 20266 18656 20272
rect 18616 20233 18644 20266
rect 19064 20256 19116 20262
rect 18602 20224 18658 20233
rect 19064 20198 19116 20204
rect 18602 20159 18658 20168
rect 19076 19718 19104 20198
rect 19064 19712 19116 19718
rect 19062 19680 19064 19689
rect 19116 19680 19118 19689
rect 19062 19615 19118 19624
rect 18972 19304 19024 19310
rect 19260 19258 19288 22063
rect 19352 21418 19380 22918
rect 19536 22166 19564 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 20088 25498 20116 27520
rect 20076 25492 20128 25498
rect 20076 25434 20128 25440
rect 20640 25226 20668 27520
rect 21088 25356 21140 25362
rect 21088 25298 21140 25304
rect 20628 25220 20680 25226
rect 20628 25162 20680 25168
rect 20168 25152 20220 25158
rect 20168 25094 20220 25100
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19800 24200 19852 24206
rect 19800 24142 19852 24148
rect 19812 23769 19840 24142
rect 19798 23760 19854 23769
rect 19798 23695 19854 23704
rect 19984 23520 20036 23526
rect 19984 23462 20036 23468
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19996 23304 20024 23462
rect 19904 23276 20024 23304
rect 19800 23248 19852 23254
rect 19798 23216 19800 23225
rect 19852 23216 19854 23225
rect 19798 23151 19854 23160
rect 19812 22710 19840 23151
rect 19800 22704 19852 22710
rect 19904 22681 19932 23276
rect 20076 23112 20128 23118
rect 20076 23054 20128 23060
rect 19984 23044 20036 23050
rect 19984 22986 20036 22992
rect 19800 22646 19852 22652
rect 19890 22672 19946 22681
rect 19890 22607 19946 22616
rect 19996 22438 20024 22986
rect 19984 22432 20036 22438
rect 19984 22374 20036 22380
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19996 22166 20024 22374
rect 20088 22234 20116 23054
rect 20180 22250 20208 25094
rect 21100 24886 21128 25298
rect 21088 24880 21140 24886
rect 20810 24848 20866 24857
rect 21192 24857 21220 27520
rect 21088 24822 21140 24828
rect 21178 24848 21234 24857
rect 20810 24783 20866 24792
rect 21178 24783 21234 24792
rect 20628 24744 20680 24750
rect 20628 24686 20680 24692
rect 20536 24676 20588 24682
rect 20536 24618 20588 24624
rect 20548 24585 20576 24618
rect 20534 24576 20590 24585
rect 20534 24511 20590 24520
rect 20444 24132 20496 24138
rect 20444 24074 20496 24080
rect 20352 24064 20404 24070
rect 20352 24006 20404 24012
rect 20364 23594 20392 24006
rect 20352 23588 20404 23594
rect 20352 23530 20404 23536
rect 20364 23254 20392 23530
rect 20352 23248 20404 23254
rect 20352 23190 20404 23196
rect 20076 22228 20128 22234
rect 20180 22222 20300 22250
rect 20076 22170 20128 22176
rect 19524 22160 19576 22166
rect 19524 22102 19576 22108
rect 19984 22160 20036 22166
rect 19984 22102 20036 22108
rect 20088 22114 20116 22170
rect 19432 22092 19484 22098
rect 20088 22086 20208 22114
rect 19432 22034 19484 22040
rect 19444 21978 19472 22034
rect 19892 22024 19944 22030
rect 19444 21950 19564 21978
rect 19892 21966 19944 21972
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 19340 21412 19392 21418
rect 19340 21354 19392 21360
rect 19338 21176 19394 21185
rect 19338 21111 19394 21120
rect 19352 21010 19380 21111
rect 19444 21026 19472 21830
rect 19536 21146 19564 21950
rect 19904 21690 19932 21966
rect 19892 21684 19944 21690
rect 19892 21626 19944 21632
rect 19984 21616 20036 21622
rect 19984 21558 20036 21564
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19524 21140 19576 21146
rect 19524 21082 19576 21088
rect 19340 21004 19392 21010
rect 19444 20998 19564 21026
rect 19340 20946 19392 20952
rect 19352 19990 19380 20946
rect 19340 19984 19392 19990
rect 19340 19926 19392 19932
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 18972 19246 19024 19252
rect 18602 19136 18658 19145
rect 18602 19071 18658 19080
rect 18616 18970 18644 19071
rect 18604 18964 18656 18970
rect 18604 18906 18656 18912
rect 18604 18080 18656 18086
rect 18602 18048 18604 18057
rect 18656 18048 18658 18057
rect 18602 17983 18658 17992
rect 18984 17882 19012 19246
rect 19168 19230 19288 19258
rect 18972 17876 19024 17882
rect 18972 17818 19024 17824
rect 18418 17232 18474 17241
rect 18418 17167 18474 17176
rect 18328 16720 18380 16726
rect 18328 16662 18380 16668
rect 18340 16425 18368 16662
rect 18326 16416 18382 16425
rect 18326 16351 18382 16360
rect 18340 16250 18368 16351
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 18432 16096 18460 17167
rect 19168 16794 19196 19230
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 19260 17513 19288 19110
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 19352 18290 19380 18702
rect 19444 18426 19472 19314
rect 19536 19242 19564 20998
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19996 19310 20024 21558
rect 20076 21548 20128 21554
rect 20076 21490 20128 21496
rect 20088 21321 20116 21490
rect 20074 21312 20130 21321
rect 20074 21247 20130 21256
rect 20180 21010 20208 22086
rect 20272 22030 20300 22222
rect 20260 22024 20312 22030
rect 20260 21966 20312 21972
rect 20364 21486 20392 23190
rect 20456 22420 20484 24074
rect 20536 23724 20588 23730
rect 20536 23666 20588 23672
rect 20548 23361 20576 23666
rect 20534 23352 20590 23361
rect 20534 23287 20590 23296
rect 20536 22976 20588 22982
rect 20536 22918 20588 22924
rect 20548 22574 20576 22918
rect 20536 22568 20588 22574
rect 20536 22510 20588 22516
rect 20456 22392 20576 22420
rect 20352 21480 20404 21486
rect 20352 21422 20404 21428
rect 20442 21448 20498 21457
rect 20442 21383 20444 21392
rect 20496 21383 20498 21392
rect 20444 21354 20496 21360
rect 20260 21344 20312 21350
rect 20260 21286 20312 21292
rect 20272 21049 20300 21286
rect 20456 21146 20484 21354
rect 20444 21140 20496 21146
rect 20444 21082 20496 21088
rect 20258 21040 20314 21049
rect 20168 21004 20220 21010
rect 20258 20975 20314 20984
rect 20168 20946 20220 20952
rect 20260 20256 20312 20262
rect 20260 20198 20312 20204
rect 20168 19712 20220 19718
rect 20168 19654 20220 19660
rect 20180 19310 20208 19654
rect 20272 19514 20300 20198
rect 20548 20058 20576 22392
rect 20640 22098 20668 24686
rect 20824 24614 20852 24783
rect 20812 24608 20864 24614
rect 20812 24550 20864 24556
rect 21652 24449 21680 27520
rect 21732 25764 21784 25770
rect 21732 25706 21784 25712
rect 21638 24440 21694 24449
rect 21638 24375 21694 24384
rect 21454 23896 21510 23905
rect 21454 23831 21456 23840
rect 21508 23831 21510 23840
rect 21456 23802 21508 23808
rect 21548 23180 21600 23186
rect 21548 23122 21600 23128
rect 20810 23080 20866 23089
rect 20810 23015 20866 23024
rect 20824 22273 20852 23015
rect 21270 22808 21326 22817
rect 21270 22743 21326 22752
rect 21454 22808 21510 22817
rect 21454 22743 21510 22752
rect 20810 22264 20866 22273
rect 20810 22199 20866 22208
rect 21178 22128 21234 22137
rect 20628 22092 20680 22098
rect 20628 22034 20680 22040
rect 20904 22092 20956 22098
rect 21178 22063 21234 22072
rect 20904 22034 20956 22040
rect 20720 21888 20772 21894
rect 20720 21830 20772 21836
rect 20732 21554 20760 21830
rect 20720 21548 20772 21554
rect 20720 21490 20772 21496
rect 20916 21078 20944 22034
rect 21088 21888 21140 21894
rect 21086 21856 21088 21865
rect 21140 21856 21142 21865
rect 21086 21791 21142 21800
rect 20904 21072 20956 21078
rect 20904 21014 20956 21020
rect 20996 21004 21048 21010
rect 20996 20946 21048 20952
rect 20904 20936 20956 20942
rect 20904 20878 20956 20884
rect 20628 20324 20680 20330
rect 20680 20284 20760 20312
rect 20628 20266 20680 20272
rect 20536 20052 20588 20058
rect 20536 19994 20588 20000
rect 20260 19508 20312 19514
rect 20260 19450 20312 19456
rect 19984 19304 20036 19310
rect 19984 19246 20036 19252
rect 20168 19304 20220 19310
rect 20168 19246 20220 19252
rect 19524 19236 19576 19242
rect 19524 19178 19576 19184
rect 20076 19236 20128 19242
rect 20076 19178 20128 19184
rect 19536 18737 19564 19178
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19522 18728 19578 18737
rect 19522 18663 19578 18672
rect 19524 18624 19576 18630
rect 19524 18566 19576 18572
rect 19432 18420 19484 18426
rect 19432 18362 19484 18368
rect 19340 18284 19392 18290
rect 19340 18226 19392 18232
rect 19432 18148 19484 18154
rect 19536 18136 19564 18566
rect 19484 18108 19564 18136
rect 19432 18090 19484 18096
rect 19246 17504 19302 17513
rect 19246 17439 19302 17448
rect 19444 16998 19472 18090
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19524 17876 19576 17882
rect 19524 17818 19576 17824
rect 19536 17338 19564 17818
rect 19616 17808 19668 17814
rect 19614 17776 19616 17785
rect 19668 17776 19670 17785
rect 19614 17711 19670 17720
rect 19524 17332 19576 17338
rect 19524 17274 19576 17280
rect 19432 16992 19484 16998
rect 19432 16934 19484 16940
rect 19156 16788 19208 16794
rect 19156 16730 19208 16736
rect 18696 16652 18748 16658
rect 18696 16594 18748 16600
rect 18340 16068 18460 16096
rect 18234 14784 18290 14793
rect 18234 14719 18290 14728
rect 18340 14634 18368 16068
rect 18604 15904 18656 15910
rect 18602 15872 18604 15881
rect 18656 15872 18658 15881
rect 18602 15807 18658 15816
rect 18248 14606 18368 14634
rect 18420 14612 18472 14618
rect 17868 14544 17920 14550
rect 17868 14486 17920 14492
rect 17776 14000 17828 14006
rect 17776 13942 17828 13948
rect 17590 13560 17646 13569
rect 17590 13495 17646 13504
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17774 13152 17830 13161
rect 17604 12782 17632 13126
rect 17774 13087 17830 13096
rect 17592 12776 17644 12782
rect 17592 12718 17644 12724
rect 17236 12396 17356 12424
rect 16764 12378 16816 12384
rect 17224 12232 17276 12238
rect 17224 12174 17276 12180
rect 17236 11558 17264 12174
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 17224 11552 17276 11558
rect 17224 11494 17276 11500
rect 16684 11150 16712 11494
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16684 10810 16712 11086
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 16684 9722 16712 10746
rect 16960 10538 16988 11154
rect 16948 10532 17000 10538
rect 16948 10474 17000 10480
rect 16960 10198 16988 10474
rect 16948 10192 17000 10198
rect 16948 10134 17000 10140
rect 16672 9716 16724 9722
rect 16672 9658 16724 9664
rect 17224 9444 17276 9450
rect 17224 9386 17276 9392
rect 17236 9178 17264 9386
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 17328 8974 17356 12396
rect 17604 12374 17632 12718
rect 17788 12481 17816 13087
rect 17774 12472 17830 12481
rect 17774 12407 17830 12416
rect 17592 12368 17644 12374
rect 17592 12310 17644 12316
rect 17604 11898 17632 12310
rect 17960 12096 18012 12102
rect 17960 12038 18012 12044
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 17684 10600 17736 10606
rect 17684 10542 17736 10548
rect 17696 10198 17724 10542
rect 17868 10532 17920 10538
rect 17972 10520 18000 12038
rect 18052 10736 18104 10742
rect 18052 10678 18104 10684
rect 17920 10492 18000 10520
rect 17868 10474 17920 10480
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 17684 10192 17736 10198
rect 17684 10134 17736 10140
rect 17500 10056 17552 10062
rect 17500 9998 17552 10004
rect 17512 9722 17540 9998
rect 17500 9716 17552 9722
rect 17500 9658 17552 9664
rect 17696 9178 17724 10134
rect 17788 9586 17816 10406
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 17684 9172 17736 9178
rect 17684 9114 17736 9120
rect 17972 9042 18000 10492
rect 18064 9450 18092 10678
rect 18144 9648 18196 9654
rect 18144 9590 18196 9596
rect 18052 9444 18104 9450
rect 18052 9386 18104 9392
rect 17960 9036 18012 9042
rect 17960 8978 18012 8984
rect 17316 8968 17368 8974
rect 17316 8910 17368 8916
rect 18156 8430 18184 9590
rect 18144 8424 18196 8430
rect 16500 8350 16620 8378
rect 18248 8401 18276 14606
rect 18420 14554 18472 14560
rect 18432 13870 18460 14554
rect 18708 13977 18736 16594
rect 18970 16280 19026 16289
rect 18970 16215 19026 16224
rect 18880 16176 18932 16182
rect 18880 16118 18932 16124
rect 18892 15638 18920 16118
rect 18880 15632 18932 15638
rect 18880 15574 18932 15580
rect 18880 15428 18932 15434
rect 18880 15370 18932 15376
rect 18892 14618 18920 15370
rect 18880 14612 18932 14618
rect 18880 14554 18932 14560
rect 18694 13968 18750 13977
rect 18694 13903 18696 13912
rect 18748 13903 18750 13912
rect 18696 13874 18748 13880
rect 18420 13864 18472 13870
rect 18420 13806 18472 13812
rect 18708 13530 18736 13874
rect 18880 13796 18932 13802
rect 18880 13738 18932 13744
rect 18696 13524 18748 13530
rect 18696 13466 18748 13472
rect 18604 12708 18656 12714
rect 18604 12650 18656 12656
rect 18616 11898 18644 12650
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 18788 11620 18840 11626
rect 18788 11562 18840 11568
rect 18604 11552 18656 11558
rect 18602 11520 18604 11529
rect 18656 11520 18658 11529
rect 18602 11455 18658 11464
rect 18800 11393 18828 11562
rect 18786 11384 18842 11393
rect 18786 11319 18788 11328
rect 18840 11319 18842 11328
rect 18892 11336 18920 13738
rect 18984 11506 19012 16215
rect 19168 16046 19196 16730
rect 19444 16561 19472 16934
rect 19536 16794 19564 17274
rect 19628 17270 19656 17711
rect 19984 17672 20036 17678
rect 19982 17640 19984 17649
rect 20036 17640 20038 17649
rect 19982 17575 20038 17584
rect 19616 17264 19668 17270
rect 19616 17206 19668 17212
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19524 16788 19576 16794
rect 19524 16730 19576 16736
rect 19996 16726 20024 17575
rect 19984 16720 20036 16726
rect 19984 16662 20036 16668
rect 19430 16552 19486 16561
rect 19430 16487 19486 16496
rect 19156 16040 19208 16046
rect 20088 16017 20116 19178
rect 20180 18426 20208 19246
rect 20732 19174 20760 20284
rect 20916 20262 20944 20878
rect 21008 20602 21036 20946
rect 20996 20596 21048 20602
rect 20996 20538 21048 20544
rect 20904 20256 20956 20262
rect 20904 20198 20956 20204
rect 21008 19990 21036 20538
rect 21192 20058 21220 22063
rect 21180 20052 21232 20058
rect 21180 19994 21232 20000
rect 20996 19984 21048 19990
rect 20996 19926 21048 19932
rect 20812 19848 20864 19854
rect 20812 19790 20864 19796
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20824 18970 20852 19790
rect 20812 18964 20864 18970
rect 20812 18906 20864 18912
rect 21178 18864 21234 18873
rect 21178 18799 21180 18808
rect 21232 18799 21234 18808
rect 21180 18770 21232 18776
rect 20168 18420 20220 18426
rect 20168 18362 20220 18368
rect 20180 18329 20208 18362
rect 20166 18320 20222 18329
rect 20166 18255 20222 18264
rect 21192 17882 21220 18770
rect 21180 17876 21232 17882
rect 21180 17818 21232 17824
rect 20168 17536 20220 17542
rect 20168 17478 20220 17484
rect 19156 15982 19208 15988
rect 20074 16008 20130 16017
rect 19168 15586 19196 15982
rect 19984 15972 20036 15978
rect 20074 15943 20130 15952
rect 19984 15914 20036 15920
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19076 15558 19196 15586
rect 19076 13326 19104 15558
rect 19996 15502 20024 15914
rect 19156 15496 19208 15502
rect 19156 15438 19208 15444
rect 19984 15496 20036 15502
rect 19984 15438 20036 15444
rect 19168 14822 19196 15438
rect 19248 15360 19300 15366
rect 19248 15302 19300 15308
rect 19156 14816 19208 14822
rect 19156 14758 19208 14764
rect 19168 14550 19196 14758
rect 19260 14634 19288 15302
rect 19996 15162 20024 15438
rect 19984 15156 20036 15162
rect 19984 15098 20036 15104
rect 19984 14952 20036 14958
rect 19984 14894 20036 14900
rect 19524 14884 19576 14890
rect 19524 14826 19576 14832
rect 19260 14618 19380 14634
rect 19260 14612 19392 14618
rect 19260 14606 19340 14612
rect 19156 14544 19208 14550
rect 19156 14486 19208 14492
rect 19260 13530 19288 14606
rect 19340 14554 19392 14560
rect 19340 14476 19392 14482
rect 19340 14418 19392 14424
rect 19248 13524 19300 13530
rect 19248 13466 19300 13472
rect 19352 13462 19380 14418
rect 19536 14006 19564 14826
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19892 14408 19944 14414
rect 19892 14350 19944 14356
rect 19904 14074 19932 14350
rect 19892 14068 19944 14074
rect 19892 14010 19944 14016
rect 19524 14000 19576 14006
rect 19524 13942 19576 13948
rect 19996 13802 20024 14894
rect 19984 13796 20036 13802
rect 19984 13738 20036 13744
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19430 13560 19486 13569
rect 19622 13552 19918 13572
rect 19486 13518 19564 13546
rect 19996 13530 20024 13738
rect 19430 13495 19486 13504
rect 19340 13456 19392 13462
rect 19340 13398 19392 13404
rect 19432 13388 19484 13394
rect 19432 13330 19484 13336
rect 19064 13320 19116 13326
rect 19064 13262 19116 13268
rect 19076 12986 19104 13262
rect 19338 13016 19394 13025
rect 19064 12980 19116 12986
rect 19338 12951 19340 12960
rect 19064 12922 19116 12928
rect 19392 12951 19394 12960
rect 19340 12922 19392 12928
rect 19444 12306 19472 13330
rect 19536 13025 19564 13518
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 19708 13456 19760 13462
rect 19708 13398 19760 13404
rect 19522 13016 19578 13025
rect 19720 12986 19748 13398
rect 19800 13184 19852 13190
rect 19800 13126 19852 13132
rect 19522 12951 19578 12960
rect 19708 12980 19760 12986
rect 19708 12922 19760 12928
rect 19524 12912 19576 12918
rect 19524 12854 19576 12860
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19444 11762 19472 12242
rect 19432 11756 19484 11762
rect 19432 11698 19484 11704
rect 19430 11656 19486 11665
rect 19430 11591 19486 11600
rect 18984 11478 19104 11506
rect 18892 11308 19012 11336
rect 18788 11290 18840 11296
rect 18880 11076 18932 11082
rect 18880 11018 18932 11024
rect 18604 10464 18656 10470
rect 18604 10406 18656 10412
rect 18616 10266 18644 10406
rect 18786 10296 18842 10305
rect 18604 10260 18656 10266
rect 18786 10231 18788 10240
rect 18604 10202 18656 10208
rect 18840 10231 18842 10240
rect 18788 10202 18840 10208
rect 18616 8906 18644 10202
rect 18800 9586 18828 10202
rect 18788 9580 18840 9586
rect 18708 9540 18788 9568
rect 18708 9178 18736 9540
rect 18788 9522 18840 9528
rect 18892 9382 18920 11018
rect 18984 10169 19012 11308
rect 18970 10160 19026 10169
rect 18970 10095 19026 10104
rect 18880 9376 18932 9382
rect 18880 9318 18932 9324
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 18788 9104 18840 9110
rect 18788 9046 18840 9052
rect 18604 8900 18656 8906
rect 18604 8842 18656 8848
rect 18800 8634 18828 9046
rect 18880 8968 18932 8974
rect 18880 8910 18932 8916
rect 18788 8628 18840 8634
rect 18788 8570 18840 8576
rect 18144 8366 18196 8372
rect 18234 8392 18290 8401
rect 14554 8327 14556 8336
rect 14608 8327 14610 8336
rect 14556 8298 14608 8304
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 16592 7954 16620 8350
rect 18234 8327 18290 8336
rect 18510 8392 18566 8401
rect 18510 8327 18512 8336
rect 18564 8327 18566 8336
rect 18512 8298 18564 8304
rect 18892 8090 18920 8910
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 14016 7546 14044 7822
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 16960 7546 16988 7890
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 13912 7540 13964 7546
rect 13912 7482 13964 7488
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 13832 7398 14044 7426
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9956 6996 10008 7002
rect 9956 6938 10008 6944
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 9600 6458 9720 6474
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 4988 6452 5040 6458
rect 4988 6394 5040 6400
rect 9588 6452 9720 6458
rect 9640 6446 9720 6452
rect 9588 6394 9640 6400
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 8114 3088 8170 3097
rect 8114 3023 8170 3032
rect 8128 2990 8156 3023
rect 8116 2984 8168 2990
rect 8116 2926 8168 2932
rect 8208 2916 8260 2922
rect 8208 2858 8260 2864
rect 8220 2650 8248 2858
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 7564 2304 7616 2310
rect 7564 2246 7616 2252
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 7576 1465 7604 2246
rect 8864 1601 8892 6054
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 8850 1592 8906 1601
rect 8850 1527 8906 1536
rect 7562 1456 7618 1465
rect 7562 1391 7618 1400
rect 14016 480 14044 7398
rect 17236 7342 17264 7822
rect 17224 7336 17276 7342
rect 17224 7278 17276 7284
rect 18234 7304 18290 7313
rect 18234 7239 18290 7248
rect 18248 7206 18276 7239
rect 18236 7200 18288 7206
rect 18236 7142 18288 7148
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 19076 5817 19104 11478
rect 19340 11280 19392 11286
rect 19340 11222 19392 11228
rect 19154 9752 19210 9761
rect 19352 9738 19380 11222
rect 19444 11150 19472 11591
rect 19536 11558 19564 12854
rect 19812 12782 19840 13126
rect 19800 12776 19852 12782
rect 19852 12736 20024 12764
rect 19800 12718 19852 12724
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19996 12442 20024 12736
rect 20076 12708 20128 12714
rect 20076 12650 20128 12656
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 20088 12102 20116 12650
rect 20076 12096 20128 12102
rect 20076 12038 20128 12044
rect 19524 11552 19576 11558
rect 19524 11494 19576 11500
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19524 11212 19576 11218
rect 19524 11154 19576 11160
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19210 9710 19380 9738
rect 19154 9687 19210 9696
rect 19168 9654 19196 9687
rect 19444 9654 19472 11086
rect 19536 11014 19564 11154
rect 19524 11008 19576 11014
rect 19524 10950 19576 10956
rect 19536 10538 19564 10950
rect 19614 10840 19670 10849
rect 19614 10775 19616 10784
rect 19668 10775 19670 10784
rect 19616 10746 19668 10752
rect 19628 10538 19656 10746
rect 20088 10606 20116 12038
rect 20076 10600 20128 10606
rect 20076 10542 20128 10548
rect 19524 10532 19576 10538
rect 19524 10474 19576 10480
rect 19616 10532 19668 10538
rect 19616 10474 19668 10480
rect 19984 10532 20036 10538
rect 19984 10474 20036 10480
rect 19536 10266 19564 10474
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19524 10260 19576 10266
rect 19524 10202 19576 10208
rect 19892 9920 19944 9926
rect 19996 9908 20024 10474
rect 19944 9880 20024 9908
rect 19892 9862 19944 9868
rect 19156 9648 19208 9654
rect 19156 9590 19208 9596
rect 19432 9648 19484 9654
rect 19904 9625 19932 9862
rect 19432 9590 19484 9596
rect 19890 9616 19946 9625
rect 19890 9551 19946 9560
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 20180 9217 20208 17478
rect 20352 17264 20404 17270
rect 20352 17206 20404 17212
rect 20258 13424 20314 13433
rect 20258 13359 20314 13368
rect 20272 13161 20300 13359
rect 20258 13152 20314 13161
rect 20258 13087 20314 13096
rect 20260 10464 20312 10470
rect 20260 10406 20312 10412
rect 20272 9897 20300 10406
rect 20258 9888 20314 9897
rect 20258 9823 20314 9832
rect 20364 9353 20392 17206
rect 20994 17096 21050 17105
rect 20994 17031 20996 17040
rect 21048 17031 21050 17040
rect 20996 17002 21048 17008
rect 20904 16040 20956 16046
rect 20904 15982 20956 15988
rect 20916 15910 20944 15982
rect 21088 15972 21140 15978
rect 21088 15914 21140 15920
rect 20904 15904 20956 15910
rect 20904 15846 20956 15852
rect 20812 15564 20864 15570
rect 20812 15506 20864 15512
rect 20720 15360 20772 15366
rect 20720 15302 20772 15308
rect 20628 15088 20680 15094
rect 20628 15030 20680 15036
rect 20640 14482 20668 15030
rect 20732 14890 20760 15302
rect 20824 15162 20852 15506
rect 20812 15156 20864 15162
rect 20812 15098 20864 15104
rect 20720 14884 20772 14890
rect 20720 14826 20772 14832
rect 20628 14476 20680 14482
rect 20628 14418 20680 14424
rect 20916 14414 20944 15846
rect 21100 15609 21128 15914
rect 21284 15706 21312 22743
rect 21364 21548 21416 21554
rect 21364 21490 21416 21496
rect 21376 18902 21404 21490
rect 21468 18970 21496 22743
rect 21560 22506 21588 23122
rect 21638 22944 21694 22953
rect 21638 22879 21694 22888
rect 21652 22778 21680 22879
rect 21640 22772 21692 22778
rect 21640 22714 21692 22720
rect 21548 22500 21600 22506
rect 21548 22442 21600 22448
rect 21560 22166 21588 22442
rect 21548 22160 21600 22166
rect 21548 22102 21600 22108
rect 21744 19922 21772 25706
rect 22204 25498 22232 27520
rect 22192 25492 22244 25498
rect 22192 25434 22244 25440
rect 22652 25356 22704 25362
rect 22652 25298 22704 25304
rect 22664 24954 22692 25298
rect 22652 24948 22704 24954
rect 22652 24890 22704 24896
rect 21914 24712 21970 24721
rect 21914 24647 21970 24656
rect 21928 24614 21956 24647
rect 21916 24608 21968 24614
rect 21916 24550 21968 24556
rect 21916 24268 21968 24274
rect 21916 24210 21968 24216
rect 21928 23905 21956 24210
rect 22100 24200 22152 24206
rect 22100 24142 22152 24148
rect 21914 23896 21970 23905
rect 21914 23831 21970 23840
rect 21824 23656 21876 23662
rect 21822 23624 21824 23633
rect 21876 23624 21878 23633
rect 21822 23559 21878 23568
rect 22008 23588 22060 23594
rect 21836 23526 21864 23559
rect 22008 23530 22060 23536
rect 21824 23520 21876 23526
rect 21824 23462 21876 23468
rect 21916 22092 21968 22098
rect 21916 22034 21968 22040
rect 21928 21690 21956 22034
rect 21916 21684 21968 21690
rect 21916 21626 21968 21632
rect 22020 21418 22048 23530
rect 22008 21412 22060 21418
rect 22008 21354 22060 21360
rect 22112 20398 22140 24142
rect 22284 23248 22336 23254
rect 22284 23190 22336 23196
rect 22296 22438 22324 23190
rect 22284 22432 22336 22438
rect 22284 22374 22336 22380
rect 22192 21548 22244 21554
rect 22192 21490 22244 21496
rect 22204 20602 22232 21490
rect 22296 21146 22324 22374
rect 22756 22137 22784 27520
rect 23308 24721 23336 27520
rect 23584 26382 23612 27639
rect 23846 27520 23902 28000
rect 24398 27520 24454 28000
rect 24858 27520 24914 28000
rect 25410 27520 25466 28000
rect 25962 27520 26018 28000
rect 26514 27520 26570 28000
rect 27066 27520 27122 28000
rect 27618 27520 27674 28000
rect 23572 26376 23624 26382
rect 23572 26318 23624 26324
rect 23480 25424 23532 25430
rect 23480 25366 23532 25372
rect 23492 24818 23520 25366
rect 23860 24970 23888 27520
rect 24306 26616 24362 26625
rect 24306 26551 24362 26560
rect 24320 26314 24348 26551
rect 24308 26308 24360 26314
rect 24308 26250 24360 26256
rect 23938 25528 23994 25537
rect 23938 25463 23994 25472
rect 23768 24942 23888 24970
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 23294 24712 23350 24721
rect 23294 24647 23350 24656
rect 23112 24336 23164 24342
rect 23112 24278 23164 24284
rect 22928 24064 22980 24070
rect 23124 24041 23152 24278
rect 23572 24200 23624 24206
rect 23572 24142 23624 24148
rect 23388 24064 23440 24070
rect 22928 24006 22980 24012
rect 23110 24032 23166 24041
rect 22940 23594 22968 24006
rect 23388 24006 23440 24012
rect 23110 23967 23166 23976
rect 23124 23866 23152 23967
rect 23112 23860 23164 23866
rect 23112 23802 23164 23808
rect 23020 23792 23072 23798
rect 23020 23734 23072 23740
rect 22928 23588 22980 23594
rect 22928 23530 22980 23536
rect 23032 23186 23060 23734
rect 23400 23338 23428 24006
rect 23400 23310 23520 23338
rect 23584 23322 23612 24142
rect 23492 23254 23520 23310
rect 23572 23316 23624 23322
rect 23572 23258 23624 23264
rect 23388 23248 23440 23254
rect 23388 23190 23440 23196
rect 23480 23248 23532 23254
rect 23480 23190 23532 23196
rect 23020 23180 23072 23186
rect 23020 23122 23072 23128
rect 22834 23080 22890 23089
rect 22834 23015 22890 23024
rect 22742 22128 22798 22137
rect 22742 22063 22798 22072
rect 22652 21888 22704 21894
rect 22652 21830 22704 21836
rect 22664 21486 22692 21830
rect 22652 21480 22704 21486
rect 22652 21422 22704 21428
rect 22560 21344 22612 21350
rect 22560 21286 22612 21292
rect 22572 21146 22600 21286
rect 22284 21140 22336 21146
rect 22284 21082 22336 21088
rect 22560 21140 22612 21146
rect 22560 21082 22612 21088
rect 22192 20596 22244 20602
rect 22192 20538 22244 20544
rect 22664 20466 22692 21422
rect 22848 20602 22876 23015
rect 23032 22778 23060 23122
rect 23020 22772 23072 22778
rect 23020 22714 23072 22720
rect 23294 22672 23350 22681
rect 23294 22607 23350 22616
rect 23202 22536 23258 22545
rect 23202 22471 23258 22480
rect 23110 22400 23166 22409
rect 23110 22335 23166 22344
rect 23124 22234 23152 22335
rect 23112 22228 23164 22234
rect 23112 22170 23164 22176
rect 23020 22024 23072 22030
rect 23020 21966 23072 21972
rect 22928 21888 22980 21894
rect 22928 21830 22980 21836
rect 22836 20596 22888 20602
rect 22836 20538 22888 20544
rect 22652 20460 22704 20466
rect 22652 20402 22704 20408
rect 22100 20392 22152 20398
rect 22100 20334 22152 20340
rect 22112 20058 22140 20334
rect 22376 20256 22428 20262
rect 22376 20198 22428 20204
rect 22100 20052 22152 20058
rect 22100 19994 22152 20000
rect 22388 19922 22416 20198
rect 21732 19916 21784 19922
rect 21732 19858 21784 19864
rect 22376 19916 22428 19922
rect 22376 19858 22428 19864
rect 22388 19514 22416 19858
rect 22376 19508 22428 19514
rect 22376 19450 22428 19456
rect 21546 19272 21602 19281
rect 21546 19207 21602 19216
rect 21456 18964 21508 18970
rect 21456 18906 21508 18912
rect 21364 18896 21416 18902
rect 21364 18838 21416 18844
rect 21376 18426 21404 18838
rect 21364 18420 21416 18426
rect 21364 18362 21416 18368
rect 21456 17740 21508 17746
rect 21456 17682 21508 17688
rect 21468 17338 21496 17682
rect 21456 17332 21508 17338
rect 21456 17274 21508 17280
rect 21272 15700 21324 15706
rect 21272 15642 21324 15648
rect 21086 15600 21142 15609
rect 21086 15535 21142 15544
rect 20996 15428 21048 15434
rect 20996 15370 21048 15376
rect 21008 15026 21036 15370
rect 21284 15162 21312 15642
rect 21272 15156 21324 15162
rect 21272 15098 21324 15104
rect 20996 15020 21048 15026
rect 20996 14962 21048 14968
rect 21180 14884 21232 14890
rect 21180 14826 21232 14832
rect 21192 14618 21220 14826
rect 21180 14612 21232 14618
rect 21180 14554 21232 14560
rect 20996 14476 21048 14482
rect 20996 14418 21048 14424
rect 20904 14408 20956 14414
rect 20904 14350 20956 14356
rect 20536 14272 20588 14278
rect 20536 14214 20588 14220
rect 20444 10532 20496 10538
rect 20444 10474 20496 10480
rect 20456 9654 20484 10474
rect 20444 9648 20496 9654
rect 20444 9590 20496 9596
rect 20350 9344 20406 9353
rect 20350 9279 20406 9288
rect 20166 9208 20222 9217
rect 20166 9143 20222 9152
rect 19156 8900 19208 8906
rect 19156 8842 19208 8848
rect 19168 8362 19196 8842
rect 19156 8356 19208 8362
rect 19156 8298 19208 8304
rect 19168 7449 19196 8298
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 20548 7732 20576 14214
rect 20916 13870 20944 14350
rect 21008 14074 21036 14418
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 20904 13864 20956 13870
rect 20904 13806 20956 13812
rect 20812 12640 20864 12646
rect 20812 12582 20864 12588
rect 20824 12345 20852 12582
rect 20810 12336 20866 12345
rect 20810 12271 20866 12280
rect 20916 12238 20944 13806
rect 21008 13530 21036 14010
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 21456 13184 21508 13190
rect 21456 13126 21508 13132
rect 21088 12912 21140 12918
rect 21088 12854 21140 12860
rect 20994 12336 21050 12345
rect 20994 12271 21050 12280
rect 20904 12232 20956 12238
rect 20904 12174 20956 12180
rect 20812 11824 20864 11830
rect 20812 11766 20864 11772
rect 20824 10810 20852 11766
rect 21008 10985 21036 12271
rect 21100 11762 21128 12854
rect 21468 12850 21496 13126
rect 21456 12844 21508 12850
rect 21456 12786 21508 12792
rect 21560 12714 21588 19207
rect 22388 18834 22416 19450
rect 22560 19168 22612 19174
rect 22560 19110 22612 19116
rect 22466 18864 22522 18873
rect 22376 18828 22428 18834
rect 22466 18799 22522 18808
rect 22376 18770 22428 18776
rect 22100 18624 22152 18630
rect 22100 18566 22152 18572
rect 22112 18222 22140 18566
rect 22388 18358 22416 18770
rect 22192 18352 22244 18358
rect 22192 18294 22244 18300
rect 22376 18352 22428 18358
rect 22376 18294 22428 18300
rect 22100 18216 22152 18222
rect 22100 18158 22152 18164
rect 22100 18080 22152 18086
rect 22100 18022 22152 18028
rect 22112 17882 22140 18022
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 22204 17678 22232 18294
rect 22192 17672 22244 17678
rect 22192 17614 22244 17620
rect 22204 17338 22232 17614
rect 22192 17332 22244 17338
rect 22192 17274 22244 17280
rect 21824 16992 21876 16998
rect 21824 16934 21876 16940
rect 21836 16794 21864 16934
rect 21824 16788 21876 16794
rect 21824 16730 21876 16736
rect 22376 16788 22428 16794
rect 22376 16730 22428 16736
rect 22284 16720 22336 16726
rect 22284 16662 22336 16668
rect 21824 16448 21876 16454
rect 21824 16390 21876 16396
rect 21640 15156 21692 15162
rect 21640 15098 21692 15104
rect 21548 12708 21600 12714
rect 21548 12650 21600 12656
rect 21180 12300 21232 12306
rect 21180 12242 21232 12248
rect 21192 12209 21220 12242
rect 21178 12200 21234 12209
rect 21178 12135 21234 12144
rect 21192 11898 21220 12135
rect 21180 11892 21232 11898
rect 21180 11834 21232 11840
rect 21088 11756 21140 11762
rect 21088 11698 21140 11704
rect 21652 11665 21680 15098
rect 21836 15065 21864 16390
rect 22296 15978 22324 16662
rect 22284 15972 22336 15978
rect 22284 15914 22336 15920
rect 21916 15904 21968 15910
rect 21916 15846 21968 15852
rect 21928 15502 21956 15846
rect 22296 15706 22324 15914
rect 22284 15700 22336 15706
rect 22284 15642 22336 15648
rect 22008 15564 22060 15570
rect 22008 15506 22060 15512
rect 21916 15496 21968 15502
rect 21916 15438 21968 15444
rect 21928 15162 21956 15438
rect 21916 15156 21968 15162
rect 21916 15098 21968 15104
rect 21822 15056 21878 15065
rect 22020 15042 22048 15506
rect 22020 15026 22140 15042
rect 22020 15020 22152 15026
rect 22020 15014 22100 15020
rect 21822 14991 21878 15000
rect 22100 14962 22152 14968
rect 22100 14816 22152 14822
rect 22100 14758 22152 14764
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 22020 12424 22048 12786
rect 22112 12782 22140 14758
rect 22284 14272 22336 14278
rect 22284 14214 22336 14220
rect 22296 13977 22324 14214
rect 22282 13968 22338 13977
rect 22282 13903 22338 13912
rect 22190 13016 22246 13025
rect 22190 12951 22192 12960
rect 22244 12951 22246 12960
rect 22192 12922 22244 12928
rect 22100 12776 22152 12782
rect 22100 12718 22152 12724
rect 22100 12436 22152 12442
rect 22020 12396 22100 12424
rect 22100 12378 22152 12384
rect 21824 12096 21876 12102
rect 21824 12038 21876 12044
rect 21836 11830 21864 12038
rect 21824 11824 21876 11830
rect 21824 11766 21876 11772
rect 21638 11656 21694 11665
rect 21364 11620 21416 11626
rect 21638 11591 21694 11600
rect 21364 11562 21416 11568
rect 21088 11552 21140 11558
rect 21088 11494 21140 11500
rect 21100 11354 21128 11494
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 21376 11218 21404 11562
rect 21836 11558 21864 11766
rect 21824 11552 21876 11558
rect 21824 11494 21876 11500
rect 21364 11212 21416 11218
rect 21364 11154 21416 11160
rect 21836 11150 21864 11494
rect 22100 11348 22152 11354
rect 22020 11308 22100 11336
rect 21824 11144 21876 11150
rect 21824 11086 21876 11092
rect 21456 11008 21508 11014
rect 20994 10976 21050 10985
rect 21456 10950 21508 10956
rect 20994 10911 21050 10920
rect 20812 10804 20864 10810
rect 20812 10746 20864 10752
rect 20628 10736 20680 10742
rect 20628 10678 20680 10684
rect 20720 10736 20772 10742
rect 20720 10678 20772 10684
rect 20640 9602 20668 10678
rect 20732 10062 20760 10678
rect 20824 10470 20852 10746
rect 21468 10538 21496 10950
rect 21836 10810 21864 11086
rect 21824 10804 21876 10810
rect 21824 10746 21876 10752
rect 21916 10736 21968 10742
rect 21916 10678 21968 10684
rect 20904 10532 20956 10538
rect 20904 10474 20956 10480
rect 21456 10532 21508 10538
rect 21456 10474 21508 10480
rect 20812 10464 20864 10470
rect 20812 10406 20864 10412
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20732 9722 20760 9998
rect 20916 9722 20944 10474
rect 21732 10124 21784 10130
rect 21732 10066 21784 10072
rect 20720 9716 20772 9722
rect 20720 9658 20772 9664
rect 20904 9716 20956 9722
rect 20904 9658 20956 9664
rect 21744 9654 21772 10066
rect 21928 9761 21956 10678
rect 22020 10674 22048 11308
rect 22100 11290 22152 11296
rect 22100 11212 22152 11218
rect 22100 11154 22152 11160
rect 22008 10668 22060 10674
rect 22008 10610 22060 10616
rect 22112 10470 22140 11154
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 22112 9926 22140 10406
rect 22100 9920 22152 9926
rect 22020 9868 22100 9874
rect 22020 9862 22152 9868
rect 22020 9846 22140 9862
rect 21914 9752 21970 9761
rect 21914 9687 21970 9696
rect 21732 9648 21784 9654
rect 20640 9574 20760 9602
rect 21732 9590 21784 9596
rect 20732 9518 20760 9574
rect 20720 9512 20772 9518
rect 20720 9454 20772 9460
rect 21546 9480 21602 9489
rect 21546 9415 21602 9424
rect 21088 9376 21140 9382
rect 21088 9318 21140 9324
rect 21100 8906 21128 9318
rect 21560 9110 21588 9415
rect 21548 9104 21600 9110
rect 21362 9072 21418 9081
rect 21548 9046 21600 9052
rect 21362 9007 21364 9016
rect 21416 9007 21418 9016
rect 21364 8978 21416 8984
rect 21088 8900 21140 8906
rect 21088 8842 21140 8848
rect 21376 8498 21404 8978
rect 21560 8634 21588 9046
rect 21744 8974 21772 9590
rect 22020 9586 22048 9846
rect 22008 9580 22060 9586
rect 22008 9522 22060 9528
rect 21732 8968 21784 8974
rect 21732 8910 21784 8916
rect 21744 8634 21772 8910
rect 21548 8628 21600 8634
rect 21548 8570 21600 8576
rect 21732 8628 21784 8634
rect 21732 8570 21784 8576
rect 21364 8492 21416 8498
rect 21364 8434 21416 8440
rect 20548 7704 20760 7732
rect 19154 7440 19210 7449
rect 19154 7375 19210 7384
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19062 5808 19118 5817
rect 20732 5778 20760 7704
rect 21376 6089 21404 8434
rect 22204 6905 22232 12922
rect 22388 9874 22416 16730
rect 22480 16590 22508 18799
rect 22572 18290 22600 19110
rect 22650 18456 22706 18465
rect 22650 18391 22706 18400
rect 22560 18284 22612 18290
rect 22560 18226 22612 18232
rect 22560 17196 22612 17202
rect 22560 17138 22612 17144
rect 22572 16726 22600 17138
rect 22560 16720 22612 16726
rect 22560 16662 22612 16668
rect 22468 16584 22520 16590
rect 22468 16526 22520 16532
rect 22480 16425 22508 16526
rect 22466 16416 22522 16425
rect 22466 16351 22522 16360
rect 22480 15706 22508 16351
rect 22468 15700 22520 15706
rect 22468 15642 22520 15648
rect 22664 15638 22692 18391
rect 22836 17264 22888 17270
rect 22836 17206 22888 17212
rect 22744 17060 22796 17066
rect 22744 17002 22796 17008
rect 22756 16658 22784 17002
rect 22744 16652 22796 16658
rect 22744 16594 22796 16600
rect 22652 15632 22704 15638
rect 22652 15574 22704 15580
rect 22664 15162 22692 15574
rect 22652 15156 22704 15162
rect 22652 15098 22704 15104
rect 22560 13456 22612 13462
rect 22560 13398 22612 13404
rect 22468 13388 22520 13394
rect 22468 13330 22520 13336
rect 22480 12918 22508 13330
rect 22572 12986 22600 13398
rect 22560 12980 22612 12986
rect 22560 12922 22612 12928
rect 22468 12912 22520 12918
rect 22664 12866 22692 15098
rect 22756 14498 22784 16594
rect 22848 14890 22876 17206
rect 22836 14884 22888 14890
rect 22836 14826 22888 14832
rect 22848 14618 22876 14826
rect 22836 14612 22888 14618
rect 22836 14554 22888 14560
rect 22756 14470 22876 14498
rect 22848 14278 22876 14470
rect 22836 14272 22888 14278
rect 22836 14214 22888 14220
rect 22848 13462 22876 14214
rect 22940 13546 22968 21830
rect 23032 21457 23060 21966
rect 23124 21690 23152 22170
rect 23112 21684 23164 21690
rect 23112 21626 23164 21632
rect 23018 21448 23074 21457
rect 23018 21383 23020 21392
rect 23072 21383 23074 21392
rect 23020 21354 23072 21360
rect 23032 21323 23060 21354
rect 23020 19916 23072 19922
rect 23020 19858 23072 19864
rect 23032 19514 23060 19858
rect 23020 19508 23072 19514
rect 23020 19450 23072 19456
rect 23110 19000 23166 19009
rect 23110 18935 23166 18944
rect 23020 17332 23072 17338
rect 23020 17274 23072 17280
rect 23032 16590 23060 17274
rect 23020 16584 23072 16590
rect 23020 16526 23072 16532
rect 23032 16250 23060 16526
rect 23124 16436 23152 18935
rect 23216 16561 23244 22471
rect 23308 22098 23336 22607
rect 23400 22114 23428 23190
rect 23492 22234 23520 23190
rect 23572 22976 23624 22982
rect 23572 22918 23624 22924
rect 23480 22228 23532 22234
rect 23480 22170 23532 22176
rect 23296 22092 23348 22098
rect 23400 22086 23520 22114
rect 23296 22034 23348 22040
rect 23308 21894 23336 22034
rect 23296 21888 23348 21894
rect 23296 21830 23348 21836
rect 23296 21616 23348 21622
rect 23492 21593 23520 22086
rect 23296 21558 23348 21564
rect 23478 21584 23534 21593
rect 23308 21049 23336 21558
rect 23478 21519 23534 21528
rect 23584 21162 23612 22918
rect 23768 22817 23796 24942
rect 23846 24848 23902 24857
rect 23846 24783 23902 24792
rect 23860 24614 23888 24783
rect 23848 24608 23900 24614
rect 23848 24550 23900 24556
rect 23754 22808 23810 22817
rect 23754 22743 23810 22752
rect 23756 22704 23808 22710
rect 23756 22646 23808 22652
rect 23664 22500 23716 22506
rect 23664 22442 23716 22448
rect 23676 21962 23704 22442
rect 23664 21956 23716 21962
rect 23664 21898 23716 21904
rect 23664 21616 23716 21622
rect 23664 21558 23716 21564
rect 23400 21146 23612 21162
rect 23388 21140 23612 21146
rect 23440 21134 23612 21140
rect 23388 21082 23440 21088
rect 23294 21040 23350 21049
rect 23294 20975 23350 20984
rect 23480 20800 23532 20806
rect 23480 20742 23532 20748
rect 23388 19712 23440 19718
rect 23388 19654 23440 19660
rect 23400 18902 23428 19654
rect 23388 18896 23440 18902
rect 23388 18838 23440 18844
rect 23388 18692 23440 18698
rect 23388 18634 23440 18640
rect 23400 17626 23428 18634
rect 23492 18426 23520 20742
rect 23572 18624 23624 18630
rect 23572 18566 23624 18572
rect 23480 18420 23532 18426
rect 23480 18362 23532 18368
rect 23480 17808 23532 17814
rect 23478 17776 23480 17785
rect 23532 17776 23534 17785
rect 23584 17746 23612 18566
rect 23478 17711 23534 17720
rect 23572 17740 23624 17746
rect 23572 17682 23624 17688
rect 23400 17598 23520 17626
rect 23388 17536 23440 17542
rect 23388 17478 23440 17484
rect 23400 16998 23428 17478
rect 23388 16992 23440 16998
rect 23388 16934 23440 16940
rect 23400 16794 23428 16934
rect 23388 16788 23440 16794
rect 23388 16730 23440 16736
rect 23296 16720 23348 16726
rect 23296 16662 23348 16668
rect 23202 16552 23258 16561
rect 23202 16487 23258 16496
rect 23124 16408 23244 16436
rect 23020 16244 23072 16250
rect 23020 16186 23072 16192
rect 23032 16046 23060 16186
rect 23020 16040 23072 16046
rect 23020 15982 23072 15988
rect 23110 15872 23166 15881
rect 23110 15807 23166 15816
rect 23020 15632 23072 15638
rect 23020 15574 23072 15580
rect 23032 14822 23060 15574
rect 23020 14816 23072 14822
rect 23020 14758 23072 14764
rect 23018 13560 23074 13569
rect 22940 13518 23018 13546
rect 23018 13495 23074 13504
rect 22836 13456 22888 13462
rect 22836 13398 22888 13404
rect 22848 12986 22876 13398
rect 22836 12980 22888 12986
rect 22836 12922 22888 12928
rect 22468 12854 22520 12860
rect 22572 12838 22692 12866
rect 22388 9846 22508 9874
rect 22374 9616 22430 9625
rect 22374 9551 22376 9560
rect 22428 9551 22430 9560
rect 22376 9522 22428 9528
rect 22480 8634 22508 9846
rect 22468 8628 22520 8634
rect 22468 8570 22520 8576
rect 22190 6896 22246 6905
rect 22190 6831 22246 6840
rect 21362 6080 21418 6089
rect 21362 6015 21418 6024
rect 19062 5743 19118 5752
rect 20720 5772 20772 5778
rect 20720 5714 20772 5720
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 20732 5370 20760 5714
rect 21088 5704 21140 5710
rect 21088 5646 21140 5652
rect 20720 5364 20772 5370
rect 20720 5306 20772 5312
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 21100 4690 21128 5646
rect 22572 5273 22600 12838
rect 22652 12776 22704 12782
rect 22652 12718 22704 12724
rect 22664 10033 22692 12718
rect 23032 10198 23060 13495
rect 23124 12782 23152 15807
rect 23216 15638 23244 16408
rect 23204 15632 23256 15638
rect 23204 15574 23256 15580
rect 23308 15484 23336 16662
rect 23492 15910 23520 17598
rect 23584 16114 23612 17682
rect 23676 16969 23704 21558
rect 23768 21554 23796 22646
rect 23848 22160 23900 22166
rect 23848 22102 23900 22108
rect 23756 21548 23808 21554
rect 23756 21490 23808 21496
rect 23860 21400 23888 22102
rect 23952 21622 23980 25463
rect 24032 25356 24084 25362
rect 24032 25298 24084 25304
rect 24044 24614 24072 25298
rect 24412 25242 24440 27520
rect 24766 27160 24822 27169
rect 24766 27095 24822 27104
rect 24780 26450 24808 27095
rect 24768 26444 24820 26450
rect 24768 26386 24820 26392
rect 24766 26072 24822 26081
rect 24766 26007 24822 26016
rect 24412 25214 24716 25242
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24032 24608 24084 24614
rect 24032 24550 24084 24556
rect 24214 24576 24270 24585
rect 24044 23225 24072 24550
rect 24214 24511 24270 24520
rect 24228 24274 24256 24511
rect 24216 24268 24268 24274
rect 24216 24210 24268 24216
rect 24122 24168 24178 24177
rect 24122 24103 24178 24112
rect 24030 23216 24086 23225
rect 24030 23151 24086 23160
rect 24032 23112 24084 23118
rect 24032 23054 24084 23060
rect 24044 22574 24072 23054
rect 24032 22568 24084 22574
rect 24032 22510 24084 22516
rect 24044 22166 24072 22510
rect 24032 22160 24084 22166
rect 24032 22102 24084 22108
rect 24032 21888 24084 21894
rect 24032 21830 24084 21836
rect 23940 21616 23992 21622
rect 23940 21558 23992 21564
rect 23940 21412 23992 21418
rect 23860 21372 23940 21400
rect 23940 21354 23992 21360
rect 23756 21344 23808 21350
rect 23756 21286 23808 21292
rect 23768 20398 23796 21286
rect 23846 21176 23902 21185
rect 23846 21111 23902 21120
rect 23756 20392 23808 20398
rect 23756 20334 23808 20340
rect 23768 19990 23796 20334
rect 23756 19984 23808 19990
rect 23756 19926 23808 19932
rect 23860 18698 23888 21111
rect 23952 19802 23980 21354
rect 24044 21010 24072 21830
rect 24136 21486 24164 24103
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24216 22976 24268 22982
rect 24216 22918 24268 22924
rect 24228 22506 24256 22918
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24688 22760 24716 25214
rect 24780 24886 24808 26007
rect 24768 24880 24820 24886
rect 24768 24822 24820 24828
rect 24872 24834 24900 27520
rect 25424 25498 25452 27520
rect 25976 25702 26004 27520
rect 25964 25696 26016 25702
rect 25964 25638 26016 25644
rect 25412 25492 25464 25498
rect 25412 25434 25464 25440
rect 25688 25356 25740 25362
rect 25688 25298 25740 25304
rect 24872 24806 25176 24834
rect 24768 24744 24820 24750
rect 24768 24686 24820 24692
rect 24950 24712 25006 24721
rect 24780 24313 24808 24686
rect 24950 24647 25006 24656
rect 24964 24614 24992 24647
rect 24952 24608 25004 24614
rect 24952 24550 25004 24556
rect 24858 24440 24914 24449
rect 24858 24375 24860 24384
rect 24912 24375 24914 24384
rect 24860 24346 24912 24352
rect 24766 24304 24822 24313
rect 24766 24239 24822 24248
rect 24952 24268 25004 24274
rect 24952 24210 25004 24216
rect 24766 23896 24822 23905
rect 24766 23831 24822 23840
rect 24780 23576 24808 23831
rect 24780 23548 24900 23576
rect 24596 22732 24716 22760
rect 24216 22500 24268 22506
rect 24216 22442 24268 22448
rect 24596 22166 24624 22732
rect 24676 22636 24728 22642
rect 24676 22578 24728 22584
rect 24216 22160 24268 22166
rect 24216 22102 24268 22108
rect 24584 22160 24636 22166
rect 24584 22102 24636 22108
rect 24228 21690 24256 22102
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24688 21690 24716 22578
rect 24768 22160 24820 22166
rect 24768 22102 24820 22108
rect 24216 21684 24268 21690
rect 24216 21626 24268 21632
rect 24676 21684 24728 21690
rect 24676 21626 24728 21632
rect 24214 21584 24270 21593
rect 24214 21519 24270 21528
rect 24124 21480 24176 21486
rect 24124 21422 24176 21428
rect 24124 21344 24176 21350
rect 24124 21286 24176 21292
rect 24032 21004 24084 21010
rect 24032 20946 24084 20952
rect 24044 20398 24072 20946
rect 24032 20392 24084 20398
rect 24032 20334 24084 20340
rect 24044 19990 24072 20334
rect 24032 19984 24084 19990
rect 24032 19926 24084 19932
rect 23952 19774 24072 19802
rect 24044 19310 24072 19774
rect 24032 19304 24084 19310
rect 24136 19281 24164 21286
rect 24228 21185 24256 21519
rect 24676 21480 24728 21486
rect 24676 21422 24728 21428
rect 24214 21176 24270 21185
rect 24214 21111 24270 21120
rect 24216 21072 24268 21078
rect 24216 21014 24268 21020
rect 24688 21026 24716 21422
rect 24780 21162 24808 22102
rect 24872 21486 24900 23548
rect 24964 23322 24992 24210
rect 25044 23520 25096 23526
rect 25044 23462 25096 23468
rect 24952 23316 25004 23322
rect 24952 23258 25004 23264
rect 24952 23180 25004 23186
rect 24952 23122 25004 23128
rect 24964 22778 24992 23122
rect 24952 22772 25004 22778
rect 24952 22714 25004 22720
rect 25056 22506 25084 23462
rect 25148 23089 25176 24806
rect 25700 24614 25728 25298
rect 25778 24984 25834 24993
rect 25778 24919 25834 24928
rect 25688 24608 25740 24614
rect 25688 24550 25740 24556
rect 25412 23860 25464 23866
rect 25412 23802 25464 23808
rect 25226 23488 25282 23497
rect 25226 23423 25282 23432
rect 25134 23080 25190 23089
rect 25134 23015 25190 23024
rect 25240 22658 25268 23423
rect 25320 22772 25372 22778
rect 25320 22714 25372 22720
rect 25148 22630 25268 22658
rect 25044 22500 25096 22506
rect 25044 22442 25096 22448
rect 24860 21480 24912 21486
rect 24860 21422 24912 21428
rect 25042 21448 25098 21457
rect 24872 21298 24900 21422
rect 25042 21383 25044 21392
rect 25096 21383 25098 21392
rect 25044 21354 25096 21360
rect 24872 21270 24992 21298
rect 24780 21146 24900 21162
rect 24780 21140 24912 21146
rect 24780 21134 24860 21140
rect 24860 21082 24912 21088
rect 24964 21078 24992 21270
rect 25056 21162 25084 21354
rect 25148 21350 25176 22630
rect 25226 21992 25282 22001
rect 25226 21927 25282 21936
rect 25136 21344 25188 21350
rect 25136 21286 25188 21292
rect 25056 21134 25176 21162
rect 24952 21072 25004 21078
rect 24228 20058 24256 21014
rect 24688 20998 24808 21026
rect 24952 21014 25004 21020
rect 24676 20936 24728 20942
rect 24676 20878 24728 20884
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24216 20052 24268 20058
rect 24216 19994 24268 20000
rect 24228 19514 24256 19994
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24216 19508 24268 19514
rect 24216 19450 24268 19456
rect 24688 19394 24716 20878
rect 24228 19366 24716 19394
rect 24032 19246 24084 19252
rect 24122 19272 24178 19281
rect 24044 19174 24072 19246
rect 24122 19207 24178 19216
rect 24032 19168 24084 19174
rect 23938 19136 23994 19145
rect 24032 19110 24084 19116
rect 23938 19071 23994 19080
rect 23848 18692 23900 18698
rect 23848 18634 23900 18640
rect 23846 18320 23902 18329
rect 23846 18255 23848 18264
rect 23900 18255 23902 18264
rect 23848 18226 23900 18232
rect 23860 18086 23888 18226
rect 23848 18080 23900 18086
rect 23848 18022 23900 18028
rect 23662 16960 23718 16969
rect 23662 16895 23718 16904
rect 23664 16788 23716 16794
rect 23664 16730 23716 16736
rect 23572 16108 23624 16114
rect 23572 16050 23624 16056
rect 23480 15904 23532 15910
rect 23480 15846 23532 15852
rect 23492 15745 23520 15846
rect 23478 15736 23534 15745
rect 23478 15671 23480 15680
rect 23532 15671 23534 15680
rect 23480 15642 23532 15648
rect 23492 15611 23520 15642
rect 23676 15609 23704 16730
rect 23662 15600 23718 15609
rect 23480 15564 23532 15570
rect 23662 15535 23718 15544
rect 23480 15506 23532 15512
rect 23216 15456 23336 15484
rect 23112 12776 23164 12782
rect 23112 12718 23164 12724
rect 23112 12368 23164 12374
rect 23112 12310 23164 12316
rect 23124 11898 23152 12310
rect 23112 11892 23164 11898
rect 23112 11834 23164 11840
rect 23216 11121 23244 15456
rect 23386 15192 23442 15201
rect 23492 15162 23520 15506
rect 23386 15127 23442 15136
rect 23480 15156 23532 15162
rect 23400 14550 23428 15127
rect 23480 15098 23532 15104
rect 23388 14544 23440 14550
rect 23308 14504 23388 14532
rect 23308 13530 23336 14504
rect 23388 14486 23440 14492
rect 23388 14408 23440 14414
rect 23388 14350 23440 14356
rect 23400 13870 23428 14350
rect 23388 13864 23440 13870
rect 23388 13806 23440 13812
rect 23676 13682 23704 15535
rect 23756 15088 23808 15094
rect 23756 15030 23808 15036
rect 23492 13654 23704 13682
rect 23296 13524 23348 13530
rect 23296 13466 23348 13472
rect 23492 12730 23520 13654
rect 23572 13524 23624 13530
rect 23572 13466 23624 13472
rect 23308 12702 23520 12730
rect 23202 11112 23258 11121
rect 23202 11047 23258 11056
rect 23308 10266 23336 12702
rect 23388 12640 23440 12646
rect 23388 12582 23440 12588
rect 23584 12594 23612 13466
rect 23664 13252 23716 13258
rect 23664 13194 23716 13200
rect 23676 12782 23704 13194
rect 23664 12776 23716 12782
rect 23664 12718 23716 12724
rect 23768 12646 23796 15030
rect 23756 12640 23808 12646
rect 23400 11218 23428 12582
rect 23584 12566 23704 12594
rect 23756 12582 23808 12588
rect 23388 11212 23440 11218
rect 23388 11154 23440 11160
rect 23478 11112 23534 11121
rect 23478 11047 23534 11056
rect 23296 10260 23348 10266
rect 23296 10202 23348 10208
rect 23020 10192 23072 10198
rect 23020 10134 23072 10140
rect 22650 10024 22706 10033
rect 22650 9959 22706 9968
rect 22928 9920 22980 9926
rect 22928 9862 22980 9868
rect 22940 9450 22968 9862
rect 23032 9654 23060 10134
rect 23308 9722 23336 10202
rect 23492 9994 23520 11047
rect 23572 10260 23624 10266
rect 23572 10202 23624 10208
rect 23480 9988 23532 9994
rect 23480 9930 23532 9936
rect 23584 9722 23612 10202
rect 23676 10130 23704 12566
rect 23768 12442 23796 12582
rect 23756 12436 23808 12442
rect 23756 12378 23808 12384
rect 23860 12322 23888 18022
rect 23952 17377 23980 19071
rect 24044 18154 24072 19110
rect 24032 18148 24084 18154
rect 24032 18090 24084 18096
rect 24032 17604 24084 17610
rect 24032 17546 24084 17552
rect 24044 17513 24072 17546
rect 24030 17504 24086 17513
rect 24086 17462 24164 17490
rect 24030 17439 24086 17448
rect 23938 17368 23994 17377
rect 23938 17303 23994 17312
rect 23940 17264 23992 17270
rect 23940 17206 23992 17212
rect 23952 12442 23980 17206
rect 24136 17066 24164 17462
rect 24032 17060 24084 17066
rect 24032 17002 24084 17008
rect 24124 17060 24176 17066
rect 24124 17002 24176 17008
rect 24044 16658 24072 17002
rect 24122 16960 24178 16969
rect 24122 16895 24178 16904
rect 24032 16652 24084 16658
rect 24032 16594 24084 16600
rect 24044 16250 24072 16594
rect 24032 16244 24084 16250
rect 24032 16186 24084 16192
rect 24030 15056 24086 15065
rect 24030 14991 24086 15000
rect 24044 14958 24072 14991
rect 24032 14952 24084 14958
rect 24032 14894 24084 14900
rect 24044 14618 24072 14894
rect 24032 14612 24084 14618
rect 24032 14554 24084 14560
rect 24136 14498 24164 16895
rect 24228 16046 24256 19366
rect 24780 19258 24808 20998
rect 24860 20868 24912 20874
rect 24860 20810 24912 20816
rect 24872 19990 24900 20810
rect 25148 20806 25176 21134
rect 25240 21010 25268 21927
rect 25228 21004 25280 21010
rect 25228 20946 25280 20952
rect 25136 20800 25188 20806
rect 25136 20742 25188 20748
rect 24860 19984 24912 19990
rect 24860 19926 24912 19932
rect 24872 19514 24900 19926
rect 24860 19508 24912 19514
rect 24860 19450 24912 19456
rect 24676 19236 24728 19242
rect 24780 19230 24900 19258
rect 24676 19178 24728 19184
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24584 18080 24636 18086
rect 24584 18022 24636 18028
rect 24596 17814 24624 18022
rect 24584 17808 24636 17814
rect 24584 17750 24636 17756
rect 24688 17610 24716 19178
rect 24768 19168 24820 19174
rect 24768 19110 24820 19116
rect 24780 18698 24808 19110
rect 24872 19009 24900 19230
rect 24858 19000 24914 19009
rect 24858 18935 24914 18944
rect 25042 19000 25098 19009
rect 25042 18935 25098 18944
rect 25056 18902 25084 18935
rect 25044 18896 25096 18902
rect 25044 18838 25096 18844
rect 24768 18692 24820 18698
rect 24768 18634 24820 18640
rect 25056 18426 25084 18838
rect 25148 18766 25176 20742
rect 25240 20602 25268 20946
rect 25228 20596 25280 20602
rect 25228 20538 25280 20544
rect 25332 20505 25360 22714
rect 25424 22098 25452 23802
rect 25594 23352 25650 23361
rect 25594 23287 25650 23296
rect 25608 22642 25636 23287
rect 25700 23254 25728 24550
rect 25688 23248 25740 23254
rect 25688 23190 25740 23196
rect 25596 22636 25648 22642
rect 25596 22578 25648 22584
rect 25412 22092 25464 22098
rect 25412 22034 25464 22040
rect 25410 21040 25466 21049
rect 25410 20975 25466 20984
rect 25318 20496 25374 20505
rect 25318 20431 25374 20440
rect 25424 20058 25452 20975
rect 25504 20256 25556 20262
rect 25504 20198 25556 20204
rect 25412 20052 25464 20058
rect 25412 19994 25464 20000
rect 25424 19378 25452 19994
rect 25516 19854 25544 20198
rect 25504 19848 25556 19854
rect 25504 19790 25556 19796
rect 25516 19446 25544 19790
rect 25504 19440 25556 19446
rect 25504 19382 25556 19388
rect 25412 19372 25464 19378
rect 25412 19314 25464 19320
rect 25226 18864 25282 18873
rect 25792 18834 25820 24919
rect 26528 24834 26556 27520
rect 26252 24806 26556 24834
rect 25872 19712 25924 19718
rect 25872 19654 25924 19660
rect 25226 18799 25228 18808
rect 25280 18799 25282 18808
rect 25780 18828 25832 18834
rect 25228 18770 25280 18776
rect 25780 18770 25832 18776
rect 25136 18760 25188 18766
rect 25136 18702 25188 18708
rect 25504 18760 25556 18766
rect 25504 18702 25556 18708
rect 25044 18420 25096 18426
rect 25044 18362 25096 18368
rect 25516 18086 25544 18702
rect 25792 18426 25820 18770
rect 25780 18420 25832 18426
rect 25780 18362 25832 18368
rect 25504 18080 25556 18086
rect 25504 18022 25556 18028
rect 24952 17808 25004 17814
rect 24952 17750 25004 17756
rect 25044 17808 25096 17814
rect 25044 17750 25096 17756
rect 25226 17776 25282 17785
rect 24676 17604 24728 17610
rect 24676 17546 24728 17552
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24398 16144 24454 16153
rect 24398 16079 24454 16088
rect 24860 16108 24912 16114
rect 24216 16040 24268 16046
rect 24216 15982 24268 15988
rect 24412 15638 24440 16079
rect 24860 16050 24912 16056
rect 24676 16040 24728 16046
rect 24676 15982 24728 15988
rect 24400 15632 24452 15638
rect 24688 15586 24716 15982
rect 24452 15580 24716 15586
rect 24400 15574 24716 15580
rect 24412 15558 24716 15574
rect 24872 15570 24900 16050
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24688 15162 24716 15558
rect 24860 15564 24912 15570
rect 24860 15506 24912 15512
rect 24768 15360 24820 15366
rect 24768 15302 24820 15308
rect 24676 15156 24728 15162
rect 24676 15098 24728 15104
rect 24044 14470 24164 14498
rect 23940 12436 23992 12442
rect 23940 12378 23992 12384
rect 23860 12294 23980 12322
rect 23848 12232 23900 12238
rect 23848 12174 23900 12180
rect 23860 11830 23888 12174
rect 23848 11824 23900 11830
rect 23848 11766 23900 11772
rect 23756 11348 23808 11354
rect 23756 11290 23808 11296
rect 23768 10606 23796 11290
rect 23756 10600 23808 10606
rect 23756 10542 23808 10548
rect 23846 10296 23902 10305
rect 23846 10231 23848 10240
rect 23900 10231 23902 10240
rect 23848 10202 23900 10208
rect 23664 10124 23716 10130
rect 23664 10066 23716 10072
rect 23848 9988 23900 9994
rect 23848 9930 23900 9936
rect 23662 9752 23718 9761
rect 23296 9716 23348 9722
rect 23296 9658 23348 9664
rect 23572 9716 23624 9722
rect 23662 9687 23718 9696
rect 23572 9658 23624 9664
rect 23020 9648 23072 9654
rect 23020 9590 23072 9596
rect 22928 9444 22980 9450
rect 22928 9386 22980 9392
rect 22940 8906 22968 9386
rect 23112 9376 23164 9382
rect 23112 9318 23164 9324
rect 23124 9178 23152 9318
rect 23570 9208 23626 9217
rect 23112 9172 23164 9178
rect 23570 9143 23626 9152
rect 23112 9114 23164 9120
rect 23584 9110 23612 9143
rect 23572 9104 23624 9110
rect 23572 9046 23624 9052
rect 23020 9036 23072 9042
rect 23020 8978 23072 8984
rect 22928 8900 22980 8906
rect 22928 8842 22980 8848
rect 23032 8566 23060 8978
rect 23020 8560 23072 8566
rect 23020 8502 23072 8508
rect 23584 8378 23612 9046
rect 23676 8430 23704 9687
rect 23756 9648 23808 9654
rect 23756 9590 23808 9596
rect 23400 8350 23612 8378
rect 23664 8424 23716 8430
rect 23664 8366 23716 8372
rect 23400 8090 23428 8350
rect 23388 8084 23440 8090
rect 23388 8026 23440 8032
rect 23664 7744 23716 7750
rect 23664 7686 23716 7692
rect 22558 5264 22614 5273
rect 22558 5199 22614 5208
rect 21270 4856 21326 4865
rect 21270 4791 21272 4800
rect 21324 4791 21326 4800
rect 21272 4762 21324 4768
rect 21088 4684 21140 4690
rect 21088 4626 21140 4632
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 21100 4282 21128 4626
rect 21088 4276 21140 4282
rect 21088 4218 21140 4224
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 23020 2304 23072 2310
rect 23020 2246 23072 2252
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 23032 649 23060 2246
rect 23676 1193 23704 7686
rect 23768 3602 23796 9590
rect 23860 9489 23888 9930
rect 23846 9480 23902 9489
rect 23846 9415 23902 9424
rect 23848 8968 23900 8974
rect 23848 8910 23900 8916
rect 23860 8634 23888 8910
rect 23848 8628 23900 8634
rect 23848 8570 23900 8576
rect 23952 8514 23980 12294
rect 24044 9994 24072 14470
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24214 13832 24270 13841
rect 24214 13767 24270 13776
rect 24124 13456 24176 13462
rect 24124 13398 24176 13404
rect 24136 12986 24164 13398
rect 24124 12980 24176 12986
rect 24124 12922 24176 12928
rect 24136 11150 24164 12922
rect 24228 12889 24256 13767
rect 24674 13288 24730 13297
rect 24674 13223 24730 13232
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24214 12880 24270 12889
rect 24214 12815 24270 12824
rect 24688 12782 24716 13223
rect 24216 12776 24268 12782
rect 24676 12776 24728 12782
rect 24216 12718 24268 12724
rect 24504 12736 24676 12764
rect 24228 11694 24256 12718
rect 24504 12084 24532 12736
rect 24676 12718 24728 12724
rect 24780 12481 24808 15302
rect 24964 14958 24992 17750
rect 25056 16998 25084 17750
rect 25226 17711 25282 17720
rect 25136 17672 25188 17678
rect 25136 17614 25188 17620
rect 25148 17066 25176 17614
rect 25240 17202 25268 17711
rect 25516 17678 25544 18022
rect 25504 17672 25556 17678
rect 25504 17614 25556 17620
rect 25228 17196 25280 17202
rect 25228 17138 25280 17144
rect 25136 17060 25188 17066
rect 25136 17002 25188 17008
rect 25044 16992 25096 16998
rect 25042 16960 25044 16969
rect 25096 16960 25098 16969
rect 25042 16895 25098 16904
rect 25148 15638 25176 17002
rect 25516 16998 25544 17614
rect 25504 16992 25556 16998
rect 25504 16934 25556 16940
rect 25136 15632 25188 15638
rect 25136 15574 25188 15580
rect 24952 14952 25004 14958
rect 24952 14894 25004 14900
rect 25044 14884 25096 14890
rect 25044 14826 25096 14832
rect 24952 14272 25004 14278
rect 24952 14214 25004 14220
rect 24964 13870 24992 14214
rect 25056 14074 25084 14826
rect 25044 14068 25096 14074
rect 25044 14010 25096 14016
rect 24952 13864 25004 13870
rect 24952 13806 25004 13812
rect 24860 13456 24912 13462
rect 24860 13398 24912 13404
rect 24766 12472 24822 12481
rect 24676 12436 24728 12442
rect 24766 12407 24822 12416
rect 24676 12378 24728 12384
rect 24688 12322 24716 12378
rect 24872 12374 24900 13398
rect 24860 12368 24912 12374
rect 24688 12294 24808 12322
rect 24860 12310 24912 12316
rect 24504 12056 24716 12084
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24216 11688 24268 11694
rect 24216 11630 24268 11636
rect 24228 11354 24256 11630
rect 24216 11348 24268 11354
rect 24216 11290 24268 11296
rect 24688 11286 24716 12056
rect 24676 11280 24728 11286
rect 24676 11222 24728 11228
rect 24216 11212 24268 11218
rect 24216 11154 24268 11160
rect 24124 11144 24176 11150
rect 24124 11086 24176 11092
rect 24124 10124 24176 10130
rect 24124 10066 24176 10072
rect 24032 9988 24084 9994
rect 24032 9930 24084 9936
rect 24030 9888 24086 9897
rect 24030 9823 24086 9832
rect 24044 8616 24072 9823
rect 24136 9178 24164 10066
rect 24124 9172 24176 9178
rect 24124 9114 24176 9120
rect 24044 8588 24164 8616
rect 23952 8486 24072 8514
rect 23940 8356 23992 8362
rect 23940 8298 23992 8304
rect 23952 7954 23980 8298
rect 24044 7954 24072 8486
rect 23940 7948 23992 7954
rect 23940 7890 23992 7896
rect 24032 7948 24084 7954
rect 24032 7890 24084 7896
rect 23848 7744 23900 7750
rect 23848 7686 23900 7692
rect 23860 7342 23888 7686
rect 23952 7546 23980 7890
rect 24044 7546 24072 7890
rect 24136 7750 24164 8588
rect 24124 7744 24176 7750
rect 24124 7686 24176 7692
rect 24228 7562 24256 11154
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24688 10266 24716 11222
rect 24676 10260 24728 10266
rect 24676 10202 24728 10208
rect 24674 10024 24730 10033
rect 24674 9959 24730 9968
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24688 9110 24716 9959
rect 24780 9450 24808 12294
rect 24858 12200 24914 12209
rect 24858 12135 24914 12144
rect 24872 11898 24900 12135
rect 24860 11892 24912 11898
rect 24860 11834 24912 11840
rect 24964 11286 24992 13806
rect 25056 13462 25084 14010
rect 25044 13456 25096 13462
rect 25044 13398 25096 13404
rect 25044 13320 25096 13326
rect 25044 13262 25096 13268
rect 25056 12986 25084 13262
rect 25044 12980 25096 12986
rect 25044 12922 25096 12928
rect 25042 11656 25098 11665
rect 25042 11591 25098 11600
rect 24860 11280 24912 11286
rect 24860 11222 24912 11228
rect 24952 11280 25004 11286
rect 24952 11222 25004 11228
rect 24872 9926 24900 11222
rect 24964 10742 24992 11222
rect 24952 10736 25004 10742
rect 24952 10678 25004 10684
rect 24950 10160 25006 10169
rect 24950 10095 24952 10104
rect 25004 10095 25006 10104
rect 24952 10066 25004 10072
rect 24860 9920 24912 9926
rect 24860 9862 24912 9868
rect 24964 9722 24992 10066
rect 24952 9716 25004 9722
rect 24952 9658 25004 9664
rect 24950 9616 25006 9625
rect 24950 9551 25006 9560
rect 24768 9444 24820 9450
rect 24768 9386 24820 9392
rect 24766 9344 24822 9353
rect 24766 9279 24822 9288
rect 24676 9104 24728 9110
rect 24676 9046 24728 9052
rect 24780 9042 24808 9279
rect 24964 9178 24992 9551
rect 25056 9518 25084 11591
rect 25148 11354 25176 15574
rect 25412 12640 25464 12646
rect 25412 12582 25464 12588
rect 25228 12096 25280 12102
rect 25228 12038 25280 12044
rect 25240 11694 25268 12038
rect 25228 11688 25280 11694
rect 25228 11630 25280 11636
rect 25136 11348 25188 11354
rect 25136 11290 25188 11296
rect 25134 10704 25190 10713
rect 25134 10639 25190 10648
rect 25148 10266 25176 10639
rect 25136 10260 25188 10266
rect 25136 10202 25188 10208
rect 25228 9920 25280 9926
rect 25228 9862 25280 9868
rect 25044 9512 25096 9518
rect 25044 9454 25096 9460
rect 25134 9208 25190 9217
rect 24952 9172 25004 9178
rect 25134 9143 25190 9152
rect 24952 9114 25004 9120
rect 24768 9036 24820 9042
rect 24768 8978 24820 8984
rect 24780 8922 24808 8978
rect 24780 8894 24900 8922
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24766 8664 24822 8673
rect 24872 8634 24900 8894
rect 25148 8634 25176 9143
rect 24766 8599 24822 8608
rect 24860 8628 24912 8634
rect 24674 8120 24730 8129
rect 24780 8090 24808 8599
rect 24860 8570 24912 8576
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 24952 8424 25004 8430
rect 24950 8392 24952 8401
rect 25004 8392 25006 8401
rect 24950 8327 25006 8336
rect 24674 8055 24730 8064
rect 24768 8084 24820 8090
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 23940 7540 23992 7546
rect 23940 7482 23992 7488
rect 24032 7540 24084 7546
rect 24032 7482 24084 7488
rect 24136 7534 24256 7562
rect 24688 7546 24716 8055
rect 24768 8026 24820 8032
rect 24766 7576 24822 7585
rect 24676 7540 24728 7546
rect 23848 7336 23900 7342
rect 23848 7278 23900 7284
rect 23756 3596 23808 3602
rect 23756 3538 23808 3544
rect 23768 3194 23796 3538
rect 23756 3188 23808 3194
rect 23756 3130 23808 3136
rect 23846 3088 23902 3097
rect 23846 3023 23902 3032
rect 23860 2990 23888 3023
rect 23848 2984 23900 2990
rect 23848 2926 23900 2932
rect 24136 2514 24164 7534
rect 24766 7511 24822 7520
rect 24676 7482 24728 7488
rect 24214 7440 24270 7449
rect 24214 7375 24270 7384
rect 24228 6254 24256 7375
rect 24780 7002 24808 7511
rect 24768 6996 24820 7002
rect 24768 6938 24820 6944
rect 24582 6896 24638 6905
rect 24582 6831 24584 6840
rect 24636 6831 24638 6840
rect 24584 6802 24636 6808
rect 24596 6746 24624 6802
rect 24596 6718 24716 6746
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24688 6390 24716 6718
rect 24766 6488 24822 6497
rect 24766 6423 24768 6432
rect 24820 6423 24822 6432
rect 24768 6394 24820 6400
rect 24676 6384 24728 6390
rect 24676 6326 24728 6332
rect 24216 6248 24268 6254
rect 24216 6190 24268 6196
rect 24858 6080 24914 6089
rect 24858 6015 24914 6024
rect 24766 5944 24822 5953
rect 24766 5879 24768 5888
rect 24820 5879 24822 5888
rect 24768 5850 24820 5856
rect 24582 5808 24638 5817
rect 24582 5743 24584 5752
rect 24636 5743 24638 5752
rect 24584 5714 24636 5720
rect 24596 5658 24624 5714
rect 24596 5630 24716 5658
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24688 5302 24716 5630
rect 24766 5400 24822 5409
rect 24766 5335 24768 5344
rect 24820 5335 24822 5344
rect 24768 5306 24820 5312
rect 24676 5296 24728 5302
rect 24582 5264 24638 5273
rect 24676 5238 24728 5244
rect 24582 5199 24638 5208
rect 24596 5166 24624 5199
rect 24584 5160 24636 5166
rect 24584 5102 24636 5108
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24872 3602 24900 6015
rect 24860 3596 24912 3602
rect 24860 3538 24912 3544
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24872 3194 24900 3538
rect 25136 3528 25188 3534
rect 25136 3470 25188 3476
rect 25044 3392 25096 3398
rect 25042 3360 25044 3369
rect 25096 3360 25098 3369
rect 25042 3295 25098 3304
rect 24860 3188 24912 3194
rect 24860 3130 24912 3136
rect 25148 2990 25176 3470
rect 24860 2984 24912 2990
rect 24860 2926 24912 2932
rect 25136 2984 25188 2990
rect 25136 2926 25188 2932
rect 24872 2514 24900 2926
rect 24124 2508 24176 2514
rect 24124 2450 24176 2456
rect 24860 2508 24912 2514
rect 24860 2450 24912 2456
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 23662 1184 23718 1193
rect 23662 1119 23718 1128
rect 23018 640 23074 649
rect 23018 575 23074 584
rect 3514 368 3570 377
rect 3514 303 3570 312
rect 14002 0 14058 480
rect 25240 241 25268 9862
rect 25320 2848 25372 2854
rect 25318 2816 25320 2825
rect 25372 2816 25374 2825
rect 25318 2751 25374 2760
rect 25424 2281 25452 12582
rect 25516 10810 25544 16934
rect 25688 15904 25740 15910
rect 25688 15846 25740 15852
rect 25596 14816 25648 14822
rect 25596 14758 25648 14764
rect 25504 10804 25556 10810
rect 25504 10746 25556 10752
rect 25502 10160 25558 10169
rect 25502 10095 25558 10104
rect 25516 9654 25544 10095
rect 25504 9648 25556 9654
rect 25504 9590 25556 9596
rect 25608 3913 25636 14758
rect 25700 4457 25728 15846
rect 25686 4448 25742 4457
rect 25686 4383 25742 4392
rect 25594 3904 25650 3913
rect 25594 3839 25650 3848
rect 25884 3097 25912 19654
rect 26252 15881 26280 24806
rect 27080 22273 27108 27520
rect 27632 23866 27660 27520
rect 27620 23860 27672 23866
rect 27620 23802 27672 23808
rect 27066 22264 27122 22273
rect 27066 22199 27122 22208
rect 26238 15872 26294 15881
rect 26238 15807 26294 15816
rect 25870 3088 25926 3097
rect 25870 3023 25926 3032
rect 25504 2304 25556 2310
rect 25410 2272 25466 2281
rect 25504 2246 25556 2252
rect 25410 2207 25466 2216
rect 25516 1737 25544 2246
rect 25502 1728 25558 1737
rect 25502 1663 25558 1672
rect 25226 232 25282 241
rect 25226 167 25282 176
<< via2 >>
rect 1306 27648 1362 27704
rect 1214 24792 1270 24848
rect 570 22344 626 22400
rect 202 22072 258 22128
rect 23570 27648 23626 27704
rect 1582 26968 1638 27024
rect 1766 23704 1822 23760
rect 1950 22480 2006 22536
rect 1674 21392 1730 21448
rect 1766 21120 1822 21176
rect 1306 18808 1362 18864
rect 1490 18264 1546 18320
rect 1398 11464 1454 11520
rect 1398 11212 1454 11248
rect 1398 11192 1400 11212
rect 1400 11192 1452 11212
rect 1452 11192 1454 11212
rect 1398 10124 1454 10160
rect 1398 10104 1400 10124
rect 1400 10104 1452 10124
rect 1452 10104 1454 10124
rect 1766 18128 1822 18184
rect 2410 24520 2466 24576
rect 3790 26288 3846 26344
rect 3698 24792 3754 24848
rect 2410 21936 2466 21992
rect 2962 22516 2964 22536
rect 2964 22516 3016 22536
rect 3016 22516 3018 22536
rect 2962 22480 3018 22516
rect 3054 22208 3110 22264
rect 2962 22072 3018 22128
rect 2318 19216 2374 19272
rect 2778 18536 2834 18592
rect 2134 16652 2190 16688
rect 2134 16632 2136 16652
rect 2136 16632 2188 16652
rect 2188 16632 2190 16652
rect 3238 23568 3294 23624
rect 3514 23180 3570 23216
rect 3514 23160 3516 23180
rect 3516 23160 3568 23180
rect 3568 23160 3570 23180
rect 3698 22480 3754 22536
rect 3790 22208 3846 22264
rect 3974 25608 4030 25664
rect 4066 25064 4122 25120
rect 3974 22616 4030 22672
rect 3974 22072 4030 22128
rect 4342 21936 4398 21992
rect 3882 20168 3938 20224
rect 3790 19216 3846 19272
rect 3330 18400 3386 18456
rect 2226 15272 2282 15328
rect 1766 13912 1822 13968
rect 1582 9424 1638 9480
rect 1398 7792 1454 7848
rect 1582 8744 1638 8800
rect 1582 8084 1638 8120
rect 1582 8064 1584 8084
rect 1584 8064 1636 8084
rect 1636 8064 1638 8084
rect 1582 7420 1584 7440
rect 1584 7420 1636 7440
rect 1636 7420 1638 7440
rect 1582 7384 1638 7420
rect 1674 4800 1730 4856
rect 1490 4120 1546 4176
rect 1582 3460 1638 3496
rect 1582 3440 1584 3460
rect 1584 3440 1636 3460
rect 1636 3440 1638 3460
rect 3606 18028 3608 18048
rect 3608 18028 3660 18048
rect 3660 18028 3662 18048
rect 3606 17992 3662 18028
rect 3974 17856 4030 17912
rect 3974 15952 4030 16008
rect 4158 16088 4214 16144
rect 4066 15816 4122 15872
rect 3606 15408 3662 15464
rect 3514 15000 3570 15056
rect 2502 14320 2558 14376
rect 2502 12688 2558 12744
rect 2042 10240 2098 10296
rect 2042 8880 2098 8936
rect 2042 8064 2098 8120
rect 2226 7928 2282 7984
rect 2318 7384 2374 7440
rect 2962 13404 2964 13424
rect 2964 13404 3016 13424
rect 3016 13404 3018 13424
rect 2962 13368 3018 13404
rect 2870 11620 2926 11656
rect 2870 11600 2872 11620
rect 2872 11600 2924 11620
rect 2924 11600 2926 11620
rect 2686 10684 2688 10704
rect 2688 10684 2740 10704
rect 2740 10684 2742 10704
rect 2686 10648 2742 10684
rect 2686 9988 2742 10024
rect 2686 9968 2688 9988
rect 2688 9968 2740 9988
rect 2740 9968 2742 9988
rect 2870 9968 2926 10024
rect 2870 9444 2926 9480
rect 2870 9424 2872 9444
rect 2872 9424 2924 9444
rect 2924 9424 2926 9444
rect 3238 14728 3294 14784
rect 3330 12164 3386 12200
rect 3330 12144 3332 12164
rect 3332 12144 3384 12164
rect 3384 12144 3386 12164
rect 3698 14592 3754 14648
rect 3974 13640 4030 13696
rect 3790 13232 3846 13288
rect 3698 12824 3754 12880
rect 3974 12008 4030 12064
rect 3790 11328 3846 11384
rect 3514 11192 3570 11248
rect 4342 14728 4398 14784
rect 4986 24792 5042 24848
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 4802 24384 4858 24440
rect 4526 23432 4582 23488
rect 4526 22480 4582 22536
rect 4526 22072 4582 22128
rect 4618 21972 4620 21992
rect 4620 21972 4672 21992
rect 4672 21972 4674 21992
rect 4618 21936 4674 21972
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5998 23296 6054 23352
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5446 22516 5448 22536
rect 5448 22516 5500 22536
rect 5500 22516 5502 22536
rect 5446 22480 5502 22516
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 4986 20304 5042 20360
rect 4802 20032 4858 20088
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 4986 19236 5042 19272
rect 4986 19216 4988 19236
rect 4988 19216 5040 19236
rect 5040 19216 5042 19236
rect 4710 18944 4766 19000
rect 4986 18808 5042 18864
rect 5262 18844 5264 18864
rect 5264 18844 5316 18864
rect 5316 18844 5318 18864
rect 4802 18692 4858 18728
rect 4802 18672 4804 18692
rect 4804 18672 4856 18692
rect 4856 18672 4858 18692
rect 4802 18400 4858 18456
rect 4710 13252 4766 13288
rect 4710 13232 4712 13252
rect 4712 13232 4764 13252
rect 4764 13232 4766 13252
rect 4250 11736 4306 11792
rect 4434 11464 4490 11520
rect 3238 8472 3294 8528
rect 3146 6704 3202 6760
rect 2962 5480 3018 5536
rect 1858 3032 1914 3088
rect 1766 2896 1822 2952
rect 1582 2252 1584 2272
rect 1584 2252 1636 2272
rect 1636 2252 1638 2272
rect 1582 2216 1638 2252
rect 4526 10412 4528 10432
rect 4528 10412 4580 10432
rect 4580 10412 4582 10432
rect 4526 10376 4582 10412
rect 4250 6160 4306 6216
rect 5262 18808 5318 18844
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5538 18128 5594 18184
rect 5446 17720 5502 17776
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 6274 23160 6330 23216
rect 6090 16632 6146 16688
rect 5998 15816 6054 15872
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 7010 21392 7066 21448
rect 7102 18672 7158 18728
rect 6734 18264 6790 18320
rect 7286 23296 7342 23352
rect 7930 24284 7932 24304
rect 7932 24284 7984 24304
rect 7984 24284 7986 24304
rect 7930 24248 7986 24284
rect 8114 22652 8116 22672
rect 8116 22652 8168 22672
rect 8168 22652 8170 22672
rect 8114 22616 8170 22652
rect 7838 22208 7894 22264
rect 7010 15852 7012 15872
rect 7012 15852 7064 15872
rect 7064 15852 7066 15872
rect 7010 15816 7066 15852
rect 6550 14592 6606 14648
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5630 13776 5686 13832
rect 5630 13676 5632 13696
rect 5632 13676 5684 13696
rect 5684 13676 5686 13696
rect 5630 13640 5686 13676
rect 5814 13504 5870 13560
rect 5170 12688 5226 12744
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5538 12280 5594 12336
rect 5998 12180 6000 12200
rect 6000 12180 6052 12200
rect 6052 12180 6054 12200
rect 5998 12144 6054 12180
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5354 11500 5356 11520
rect 5356 11500 5408 11520
rect 5408 11500 5410 11520
rect 5354 11464 5410 11500
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 4710 9594 4766 9650
rect 6734 12008 6790 12064
rect 4894 9560 4950 9616
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 6458 9696 6514 9752
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 7378 16224 7434 16280
rect 7286 15000 7342 15056
rect 7562 20440 7618 20496
rect 7562 19896 7618 19952
rect 7470 15136 7526 15192
rect 7378 14728 7434 14784
rect 7654 17040 7710 17096
rect 7194 11872 7250 11928
rect 8390 24792 8446 24848
rect 8390 23976 8446 24032
rect 8482 23704 8538 23760
rect 8574 22888 8630 22944
rect 7838 20848 7894 20904
rect 7838 17756 7840 17776
rect 7840 17756 7892 17776
rect 7892 17756 7894 17776
rect 7838 17720 7894 17756
rect 7102 11464 7158 11520
rect 7010 10920 7066 10976
rect 8206 21800 8262 21856
rect 8666 21800 8722 21856
rect 9494 23196 9496 23216
rect 9496 23196 9548 23216
rect 9548 23196 9550 23216
rect 9494 23160 9550 23196
rect 9494 22092 9550 22128
rect 9494 22072 9496 22092
rect 9496 22072 9548 22092
rect 9548 22072 9550 22092
rect 8390 21020 8392 21040
rect 8392 21020 8444 21040
rect 8444 21020 8446 21040
rect 8390 20984 8446 21020
rect 8206 20848 8262 20904
rect 9494 21664 9550 21720
rect 9402 20440 9458 20496
rect 8758 20168 8814 20224
rect 8390 19488 8446 19544
rect 8482 18400 8538 18456
rect 9586 20204 9588 20224
rect 9588 20204 9640 20224
rect 9640 20204 9642 20224
rect 9586 20168 9642 20204
rect 9954 24520 10010 24576
rect 10046 24248 10102 24304
rect 9954 24112 10010 24168
rect 9954 23432 10010 23488
rect 10046 22208 10102 22264
rect 9954 21800 10010 21856
rect 9770 20052 9826 20088
rect 9770 20032 9772 20052
rect 9772 20032 9824 20052
rect 9824 20032 9826 20052
rect 9126 17720 9182 17776
rect 8298 16360 8354 16416
rect 8206 16224 8262 16280
rect 8114 15272 8170 15328
rect 8390 15544 8446 15600
rect 8298 14884 8354 14920
rect 8298 14864 8300 14884
rect 8300 14864 8352 14884
rect 8352 14864 8354 14884
rect 8390 14612 8446 14648
rect 8390 14592 8392 14612
rect 8392 14592 8444 14612
rect 8444 14592 8446 14612
rect 8206 14048 8262 14104
rect 8022 12860 8024 12880
rect 8024 12860 8076 12880
rect 8076 12860 8078 12880
rect 8022 12824 8078 12860
rect 6918 9968 6974 10024
rect 7654 10784 7710 10840
rect 7654 10376 7710 10432
rect 7562 9968 7618 10024
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 8390 13640 8446 13696
rect 8574 14320 8630 14376
rect 8574 13232 8630 13288
rect 8942 16496 8998 16552
rect 8758 15000 8814 15056
rect 9862 18944 9918 19000
rect 9126 16496 9182 16552
rect 9126 16224 9182 16280
rect 8942 14456 8998 14512
rect 9034 13504 9090 13560
rect 8390 12144 8446 12200
rect 7746 8880 7802 8936
rect 8206 9560 8262 9616
rect 7102 7792 7158 7848
rect 9402 16224 9458 16280
rect 9954 16224 10010 16280
rect 9862 15272 9918 15328
rect 9310 12688 9366 12744
rect 9770 12688 9826 12744
rect 9678 12044 9680 12064
rect 9680 12044 9732 12064
rect 9732 12044 9734 12064
rect 9678 12008 9734 12044
rect 9678 10920 9734 10976
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 11334 25200 11390 25256
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10414 21800 10470 21856
rect 10966 23296 11022 23352
rect 11058 23160 11114 23216
rect 11242 23024 11298 23080
rect 11242 22344 11298 22400
rect 11334 22072 11390 22128
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10322 20576 10378 20632
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10782 19216 10838 19272
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10690 18148 10746 18184
rect 10690 18128 10692 18148
rect 10692 18128 10744 18148
rect 10744 18128 10746 18148
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10138 15156 10194 15192
rect 10138 15136 10140 15156
rect 10140 15136 10192 15156
rect 10192 15136 10194 15156
rect 10782 15272 10838 15328
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10230 14048 10286 14104
rect 10782 13640 10838 13696
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 9218 9696 9274 9752
rect 8666 7828 8668 7848
rect 8668 7828 8720 7848
rect 8720 7828 8722 7848
rect 8666 7792 8722 7828
rect 10782 13096 10838 13152
rect 11242 21392 11298 21448
rect 11242 20848 11298 20904
rect 11058 20304 11114 20360
rect 11150 20032 11206 20088
rect 11058 19760 11114 19816
rect 11150 19624 11206 19680
rect 10966 19352 11022 19408
rect 11058 19216 11114 19272
rect 11058 18264 11114 18320
rect 11518 23468 11520 23488
rect 11520 23468 11572 23488
rect 11572 23468 11574 23488
rect 11518 23432 11574 23468
rect 11610 22752 11666 22808
rect 11702 18844 11704 18864
rect 11704 18844 11756 18864
rect 11756 18844 11758 18864
rect 11702 18808 11758 18844
rect 11518 17856 11574 17912
rect 11702 17720 11758 17776
rect 11518 15544 11574 15600
rect 10966 14728 11022 14784
rect 11150 15000 11206 15056
rect 11334 15000 11390 15056
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10690 11600 10746 11656
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10874 12416 10930 12472
rect 10966 12144 11022 12200
rect 9954 10512 10010 10568
rect 10230 11056 10286 11112
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 9862 9016 9918 9072
rect 9770 7928 9826 7984
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 10598 9832 10654 9888
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 12346 23976 12402 24032
rect 12162 23604 12164 23624
rect 12164 23604 12216 23624
rect 12216 23604 12218 23624
rect 12162 23568 12218 23604
rect 12346 23568 12402 23624
rect 12254 22636 12310 22672
rect 12254 22616 12256 22636
rect 12256 22616 12308 22636
rect 12308 22616 12310 22636
rect 12346 22480 12402 22536
rect 12070 21800 12126 21856
rect 12714 24792 12770 24848
rect 12622 24112 12678 24168
rect 12990 24112 13046 24168
rect 12622 22480 12678 22536
rect 12438 21392 12494 21448
rect 11794 13504 11850 13560
rect 12990 22888 13046 22944
rect 12714 19760 12770 19816
rect 12714 19488 12770 19544
rect 12162 17720 12218 17776
rect 11978 16768 12034 16824
rect 12806 17584 12862 17640
rect 12254 15272 12310 15328
rect 11610 12280 11666 12336
rect 12070 12280 12126 12336
rect 11794 11892 11850 11928
rect 11794 11872 11796 11892
rect 11796 11872 11848 11892
rect 11848 11872 11850 11892
rect 11518 11192 11574 11248
rect 11242 10240 11298 10296
rect 11242 9968 11298 10024
rect 11610 9560 11666 9616
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 11886 10784 11942 10840
rect 12162 10376 12218 10432
rect 12162 9696 12218 9752
rect 12714 15816 12770 15872
rect 13082 17040 13138 17096
rect 13082 16768 13138 16824
rect 13266 21392 13322 21448
rect 13726 23160 13782 23216
rect 14002 22888 14058 22944
rect 13634 21528 13690 21584
rect 13266 20848 13322 20904
rect 13358 19216 13414 19272
rect 13818 21800 13874 21856
rect 13542 19116 13544 19136
rect 13544 19116 13596 19136
rect 13596 19116 13598 19136
rect 13542 19080 13598 19116
rect 14002 20576 14058 20632
rect 14278 23468 14280 23488
rect 14280 23468 14332 23488
rect 14332 23468 14334 23488
rect 14278 23432 14334 23468
rect 13910 20304 13966 20360
rect 13450 18264 13506 18320
rect 13266 17992 13322 18048
rect 13542 18128 13598 18184
rect 13450 17856 13506 17912
rect 13266 17040 13322 17096
rect 13174 15988 13176 16008
rect 13176 15988 13228 16008
rect 13228 15988 13230 16008
rect 13174 15952 13230 15988
rect 12898 14864 12954 14920
rect 12714 13368 12770 13424
rect 13358 15000 13414 15056
rect 14278 20440 14334 20496
rect 13634 15680 13690 15736
rect 13818 16088 13874 16144
rect 14094 16360 14150 16416
rect 13542 14864 13598 14920
rect 13450 14592 13506 14648
rect 13450 14476 13506 14512
rect 13450 14456 13452 14476
rect 13452 14456 13504 14476
rect 13504 14456 13506 14476
rect 12622 12416 12678 12472
rect 13266 12416 13322 12472
rect 12254 9016 12310 9072
rect 12254 8880 12310 8936
rect 11794 7792 11850 7848
rect 11978 7384 12034 7440
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 13266 11500 13268 11520
rect 13268 11500 13320 11520
rect 13320 11500 13322 11520
rect 13266 11464 13322 11500
rect 13174 11328 13230 11384
rect 13082 10376 13138 10432
rect 13910 15020 13966 15056
rect 13910 15000 13912 15020
rect 13912 15000 13964 15020
rect 13964 15000 13966 15020
rect 14278 13776 14334 13832
rect 14002 12824 14058 12880
rect 13818 9596 13820 9616
rect 13820 9596 13872 9616
rect 13872 9596 13874 9616
rect 13818 9560 13874 9596
rect 13634 8472 13690 8528
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 15382 24792 15438 24848
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 15290 23160 15346 23216
rect 14462 21256 14518 21312
rect 14462 20712 14518 20768
rect 14646 20204 14648 20224
rect 14648 20204 14700 20224
rect 14700 20204 14702 20224
rect 14646 20168 14702 20204
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 15474 22752 15530 22808
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 15382 21528 15438 21584
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 15290 20168 15346 20224
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14922 19216 14978 19272
rect 15474 20168 15530 20224
rect 15474 20032 15530 20088
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14554 16224 14610 16280
rect 15382 17992 15438 18048
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 16486 24656 16542 24712
rect 15750 23296 15806 23352
rect 15750 22344 15806 22400
rect 15842 21120 15898 21176
rect 15842 20712 15898 20768
rect 15750 20204 15752 20224
rect 15752 20204 15804 20224
rect 15804 20204 15806 20224
rect 15750 20168 15806 20204
rect 15750 19624 15806 19680
rect 15750 15700 15806 15736
rect 15750 15680 15752 15700
rect 15752 15680 15804 15700
rect 15804 15680 15806 15700
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14554 14864 14610 14920
rect 15106 14320 15162 14376
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 15474 13504 15530 13560
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 15566 13404 15568 13424
rect 15568 13404 15620 13424
rect 15620 13404 15622 13424
rect 15566 13368 15622 13404
rect 15474 12960 15530 13016
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14370 11056 14426 11112
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14186 10240 14242 10296
rect 14646 10260 14702 10296
rect 14646 10240 14648 10260
rect 14648 10240 14700 10260
rect 14700 10240 14702 10260
rect 14186 9968 14242 10024
rect 14094 9424 14150 9480
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 15382 9696 15438 9752
rect 15750 11600 15806 11656
rect 15750 10920 15806 10976
rect 17222 25236 17224 25256
rect 17224 25236 17276 25256
rect 17276 25236 17278 25256
rect 17222 25200 17278 25236
rect 17866 24792 17922 24848
rect 18050 24692 18052 24712
rect 18052 24692 18104 24712
rect 18104 24692 18106 24712
rect 18050 24656 18106 24692
rect 18418 24656 18474 24712
rect 17498 24148 17500 24168
rect 17500 24148 17552 24168
rect 17552 24148 17554 24168
rect 17498 24112 17554 24148
rect 16762 22480 16818 22536
rect 16394 21256 16450 21312
rect 16026 21120 16082 21176
rect 16394 20168 16450 20224
rect 16210 17992 16266 18048
rect 16026 17312 16082 17368
rect 17406 22888 17462 22944
rect 17682 23704 17738 23760
rect 17498 20712 17554 20768
rect 18234 23296 18290 23352
rect 16302 16632 16358 16688
rect 17222 19896 17278 19952
rect 16946 18536 17002 18592
rect 17038 18264 17094 18320
rect 16854 16496 16910 16552
rect 17038 16496 17094 16552
rect 16762 14320 16818 14376
rect 16946 15408 17002 15464
rect 17038 14320 17094 14376
rect 16026 13912 16082 13968
rect 16118 12280 16174 12336
rect 15934 10784 15990 10840
rect 15842 10512 15898 10568
rect 15750 10104 15806 10160
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14554 8356 14610 8392
rect 14554 8336 14556 8356
rect 14556 8336 14608 8356
rect 14608 8336 14610 8356
rect 17038 13640 17094 13696
rect 18142 21256 18198 21312
rect 18142 20576 18198 20632
rect 18234 20440 18290 20496
rect 17774 14592 17830 14648
rect 18142 16244 18198 16280
rect 18142 16224 18144 16244
rect 18144 16224 18196 16244
rect 18196 16224 18198 16244
rect 18326 19760 18382 19816
rect 19338 24112 19394 24168
rect 19338 23160 19394 23216
rect 19246 22072 19302 22128
rect 19154 21800 19210 21856
rect 18602 20168 18658 20224
rect 19062 19660 19064 19680
rect 19064 19660 19116 19680
rect 19116 19660 19118 19680
rect 19062 19624 19118 19660
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19798 23704 19854 23760
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19798 23196 19800 23216
rect 19800 23196 19852 23216
rect 19852 23196 19854 23216
rect 19798 23160 19854 23196
rect 19890 22616 19946 22672
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 20810 24792 20866 24848
rect 21178 24792 21234 24848
rect 20534 24520 20590 24576
rect 19338 21120 19394 21176
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 18602 19080 18658 19136
rect 18602 18028 18604 18048
rect 18604 18028 18656 18048
rect 18656 18028 18658 18048
rect 18602 17992 18658 18028
rect 18418 17176 18474 17232
rect 18326 16360 18382 16416
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 20074 21256 20130 21312
rect 20534 23296 20590 23352
rect 20442 21412 20498 21448
rect 20442 21392 20444 21412
rect 20444 21392 20496 21412
rect 20496 21392 20498 21412
rect 20258 20984 20314 21040
rect 21638 24384 21694 24440
rect 21454 23860 21510 23896
rect 21454 23840 21456 23860
rect 21456 23840 21508 23860
rect 21508 23840 21510 23860
rect 20810 23024 20866 23080
rect 21270 22752 21326 22808
rect 21454 22752 21510 22808
rect 20810 22208 20866 22264
rect 21178 22072 21234 22128
rect 21086 21836 21088 21856
rect 21088 21836 21140 21856
rect 21140 21836 21142 21856
rect 21086 21800 21142 21836
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19522 18672 19578 18728
rect 19246 17448 19302 17504
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19614 17756 19616 17776
rect 19616 17756 19668 17776
rect 19668 17756 19670 17776
rect 19614 17720 19670 17756
rect 18234 14728 18290 14784
rect 18602 15852 18604 15872
rect 18604 15852 18656 15872
rect 18656 15852 18658 15872
rect 18602 15816 18658 15852
rect 17590 13504 17646 13560
rect 17774 13096 17830 13152
rect 17774 12416 17830 12472
rect 18970 16224 19026 16280
rect 18694 13932 18750 13968
rect 18694 13912 18696 13932
rect 18696 13912 18748 13932
rect 18748 13912 18750 13932
rect 18602 11500 18604 11520
rect 18604 11500 18656 11520
rect 18656 11500 18658 11520
rect 18602 11464 18658 11500
rect 18786 11348 18842 11384
rect 18786 11328 18788 11348
rect 18788 11328 18840 11348
rect 18840 11328 18842 11348
rect 19982 17620 19984 17640
rect 19984 17620 20036 17640
rect 20036 17620 20038 17640
rect 19982 17584 20038 17620
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19430 16496 19486 16552
rect 21178 18828 21234 18864
rect 21178 18808 21180 18828
rect 21180 18808 21232 18828
rect 21232 18808 21234 18828
rect 20166 18264 20222 18320
rect 20074 15952 20130 16008
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19430 13504 19486 13560
rect 19338 12980 19394 13016
rect 19338 12960 19340 12980
rect 19340 12960 19392 12980
rect 19392 12960 19394 12980
rect 19522 12960 19578 13016
rect 19430 11600 19486 11656
rect 18786 10260 18842 10296
rect 18786 10240 18788 10260
rect 18788 10240 18840 10260
rect 18840 10240 18842 10260
rect 18970 10104 19026 10160
rect 18234 8336 18290 8392
rect 18510 8356 18566 8392
rect 18510 8336 18512 8356
rect 18512 8336 18564 8356
rect 18564 8336 18566 8356
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 8114 3032 8170 3088
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 8850 1536 8906 1592
rect 7562 1400 7618 1456
rect 18234 7248 18290 7304
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 19154 9696 19210 9752
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19614 10804 19670 10840
rect 19614 10784 19616 10804
rect 19616 10784 19668 10804
rect 19668 10784 19670 10804
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19890 9560 19946 9616
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 20258 13368 20314 13424
rect 20258 13096 20314 13152
rect 20258 9832 20314 9888
rect 20994 17060 21050 17096
rect 20994 17040 20996 17060
rect 20996 17040 21048 17060
rect 21048 17040 21050 17060
rect 21638 22888 21694 22944
rect 21914 24656 21970 24712
rect 21914 23840 21970 23896
rect 21822 23604 21824 23624
rect 21824 23604 21876 23624
rect 21876 23604 21878 23624
rect 21822 23568 21878 23604
rect 24306 26560 24362 26616
rect 23938 25472 23994 25528
rect 23294 24656 23350 24712
rect 23110 23976 23166 24032
rect 22834 23024 22890 23080
rect 22742 22072 22798 22128
rect 23294 22616 23350 22672
rect 23202 22480 23258 22536
rect 23110 22344 23166 22400
rect 21546 19216 21602 19272
rect 21086 15544 21142 15600
rect 20350 9288 20406 9344
rect 20166 9152 20222 9208
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 20810 12280 20866 12336
rect 20994 12280 21050 12336
rect 22466 18808 22522 18864
rect 21178 12144 21234 12200
rect 21822 15000 21878 15056
rect 22282 13912 22338 13968
rect 22190 12980 22246 13016
rect 22190 12960 22192 12980
rect 22192 12960 22244 12980
rect 22244 12960 22246 12980
rect 21638 11600 21694 11656
rect 20994 10920 21050 10976
rect 21914 9696 21970 9752
rect 21546 9424 21602 9480
rect 21362 9036 21418 9072
rect 21362 9016 21364 9036
rect 21364 9016 21416 9036
rect 21416 9016 21418 9036
rect 19154 7384 19210 7440
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19062 5752 19118 5808
rect 22650 18400 22706 18456
rect 22466 16360 22522 16416
rect 23018 21412 23074 21448
rect 23018 21392 23020 21412
rect 23020 21392 23072 21412
rect 23072 21392 23074 21412
rect 23110 18944 23166 19000
rect 23478 21528 23534 21584
rect 23846 24792 23902 24848
rect 23754 22752 23810 22808
rect 23294 20984 23350 21040
rect 23478 17756 23480 17776
rect 23480 17756 23532 17776
rect 23532 17756 23534 17776
rect 23478 17720 23534 17756
rect 23202 16496 23258 16552
rect 23110 15816 23166 15872
rect 23018 13504 23074 13560
rect 22374 9580 22430 9616
rect 22374 9560 22376 9580
rect 22376 9560 22428 9580
rect 22428 9560 22430 9580
rect 22190 6840 22246 6896
rect 21362 6024 21418 6080
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 24766 27104 24822 27160
rect 24766 26016 24822 26072
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24214 24520 24270 24576
rect 24122 24112 24178 24168
rect 24030 23160 24086 23216
rect 23846 21120 23902 21176
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24950 24656 25006 24712
rect 24858 24404 24914 24440
rect 24858 24384 24860 24404
rect 24860 24384 24912 24404
rect 24912 24384 24914 24404
rect 24766 24248 24822 24304
rect 24766 23840 24822 23896
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24214 21528 24270 21584
rect 24214 21120 24270 21176
rect 25778 24928 25834 24984
rect 25226 23432 25282 23488
rect 25134 23024 25190 23080
rect 25042 21412 25098 21448
rect 25042 21392 25044 21412
rect 25044 21392 25096 21412
rect 25096 21392 25098 21412
rect 25226 21936 25282 21992
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24122 19216 24178 19272
rect 23938 19080 23994 19136
rect 23846 18284 23902 18320
rect 23846 18264 23848 18284
rect 23848 18264 23900 18284
rect 23900 18264 23902 18284
rect 23662 16904 23718 16960
rect 23478 15700 23534 15736
rect 23478 15680 23480 15700
rect 23480 15680 23532 15700
rect 23532 15680 23534 15700
rect 23662 15544 23718 15600
rect 23386 15136 23442 15192
rect 23202 11056 23258 11112
rect 23478 11056 23534 11112
rect 22650 9968 22706 10024
rect 24030 17448 24086 17504
rect 23938 17312 23994 17368
rect 24122 16904 24178 16960
rect 24030 15000 24086 15056
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24858 18944 24914 19000
rect 25042 18944 25098 19000
rect 25594 23296 25650 23352
rect 25410 20984 25466 21040
rect 25318 20440 25374 20496
rect 25226 18828 25282 18864
rect 25226 18808 25228 18828
rect 25228 18808 25280 18828
rect 25280 18808 25282 18828
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24398 16088 24454 16144
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 23846 10260 23902 10296
rect 23846 10240 23848 10260
rect 23848 10240 23900 10260
rect 23900 10240 23902 10260
rect 23662 9696 23718 9752
rect 23570 9152 23626 9208
rect 22558 5208 22614 5264
rect 21270 4820 21326 4856
rect 21270 4800 21272 4820
rect 21272 4800 21324 4820
rect 21324 4800 21326 4820
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 23846 9424 23902 9480
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24214 13776 24270 13832
rect 24674 13232 24730 13288
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24214 12824 24270 12880
rect 25226 17720 25282 17776
rect 25042 16940 25044 16960
rect 25044 16940 25096 16960
rect 25096 16940 25098 16960
rect 25042 16904 25098 16940
rect 24766 12416 24822 12472
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24030 9832 24086 9888
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24674 9968 24730 10024
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24858 12144 24914 12200
rect 25042 11600 25098 11656
rect 24950 10124 25006 10160
rect 24950 10104 24952 10124
rect 24952 10104 25004 10124
rect 25004 10104 25006 10124
rect 24950 9560 25006 9616
rect 24766 9288 24822 9344
rect 25134 10648 25190 10704
rect 25134 9152 25190 9208
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24766 8608 24822 8664
rect 24674 8064 24730 8120
rect 24950 8372 24952 8392
rect 24952 8372 25004 8392
rect 25004 8372 25006 8392
rect 24950 8336 25006 8372
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 23846 3032 23902 3088
rect 24766 7520 24822 7576
rect 24214 7384 24270 7440
rect 24582 6860 24638 6896
rect 24582 6840 24584 6860
rect 24584 6840 24636 6860
rect 24636 6840 24638 6860
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24766 6452 24822 6488
rect 24766 6432 24768 6452
rect 24768 6432 24820 6452
rect 24820 6432 24822 6452
rect 24858 6024 24914 6080
rect 24766 5908 24822 5944
rect 24766 5888 24768 5908
rect 24768 5888 24820 5908
rect 24820 5888 24822 5908
rect 24582 5772 24638 5808
rect 24582 5752 24584 5772
rect 24584 5752 24636 5772
rect 24636 5752 24638 5772
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24766 5364 24822 5400
rect 24766 5344 24768 5364
rect 24768 5344 24820 5364
rect 24820 5344 24822 5364
rect 24582 5208 24638 5264
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 25042 3340 25044 3360
rect 25044 3340 25096 3360
rect 25096 3340 25098 3360
rect 25042 3304 25098 3340
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 23662 1128 23718 1184
rect 23018 584 23074 640
rect 3514 312 3570 368
rect 25318 2796 25320 2816
rect 25320 2796 25372 2816
rect 25372 2796 25374 2816
rect 25318 2760 25374 2796
rect 25502 10104 25558 10160
rect 25686 4392 25742 4448
rect 25594 3848 25650 3904
rect 27066 22208 27122 22264
rect 26238 15816 26294 15872
rect 25870 3032 25926 3088
rect 25410 2216 25466 2272
rect 25502 1672 25558 1728
rect 25226 176 25282 232
<< metal3 >>
rect 0 27706 480 27736
rect 1301 27706 1367 27709
rect 0 27704 1367 27706
rect 0 27648 1306 27704
rect 1362 27648 1367 27704
rect 0 27646 1367 27648
rect 0 27616 480 27646
rect 1301 27643 1367 27646
rect 23565 27706 23631 27709
rect 27520 27706 28000 27736
rect 23565 27704 28000 27706
rect 23565 27648 23570 27704
rect 23626 27648 28000 27704
rect 23565 27646 28000 27648
rect 23565 27643 23631 27646
rect 27520 27616 28000 27646
rect 24761 27162 24827 27165
rect 27520 27162 28000 27192
rect 24761 27160 28000 27162
rect 24761 27104 24766 27160
rect 24822 27104 28000 27160
rect 24761 27102 28000 27104
rect 24761 27099 24827 27102
rect 27520 27072 28000 27102
rect 0 27026 480 27056
rect 1577 27026 1643 27029
rect 0 27024 1643 27026
rect 0 26968 1582 27024
rect 1638 26968 1643 27024
rect 0 26966 1643 26968
rect 0 26936 480 26966
rect 1577 26963 1643 26966
rect 24301 26618 24367 26621
rect 27520 26618 28000 26648
rect 24301 26616 28000 26618
rect 24301 26560 24306 26616
rect 24362 26560 28000 26616
rect 24301 26558 28000 26560
rect 24301 26555 24367 26558
rect 27520 26528 28000 26558
rect 0 26346 480 26376
rect 3785 26346 3851 26349
rect 0 26344 3851 26346
rect 0 26288 3790 26344
rect 3846 26288 3851 26344
rect 0 26286 3851 26288
rect 0 26256 480 26286
rect 3785 26283 3851 26286
rect 24761 26074 24827 26077
rect 27520 26074 28000 26104
rect 24761 26072 28000 26074
rect 24761 26016 24766 26072
rect 24822 26016 28000 26072
rect 24761 26014 28000 26016
rect 24761 26011 24827 26014
rect 27520 25984 28000 26014
rect 0 25666 480 25696
rect 3969 25666 4035 25669
rect 0 25664 4035 25666
rect 0 25608 3974 25664
rect 4030 25608 4035 25664
rect 0 25606 4035 25608
rect 0 25576 480 25606
rect 3969 25603 4035 25606
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 23933 25530 23999 25533
rect 27520 25530 28000 25560
rect 23933 25528 28000 25530
rect 23933 25472 23938 25528
rect 23994 25472 28000 25528
rect 23933 25470 28000 25472
rect 23933 25467 23999 25470
rect 27520 25440 28000 25470
rect 11329 25258 11395 25261
rect 17217 25258 17283 25261
rect 11329 25256 17283 25258
rect 11329 25200 11334 25256
rect 11390 25200 17222 25256
rect 17278 25200 17283 25256
rect 11329 25198 17283 25200
rect 11329 25195 11395 25198
rect 17217 25195 17283 25198
rect 0 25122 480 25152
rect 4061 25122 4127 25125
rect 0 25120 4127 25122
rect 0 25064 4066 25120
rect 4122 25064 4127 25120
rect 0 25062 4127 25064
rect 0 25032 480 25062
rect 4061 25059 4127 25062
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 25773 24986 25839 24989
rect 27520 24986 28000 25016
rect 25773 24984 28000 24986
rect 25773 24928 25778 24984
rect 25834 24928 28000 24984
rect 25773 24926 28000 24928
rect 25773 24923 25839 24926
rect 27520 24896 28000 24926
rect 1209 24850 1275 24853
rect 3693 24850 3759 24853
rect 1209 24848 3759 24850
rect 1209 24792 1214 24848
rect 1270 24792 3698 24848
rect 3754 24792 3759 24848
rect 1209 24790 3759 24792
rect 1209 24787 1275 24790
rect 3693 24787 3759 24790
rect 4981 24850 5047 24853
rect 8385 24850 8451 24853
rect 4981 24848 8451 24850
rect 4981 24792 4986 24848
rect 5042 24792 8390 24848
rect 8446 24792 8451 24848
rect 4981 24790 8451 24792
rect 4981 24787 5047 24790
rect 8385 24787 8451 24790
rect 12709 24850 12775 24853
rect 15377 24850 15443 24853
rect 12709 24848 15443 24850
rect 12709 24792 12714 24848
rect 12770 24792 15382 24848
rect 15438 24792 15443 24848
rect 12709 24790 15443 24792
rect 12709 24787 12775 24790
rect 15377 24787 15443 24790
rect 17861 24850 17927 24853
rect 20805 24850 20871 24853
rect 17861 24848 20871 24850
rect 17861 24792 17866 24848
rect 17922 24792 20810 24848
rect 20866 24792 20871 24848
rect 17861 24790 20871 24792
rect 17861 24787 17927 24790
rect 20805 24787 20871 24790
rect 21173 24850 21239 24853
rect 23841 24850 23907 24853
rect 21173 24848 23907 24850
rect 21173 24792 21178 24848
rect 21234 24792 23846 24848
rect 23902 24792 23907 24848
rect 21173 24790 23907 24792
rect 21173 24787 21239 24790
rect 23841 24787 23907 24790
rect 16481 24714 16547 24717
rect 18045 24714 18111 24717
rect 16481 24712 18111 24714
rect 16481 24656 16486 24712
rect 16542 24656 18050 24712
rect 18106 24656 18111 24712
rect 16481 24654 18111 24656
rect 16481 24651 16547 24654
rect 18045 24651 18111 24654
rect 18413 24714 18479 24717
rect 21909 24714 21975 24717
rect 18413 24712 21975 24714
rect 18413 24656 18418 24712
rect 18474 24656 21914 24712
rect 21970 24656 21975 24712
rect 18413 24654 21975 24656
rect 18413 24651 18479 24654
rect 21909 24651 21975 24654
rect 23289 24714 23355 24717
rect 24945 24714 25011 24717
rect 23289 24712 25011 24714
rect 23289 24656 23294 24712
rect 23350 24656 24950 24712
rect 25006 24656 25011 24712
rect 23289 24654 25011 24656
rect 23289 24651 23355 24654
rect 24945 24651 25011 24654
rect 2405 24578 2471 24581
rect 9949 24578 10015 24581
rect 2405 24576 10015 24578
rect 2405 24520 2410 24576
rect 2466 24520 9954 24576
rect 10010 24520 10015 24576
rect 2405 24518 10015 24520
rect 2405 24515 2471 24518
rect 9949 24515 10015 24518
rect 20529 24578 20595 24581
rect 24209 24578 24275 24581
rect 20529 24576 24275 24578
rect 20529 24520 20534 24576
rect 20590 24520 24214 24576
rect 24270 24520 24275 24576
rect 20529 24518 24275 24520
rect 20529 24515 20595 24518
rect 24209 24515 24275 24518
rect 10277 24512 10597 24513
rect 0 24442 480 24472
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 4797 24442 4863 24445
rect 0 24440 4863 24442
rect 0 24384 4802 24440
rect 4858 24384 4863 24440
rect 0 24382 4863 24384
rect 0 24352 480 24382
rect 4797 24379 4863 24382
rect 21633 24442 21699 24445
rect 24853 24442 24919 24445
rect 27520 24442 28000 24472
rect 21633 24440 24919 24442
rect 21633 24384 21638 24440
rect 21694 24384 24858 24440
rect 24914 24384 24919 24440
rect 21633 24382 24919 24384
rect 21633 24379 21699 24382
rect 24853 24379 24919 24382
rect 25454 24382 28000 24442
rect 7925 24306 7991 24309
rect 10041 24306 10107 24309
rect 19382 24306 19626 24340
rect 24761 24306 24827 24309
rect 7925 24304 10107 24306
rect 7925 24248 7930 24304
rect 7986 24248 10046 24304
rect 10102 24248 10107 24304
rect 7925 24246 10107 24248
rect 7925 24243 7991 24246
rect 10041 24243 10107 24246
rect 10182 24304 24827 24306
rect 10182 24280 24766 24304
rect 10182 24246 19442 24280
rect 19566 24248 24766 24280
rect 24822 24248 24827 24304
rect 19566 24246 24827 24248
rect 9949 24170 10015 24173
rect 10182 24170 10242 24246
rect 24761 24243 24827 24246
rect 9949 24168 10242 24170
rect 9949 24112 9954 24168
rect 10010 24112 10242 24168
rect 9949 24110 10242 24112
rect 12617 24170 12683 24173
rect 12985 24170 13051 24173
rect 17493 24170 17559 24173
rect 19333 24170 19399 24173
rect 12617 24168 15394 24170
rect 12617 24112 12622 24168
rect 12678 24112 12990 24168
rect 13046 24112 15394 24168
rect 12617 24110 15394 24112
rect 9949 24107 10015 24110
rect 12617 24107 12683 24110
rect 12985 24107 13051 24110
rect 8385 24034 8451 24037
rect 12341 24034 12407 24037
rect 8385 24032 12407 24034
rect 8385 23976 8390 24032
rect 8446 23976 12346 24032
rect 12402 23976 12407 24032
rect 8385 23974 12407 23976
rect 15334 24034 15394 24110
rect 17493 24168 19399 24170
rect 17493 24112 17498 24168
rect 17554 24112 19338 24168
rect 19394 24112 19399 24168
rect 17493 24110 19399 24112
rect 17493 24107 17559 24110
rect 19333 24107 19399 24110
rect 24117 24170 24183 24173
rect 25454 24170 25514 24382
rect 27520 24352 28000 24382
rect 24117 24168 25514 24170
rect 24117 24112 24122 24168
rect 24178 24112 25514 24168
rect 24117 24110 25514 24112
rect 24117 24107 24183 24110
rect 23105 24034 23171 24037
rect 15334 24032 23171 24034
rect 15334 23976 23110 24032
rect 23166 23976 23171 24032
rect 15334 23974 23171 23976
rect 8385 23971 8451 23974
rect 12341 23971 12407 23974
rect 23105 23971 23171 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 21449 23898 21515 23901
rect 17542 23896 21515 23898
rect 17542 23840 21454 23896
rect 21510 23840 21515 23896
rect 17542 23838 21515 23840
rect 0 23762 480 23792
rect 1761 23762 1827 23765
rect 0 23760 1827 23762
rect 0 23704 1766 23760
rect 1822 23704 1827 23760
rect 0 23702 1827 23704
rect 0 23672 480 23702
rect 1761 23699 1827 23702
rect 8477 23762 8543 23765
rect 17542 23762 17602 23838
rect 21449 23835 21515 23838
rect 21766 23836 21772 23900
rect 21836 23898 21842 23900
rect 21909 23898 21975 23901
rect 21836 23896 21975 23898
rect 21836 23840 21914 23896
rect 21970 23840 21975 23896
rect 21836 23838 21975 23840
rect 21836 23836 21842 23838
rect 21909 23835 21975 23838
rect 24761 23898 24827 23901
rect 27520 23898 28000 23928
rect 24761 23896 28000 23898
rect 24761 23840 24766 23896
rect 24822 23840 28000 23896
rect 24761 23838 28000 23840
rect 24761 23835 24827 23838
rect 27520 23808 28000 23838
rect 8477 23760 17602 23762
rect 8477 23704 8482 23760
rect 8538 23704 17602 23760
rect 8477 23702 17602 23704
rect 17677 23762 17743 23765
rect 19793 23762 19859 23765
rect 17677 23760 19859 23762
rect 17677 23704 17682 23760
rect 17738 23704 19798 23760
rect 19854 23704 19859 23760
rect 17677 23702 19859 23704
rect 8477 23699 8543 23702
rect 17677 23699 17743 23702
rect 19793 23699 19859 23702
rect 3233 23626 3299 23629
rect 12157 23626 12223 23629
rect 3233 23624 12223 23626
rect 3233 23568 3238 23624
rect 3294 23568 12162 23624
rect 12218 23568 12223 23624
rect 3233 23566 12223 23568
rect 3233 23563 3299 23566
rect 12157 23563 12223 23566
rect 12341 23626 12407 23629
rect 21817 23626 21883 23629
rect 12341 23624 21883 23626
rect 12341 23568 12346 23624
rect 12402 23568 21822 23624
rect 21878 23568 21883 23624
rect 12341 23566 21883 23568
rect 12341 23563 12407 23566
rect 21817 23563 21883 23566
rect 4521 23490 4587 23493
rect 9949 23490 10015 23493
rect 4521 23488 10015 23490
rect 4521 23432 4526 23488
rect 4582 23432 9954 23488
rect 10010 23432 10015 23488
rect 4521 23430 10015 23432
rect 4521 23427 4587 23430
rect 9949 23427 10015 23430
rect 11513 23490 11579 23493
rect 14273 23490 14339 23493
rect 11513 23488 14339 23490
rect 11513 23432 11518 23488
rect 11574 23432 14278 23488
rect 14334 23432 14339 23488
rect 11513 23430 14339 23432
rect 11513 23427 11579 23430
rect 14273 23427 14339 23430
rect 25221 23490 25287 23493
rect 27520 23490 28000 23520
rect 25221 23488 28000 23490
rect 25221 23432 25226 23488
rect 25282 23432 28000 23488
rect 25221 23430 28000 23432
rect 25221 23427 25287 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 27520 23400 28000 23430
rect 19610 23359 19930 23360
rect 5993 23354 6059 23357
rect 7281 23354 7347 23357
rect 5993 23352 7347 23354
rect 5993 23296 5998 23352
rect 6054 23296 7286 23352
rect 7342 23296 7347 23352
rect 5993 23294 7347 23296
rect 5993 23291 6059 23294
rect 7281 23291 7347 23294
rect 10961 23354 11027 23357
rect 15745 23354 15811 23357
rect 18229 23354 18295 23357
rect 10961 23352 15578 23354
rect 10961 23296 10966 23352
rect 11022 23296 15578 23352
rect 10961 23294 15578 23296
rect 10961 23291 11027 23294
rect 3509 23218 3575 23221
rect 6269 23218 6335 23221
rect 3509 23216 6335 23218
rect 3509 23160 3514 23216
rect 3570 23160 6274 23216
rect 6330 23160 6335 23216
rect 3509 23158 6335 23160
rect 3509 23155 3575 23158
rect 6269 23155 6335 23158
rect 9489 23218 9555 23221
rect 11053 23218 11119 23221
rect 9489 23216 11119 23218
rect 9489 23160 9494 23216
rect 9550 23160 11058 23216
rect 11114 23160 11119 23216
rect 9489 23158 11119 23160
rect 9489 23155 9555 23158
rect 11053 23155 11119 23158
rect 13721 23218 13787 23221
rect 15285 23218 15351 23221
rect 13721 23216 15351 23218
rect 13721 23160 13726 23216
rect 13782 23160 15290 23216
rect 15346 23160 15351 23216
rect 13721 23158 15351 23160
rect 15518 23218 15578 23294
rect 15745 23352 18295 23354
rect 15745 23296 15750 23352
rect 15806 23296 18234 23352
rect 18290 23296 18295 23352
rect 15745 23294 18295 23296
rect 15745 23291 15811 23294
rect 18229 23291 18295 23294
rect 20529 23354 20595 23357
rect 25589 23354 25655 23357
rect 20529 23352 25655 23354
rect 20529 23296 20534 23352
rect 20590 23296 25594 23352
rect 25650 23296 25655 23352
rect 20529 23294 25655 23296
rect 20529 23291 20595 23294
rect 25589 23291 25655 23294
rect 19333 23218 19399 23221
rect 15518 23216 19399 23218
rect 15518 23160 19338 23216
rect 19394 23160 19399 23216
rect 15518 23158 19399 23160
rect 13721 23155 13787 23158
rect 15285 23155 15351 23158
rect 19333 23155 19399 23158
rect 19793 23218 19859 23221
rect 24025 23218 24091 23221
rect 19793 23216 24091 23218
rect 19793 23160 19798 23216
rect 19854 23160 24030 23216
rect 24086 23160 24091 23216
rect 19793 23158 24091 23160
rect 19793 23155 19859 23158
rect 24025 23155 24091 23158
rect 0 23082 480 23112
rect 11237 23082 11303 23085
rect 20805 23082 20871 23085
rect 0 23080 11303 23082
rect 0 23024 11242 23080
rect 11298 23024 11303 23080
rect 0 23022 11303 23024
rect 0 22992 480 23022
rect 11237 23019 11303 23022
rect 14046 23080 20871 23082
rect 14046 23024 20810 23080
rect 20866 23024 20871 23080
rect 14046 23022 20871 23024
rect 14046 22949 14106 23022
rect 20805 23019 20871 23022
rect 22829 23082 22895 23085
rect 25129 23082 25195 23085
rect 22829 23080 25195 23082
rect 22829 23024 22834 23080
rect 22890 23024 25134 23080
rect 25190 23024 25195 23080
rect 22829 23022 25195 23024
rect 22829 23019 22895 23022
rect 25129 23019 25195 23022
rect 8569 22946 8635 22949
rect 12985 22946 13051 22949
rect 8569 22944 13051 22946
rect 8569 22888 8574 22944
rect 8630 22888 12990 22944
rect 13046 22888 13051 22944
rect 8569 22886 13051 22888
rect 8569 22883 8635 22886
rect 12985 22883 13051 22886
rect 13997 22944 14106 22949
rect 13997 22888 14002 22944
rect 14058 22888 14106 22944
rect 13997 22886 14106 22888
rect 17401 22946 17467 22949
rect 21633 22946 21699 22949
rect 27520 22946 28000 22976
rect 17401 22944 21699 22946
rect 17401 22888 17406 22944
rect 17462 22888 21638 22944
rect 21694 22888 21699 22944
rect 17401 22886 21699 22888
rect 13997 22883 14063 22886
rect 17401 22883 17467 22886
rect 21633 22883 21699 22886
rect 25086 22886 28000 22946
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 11605 22810 11671 22813
rect 7790 22808 11671 22810
rect 7790 22752 11610 22808
rect 11666 22752 11671 22808
rect 7790 22750 11671 22752
rect 3969 22674 4035 22677
rect 7790 22674 7850 22750
rect 11605 22747 11671 22750
rect 15469 22810 15535 22813
rect 21265 22810 21331 22813
rect 15469 22808 21331 22810
rect 15469 22752 15474 22808
rect 15530 22752 21270 22808
rect 21326 22752 21331 22808
rect 15469 22750 21331 22752
rect 15469 22747 15535 22750
rect 21265 22747 21331 22750
rect 21449 22810 21515 22813
rect 23749 22810 23815 22813
rect 21449 22808 23815 22810
rect 21449 22752 21454 22808
rect 21510 22752 23754 22808
rect 23810 22752 23815 22808
rect 21449 22750 23815 22752
rect 21449 22747 21515 22750
rect 23749 22747 23815 22750
rect 8109 22676 8175 22677
rect 8109 22674 8156 22676
rect 3969 22672 7850 22674
rect 3969 22616 3974 22672
rect 4030 22616 7850 22672
rect 3969 22614 7850 22616
rect 8028 22672 8156 22674
rect 8220 22674 8226 22676
rect 12249 22674 12315 22677
rect 8220 22672 12315 22674
rect 8028 22616 8114 22672
rect 8220 22616 12254 22672
rect 12310 22616 12315 22672
rect 8028 22614 8156 22616
rect 3969 22611 4035 22614
rect 8109 22612 8156 22614
rect 8220 22614 12315 22616
rect 8220 22612 8226 22614
rect 8109 22611 8175 22612
rect 12249 22611 12315 22614
rect 19374 22612 19380 22676
rect 19444 22674 19450 22676
rect 19885 22674 19951 22677
rect 19444 22672 19951 22674
rect 19444 22616 19890 22672
rect 19946 22616 19951 22672
rect 19444 22614 19951 22616
rect 19444 22612 19450 22614
rect 19885 22611 19951 22614
rect 23289 22674 23355 22677
rect 25086 22674 25146 22886
rect 27520 22856 28000 22886
rect 23289 22672 25146 22674
rect 23289 22616 23294 22672
rect 23350 22616 25146 22672
rect 23289 22614 25146 22616
rect 23289 22611 23355 22614
rect 1945 22538 2011 22541
rect 2957 22538 3023 22541
rect 1945 22536 3023 22538
rect 1945 22480 1950 22536
rect 2006 22480 2962 22536
rect 3018 22480 3023 22536
rect 1945 22478 3023 22480
rect 1945 22475 2011 22478
rect 2957 22475 3023 22478
rect 3693 22538 3759 22541
rect 4521 22538 4587 22541
rect 3693 22536 4587 22538
rect 3693 22480 3698 22536
rect 3754 22480 4526 22536
rect 4582 22480 4587 22536
rect 3693 22478 4587 22480
rect 3693 22475 3759 22478
rect 4521 22475 4587 22478
rect 5441 22538 5507 22541
rect 12341 22538 12407 22541
rect 5441 22536 12407 22538
rect 5441 22480 5446 22536
rect 5502 22480 12346 22536
rect 12402 22480 12407 22536
rect 5441 22478 12407 22480
rect 5441 22475 5507 22478
rect 12341 22475 12407 22478
rect 12617 22538 12683 22541
rect 16757 22538 16823 22541
rect 23197 22538 23263 22541
rect 12617 22536 23263 22538
rect 12617 22480 12622 22536
rect 12678 22480 16762 22536
rect 16818 22480 23202 22536
rect 23258 22480 23263 22536
rect 12617 22478 23263 22480
rect 12617 22475 12683 22478
rect 16757 22475 16823 22478
rect 23197 22475 23263 22478
rect 0 22402 480 22432
rect 565 22402 631 22405
rect 0 22400 631 22402
rect 0 22344 570 22400
rect 626 22344 631 22400
rect 0 22342 631 22344
rect 0 22312 480 22342
rect 565 22339 631 22342
rect 11237 22402 11303 22405
rect 15745 22402 15811 22405
rect 23105 22402 23171 22405
rect 27520 22402 28000 22432
rect 11237 22400 15811 22402
rect 11237 22344 11242 22400
rect 11298 22344 15750 22400
rect 15806 22344 15811 22400
rect 11237 22342 15811 22344
rect 11237 22339 11303 22342
rect 15745 22339 15811 22342
rect 20118 22400 28000 22402
rect 20118 22344 23110 22400
rect 23166 22344 28000 22400
rect 20118 22342 28000 22344
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 3049 22266 3115 22269
rect 3785 22266 3851 22269
rect 7833 22266 7899 22269
rect 10041 22266 10107 22269
rect 3049 22264 7899 22266
rect 3049 22208 3054 22264
rect 3110 22208 3790 22264
rect 3846 22208 7838 22264
rect 7894 22208 7899 22264
rect 3049 22206 7899 22208
rect 3049 22203 3115 22206
rect 3785 22203 3851 22206
rect 7833 22203 7899 22206
rect 7974 22264 10107 22266
rect 7974 22208 10046 22264
rect 10102 22208 10107 22264
rect 7974 22206 10107 22208
rect 197 22130 263 22133
rect 2957 22130 3023 22133
rect 3969 22130 4035 22133
rect 197 22128 4035 22130
rect 197 22072 202 22128
rect 258 22072 2962 22128
rect 3018 22072 3974 22128
rect 4030 22072 4035 22128
rect 197 22070 4035 22072
rect 197 22067 263 22070
rect 2957 22067 3023 22070
rect 3969 22067 4035 22070
rect 4521 22130 4587 22133
rect 7974 22130 8034 22206
rect 10041 22203 10107 22206
rect 4521 22128 8034 22130
rect 4521 22072 4526 22128
rect 4582 22072 8034 22128
rect 4521 22070 8034 22072
rect 9489 22130 9555 22133
rect 11329 22130 11395 22133
rect 9489 22128 11395 22130
rect 9489 22072 9494 22128
rect 9550 22072 11334 22128
rect 11390 22072 11395 22128
rect 9489 22070 11395 22072
rect 4521 22067 4587 22070
rect 9489 22067 9555 22070
rect 11329 22067 11395 22070
rect 19241 22130 19307 22133
rect 20118 22130 20178 22342
rect 23105 22339 23171 22342
rect 27520 22312 28000 22342
rect 20805 22266 20871 22269
rect 27061 22266 27127 22269
rect 20805 22264 27127 22266
rect 20805 22208 20810 22264
rect 20866 22208 27066 22264
rect 27122 22208 27127 22264
rect 20805 22206 27127 22208
rect 20805 22203 20871 22206
rect 27061 22203 27127 22206
rect 19241 22128 20178 22130
rect 19241 22072 19246 22128
rect 19302 22072 20178 22128
rect 19241 22070 20178 22072
rect 21173 22130 21239 22133
rect 22737 22130 22803 22133
rect 21173 22128 22803 22130
rect 21173 22072 21178 22128
rect 21234 22072 22742 22128
rect 22798 22072 22803 22128
rect 21173 22070 22803 22072
rect 19241 22067 19307 22070
rect 21173 22067 21239 22070
rect 22737 22067 22803 22070
rect 2405 21994 2471 21997
rect 4337 21994 4403 21997
rect 2405 21992 4403 21994
rect 2405 21936 2410 21992
rect 2466 21936 4342 21992
rect 4398 21936 4403 21992
rect 2405 21934 4403 21936
rect 2405 21931 2471 21934
rect 4337 21931 4403 21934
rect 4613 21994 4679 21997
rect 25221 21994 25287 21997
rect 4613 21992 25287 21994
rect 4613 21936 4618 21992
rect 4674 21936 25226 21992
rect 25282 21936 25287 21992
rect 4613 21934 25287 21936
rect 4613 21931 4679 21934
rect 25221 21931 25287 21934
rect 0 21858 480 21888
rect 8201 21858 8267 21861
rect 8661 21858 8727 21861
rect 9949 21858 10015 21861
rect 0 21798 4906 21858
rect 0 21768 480 21798
rect 4846 21586 4906 21798
rect 8201 21856 10015 21858
rect 8201 21800 8206 21856
rect 8262 21800 8666 21856
rect 8722 21800 9954 21856
rect 10010 21800 10015 21856
rect 8201 21798 10015 21800
rect 8201 21795 8267 21798
rect 8661 21795 8727 21798
rect 9949 21795 10015 21798
rect 10409 21858 10475 21861
rect 12065 21858 12131 21861
rect 13813 21858 13879 21861
rect 10409 21856 13879 21858
rect 10409 21800 10414 21856
rect 10470 21800 12070 21856
rect 12126 21800 13818 21856
rect 13874 21800 13879 21856
rect 10409 21798 13879 21800
rect 10409 21795 10475 21798
rect 12065 21795 12131 21798
rect 13813 21795 13879 21798
rect 19149 21858 19215 21861
rect 21081 21858 21147 21861
rect 27520 21858 28000 21888
rect 19149 21856 21147 21858
rect 19149 21800 19154 21856
rect 19210 21800 21086 21856
rect 21142 21800 21147 21856
rect 19149 21798 21147 21800
rect 19149 21795 19215 21798
rect 21081 21795 21147 21798
rect 24718 21798 28000 21858
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 9489 21722 9555 21725
rect 9489 21720 13554 21722
rect 9489 21664 9494 21720
rect 9550 21664 13554 21720
rect 9489 21662 13554 21664
rect 9489 21659 9555 21662
rect 4846 21526 10794 21586
rect 1669 21450 1735 21453
rect 7005 21450 7071 21453
rect 1669 21448 7071 21450
rect 1669 21392 1674 21448
rect 1730 21392 7010 21448
rect 7066 21392 7071 21448
rect 1669 21390 7071 21392
rect 1669 21387 1735 21390
rect 7005 21387 7071 21390
rect 10734 21314 10794 21526
rect 11237 21450 11303 21453
rect 12433 21450 12499 21453
rect 13261 21450 13327 21453
rect 11237 21448 13327 21450
rect 11237 21392 11242 21448
rect 11298 21392 12438 21448
rect 12494 21392 13266 21448
rect 13322 21392 13327 21448
rect 11237 21390 13327 21392
rect 13494 21450 13554 21662
rect 13629 21586 13695 21589
rect 15377 21586 15443 21589
rect 13629 21584 15443 21586
rect 13629 21528 13634 21584
rect 13690 21528 15382 21584
rect 15438 21528 15443 21584
rect 13629 21526 15443 21528
rect 13629 21523 13695 21526
rect 15377 21523 15443 21526
rect 23473 21586 23539 21589
rect 24209 21586 24275 21589
rect 24718 21586 24778 21798
rect 27520 21768 28000 21798
rect 23473 21584 24778 21586
rect 23473 21528 23478 21584
rect 23534 21528 24214 21584
rect 24270 21528 24778 21584
rect 23473 21526 24778 21528
rect 23473 21523 23539 21526
rect 24209 21523 24275 21526
rect 20437 21450 20503 21453
rect 13494 21448 20503 21450
rect 13494 21392 20442 21448
rect 20498 21392 20503 21448
rect 13494 21390 20503 21392
rect 11237 21387 11303 21390
rect 12433 21387 12499 21390
rect 13261 21387 13327 21390
rect 20437 21387 20503 21390
rect 23013 21450 23079 21453
rect 25037 21450 25103 21453
rect 23013 21448 25103 21450
rect 23013 21392 23018 21448
rect 23074 21392 25042 21448
rect 25098 21392 25103 21448
rect 23013 21390 25103 21392
rect 23013 21387 23079 21390
rect 25037 21387 25103 21390
rect 14457 21314 14523 21317
rect 16389 21314 16455 21317
rect 18137 21314 18203 21317
rect 10734 21254 14290 21314
rect 10277 21248 10597 21249
rect 0 21178 480 21208
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 1761 21178 1827 21181
rect 0 21176 1827 21178
rect 0 21120 1766 21176
rect 1822 21120 1827 21176
rect 0 21118 1827 21120
rect 14230 21178 14290 21254
rect 14457 21312 18203 21314
rect 14457 21256 14462 21312
rect 14518 21256 16394 21312
rect 16450 21256 18142 21312
rect 18198 21256 18203 21312
rect 14457 21254 18203 21256
rect 14457 21251 14523 21254
rect 16389 21251 16455 21254
rect 18137 21251 18203 21254
rect 20069 21314 20135 21317
rect 27520 21314 28000 21344
rect 20069 21312 28000 21314
rect 20069 21256 20074 21312
rect 20130 21256 28000 21312
rect 20069 21254 28000 21256
rect 20069 21251 20135 21254
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 27520 21224 28000 21254
rect 19610 21183 19930 21184
rect 15837 21178 15903 21181
rect 14230 21176 15903 21178
rect 14230 21120 15842 21176
rect 15898 21120 15903 21176
rect 14230 21118 15903 21120
rect 0 21088 480 21118
rect 1761 21115 1827 21118
rect 15837 21115 15903 21118
rect 16021 21178 16087 21181
rect 19333 21178 19399 21181
rect 16021 21176 19399 21178
rect 16021 21120 16026 21176
rect 16082 21120 19338 21176
rect 19394 21120 19399 21176
rect 16021 21118 19399 21120
rect 16021 21115 16087 21118
rect 19333 21115 19399 21118
rect 23841 21178 23907 21181
rect 24209 21178 24275 21181
rect 23841 21176 24275 21178
rect 23841 21120 23846 21176
rect 23902 21120 24214 21176
rect 24270 21120 24275 21176
rect 23841 21118 24275 21120
rect 23841 21115 23907 21118
rect 24209 21115 24275 21118
rect 8385 21042 8451 21045
rect 20253 21042 20319 21045
rect 8385 21040 20319 21042
rect 8385 20984 8390 21040
rect 8446 20984 20258 21040
rect 20314 20984 20319 21040
rect 8385 20982 20319 20984
rect 8385 20979 8451 20982
rect 20253 20979 20319 20982
rect 23289 21042 23355 21045
rect 25405 21042 25471 21045
rect 23289 21040 25471 21042
rect 23289 20984 23294 21040
rect 23350 20984 25410 21040
rect 25466 20984 25471 21040
rect 23289 20982 25471 20984
rect 23289 20979 23355 20982
rect 25405 20979 25471 20982
rect 7833 20904 7899 20909
rect 7833 20848 7838 20904
rect 7894 20848 7899 20904
rect 7833 20843 7899 20848
rect 8201 20906 8267 20909
rect 11237 20906 11303 20909
rect 8201 20904 11303 20906
rect 8201 20848 8206 20904
rect 8262 20848 11242 20904
rect 11298 20848 11303 20904
rect 8201 20846 11303 20848
rect 8201 20843 8267 20846
rect 11237 20843 11303 20846
rect 13261 20906 13327 20909
rect 13261 20904 24916 20906
rect 13261 20848 13266 20904
rect 13322 20848 24916 20904
rect 13261 20846 24916 20848
rect 13261 20843 13327 20846
rect 7836 20770 7896 20843
rect 14457 20770 14523 20773
rect 7836 20768 14523 20770
rect 7836 20712 14462 20768
rect 14518 20712 14523 20768
rect 7836 20710 14523 20712
rect 14457 20707 14523 20710
rect 15837 20770 15903 20773
rect 17493 20770 17559 20773
rect 15837 20768 17559 20770
rect 15837 20712 15842 20768
rect 15898 20712 17498 20768
rect 17554 20712 17559 20768
rect 15837 20710 17559 20712
rect 24856 20770 24916 20846
rect 27520 20770 28000 20800
rect 24856 20710 28000 20770
rect 15837 20707 15903 20710
rect 17493 20707 17559 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 27520 20680 28000 20710
rect 24277 20639 24597 20640
rect 10317 20634 10383 20637
rect 13997 20634 14063 20637
rect 10317 20632 14063 20634
rect 10317 20576 10322 20632
rect 10378 20576 14002 20632
rect 14058 20576 14063 20632
rect 10317 20574 14063 20576
rect 10317 20571 10383 20574
rect 13997 20571 14063 20574
rect 14222 20572 14228 20636
rect 14292 20634 14298 20636
rect 18137 20634 18203 20637
rect 19374 20634 19380 20636
rect 14292 20574 14842 20634
rect 18010 20632 19380 20634
rect 18010 20576 18142 20632
rect 18198 20576 19380 20632
rect 18010 20574 19380 20576
rect 14292 20572 14298 20574
rect 0 20498 480 20528
rect 7557 20498 7623 20501
rect 0 20496 7623 20498
rect 0 20440 7562 20496
rect 7618 20440 7623 20496
rect 0 20438 7623 20440
rect 0 20408 480 20438
rect 7557 20435 7623 20438
rect 9397 20498 9463 20501
rect 14273 20498 14339 20501
rect 9397 20496 14339 20498
rect 9397 20440 9402 20496
rect 9458 20440 14278 20496
rect 14334 20440 14339 20496
rect 9397 20438 14339 20440
rect 14782 20498 14842 20574
rect 18094 20571 18203 20574
rect 19374 20572 19380 20574
rect 19444 20572 19450 20636
rect 18094 20498 18154 20571
rect 14782 20438 18154 20498
rect 18229 20498 18295 20501
rect 25313 20498 25379 20501
rect 18229 20496 25379 20498
rect 18229 20440 18234 20496
rect 18290 20440 25318 20496
rect 25374 20440 25379 20496
rect 18229 20438 25379 20440
rect 9397 20435 9463 20438
rect 14273 20435 14339 20438
rect 18229 20435 18295 20438
rect 25313 20435 25379 20438
rect 4981 20362 5047 20365
rect 11053 20362 11119 20365
rect 13670 20362 13676 20364
rect 4981 20360 10794 20362
rect 4981 20304 4986 20360
rect 5042 20304 10794 20360
rect 4981 20302 10794 20304
rect 4981 20299 5047 20302
rect 3877 20226 3943 20229
rect 8753 20226 8819 20229
rect 9581 20226 9647 20229
rect 3877 20224 9647 20226
rect 3877 20168 3882 20224
rect 3938 20168 8758 20224
rect 8814 20168 9586 20224
rect 9642 20168 9647 20224
rect 3877 20166 9647 20168
rect 10734 20226 10794 20302
rect 11053 20360 13676 20362
rect 11053 20304 11058 20360
rect 11114 20304 13676 20360
rect 11053 20302 13676 20304
rect 11053 20299 11119 20302
rect 13670 20300 13676 20302
rect 13740 20300 13746 20364
rect 13905 20362 13971 20365
rect 13905 20360 24916 20362
rect 13905 20304 13910 20360
rect 13966 20304 24916 20360
rect 13905 20302 24916 20304
rect 13905 20299 13971 20302
rect 14641 20226 14707 20229
rect 10734 20224 14707 20226
rect 10734 20168 14646 20224
rect 14702 20168 14707 20224
rect 10734 20166 14707 20168
rect 3877 20163 3943 20166
rect 8753 20163 8819 20166
rect 9581 20163 9647 20166
rect 14641 20163 14707 20166
rect 15285 20226 15351 20229
rect 15469 20226 15535 20229
rect 15285 20224 15535 20226
rect 15285 20168 15290 20224
rect 15346 20168 15474 20224
rect 15530 20168 15535 20224
rect 15285 20166 15535 20168
rect 15285 20163 15351 20166
rect 15469 20163 15535 20166
rect 15745 20226 15811 20229
rect 15878 20226 15884 20228
rect 15745 20224 15884 20226
rect 15745 20168 15750 20224
rect 15806 20168 15884 20224
rect 15745 20166 15884 20168
rect 15745 20163 15811 20166
rect 15878 20164 15884 20166
rect 15948 20164 15954 20228
rect 16389 20226 16455 20229
rect 18597 20226 18663 20229
rect 16389 20224 18663 20226
rect 16389 20168 16394 20224
rect 16450 20168 18602 20224
rect 18658 20168 18663 20224
rect 16389 20166 18663 20168
rect 24856 20226 24916 20302
rect 27520 20226 28000 20256
rect 24856 20166 28000 20226
rect 16389 20163 16455 20166
rect 18597 20163 18663 20166
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 27520 20136 28000 20166
rect 19610 20095 19930 20096
rect 4797 20090 4863 20093
rect 9765 20090 9831 20093
rect 4797 20088 9831 20090
rect 4797 20032 4802 20088
rect 4858 20032 9770 20088
rect 9826 20032 9831 20088
rect 4797 20030 9831 20032
rect 4797 20027 4863 20030
rect 9765 20027 9831 20030
rect 11145 20090 11211 20093
rect 15469 20090 15535 20093
rect 11145 20088 15535 20090
rect 11145 20032 11150 20088
rect 11206 20032 15474 20088
rect 15530 20032 15535 20088
rect 11145 20030 15535 20032
rect 11145 20027 11211 20030
rect 15469 20027 15535 20030
rect 7557 19954 7623 19957
rect 17217 19954 17283 19957
rect 7557 19952 17283 19954
rect 7557 19896 7562 19952
rect 7618 19896 17222 19952
rect 17278 19896 17283 19952
rect 7557 19894 17283 19896
rect 7557 19891 7623 19894
rect 17217 19891 17283 19894
rect 0 19818 480 19848
rect 11053 19818 11119 19821
rect 0 19816 11119 19818
rect 0 19760 11058 19816
rect 11114 19760 11119 19816
rect 0 19758 11119 19760
rect 0 19728 480 19758
rect 11053 19755 11119 19758
rect 12709 19818 12775 19821
rect 18321 19818 18387 19821
rect 12709 19816 18387 19818
rect 12709 19760 12714 19816
rect 12770 19760 18326 19816
rect 18382 19760 18387 19816
rect 12709 19758 18387 19760
rect 12709 19755 12775 19758
rect 18321 19755 18387 19758
rect 11145 19682 11211 19685
rect 5996 19680 11211 19682
rect 5996 19624 11150 19680
rect 11206 19624 11211 19680
rect 5996 19622 11211 19624
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 5996 19410 6056 19622
rect 11145 19619 11211 19622
rect 15745 19682 15811 19685
rect 19057 19682 19123 19685
rect 27520 19682 28000 19712
rect 15745 19680 19123 19682
rect 15745 19624 15750 19680
rect 15806 19624 19062 19680
rect 19118 19624 19123 19680
rect 15745 19622 19123 19624
rect 15745 19619 15811 19622
rect 19057 19619 19123 19622
rect 24856 19622 28000 19682
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 8385 19546 8451 19549
rect 12709 19546 12775 19549
rect 8385 19544 12775 19546
rect 8385 19488 8390 19544
rect 8446 19488 12714 19544
rect 12770 19488 12775 19544
rect 8385 19486 12775 19488
rect 8385 19483 8451 19486
rect 12709 19483 12775 19486
rect 3972 19350 6056 19410
rect 10961 19410 11027 19413
rect 24856 19410 24916 19622
rect 27520 19592 28000 19622
rect 10961 19408 24916 19410
rect 10961 19352 10966 19408
rect 11022 19352 24916 19408
rect 10961 19350 24916 19352
rect 2313 19274 2379 19277
rect 3785 19274 3851 19277
rect 2313 19272 3851 19274
rect 2313 19216 2318 19272
rect 2374 19216 3790 19272
rect 3846 19216 3851 19272
rect 2313 19214 3851 19216
rect 2313 19211 2379 19214
rect 3785 19211 3851 19214
rect 0 19138 480 19168
rect 3972 19138 4032 19350
rect 10961 19347 11027 19350
rect 4981 19274 5047 19277
rect 10777 19274 10843 19277
rect 4981 19272 10843 19274
rect 4981 19216 4986 19272
rect 5042 19216 10782 19272
rect 10838 19216 10843 19272
rect 4981 19214 10843 19216
rect 4981 19211 5047 19214
rect 10777 19211 10843 19214
rect 11053 19274 11119 19277
rect 13353 19274 13419 19277
rect 11053 19272 13419 19274
rect 11053 19216 11058 19272
rect 11114 19216 13358 19272
rect 13414 19216 13419 19272
rect 11053 19214 13419 19216
rect 11053 19211 11119 19214
rect 13353 19211 13419 19214
rect 14917 19274 14983 19277
rect 21541 19274 21607 19277
rect 24117 19274 24183 19277
rect 14917 19272 20178 19274
rect 14917 19216 14922 19272
rect 14978 19216 20178 19272
rect 14917 19214 20178 19216
rect 14917 19211 14983 19214
rect 0 19078 4032 19138
rect 13537 19138 13603 19141
rect 18597 19138 18663 19141
rect 13537 19136 18663 19138
rect 13537 19080 13542 19136
rect 13598 19080 18602 19136
rect 18658 19080 18663 19136
rect 13537 19078 18663 19080
rect 20118 19138 20178 19214
rect 21541 19272 24183 19274
rect 21541 19216 21546 19272
rect 21602 19216 24122 19272
rect 24178 19216 24183 19272
rect 21541 19214 24183 19216
rect 21541 19211 21607 19214
rect 24117 19211 24183 19214
rect 23933 19138 23999 19141
rect 27520 19138 28000 19168
rect 20118 19078 22386 19138
rect 0 19048 480 19078
rect 13537 19075 13603 19078
rect 18597 19075 18663 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 4705 19002 4771 19005
rect 9857 19002 9923 19005
rect 4705 19000 9923 19002
rect 4705 18944 4710 19000
rect 4766 18944 9862 19000
rect 9918 18944 9923 19000
rect 4705 18942 9923 18944
rect 4705 18939 4771 18942
rect 9857 18939 9923 18942
rect 1301 18866 1367 18869
rect 4981 18866 5047 18869
rect 1301 18864 5047 18866
rect 1301 18808 1306 18864
rect 1362 18808 4986 18864
rect 5042 18808 5047 18864
rect 1301 18806 5047 18808
rect 1301 18803 1367 18806
rect 4981 18803 5047 18806
rect 5257 18866 5323 18869
rect 11697 18866 11763 18869
rect 21173 18866 21239 18869
rect 5257 18864 11763 18866
rect 5257 18808 5262 18864
rect 5318 18808 11702 18864
rect 11758 18808 11763 18864
rect 5257 18806 11763 18808
rect 5257 18803 5323 18806
rect 11697 18803 11763 18806
rect 11838 18864 21239 18866
rect 11838 18808 21178 18864
rect 21234 18808 21239 18864
rect 11838 18806 21239 18808
rect 4797 18730 4863 18733
rect 5390 18730 5396 18732
rect 4797 18728 5396 18730
rect 4797 18672 4802 18728
rect 4858 18672 5396 18728
rect 4797 18670 5396 18672
rect 4797 18667 4863 18670
rect 5390 18668 5396 18670
rect 5460 18668 5466 18732
rect 7097 18730 7163 18733
rect 11838 18730 11898 18806
rect 21173 18803 21239 18806
rect 19517 18730 19583 18733
rect 7097 18728 11898 18730
rect 7097 18672 7102 18728
rect 7158 18672 11898 18728
rect 7097 18670 11898 18672
rect 14414 18728 19583 18730
rect 14414 18672 19522 18728
rect 19578 18672 19583 18728
rect 14414 18670 19583 18672
rect 22326 18730 22386 19078
rect 23933 19136 28000 19138
rect 23933 19080 23938 19136
rect 23994 19080 28000 19136
rect 23933 19078 28000 19080
rect 23933 19075 23999 19078
rect 27520 19048 28000 19078
rect 23105 19002 23171 19005
rect 24853 19002 24919 19005
rect 25037 19002 25103 19005
rect 23105 19000 25103 19002
rect 23105 18944 23110 19000
rect 23166 18944 24858 19000
rect 24914 18944 25042 19000
rect 25098 18944 25103 19000
rect 23105 18942 25103 18944
rect 23105 18939 23171 18942
rect 24853 18939 24919 18942
rect 25037 18939 25103 18942
rect 22461 18866 22527 18869
rect 25221 18866 25287 18869
rect 22461 18864 25287 18866
rect 22461 18808 22466 18864
rect 22522 18808 25226 18864
rect 25282 18808 25287 18864
rect 22461 18806 25287 18808
rect 22461 18803 22527 18806
rect 25221 18803 25287 18806
rect 27520 18730 28000 18760
rect 22326 18670 28000 18730
rect 7097 18667 7163 18670
rect 0 18594 480 18624
rect 2773 18594 2839 18597
rect 0 18592 2839 18594
rect 0 18536 2778 18592
rect 2834 18536 2839 18592
rect 0 18534 2839 18536
rect 0 18504 480 18534
rect 2773 18531 2839 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 3325 18458 3391 18461
rect 4797 18458 4863 18461
rect 3325 18456 4863 18458
rect 3325 18400 3330 18456
rect 3386 18400 4802 18456
rect 4858 18400 4863 18456
rect 3325 18398 4863 18400
rect 3325 18395 3391 18398
rect 4797 18395 4863 18398
rect 8477 18458 8543 18461
rect 14414 18458 14474 18670
rect 19517 18667 19583 18670
rect 27520 18640 28000 18670
rect 16941 18594 17007 18597
rect 16941 18592 19396 18594
rect 16941 18536 16946 18592
rect 17002 18536 19396 18592
rect 16941 18534 19396 18536
rect 16941 18531 17007 18534
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 8477 18456 14474 18458
rect 8477 18400 8482 18456
rect 8538 18400 14474 18456
rect 8477 18398 14474 18400
rect 19336 18458 19396 18534
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 22645 18458 22711 18461
rect 19336 18456 22711 18458
rect 19336 18400 22650 18456
rect 22706 18400 22711 18456
rect 19336 18398 22711 18400
rect 8477 18395 8543 18398
rect 22645 18395 22711 18398
rect 1485 18322 1551 18325
rect 6729 18322 6795 18325
rect 11053 18322 11119 18325
rect 1485 18320 6795 18322
rect 1485 18264 1490 18320
rect 1546 18264 6734 18320
rect 6790 18264 6795 18320
rect 1485 18262 6795 18264
rect 1485 18259 1551 18262
rect 6729 18259 6795 18262
rect 6870 18320 11119 18322
rect 6870 18264 11058 18320
rect 11114 18264 11119 18320
rect 6870 18262 11119 18264
rect 1761 18186 1827 18189
rect 5533 18186 5599 18189
rect 1761 18184 5599 18186
rect 1761 18128 1766 18184
rect 1822 18128 5538 18184
rect 5594 18128 5599 18184
rect 1761 18126 5599 18128
rect 1761 18123 1827 18126
rect 5533 18123 5599 18126
rect 3601 18050 3667 18053
rect 6870 18050 6930 18262
rect 11053 18259 11119 18262
rect 13445 18322 13511 18325
rect 17033 18322 17099 18325
rect 20161 18322 20227 18325
rect 23841 18324 23907 18325
rect 13445 18320 15532 18322
rect 13445 18264 13450 18320
rect 13506 18264 15532 18320
rect 13445 18262 15532 18264
rect 13445 18259 13511 18262
rect 10685 18186 10751 18189
rect 13537 18186 13603 18189
rect 10685 18184 13603 18186
rect 10685 18128 10690 18184
rect 10746 18128 13542 18184
rect 13598 18128 13603 18184
rect 10685 18126 13603 18128
rect 15472 18186 15532 18262
rect 17033 18320 20227 18322
rect 17033 18264 17038 18320
rect 17094 18264 20166 18320
rect 20222 18264 20227 18320
rect 17033 18262 20227 18264
rect 17033 18259 17099 18262
rect 20161 18259 20227 18262
rect 23790 18260 23796 18324
rect 23860 18322 23907 18324
rect 23860 18320 23952 18322
rect 23902 18264 23952 18320
rect 23860 18262 23952 18264
rect 23860 18260 23907 18262
rect 23841 18259 23907 18260
rect 27520 18186 28000 18216
rect 15472 18126 28000 18186
rect 10685 18123 10751 18126
rect 13537 18123 13603 18126
rect 27520 18096 28000 18126
rect 3601 18048 6930 18050
rect 3601 17992 3606 18048
rect 3662 17992 6930 18048
rect 3601 17990 6930 17992
rect 13261 18050 13327 18053
rect 15377 18050 15443 18053
rect 13261 18048 15443 18050
rect 13261 17992 13266 18048
rect 13322 17992 15382 18048
rect 15438 17992 15443 18048
rect 13261 17990 15443 17992
rect 3601 17987 3667 17990
rect 13261 17987 13327 17990
rect 15377 17987 15443 17990
rect 16205 18050 16271 18053
rect 18597 18050 18663 18053
rect 16205 18048 18663 18050
rect 16205 17992 16210 18048
rect 16266 17992 18602 18048
rect 18658 17992 18663 18048
rect 16205 17990 18663 17992
rect 16205 17987 16271 17990
rect 18597 17987 18663 17990
rect 10277 17984 10597 17985
rect 0 17914 480 17944
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 3969 17914 4035 17917
rect 0 17912 4035 17914
rect 0 17856 3974 17912
rect 4030 17856 4035 17912
rect 0 17854 4035 17856
rect 0 17824 480 17854
rect 3969 17851 4035 17854
rect 11513 17914 11579 17917
rect 13445 17914 13511 17917
rect 11513 17912 13511 17914
rect 11513 17856 11518 17912
rect 11574 17856 13450 17912
rect 13506 17856 13511 17912
rect 11513 17854 13511 17856
rect 11513 17851 11579 17854
rect 13445 17851 13511 17854
rect 5441 17778 5507 17781
rect 7833 17778 7899 17781
rect 9121 17778 9187 17781
rect 11697 17778 11763 17781
rect 5441 17776 11763 17778
rect 5441 17720 5446 17776
rect 5502 17720 7838 17776
rect 7894 17720 9126 17776
rect 9182 17720 11702 17776
rect 11758 17720 11763 17776
rect 5441 17718 11763 17720
rect 5441 17715 5507 17718
rect 7833 17715 7899 17718
rect 9121 17715 9187 17718
rect 11697 17715 11763 17718
rect 12157 17778 12223 17781
rect 19609 17778 19675 17781
rect 23473 17778 23539 17781
rect 25221 17778 25287 17781
rect 12157 17776 19675 17778
rect 12157 17720 12162 17776
rect 12218 17720 19614 17776
rect 19670 17720 19675 17776
rect 12157 17718 19675 17720
rect 12157 17715 12223 17718
rect 19609 17715 19675 17718
rect 19750 17776 23539 17778
rect 19750 17720 23478 17776
rect 23534 17720 23539 17776
rect 19750 17718 23539 17720
rect 12801 17642 12867 17645
rect 19750 17642 19810 17718
rect 23473 17715 23539 17718
rect 23614 17776 25287 17778
rect 23614 17720 25226 17776
rect 25282 17720 25287 17776
rect 23614 17718 25287 17720
rect 2270 17640 19810 17642
rect 2270 17584 12806 17640
rect 12862 17584 19810 17640
rect 2270 17582 19810 17584
rect 19977 17642 20043 17645
rect 23614 17642 23674 17718
rect 25221 17715 25287 17718
rect 27520 17642 28000 17672
rect 19977 17640 23674 17642
rect 19977 17584 19982 17640
rect 20038 17584 23674 17640
rect 19977 17582 23674 17584
rect 24856 17582 28000 17642
rect 0 17234 480 17264
rect 2270 17234 2330 17582
rect 12801 17579 12867 17582
rect 19977 17579 20043 17582
rect 19241 17506 19307 17509
rect 24025 17506 24091 17509
rect 19241 17504 24091 17506
rect 19241 17448 19246 17504
rect 19302 17448 24030 17504
rect 24086 17448 24091 17504
rect 19241 17446 24091 17448
rect 19241 17443 19307 17446
rect 24025 17443 24091 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 16021 17370 16087 17373
rect 23933 17370 23999 17373
rect 16021 17368 23999 17370
rect 16021 17312 16026 17368
rect 16082 17312 23938 17368
rect 23994 17312 23999 17368
rect 16021 17310 23999 17312
rect 16021 17307 16087 17310
rect 23933 17307 23999 17310
rect 0 17174 2330 17234
rect 18413 17234 18479 17237
rect 24856 17234 24916 17582
rect 27520 17552 28000 17582
rect 18413 17232 24916 17234
rect 18413 17176 18418 17232
rect 18474 17176 24916 17232
rect 18413 17174 24916 17176
rect 0 17144 480 17174
rect 18413 17171 18479 17174
rect 7649 17098 7715 17101
rect 13077 17098 13143 17101
rect 7649 17096 13143 17098
rect 7649 17040 7654 17096
rect 7710 17040 13082 17096
rect 13138 17040 13143 17096
rect 7649 17038 13143 17040
rect 7649 17035 7715 17038
rect 13077 17035 13143 17038
rect 13261 17098 13327 17101
rect 20989 17098 21055 17101
rect 27520 17098 28000 17128
rect 13261 17096 21055 17098
rect 13261 17040 13266 17096
rect 13322 17040 20994 17096
rect 21050 17040 21055 17096
rect 13261 17038 21055 17040
rect 13261 17035 13327 17038
rect 20989 17035 21055 17038
rect 25270 17038 28000 17098
rect 23657 16962 23723 16965
rect 24117 16962 24183 16965
rect 25037 16962 25103 16965
rect 23657 16960 25103 16962
rect 23657 16904 23662 16960
rect 23718 16904 24122 16960
rect 24178 16904 25042 16960
rect 25098 16904 25103 16960
rect 23657 16902 25103 16904
rect 23657 16899 23723 16902
rect 24117 16899 24183 16902
rect 25037 16899 25103 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 11973 16826 12039 16829
rect 13077 16826 13143 16829
rect 11973 16824 13143 16826
rect 11973 16768 11978 16824
rect 12034 16768 13082 16824
rect 13138 16768 13143 16824
rect 11973 16766 13143 16768
rect 11973 16763 12039 16766
rect 13077 16763 13143 16766
rect 2129 16690 2195 16693
rect 6085 16690 6151 16693
rect 2129 16688 6151 16690
rect 2129 16632 2134 16688
rect 2190 16632 6090 16688
rect 6146 16632 6151 16688
rect 2129 16630 6151 16632
rect 2129 16627 2195 16630
rect 6085 16627 6151 16630
rect 16297 16690 16363 16693
rect 25270 16690 25330 17038
rect 27520 17008 28000 17038
rect 16297 16688 25330 16690
rect 16297 16632 16302 16688
rect 16358 16632 25330 16688
rect 16297 16630 25330 16632
rect 16297 16627 16363 16630
rect 0 16554 480 16584
rect 8937 16554 9003 16557
rect 0 16552 9003 16554
rect 0 16496 8942 16552
rect 8998 16496 9003 16552
rect 0 16494 9003 16496
rect 0 16464 480 16494
rect 8937 16491 9003 16494
rect 9121 16554 9187 16557
rect 16849 16554 16915 16557
rect 9121 16552 16915 16554
rect 9121 16496 9126 16552
rect 9182 16496 16854 16552
rect 16910 16496 16915 16552
rect 9121 16494 16915 16496
rect 9121 16491 9187 16494
rect 16849 16491 16915 16494
rect 17033 16554 17099 16557
rect 19425 16554 19491 16557
rect 17033 16552 19491 16554
rect 17033 16496 17038 16552
rect 17094 16496 19430 16552
rect 19486 16496 19491 16552
rect 17033 16494 19491 16496
rect 17033 16491 17099 16494
rect 19425 16491 19491 16494
rect 23197 16554 23263 16557
rect 27520 16554 28000 16584
rect 23197 16552 28000 16554
rect 23197 16496 23202 16552
rect 23258 16496 28000 16552
rect 23197 16494 28000 16496
rect 23197 16491 23263 16494
rect 27520 16464 28000 16494
rect 8293 16418 8359 16421
rect 14089 16418 14155 16421
rect 8293 16416 14155 16418
rect 8293 16360 8298 16416
rect 8354 16360 14094 16416
rect 14150 16360 14155 16416
rect 8293 16358 14155 16360
rect 8293 16355 8359 16358
rect 14089 16355 14155 16358
rect 18321 16418 18387 16421
rect 22461 16418 22527 16421
rect 18321 16416 22527 16418
rect 18321 16360 18326 16416
rect 18382 16360 22466 16416
rect 22522 16360 22527 16416
rect 18321 16358 22527 16360
rect 18321 16355 18387 16358
rect 22461 16355 22527 16358
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 7373 16282 7439 16285
rect 5996 16280 7439 16282
rect 5996 16224 7378 16280
rect 7434 16224 7439 16280
rect 5996 16222 7439 16224
rect 4153 16146 4219 16149
rect 5996 16146 6056 16222
rect 7373 16219 7439 16222
rect 8201 16282 8267 16285
rect 9121 16282 9187 16285
rect 8201 16280 9187 16282
rect 8201 16224 8206 16280
rect 8262 16224 9126 16280
rect 9182 16224 9187 16280
rect 8201 16222 9187 16224
rect 8201 16219 8267 16222
rect 9121 16219 9187 16222
rect 9397 16282 9463 16285
rect 9949 16282 10015 16285
rect 14549 16282 14615 16285
rect 9397 16280 14615 16282
rect 9397 16224 9402 16280
rect 9458 16224 9954 16280
rect 10010 16224 14554 16280
rect 14610 16224 14615 16280
rect 9397 16222 14615 16224
rect 9397 16219 9463 16222
rect 9949 16219 10015 16222
rect 14549 16219 14615 16222
rect 18137 16282 18203 16285
rect 18965 16282 19031 16285
rect 18137 16280 19031 16282
rect 18137 16224 18142 16280
rect 18198 16224 18970 16280
rect 19026 16224 19031 16280
rect 18137 16222 19031 16224
rect 18137 16219 18203 16222
rect 18965 16219 19031 16222
rect 4153 16144 6056 16146
rect 4153 16088 4158 16144
rect 4214 16088 6056 16144
rect 4153 16086 6056 16088
rect 13813 16146 13879 16149
rect 24393 16146 24459 16149
rect 13813 16144 24459 16146
rect 13813 16088 13818 16144
rect 13874 16088 24398 16144
rect 24454 16088 24459 16144
rect 13813 16086 24459 16088
rect 4153 16083 4219 16086
rect 13813 16083 13879 16086
rect 24393 16083 24459 16086
rect 3969 16010 4035 16013
rect 13169 16010 13235 16013
rect 3969 16008 13235 16010
rect 3969 15952 3974 16008
rect 4030 15952 13174 16008
rect 13230 15952 13235 16008
rect 3969 15950 13235 15952
rect 3969 15947 4035 15950
rect 13169 15947 13235 15950
rect 20069 16010 20135 16013
rect 27520 16010 28000 16040
rect 20069 16008 28000 16010
rect 20069 15952 20074 16008
rect 20130 15952 28000 16008
rect 20069 15950 28000 15952
rect 20069 15947 20135 15950
rect 27520 15920 28000 15950
rect 0 15874 480 15904
rect 4061 15874 4127 15877
rect 0 15872 4127 15874
rect 0 15816 4066 15872
rect 4122 15816 4127 15872
rect 0 15814 4127 15816
rect 0 15784 480 15814
rect 4061 15811 4127 15814
rect 5993 15874 6059 15877
rect 7005 15874 7071 15877
rect 5993 15872 7071 15874
rect 5993 15816 5998 15872
rect 6054 15816 7010 15872
rect 7066 15816 7071 15872
rect 5993 15814 7071 15816
rect 5993 15811 6059 15814
rect 7005 15811 7071 15814
rect 12709 15874 12775 15877
rect 18597 15874 18663 15877
rect 12709 15872 18663 15874
rect 12709 15816 12714 15872
rect 12770 15816 18602 15872
rect 18658 15816 18663 15872
rect 12709 15814 18663 15816
rect 12709 15811 12775 15814
rect 18597 15811 18663 15814
rect 23105 15874 23171 15877
rect 26233 15874 26299 15877
rect 23105 15872 26299 15874
rect 23105 15816 23110 15872
rect 23166 15816 26238 15872
rect 26294 15816 26299 15872
rect 23105 15814 26299 15816
rect 23105 15811 23171 15814
rect 26233 15811 26299 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 13629 15738 13695 15741
rect 15745 15738 15811 15741
rect 13629 15736 15811 15738
rect 13629 15680 13634 15736
rect 13690 15680 15750 15736
rect 15806 15680 15811 15736
rect 13629 15678 15811 15680
rect 13629 15675 13695 15678
rect 15745 15675 15811 15678
rect 23473 15738 23539 15741
rect 23790 15738 23796 15740
rect 23473 15736 23796 15738
rect 23473 15680 23478 15736
rect 23534 15680 23796 15736
rect 23473 15678 23796 15680
rect 23473 15675 23539 15678
rect 23790 15676 23796 15678
rect 23860 15676 23866 15740
rect 8385 15602 8451 15605
rect 11513 15602 11579 15605
rect 8385 15600 11579 15602
rect 8385 15544 8390 15600
rect 8446 15544 11518 15600
rect 11574 15544 11579 15600
rect 8385 15542 11579 15544
rect 8385 15539 8451 15542
rect 11513 15539 11579 15542
rect 21081 15602 21147 15605
rect 23657 15602 23723 15605
rect 21081 15600 23723 15602
rect 21081 15544 21086 15600
rect 21142 15544 23662 15600
rect 23718 15544 23723 15600
rect 21081 15542 23723 15544
rect 21081 15539 21147 15542
rect 23657 15539 23723 15542
rect 3601 15466 3667 15469
rect 16941 15466 17007 15469
rect 27520 15466 28000 15496
rect 3601 15464 28000 15466
rect 3601 15408 3606 15464
rect 3662 15408 16946 15464
rect 17002 15408 28000 15464
rect 3601 15406 28000 15408
rect 3601 15403 3667 15406
rect 16941 15403 17007 15406
rect 27520 15376 28000 15406
rect 0 15330 480 15360
rect 2221 15330 2287 15333
rect 0 15328 2287 15330
rect 0 15272 2226 15328
rect 2282 15272 2287 15328
rect 0 15270 2287 15272
rect 0 15240 480 15270
rect 2221 15267 2287 15270
rect 8109 15330 8175 15333
rect 9857 15330 9923 15333
rect 8109 15328 9923 15330
rect 8109 15272 8114 15328
rect 8170 15272 9862 15328
rect 9918 15272 9923 15328
rect 8109 15270 9923 15272
rect 8109 15267 8175 15270
rect 9857 15267 9923 15270
rect 10777 15330 10843 15333
rect 12249 15330 12315 15333
rect 10777 15328 12315 15330
rect 10777 15272 10782 15328
rect 10838 15272 12254 15328
rect 12310 15272 12315 15328
rect 10777 15270 12315 15272
rect 10777 15267 10843 15270
rect 12249 15267 12315 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 7465 15194 7531 15197
rect 10133 15194 10199 15197
rect 23381 15194 23447 15197
rect 7465 15192 10199 15194
rect 7465 15136 7470 15192
rect 7526 15136 10138 15192
rect 10194 15136 10199 15192
rect 7465 15134 10199 15136
rect 7465 15131 7531 15134
rect 10133 15131 10199 15134
rect 15380 15192 23447 15194
rect 15380 15136 23386 15192
rect 23442 15136 23447 15192
rect 15380 15134 23447 15136
rect 3509 15058 3575 15061
rect 7281 15058 7347 15061
rect 3509 15056 7347 15058
rect 3509 15000 3514 15056
rect 3570 15000 7286 15056
rect 7342 15000 7347 15056
rect 3509 14998 7347 15000
rect 3509 14995 3575 14998
rect 7281 14995 7347 14998
rect 8753 15058 8819 15061
rect 11145 15058 11211 15061
rect 8753 15056 11211 15058
rect 8753 15000 8758 15056
rect 8814 15000 11150 15056
rect 11206 15000 11211 15056
rect 8753 14998 11211 15000
rect 8753 14995 8819 14998
rect 11145 14995 11211 14998
rect 11329 15058 11395 15061
rect 13353 15058 13419 15061
rect 11329 15056 13419 15058
rect 11329 15000 11334 15056
rect 11390 15000 13358 15056
rect 13414 15000 13419 15056
rect 11329 14998 13419 15000
rect 11329 14995 11395 14998
rect 13353 14995 13419 14998
rect 13905 15058 13971 15061
rect 15380 15058 15440 15134
rect 23381 15131 23447 15134
rect 13905 15056 15440 15058
rect 13905 15000 13910 15056
rect 13966 15000 15440 15056
rect 13905 14998 15440 15000
rect 21817 15058 21883 15061
rect 24025 15058 24091 15061
rect 21817 15056 24091 15058
rect 21817 15000 21822 15056
rect 21878 15000 24030 15056
rect 24086 15000 24091 15056
rect 21817 14998 24091 15000
rect 13905 14995 13971 14998
rect 21817 14995 21883 14998
rect 24025 14995 24091 14998
rect 8293 14922 8359 14925
rect 12893 14922 12959 14925
rect 13537 14922 13603 14925
rect 7422 14920 13603 14922
rect 7422 14864 8298 14920
rect 8354 14864 12898 14920
rect 12954 14864 13542 14920
rect 13598 14864 13603 14920
rect 7422 14862 13603 14864
rect 7422 14789 7482 14862
rect 8293 14859 8359 14862
rect 12893 14859 12959 14862
rect 13537 14859 13603 14862
rect 14549 14922 14615 14925
rect 27520 14922 28000 14952
rect 14549 14920 28000 14922
rect 14549 14864 14554 14920
rect 14610 14864 28000 14920
rect 14549 14862 28000 14864
rect 14549 14859 14615 14862
rect 27520 14832 28000 14862
rect 3233 14786 3299 14789
rect 4337 14786 4403 14789
rect 3233 14784 4403 14786
rect 3233 14728 3238 14784
rect 3294 14728 4342 14784
rect 4398 14728 4403 14784
rect 3233 14726 4403 14728
rect 3233 14723 3299 14726
rect 4337 14723 4403 14726
rect 7373 14784 7482 14789
rect 7373 14728 7378 14784
rect 7434 14728 7482 14784
rect 7373 14726 7482 14728
rect 10961 14786 11027 14789
rect 18229 14786 18295 14789
rect 10961 14784 18295 14786
rect 10961 14728 10966 14784
rect 11022 14728 18234 14784
rect 18290 14728 18295 14784
rect 10961 14726 18295 14728
rect 7373 14723 7439 14726
rect 10961 14723 11027 14726
rect 18229 14723 18295 14726
rect 10277 14720 10597 14721
rect 0 14650 480 14680
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 3693 14650 3759 14653
rect 0 14648 3759 14650
rect 0 14592 3698 14648
rect 3754 14592 3759 14648
rect 0 14590 3759 14592
rect 0 14560 480 14590
rect 3693 14587 3759 14590
rect 6545 14650 6611 14653
rect 8385 14650 8451 14653
rect 6545 14648 8451 14650
rect 6545 14592 6550 14648
rect 6606 14592 8390 14648
rect 8446 14592 8451 14648
rect 6545 14590 8451 14592
rect 6545 14587 6611 14590
rect 8385 14587 8451 14590
rect 13445 14650 13511 14653
rect 17769 14650 17835 14653
rect 13445 14648 17835 14650
rect 13445 14592 13450 14648
rect 13506 14592 17774 14648
rect 17830 14592 17835 14648
rect 13445 14590 17835 14592
rect 13445 14587 13511 14590
rect 17769 14587 17835 14590
rect 8937 14514 9003 14517
rect 13445 14514 13511 14517
rect 8937 14512 13511 14514
rect 8937 14456 8942 14512
rect 8998 14456 13450 14512
rect 13506 14456 13511 14512
rect 8937 14454 13511 14456
rect 8937 14451 9003 14454
rect 13445 14451 13511 14454
rect 2497 14378 2563 14381
rect 8569 14378 8635 14381
rect 2497 14376 8635 14378
rect 2497 14320 2502 14376
rect 2558 14320 8574 14376
rect 8630 14320 8635 14376
rect 2497 14318 8635 14320
rect 2497 14315 2563 14318
rect 8569 14315 8635 14318
rect 15101 14378 15167 14381
rect 16757 14378 16823 14381
rect 15101 14376 16823 14378
rect 15101 14320 15106 14376
rect 15162 14320 16762 14376
rect 16818 14320 16823 14376
rect 15101 14318 16823 14320
rect 15101 14315 15167 14318
rect 16757 14315 16823 14318
rect 17033 14378 17099 14381
rect 27520 14378 28000 14408
rect 17033 14376 28000 14378
rect 17033 14320 17038 14376
rect 17094 14320 28000 14376
rect 17033 14318 28000 14320
rect 17033 14315 17099 14318
rect 27520 14288 28000 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 8201 14106 8267 14109
rect 10225 14106 10291 14109
rect 8201 14104 10291 14106
rect 8201 14048 8206 14104
rect 8262 14048 10230 14104
rect 10286 14048 10291 14104
rect 8201 14046 10291 14048
rect 8201 14043 8267 14046
rect 10225 14043 10291 14046
rect 0 13970 480 14000
rect 1761 13970 1827 13973
rect 0 13968 1827 13970
rect 0 13912 1766 13968
rect 1822 13912 1827 13968
rect 0 13910 1827 13912
rect 0 13880 480 13910
rect 1761 13907 1827 13910
rect 16021 13970 16087 13973
rect 18689 13970 18755 13973
rect 22277 13970 22343 13973
rect 27520 13970 28000 14000
rect 16021 13968 22343 13970
rect 16021 13912 16026 13968
rect 16082 13912 18694 13968
rect 18750 13912 22282 13968
rect 22338 13912 22343 13968
rect 16021 13910 22343 13912
rect 16021 13907 16087 13910
rect 18689 13907 18755 13910
rect 22277 13907 22343 13910
rect 24350 13910 28000 13970
rect 5625 13834 5691 13837
rect 14273 13834 14339 13837
rect 5625 13832 14339 13834
rect 5625 13776 5630 13832
rect 5686 13776 14278 13832
rect 14334 13776 14339 13832
rect 5625 13774 14339 13776
rect 5625 13771 5691 13774
rect 14273 13771 14339 13774
rect 24209 13834 24275 13837
rect 24350 13834 24410 13910
rect 27520 13880 28000 13910
rect 24209 13832 24410 13834
rect 24209 13776 24214 13832
rect 24270 13776 24410 13832
rect 24209 13774 24410 13776
rect 24209 13771 24275 13774
rect 3969 13698 4035 13701
rect 5625 13698 5691 13701
rect 8385 13698 8451 13701
rect 3969 13696 8451 13698
rect 3969 13640 3974 13696
rect 4030 13640 5630 13696
rect 5686 13640 8390 13696
rect 8446 13640 8451 13696
rect 3969 13638 8451 13640
rect 3969 13635 4035 13638
rect 5625 13635 5691 13638
rect 8385 13635 8451 13638
rect 10777 13698 10843 13701
rect 17033 13698 17099 13701
rect 10777 13696 17099 13698
rect 10777 13640 10782 13696
rect 10838 13640 17038 13696
rect 17094 13640 17099 13696
rect 10777 13638 17099 13640
rect 10777 13635 10843 13638
rect 17033 13635 17099 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 5809 13562 5875 13565
rect 9029 13562 9095 13565
rect 5809 13560 9095 13562
rect 5809 13504 5814 13560
rect 5870 13504 9034 13560
rect 9090 13504 9095 13560
rect 5809 13502 9095 13504
rect 5809 13499 5875 13502
rect 9029 13499 9095 13502
rect 11789 13562 11855 13565
rect 15469 13562 15535 13565
rect 11789 13560 15535 13562
rect 11789 13504 11794 13560
rect 11850 13504 15474 13560
rect 15530 13504 15535 13560
rect 11789 13502 15535 13504
rect 11789 13499 11855 13502
rect 15469 13499 15535 13502
rect 17585 13562 17651 13565
rect 19425 13562 19491 13565
rect 23013 13562 23079 13565
rect 17585 13560 19491 13562
rect 17585 13504 17590 13560
rect 17646 13504 19430 13560
rect 19486 13504 19491 13560
rect 17585 13502 19491 13504
rect 17585 13499 17651 13502
rect 19425 13499 19491 13502
rect 20118 13560 23079 13562
rect 20118 13504 23018 13560
rect 23074 13504 23079 13560
rect 20118 13502 23079 13504
rect 2957 13426 3023 13429
rect 12709 13426 12775 13429
rect 2957 13424 12775 13426
rect 2957 13368 2962 13424
rect 3018 13368 12714 13424
rect 12770 13368 12775 13424
rect 2957 13366 12775 13368
rect 2957 13363 3023 13366
rect 12709 13363 12775 13366
rect 15561 13426 15627 13429
rect 20118 13426 20178 13502
rect 23013 13499 23079 13502
rect 15561 13424 20178 13426
rect 15561 13368 15566 13424
rect 15622 13368 20178 13424
rect 15561 13366 20178 13368
rect 20253 13426 20319 13429
rect 27520 13426 28000 13456
rect 20253 13424 28000 13426
rect 20253 13368 20258 13424
rect 20314 13368 28000 13424
rect 20253 13366 28000 13368
rect 15561 13363 15627 13366
rect 20253 13363 20319 13366
rect 27520 13336 28000 13366
rect 0 13290 480 13320
rect 3785 13290 3851 13293
rect 0 13288 3851 13290
rect 0 13232 3790 13288
rect 3846 13232 3851 13288
rect 0 13230 3851 13232
rect 0 13200 480 13230
rect 3785 13227 3851 13230
rect 4705 13290 4771 13293
rect 8569 13290 8635 13293
rect 24669 13290 24735 13293
rect 4705 13288 6562 13290
rect 4705 13232 4710 13288
rect 4766 13232 6562 13288
rect 4705 13230 6562 13232
rect 4705 13227 4771 13230
rect 6502 13154 6562 13230
rect 8569 13288 24735 13290
rect 8569 13232 8574 13288
rect 8630 13232 24674 13288
rect 24730 13232 24735 13288
rect 8569 13230 24735 13232
rect 8569 13227 8635 13230
rect 24669 13227 24735 13230
rect 10777 13154 10843 13157
rect 6502 13152 10843 13154
rect 6502 13096 10782 13152
rect 10838 13096 10843 13152
rect 6502 13094 10843 13096
rect 10777 13091 10843 13094
rect 17769 13154 17835 13157
rect 20253 13154 20319 13157
rect 17769 13152 20319 13154
rect 17769 13096 17774 13152
rect 17830 13096 20258 13152
rect 20314 13096 20319 13152
rect 17769 13094 20319 13096
rect 17769 13091 17835 13094
rect 20253 13091 20319 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 15469 13018 15535 13021
rect 19333 13018 19399 13021
rect 15469 13016 19399 13018
rect 15469 12960 15474 13016
rect 15530 12960 19338 13016
rect 19394 12960 19399 13016
rect 15469 12958 19399 12960
rect 15469 12955 15535 12958
rect 19333 12955 19399 12958
rect 19517 13018 19583 13021
rect 22185 13018 22251 13021
rect 19517 13016 22251 13018
rect 19517 12960 19522 13016
rect 19578 12960 22190 13016
rect 22246 12960 22251 13016
rect 19517 12958 22251 12960
rect 19517 12955 19583 12958
rect 22185 12955 22251 12958
rect 3693 12882 3759 12885
rect 8017 12882 8083 12885
rect 3693 12880 8083 12882
rect 3693 12824 3698 12880
rect 3754 12824 8022 12880
rect 8078 12824 8083 12880
rect 3693 12822 8083 12824
rect 3693 12819 3759 12822
rect 8017 12819 8083 12822
rect 13997 12882 14063 12885
rect 24209 12882 24275 12885
rect 27520 12882 28000 12912
rect 13997 12880 24275 12882
rect 13997 12824 14002 12880
rect 14058 12824 24214 12880
rect 24270 12824 24275 12880
rect 13997 12822 24275 12824
rect 13997 12819 14063 12822
rect 24209 12819 24275 12822
rect 24856 12822 28000 12882
rect 0 12746 480 12776
rect 2497 12746 2563 12749
rect 0 12744 2563 12746
rect 0 12688 2502 12744
rect 2558 12688 2563 12744
rect 0 12686 2563 12688
rect 0 12656 480 12686
rect 2497 12683 2563 12686
rect 5165 12746 5231 12749
rect 9305 12746 9371 12749
rect 5165 12744 9371 12746
rect 5165 12688 5170 12744
rect 5226 12688 9310 12744
rect 9366 12688 9371 12744
rect 5165 12686 9371 12688
rect 5165 12683 5231 12686
rect 9305 12683 9371 12686
rect 9765 12746 9831 12749
rect 24856 12746 24916 12822
rect 27520 12792 28000 12822
rect 9765 12744 24916 12746
rect 9765 12688 9770 12744
rect 9826 12688 24916 12744
rect 9765 12686 24916 12688
rect 9765 12683 9831 12686
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 10869 12474 10935 12477
rect 12617 12474 12683 12477
rect 13261 12474 13327 12477
rect 17769 12474 17835 12477
rect 24761 12476 24827 12477
rect 24710 12474 24716 12476
rect 10869 12472 13327 12474
rect 10869 12416 10874 12472
rect 10930 12416 12622 12472
rect 12678 12416 13266 12472
rect 13322 12416 13327 12472
rect 10869 12414 13327 12416
rect 10869 12411 10935 12414
rect 12617 12411 12683 12414
rect 13261 12411 13327 12414
rect 13494 12472 17835 12474
rect 13494 12416 17774 12472
rect 17830 12416 17835 12472
rect 13494 12414 17835 12416
rect 24670 12414 24716 12474
rect 24780 12472 24827 12476
rect 24822 12416 24827 12472
rect 5533 12338 5599 12341
rect 11605 12338 11671 12341
rect 5533 12336 11671 12338
rect 5533 12280 5538 12336
rect 5594 12280 11610 12336
rect 11666 12280 11671 12336
rect 5533 12278 11671 12280
rect 5533 12275 5599 12278
rect 11605 12275 11671 12278
rect 12065 12338 12131 12341
rect 13494 12338 13554 12414
rect 17769 12411 17835 12414
rect 24710 12412 24716 12414
rect 24780 12412 24827 12416
rect 24761 12411 24827 12412
rect 12065 12336 13554 12338
rect 12065 12280 12070 12336
rect 12126 12280 13554 12336
rect 12065 12278 13554 12280
rect 16113 12338 16179 12341
rect 20805 12338 20871 12341
rect 16113 12336 20871 12338
rect 16113 12280 16118 12336
rect 16174 12280 20810 12336
rect 20866 12280 20871 12336
rect 16113 12278 20871 12280
rect 12065 12275 12131 12278
rect 16113 12275 16179 12278
rect 20805 12275 20871 12278
rect 20989 12338 21055 12341
rect 27520 12338 28000 12368
rect 20989 12336 28000 12338
rect 20989 12280 20994 12336
rect 21050 12280 28000 12336
rect 20989 12278 28000 12280
rect 20989 12275 21055 12278
rect 27520 12248 28000 12278
rect 3325 12202 3391 12205
rect 5993 12202 6059 12205
rect 3325 12200 6059 12202
rect 3325 12144 3330 12200
rect 3386 12144 5998 12200
rect 6054 12144 6059 12200
rect 3325 12142 6059 12144
rect 3325 12139 3391 12142
rect 5993 12139 6059 12142
rect 8385 12202 8451 12205
rect 10961 12202 11027 12205
rect 8385 12200 11027 12202
rect 8385 12144 8390 12200
rect 8446 12144 10966 12200
rect 11022 12144 11027 12200
rect 8385 12142 11027 12144
rect 8385 12139 8451 12142
rect 10961 12139 11027 12142
rect 21173 12202 21239 12205
rect 24853 12202 24919 12205
rect 21173 12200 24919 12202
rect 21173 12144 21178 12200
rect 21234 12144 24858 12200
rect 24914 12144 24919 12200
rect 21173 12142 24919 12144
rect 21173 12139 21239 12142
rect 24853 12139 24919 12142
rect 0 12066 480 12096
rect 3969 12066 4035 12069
rect 0 12064 4035 12066
rect 0 12008 3974 12064
rect 4030 12008 4035 12064
rect 0 12006 4035 12008
rect 0 11976 480 12006
rect 3969 12003 4035 12006
rect 6729 12066 6795 12069
rect 9673 12066 9739 12069
rect 6729 12064 9739 12066
rect 6729 12008 6734 12064
rect 6790 12008 9678 12064
rect 9734 12008 9739 12064
rect 6729 12006 9739 12008
rect 6729 12003 6795 12006
rect 9673 12003 9739 12006
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 7189 11930 7255 11933
rect 11789 11930 11855 11933
rect 7189 11928 11855 11930
rect 7189 11872 7194 11928
rect 7250 11872 11794 11928
rect 11850 11872 11855 11928
rect 7189 11870 11855 11872
rect 7189 11867 7255 11870
rect 11789 11867 11855 11870
rect 4245 11794 4311 11797
rect 27520 11794 28000 11824
rect 4245 11792 28000 11794
rect 4245 11736 4250 11792
rect 4306 11736 28000 11792
rect 4245 11734 28000 11736
rect 4245 11731 4311 11734
rect 27520 11704 28000 11734
rect 2865 11658 2931 11661
rect 10685 11658 10751 11661
rect 2865 11656 10751 11658
rect 2865 11600 2870 11656
rect 2926 11600 10690 11656
rect 10746 11600 10751 11656
rect 2865 11598 10751 11600
rect 2865 11595 2931 11598
rect 10685 11595 10751 11598
rect 15745 11658 15811 11661
rect 19425 11658 19491 11661
rect 15745 11656 19491 11658
rect 15745 11600 15750 11656
rect 15806 11600 19430 11656
rect 19486 11600 19491 11656
rect 15745 11598 19491 11600
rect 15745 11595 15811 11598
rect 19425 11595 19491 11598
rect 21633 11658 21699 11661
rect 25037 11658 25103 11661
rect 21633 11656 25103 11658
rect 21633 11600 21638 11656
rect 21694 11600 25042 11656
rect 25098 11600 25103 11656
rect 21633 11598 25103 11600
rect 21633 11595 21699 11598
rect 25037 11595 25103 11598
rect 1393 11522 1459 11525
rect 4429 11522 4495 11525
rect 1393 11520 4495 11522
rect 1393 11464 1398 11520
rect 1454 11464 4434 11520
rect 4490 11464 4495 11520
rect 1393 11462 4495 11464
rect 1393 11459 1459 11462
rect 4429 11459 4495 11462
rect 5349 11522 5415 11525
rect 7097 11522 7163 11525
rect 5349 11520 7163 11522
rect 5349 11464 5354 11520
rect 5410 11464 7102 11520
rect 7158 11464 7163 11520
rect 5349 11462 7163 11464
rect 5349 11459 5415 11462
rect 7097 11459 7163 11462
rect 13261 11522 13327 11525
rect 18597 11522 18663 11525
rect 13261 11520 18663 11522
rect 13261 11464 13266 11520
rect 13322 11464 18602 11520
rect 18658 11464 18663 11520
rect 13261 11462 18663 11464
rect 13261 11459 13327 11462
rect 18597 11459 18663 11462
rect 10277 11456 10597 11457
rect 0 11386 480 11416
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 3785 11386 3851 11389
rect 0 11384 3851 11386
rect 0 11328 3790 11384
rect 3846 11328 3851 11384
rect 0 11326 3851 11328
rect 0 11296 480 11326
rect 3785 11323 3851 11326
rect 13169 11386 13235 11389
rect 18781 11386 18847 11389
rect 13169 11384 18847 11386
rect 13169 11328 13174 11384
rect 13230 11328 18786 11384
rect 18842 11328 18847 11384
rect 13169 11326 18847 11328
rect 13169 11323 13235 11326
rect 18781 11323 18847 11326
rect 1393 11250 1459 11253
rect 3509 11250 3575 11253
rect 1393 11248 3575 11250
rect 1393 11192 1398 11248
rect 1454 11192 3514 11248
rect 3570 11192 3575 11248
rect 1393 11190 3575 11192
rect 1393 11187 1459 11190
rect 3509 11187 3575 11190
rect 11513 11250 11579 11253
rect 27520 11250 28000 11280
rect 11513 11248 28000 11250
rect 11513 11192 11518 11248
rect 11574 11192 28000 11248
rect 11513 11190 28000 11192
rect 11513 11187 11579 11190
rect 27520 11160 28000 11190
rect 10225 11114 10291 11117
rect 14365 11114 14431 11117
rect 10225 11112 14431 11114
rect 10225 11056 10230 11112
rect 10286 11056 14370 11112
rect 14426 11056 14431 11112
rect 10225 11054 14431 11056
rect 10225 11051 10291 11054
rect 14365 11051 14431 11054
rect 23197 11114 23263 11117
rect 23473 11114 23539 11117
rect 23197 11112 23539 11114
rect 23197 11056 23202 11112
rect 23258 11056 23478 11112
rect 23534 11056 23539 11112
rect 23197 11054 23539 11056
rect 23197 11051 23263 11054
rect 23473 11051 23539 11054
rect 7005 10978 7071 10981
rect 9673 10978 9739 10981
rect 7005 10976 9739 10978
rect 7005 10920 7010 10976
rect 7066 10920 9678 10976
rect 9734 10920 9739 10976
rect 7005 10918 9739 10920
rect 7005 10915 7071 10918
rect 9673 10915 9739 10918
rect 15745 10978 15811 10981
rect 20989 10978 21055 10981
rect 15745 10976 21055 10978
rect 15745 10920 15750 10976
rect 15806 10920 20994 10976
rect 21050 10920 21055 10976
rect 15745 10918 21055 10920
rect 15745 10915 15811 10918
rect 20989 10915 21055 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 7649 10842 7715 10845
rect 11881 10842 11947 10845
rect 7649 10840 11947 10842
rect 7649 10784 7654 10840
rect 7710 10784 11886 10840
rect 11942 10784 11947 10840
rect 7649 10782 11947 10784
rect 7649 10779 7715 10782
rect 11881 10779 11947 10782
rect 15929 10842 15995 10845
rect 19609 10842 19675 10845
rect 15929 10840 19675 10842
rect 15929 10784 15934 10840
rect 15990 10784 19614 10840
rect 19670 10784 19675 10840
rect 15929 10782 19675 10784
rect 15929 10779 15995 10782
rect 19609 10779 19675 10782
rect 0 10706 480 10736
rect 2681 10706 2747 10709
rect 0 10704 2747 10706
rect 0 10648 2686 10704
rect 2742 10648 2747 10704
rect 0 10646 2747 10648
rect 0 10616 480 10646
rect 2681 10643 2747 10646
rect 25129 10706 25195 10709
rect 27520 10706 28000 10736
rect 25129 10704 28000 10706
rect 25129 10648 25134 10704
rect 25190 10648 28000 10704
rect 25129 10646 28000 10648
rect 25129 10643 25195 10646
rect 27520 10616 28000 10646
rect 9949 10570 10015 10573
rect 15837 10570 15903 10573
rect 9949 10568 15903 10570
rect 9949 10512 9954 10568
rect 10010 10512 15842 10568
rect 15898 10512 15903 10568
rect 9949 10510 15903 10512
rect 9949 10507 10015 10510
rect 15837 10507 15903 10510
rect 4521 10434 4587 10437
rect 7649 10434 7715 10437
rect 4521 10432 7715 10434
rect 4521 10376 4526 10432
rect 4582 10376 7654 10432
rect 7710 10376 7715 10432
rect 4521 10374 7715 10376
rect 4521 10371 4587 10374
rect 7649 10371 7715 10374
rect 12157 10434 12223 10437
rect 13077 10434 13143 10437
rect 12157 10432 13143 10434
rect 12157 10376 12162 10432
rect 12218 10376 13082 10432
rect 13138 10376 13143 10432
rect 12157 10374 13143 10376
rect 12157 10371 12223 10374
rect 13077 10371 13143 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 2037 10298 2103 10301
rect 11237 10298 11303 10301
rect 14181 10298 14247 10301
rect 2037 10296 7666 10298
rect 2037 10240 2042 10296
rect 2098 10240 7666 10296
rect 2037 10238 7666 10240
rect 2037 10235 2103 10238
rect 1393 10162 1459 10165
rect 7606 10162 7666 10238
rect 11237 10296 14247 10298
rect 11237 10240 11242 10296
rect 11298 10240 14186 10296
rect 14242 10240 14247 10296
rect 11237 10238 14247 10240
rect 11237 10235 11303 10238
rect 14181 10235 14247 10238
rect 14641 10298 14707 10301
rect 18781 10298 18847 10301
rect 23841 10300 23907 10301
rect 14641 10296 18847 10298
rect 14641 10240 14646 10296
rect 14702 10240 18786 10296
rect 18842 10240 18847 10296
rect 14641 10238 18847 10240
rect 14641 10235 14707 10238
rect 18781 10235 18847 10238
rect 23790 10236 23796 10300
rect 23860 10298 23907 10300
rect 23860 10296 23952 10298
rect 23902 10240 23952 10296
rect 23860 10238 23952 10240
rect 23860 10236 23907 10238
rect 23841 10235 23907 10236
rect 15745 10162 15811 10165
rect 1393 10160 7482 10162
rect 1393 10104 1398 10160
rect 1454 10104 7482 10160
rect 1393 10102 7482 10104
rect 7606 10160 15811 10162
rect 7606 10104 15750 10160
rect 15806 10104 15811 10160
rect 7606 10102 15811 10104
rect 1393 10099 1459 10102
rect 0 10026 480 10056
rect 2681 10026 2747 10029
rect 0 10024 2747 10026
rect 0 9968 2686 10024
rect 2742 9968 2747 10024
rect 0 9966 2747 9968
rect 0 9936 480 9966
rect 2681 9963 2747 9966
rect 2865 10026 2931 10029
rect 6913 10026 6979 10029
rect 2865 10024 6979 10026
rect 2865 9968 2870 10024
rect 2926 9968 6918 10024
rect 6974 9968 6979 10024
rect 2865 9966 6979 9968
rect 2865 9963 2931 9966
rect 6913 9963 6979 9966
rect 7422 9890 7482 10102
rect 15745 10099 15811 10102
rect 18965 10162 19031 10165
rect 24945 10162 25011 10165
rect 18965 10160 25011 10162
rect 18965 10104 18970 10160
rect 19026 10104 24950 10160
rect 25006 10104 25011 10160
rect 18965 10102 25011 10104
rect 18965 10099 19031 10102
rect 24945 10099 25011 10102
rect 25497 10162 25563 10165
rect 27520 10162 28000 10192
rect 25497 10160 28000 10162
rect 25497 10104 25502 10160
rect 25558 10104 28000 10160
rect 25497 10102 28000 10104
rect 25497 10099 25563 10102
rect 27520 10072 28000 10102
rect 7557 10026 7623 10029
rect 11237 10026 11303 10029
rect 7557 10024 11303 10026
rect 7557 9968 7562 10024
rect 7618 9968 11242 10024
rect 11298 9968 11303 10024
rect 7557 9966 11303 9968
rect 7557 9963 7623 9966
rect 11237 9963 11303 9966
rect 14181 10026 14247 10029
rect 22645 10026 22711 10029
rect 24669 10028 24735 10029
rect 24669 10026 24716 10028
rect 14181 10024 22711 10026
rect 14181 9968 14186 10024
rect 14242 9968 22650 10024
rect 22706 9968 22711 10024
rect 14181 9966 22711 9968
rect 24624 10024 24716 10026
rect 24624 9968 24674 10024
rect 24624 9966 24716 9968
rect 14181 9963 14247 9966
rect 22645 9963 22711 9966
rect 24669 9964 24716 9966
rect 24780 9964 24786 10028
rect 24669 9963 24735 9964
rect 10593 9890 10659 9893
rect 7422 9888 10659 9890
rect 7422 9832 10598 9888
rect 10654 9832 10659 9888
rect 7422 9830 10659 9832
rect 10593 9827 10659 9830
rect 20253 9890 20319 9893
rect 24025 9890 24091 9893
rect 20253 9888 24091 9890
rect 20253 9832 20258 9888
rect 20314 9832 24030 9888
rect 24086 9832 24091 9888
rect 20253 9830 24091 9832
rect 20253 9827 20319 9830
rect 24025 9827 24091 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 6453 9754 6519 9757
rect 9213 9754 9279 9757
rect 12157 9754 12223 9757
rect 6453 9752 9279 9754
rect 6453 9696 6458 9752
rect 6514 9696 9218 9752
rect 9274 9696 9279 9752
rect 6453 9694 9279 9696
rect 6453 9691 6519 9694
rect 9213 9691 9279 9694
rect 9446 9752 12223 9754
rect 9446 9696 12162 9752
rect 12218 9696 12223 9752
rect 9446 9694 12223 9696
rect 4705 9652 4771 9655
rect 4705 9650 4906 9652
rect 4705 9594 4710 9650
rect 4766 9621 4906 9650
rect 4766 9616 4955 9621
rect 4766 9594 4894 9616
rect 4705 9592 4894 9594
rect 4705 9589 4771 9592
rect 4846 9560 4894 9592
rect 4950 9560 4955 9616
rect 4846 9558 4955 9560
rect 4889 9555 4955 9558
rect 8201 9618 8267 9621
rect 9446 9618 9506 9694
rect 12157 9691 12223 9694
rect 15377 9754 15443 9757
rect 19149 9754 19215 9757
rect 15377 9752 19215 9754
rect 15377 9696 15382 9752
rect 15438 9696 19154 9752
rect 19210 9696 19215 9752
rect 15377 9694 19215 9696
rect 15377 9691 15443 9694
rect 19149 9691 19215 9694
rect 21909 9754 21975 9757
rect 23657 9754 23723 9757
rect 21909 9752 23723 9754
rect 21909 9696 21914 9752
rect 21970 9696 23662 9752
rect 23718 9696 23723 9752
rect 21909 9694 23723 9696
rect 21909 9691 21975 9694
rect 23657 9691 23723 9694
rect 8201 9616 9506 9618
rect 8201 9560 8206 9616
rect 8262 9560 9506 9616
rect 8201 9558 9506 9560
rect 11605 9618 11671 9621
rect 13813 9618 13879 9621
rect 11605 9616 13879 9618
rect 11605 9560 11610 9616
rect 11666 9560 13818 9616
rect 13874 9560 13879 9616
rect 11605 9558 13879 9560
rect 8201 9555 8267 9558
rect 11605 9555 11671 9558
rect 13813 9555 13879 9558
rect 19885 9618 19951 9621
rect 22369 9618 22435 9621
rect 19885 9616 22435 9618
rect 19885 9560 19890 9616
rect 19946 9560 22374 9616
rect 22430 9560 22435 9616
rect 19885 9558 22435 9560
rect 19885 9555 19951 9558
rect 22369 9555 22435 9558
rect 24945 9618 25011 9621
rect 27520 9618 28000 9648
rect 24945 9616 28000 9618
rect 24945 9560 24950 9616
rect 25006 9560 28000 9616
rect 24945 9558 28000 9560
rect 24945 9555 25011 9558
rect 27520 9528 28000 9558
rect 0 9482 480 9512
rect 1577 9482 1643 9485
rect 0 9480 1643 9482
rect 0 9424 1582 9480
rect 1638 9424 1643 9480
rect 0 9422 1643 9424
rect 0 9392 480 9422
rect 1577 9419 1643 9422
rect 2865 9482 2931 9485
rect 14089 9482 14155 9485
rect 2865 9480 14155 9482
rect 2865 9424 2870 9480
rect 2926 9424 14094 9480
rect 14150 9424 14155 9480
rect 2865 9422 14155 9424
rect 2865 9419 2931 9422
rect 14089 9419 14155 9422
rect 21541 9482 21607 9485
rect 23841 9482 23907 9485
rect 21541 9480 23907 9482
rect 21541 9424 21546 9480
rect 21602 9424 23846 9480
rect 23902 9424 23907 9480
rect 21541 9422 23907 9424
rect 21541 9419 21607 9422
rect 23841 9419 23907 9422
rect 20345 9346 20411 9349
rect 24761 9346 24827 9349
rect 20345 9344 24827 9346
rect 20345 9288 20350 9344
rect 20406 9288 24766 9344
rect 24822 9288 24827 9344
rect 20345 9286 24827 9288
rect 20345 9283 20411 9286
rect 24761 9283 24827 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 20161 9210 20227 9213
rect 23565 9210 23631 9213
rect 20161 9208 23631 9210
rect 20161 9152 20166 9208
rect 20222 9152 23570 9208
rect 23626 9152 23631 9208
rect 20161 9150 23631 9152
rect 20161 9147 20227 9150
rect 23565 9147 23631 9150
rect 25129 9210 25195 9213
rect 27520 9210 28000 9240
rect 25129 9208 28000 9210
rect 25129 9152 25134 9208
rect 25190 9152 28000 9208
rect 25129 9150 28000 9152
rect 25129 9147 25195 9150
rect 27520 9120 28000 9150
rect 9857 9074 9923 9077
rect 7606 9072 9923 9074
rect 7606 9016 9862 9072
rect 9918 9016 9923 9072
rect 7606 9014 9923 9016
rect 2037 8938 2103 8941
rect 7606 8938 7666 9014
rect 9857 9011 9923 9014
rect 12249 9074 12315 9077
rect 21357 9074 21423 9077
rect 12249 9072 21423 9074
rect 12249 9016 12254 9072
rect 12310 9016 21362 9072
rect 21418 9016 21423 9072
rect 12249 9014 21423 9016
rect 12249 9011 12315 9014
rect 21357 9011 21423 9014
rect 2037 8936 7666 8938
rect 2037 8880 2042 8936
rect 2098 8880 7666 8936
rect 2037 8878 7666 8880
rect 7741 8938 7807 8941
rect 12249 8938 12315 8941
rect 7741 8936 12315 8938
rect 7741 8880 7746 8936
rect 7802 8880 12254 8936
rect 12310 8880 12315 8936
rect 7741 8878 12315 8880
rect 2037 8875 2103 8878
rect 7741 8875 7807 8878
rect 12249 8875 12315 8878
rect 0 8802 480 8832
rect 1577 8802 1643 8805
rect 0 8800 1643 8802
rect 0 8744 1582 8800
rect 1638 8744 1643 8800
rect 0 8742 1643 8744
rect 0 8712 480 8742
rect 1577 8739 1643 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 24761 8666 24827 8669
rect 27520 8666 28000 8696
rect 24761 8664 28000 8666
rect 24761 8608 24766 8664
rect 24822 8608 28000 8664
rect 24761 8606 28000 8608
rect 24761 8603 24827 8606
rect 27520 8576 28000 8606
rect 3233 8530 3299 8533
rect 13629 8530 13695 8533
rect 3233 8528 13695 8530
rect 3233 8472 3238 8528
rect 3294 8472 13634 8528
rect 13690 8472 13695 8528
rect 3233 8470 13695 8472
rect 3233 8467 3299 8470
rect 13629 8467 13695 8470
rect 14549 8394 14615 8397
rect 18229 8394 18295 8397
rect 14549 8392 18295 8394
rect 14549 8336 14554 8392
rect 14610 8336 18234 8392
rect 18290 8336 18295 8392
rect 14549 8334 18295 8336
rect 14549 8331 14615 8334
rect 18229 8331 18295 8334
rect 18505 8394 18571 8397
rect 24945 8394 25011 8397
rect 18505 8392 25011 8394
rect 18505 8336 18510 8392
rect 18566 8336 24950 8392
rect 25006 8336 25011 8392
rect 18505 8334 25011 8336
rect 18505 8331 18571 8334
rect 24945 8331 25011 8334
rect 10277 8192 10597 8193
rect 0 8122 480 8152
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 1577 8122 1643 8125
rect 0 8120 1643 8122
rect 0 8064 1582 8120
rect 1638 8064 1643 8120
rect 0 8062 1643 8064
rect 0 8032 480 8062
rect 1577 8059 1643 8062
rect 2037 8122 2103 8125
rect 8150 8122 8156 8124
rect 2037 8120 8156 8122
rect 2037 8064 2042 8120
rect 2098 8064 8156 8120
rect 2037 8062 8156 8064
rect 2037 8059 2103 8062
rect 8150 8060 8156 8062
rect 8220 8060 8226 8124
rect 24669 8122 24735 8125
rect 27520 8122 28000 8152
rect 24669 8120 28000 8122
rect 24669 8064 24674 8120
rect 24730 8064 28000 8120
rect 24669 8062 28000 8064
rect 24669 8059 24735 8062
rect 27520 8032 28000 8062
rect 2221 7986 2287 7989
rect 9765 7986 9831 7989
rect 2221 7984 9831 7986
rect 2221 7928 2226 7984
rect 2282 7928 9770 7984
rect 9826 7928 9831 7984
rect 2221 7926 9831 7928
rect 2221 7923 2287 7926
rect 9765 7923 9831 7926
rect 1393 7850 1459 7853
rect 7097 7850 7163 7853
rect 1393 7848 7163 7850
rect 1393 7792 1398 7848
rect 1454 7792 7102 7848
rect 7158 7792 7163 7848
rect 1393 7790 7163 7792
rect 1393 7787 1459 7790
rect 7097 7787 7163 7790
rect 8661 7850 8727 7853
rect 11789 7850 11855 7853
rect 8661 7848 11855 7850
rect 8661 7792 8666 7848
rect 8722 7792 11794 7848
rect 11850 7792 11855 7848
rect 8661 7790 11855 7792
rect 8661 7787 8727 7790
rect 11789 7787 11855 7790
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 24761 7578 24827 7581
rect 27520 7578 28000 7608
rect 24761 7576 28000 7578
rect 24761 7520 24766 7576
rect 24822 7520 28000 7576
rect 24761 7518 28000 7520
rect 24761 7515 24827 7518
rect 27520 7488 28000 7518
rect 0 7442 480 7472
rect 1577 7442 1643 7445
rect 0 7440 1643 7442
rect 0 7384 1582 7440
rect 1638 7384 1643 7440
rect 0 7382 1643 7384
rect 0 7352 480 7382
rect 1577 7379 1643 7382
rect 2313 7442 2379 7445
rect 11973 7442 12039 7445
rect 2313 7440 12039 7442
rect 2313 7384 2318 7440
rect 2374 7384 11978 7440
rect 12034 7384 12039 7440
rect 2313 7382 12039 7384
rect 2313 7379 2379 7382
rect 11973 7379 12039 7382
rect 19149 7442 19215 7445
rect 24209 7442 24275 7445
rect 19149 7440 24275 7442
rect 19149 7384 19154 7440
rect 19210 7384 24214 7440
rect 24270 7384 24275 7440
rect 19149 7382 24275 7384
rect 19149 7379 19215 7382
rect 24209 7379 24275 7382
rect 18229 7306 18295 7309
rect 18229 7304 24916 7306
rect 18229 7248 18234 7304
rect 18290 7248 24916 7304
rect 18229 7246 24916 7248
rect 18229 7243 18295 7246
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 24856 7034 24916 7246
rect 27520 7034 28000 7064
rect 24856 6974 28000 7034
rect 27520 6944 28000 6974
rect 22185 6898 22251 6901
rect 24577 6898 24643 6901
rect 22185 6896 24643 6898
rect 22185 6840 22190 6896
rect 22246 6840 24582 6896
rect 24638 6840 24643 6896
rect 22185 6838 24643 6840
rect 22185 6835 22251 6838
rect 24577 6835 24643 6838
rect 0 6762 480 6792
rect 3141 6762 3207 6765
rect 0 6760 3207 6762
rect 0 6704 3146 6760
rect 3202 6704 3207 6760
rect 0 6702 3207 6704
rect 0 6672 480 6702
rect 3141 6699 3207 6702
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 24761 6490 24827 6493
rect 27520 6490 28000 6520
rect 24761 6488 28000 6490
rect 24761 6432 24766 6488
rect 24822 6432 28000 6488
rect 24761 6430 28000 6432
rect 24761 6427 24827 6430
rect 27520 6400 28000 6430
rect 0 6218 480 6248
rect 4245 6218 4311 6221
rect 0 6216 4311 6218
rect 0 6160 4250 6216
rect 4306 6160 4311 6216
rect 0 6158 4311 6160
rect 0 6128 480 6158
rect 4245 6155 4311 6158
rect 21357 6082 21423 6085
rect 24853 6082 24919 6085
rect 21357 6080 24919 6082
rect 21357 6024 21362 6080
rect 21418 6024 24858 6080
rect 24914 6024 24919 6080
rect 21357 6022 24919 6024
rect 21357 6019 21423 6022
rect 24853 6019 24919 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 24761 5946 24827 5949
rect 27520 5946 28000 5976
rect 24761 5944 28000 5946
rect 24761 5888 24766 5944
rect 24822 5888 28000 5944
rect 24761 5886 28000 5888
rect 24761 5883 24827 5886
rect 27520 5856 28000 5886
rect 19057 5810 19123 5813
rect 24577 5810 24643 5813
rect 19057 5808 24643 5810
rect 19057 5752 19062 5808
rect 19118 5752 24582 5808
rect 24638 5752 24643 5808
rect 19057 5750 24643 5752
rect 19057 5747 19123 5750
rect 24577 5747 24643 5750
rect 0 5538 480 5568
rect 2957 5538 3023 5541
rect 0 5536 3023 5538
rect 0 5480 2962 5536
rect 3018 5480 3023 5536
rect 0 5478 3023 5480
rect 0 5448 480 5478
rect 2957 5475 3023 5478
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 24761 5402 24827 5405
rect 27520 5402 28000 5432
rect 24761 5400 28000 5402
rect 24761 5344 24766 5400
rect 24822 5344 28000 5400
rect 24761 5342 28000 5344
rect 24761 5339 24827 5342
rect 27520 5312 28000 5342
rect 22553 5266 22619 5269
rect 24577 5266 24643 5269
rect 22553 5264 24643 5266
rect 22553 5208 22558 5264
rect 22614 5208 24582 5264
rect 24638 5208 24643 5264
rect 22553 5206 24643 5208
rect 22553 5203 22619 5206
rect 24577 5203 24643 5206
rect 10277 4928 10597 4929
rect 0 4858 480 4888
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 1669 4858 1735 4861
rect 0 4856 1735 4858
rect 0 4800 1674 4856
rect 1730 4800 1735 4856
rect 0 4798 1735 4800
rect 0 4768 480 4798
rect 1669 4795 1735 4798
rect 21265 4858 21331 4861
rect 27520 4858 28000 4888
rect 21265 4856 28000 4858
rect 21265 4800 21270 4856
rect 21326 4800 28000 4856
rect 21265 4798 28000 4800
rect 21265 4795 21331 4798
rect 27520 4768 28000 4798
rect 25681 4450 25747 4453
rect 27520 4450 28000 4480
rect 25681 4448 28000 4450
rect 25681 4392 25686 4448
rect 25742 4392 28000 4448
rect 25681 4390 28000 4392
rect 25681 4387 25747 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 27520 4360 28000 4390
rect 24277 4319 24597 4320
rect 0 4178 480 4208
rect 1485 4178 1551 4181
rect 0 4176 1551 4178
rect 0 4120 1490 4176
rect 1546 4120 1551 4176
rect 0 4118 1551 4120
rect 0 4088 480 4118
rect 1485 4115 1551 4118
rect 25589 3906 25655 3909
rect 27520 3906 28000 3936
rect 25589 3904 28000 3906
rect 25589 3848 25594 3904
rect 25650 3848 28000 3904
rect 25589 3846 28000 3848
rect 25589 3843 25655 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 27520 3816 28000 3846
rect 19610 3775 19930 3776
rect 0 3498 480 3528
rect 1577 3498 1643 3501
rect 0 3496 1643 3498
rect 0 3440 1582 3496
rect 1638 3440 1643 3496
rect 0 3438 1643 3440
rect 0 3408 480 3438
rect 1577 3435 1643 3438
rect 25037 3362 25103 3365
rect 27520 3362 28000 3392
rect 25037 3360 28000 3362
rect 25037 3304 25042 3360
rect 25098 3304 28000 3360
rect 25037 3302 28000 3304
rect 25037 3299 25103 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 27520 3272 28000 3302
rect 24277 3231 24597 3232
rect 1853 3090 1919 3093
rect 8109 3090 8175 3093
rect 1853 3088 8175 3090
rect 1853 3032 1858 3088
rect 1914 3032 8114 3088
rect 8170 3032 8175 3088
rect 1853 3030 8175 3032
rect 1853 3027 1919 3030
rect 8109 3027 8175 3030
rect 23841 3090 23907 3093
rect 25865 3090 25931 3093
rect 23841 3088 25931 3090
rect 23841 3032 23846 3088
rect 23902 3032 25870 3088
rect 25926 3032 25931 3088
rect 23841 3030 25931 3032
rect 23841 3027 23907 3030
rect 25865 3027 25931 3030
rect 0 2954 480 2984
rect 1761 2954 1827 2957
rect 0 2952 1827 2954
rect 0 2896 1766 2952
rect 1822 2896 1827 2952
rect 0 2894 1827 2896
rect 0 2864 480 2894
rect 1761 2891 1827 2894
rect 25313 2818 25379 2821
rect 27520 2818 28000 2848
rect 25313 2816 28000 2818
rect 25313 2760 25318 2816
rect 25374 2760 28000 2816
rect 25313 2758 28000 2760
rect 25313 2755 25379 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 27520 2728 28000 2758
rect 19610 2687 19930 2688
rect 0 2274 480 2304
rect 1577 2274 1643 2277
rect 0 2272 1643 2274
rect 0 2216 1582 2272
rect 1638 2216 1643 2272
rect 0 2214 1643 2216
rect 0 2184 480 2214
rect 1577 2211 1643 2214
rect 25405 2274 25471 2277
rect 27520 2274 28000 2304
rect 25405 2272 28000 2274
rect 25405 2216 25410 2272
rect 25466 2216 28000 2272
rect 25405 2214 28000 2216
rect 25405 2211 25471 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 27520 2184 28000 2214
rect 24277 2143 24597 2144
rect 25497 1730 25563 1733
rect 27520 1730 28000 1760
rect 25497 1728 28000 1730
rect 25497 1672 25502 1728
rect 25558 1672 28000 1728
rect 25497 1670 28000 1672
rect 25497 1667 25563 1670
rect 27520 1640 28000 1670
rect 0 1594 480 1624
rect 8845 1594 8911 1597
rect 0 1592 8911 1594
rect 0 1536 8850 1592
rect 8906 1536 8911 1592
rect 0 1534 8911 1536
rect 0 1504 480 1534
rect 8845 1531 8911 1534
rect 7557 1458 7623 1461
rect 3374 1456 7623 1458
rect 3374 1400 7562 1456
rect 7618 1400 7623 1456
rect 3374 1398 7623 1400
rect 0 914 480 944
rect 3374 914 3434 1398
rect 7557 1395 7623 1398
rect 23657 1186 23723 1189
rect 27520 1186 28000 1216
rect 23657 1184 28000 1186
rect 23657 1128 23662 1184
rect 23718 1128 28000 1184
rect 23657 1126 28000 1128
rect 23657 1123 23723 1126
rect 27520 1096 28000 1126
rect 0 854 3434 914
rect 0 824 480 854
rect 23013 642 23079 645
rect 27520 642 28000 672
rect 23013 640 28000 642
rect 23013 584 23018 640
rect 23074 584 28000 640
rect 23013 582 28000 584
rect 23013 579 23079 582
rect 27520 552 28000 582
rect 0 370 480 400
rect 3509 370 3575 373
rect 0 368 3575 370
rect 0 312 3514 368
rect 3570 312 3575 368
rect 0 310 3575 312
rect 0 280 480 310
rect 3509 307 3575 310
rect 25221 234 25287 237
rect 27520 234 28000 264
rect 25221 232 28000 234
rect 25221 176 25226 232
rect 25282 176 28000 232
rect 25221 174 28000 176
rect 25221 171 25287 174
rect 27520 144 28000 174
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 21772 23836 21836 23900
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 8156 22672 8220 22676
rect 8156 22616 8170 22672
rect 8170 22616 8220 22672
rect 8156 22612 8220 22616
rect 19380 22612 19444 22676
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 14228 20572 14292 20636
rect 19380 20572 19444 20636
rect 13676 20300 13740 20364
rect 15884 20164 15948 20228
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5396 18668 5460 18732
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 23796 18320 23860 18324
rect 23796 18264 23846 18320
rect 23846 18264 23860 18320
rect 23796 18260 23860 18264
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 23796 15676 23860 15740
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 24716 12472 24780 12476
rect 24716 12416 24766 12472
rect 24766 12416 24780 12472
rect 24716 12412 24780 12416
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 23796 10296 23860 10300
rect 23796 10240 23846 10296
rect 23846 10240 23860 10296
rect 23796 10236 23860 10240
rect 24716 10024 24780 10028
rect 24716 9968 24730 10024
rect 24730 9968 24780 10024
rect 24716 9964 24780 9968
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 8156 8060 8220 8124
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 8155 22676 8221 22677
rect 8155 22612 8156 22676
rect 8220 22612 8221 22676
rect 8155 22611 8221 22612
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 8158 8125 8218 22611
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 21771 23900 21837 23901
rect 21771 23836 21772 23900
rect 21836 23836 21837 23900
rect 21771 23835 21837 23836
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19379 22676 19445 22677
rect 19379 22612 19380 22676
rect 19444 22612 19445 22676
rect 19379 22611 19445 22612
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 13678 20710 14290 20770
rect 13678 20365 13738 20710
rect 14230 20637 14290 20710
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14227 20636 14293 20637
rect 14227 20572 14228 20636
rect 14292 20572 14293 20636
rect 14227 20571 14293 20572
rect 13675 20364 13741 20365
rect 13675 20300 13676 20364
rect 13740 20300 13741 20364
rect 13675 20299 13741 20300
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 8155 8124 8221 8125
rect 8155 8060 8156 8124
rect 8220 8060 8221 8124
rect 8155 8059 8221 8060
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 19616 15264 20640
rect 19382 20637 19442 22611
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19379 20636 19445 20637
rect 19379 20572 19380 20636
rect 19444 20572 19445 20636
rect 19379 20571 19445 20572
rect 15883 20228 15949 20229
rect 15883 20164 15884 20228
rect 15948 20164 15949 20228
rect 15883 20163 15949 20164
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 15886 18138 15946 20163
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 21774 18818 21834 23835
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 23795 18324 23861 18325
rect 23795 18260 23796 18324
rect 23860 18260 23861 18324
rect 23795 18259 23861 18260
rect 23798 18138 23858 18259
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 23795 15740 23861 15741
rect 23795 15676 23796 15740
rect 23860 15676 23861 15740
rect 23795 15675 23861 15676
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 23798 10301 23858 15675
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24715 12476 24781 12477
rect 24715 12412 24716 12476
rect 24780 12412 24781 12476
rect 24715 12411 24781 12412
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 23795 10300 23861 10301
rect 23795 10236 23796 10300
rect 23860 10236 23861 10300
rect 23795 10235 23861 10236
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 9824 24597 10848
rect 24718 10029 24778 12411
rect 24715 10028 24781 10029
rect 24715 9964 24716 10028
rect 24780 9964 24781 10028
rect 24715 9963 24781 9964
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 5310 18732 5546 18818
rect 5310 18668 5396 18732
rect 5396 18668 5460 18732
rect 5460 18668 5546 18732
rect 5310 18582 5546 18668
rect 15798 17902 16034 18138
rect 21686 18582 21922 18818
rect 23710 17902 23946 18138
<< metal5 >>
rect 5268 18818 21964 18860
rect 5268 18582 5310 18818
rect 5546 18582 21686 18818
rect 21922 18582 21964 18818
rect 5268 18540 21964 18582
rect 15756 18138 23988 18180
rect 15756 17902 15798 18138
rect 16034 17902 23710 18138
rect 23946 17902 23988 18138
rect 15756 17860 23988 17902
use scs8hd_fill_2  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_7
timestamp 1586364061
transform 1 0 1748 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1564 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_buf_2  _083_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_1_19 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2852 0 1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_11
timestamp 1586364061
transform 1 0 2116 0 -1 2720
box -38 -48 1142 592
use scs8hd_buf_4  mux_left_track_5.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3680 0 1 2720
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_34
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_38
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_8  FILLER_1_50
timestamp 1586364061
transform 1 0 5704 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  FILLER_1_58
timestamp 1586364061
transform 1 0 6440 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_67
timestamp 1586364061
transform 1 0 7268 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_63 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _085_
timestamp 1586364061
transform 1 0 7360 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_4  mux_left_track_1.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 8096 0 1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_76
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_88
timestamp 1586364061
transform 1 0 9200 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_92
timestamp 1586364061
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_82
timestamp 1586364061
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _105_
timestamp 1586364061
transform 1 0 22816 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_244
timestamp 1586364061
transform 1 0 23552 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_240
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_4  mux_right_track_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23828 0 1 2720
box -38 -48 590 592
use scs8hd_buf_4  mux_right_track_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_253
timestamp 1586364061
transform 1 0 24380 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_255
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24748 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_265
timestamp 1586364061
transform 1 0 25484 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_260
timestamp 1586364061
transform 1 0 25024 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_259
timestamp 1586364061
transform 1 0 24932 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 24840 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _103_
timestamp 1586364061
transform 1 0 25300 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_2  _101_
timestamp 1586364061
transform 1 0 25116 0 1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use scs8hd_decap_6  FILLER_0_271
timestamp 1586364061
transform 1 0 26036 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_267
timestamp 1586364061
transform 1 0 25668 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 25668 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 25852 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_buf_2  _081_
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_7
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_19
timestamp 1586364061
transform 1 0 2852 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_buf_4  mux_right_track_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23552 0 -1 3808
box -38 -48 590 592
use scs8hd_decap_4  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_243
timestamp 1586364061
transform 1 0 23460 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_250
timestamp 1586364061
transform 1 0 24104 0 -1 3808
box -38 -48 774 592
use scs8hd_buf_2  _100_
timestamp 1586364061
transform 1 0 24840 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_262
timestamp 1586364061
transform 1 0 25208 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_2_274
timestamp 1586364061
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_buf_4  mux_left_track_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1656 0 1 3808
box -38 -48 590 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_12
timestamp 1586364061
transform 1 0 2208 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_16
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_28
timestamp 1586364061
transform 1 0 3680 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_40
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_52
timestamp 1586364061
transform 1 0 5888 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_60
timestamp 1586364061
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 21068 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_3_216
timestamp 1586364061
transform 1 0 20976 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_219
timestamp 1586364061
transform 1 0 21252 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_231
timestamp 1586364061
transform 1 0 22356 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_243
timestamp 1586364061
transform 1 0 23460 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_buf_2  _097_
timestamp 1586364061
transform 1 0 21068 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_221
timestamp 1586364061
transform 1 0 21436 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_233
timestamp 1586364061
transform 1 0 22540 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_245
timestamp 1586364061
transform 1 0 23644 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_257
timestamp 1586364061
transform 1 0 24748 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_4_269
timestamp 1586364061
transform 1 0 25852 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20884 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_214
timestamp 1586364061
transform 1 0 20792 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_217
timestamp 1586364061
transform 1 0 21068 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_229
timestamp 1586364061
transform 1 0 22172 0 1 4896
box -38 -48 1142 592
use scs8hd_buf_2  _096_
timestamp 1586364061
transform 1 0 24564 0 1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 24380 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_241
timestamp 1586364061
transform 1 0 23276 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 25116 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_259
timestamp 1586364061
transform 1 0 24932 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_263
timestamp 1586364061
transform 1 0 25300 0 1 4896
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_5_275
timestamp 1586364061
transform 1 0 26404 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_buf_2  _077_
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_31
timestamp 1586364061
transform 1 0 3956 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_36
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_40
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_44
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_56
timestamp 1586364061
transform 1 0 6256 0 1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_60
timestamp 1586364061
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 774 592
use scs8hd_buf_2  _084_
timestamp 1586364061
transform 1 0 8648 0 1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_90
timestamp 1586364061
transform 1 0 9384 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_102
timestamp 1586364061
transform 1 0 10488 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_171
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use scs8hd_buf_4  mux_right_track_16.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_221
timestamp 1586364061
transform 1 0 21436 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_233
timestamp 1586364061
transform 1 0 22540 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use scs8hd_buf_2  _094_
timestamp 1586364061
transform 1 0 24564 0 1 5984
box -38 -48 406 592
use scs8hd_buf_2  _095_
timestamp 1586364061
transform 1 0 24564 0 -1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 24380 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_245
timestamp 1586364061
transform 1 0 23644 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_253
timestamp 1586364061
transform 1 0 24380 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_259
timestamp 1586364061
transform 1 0 24932 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 25116 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_275
timestamp 1586364061
transform 1 0 26404 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_271
timestamp 1586364061
transform 1 0 26036 0 -1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_263
timestamp 1586364061
transform 1 0 25300 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_259
timestamp 1586364061
transform 1 0 24932 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 1564 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_7
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_19
timestamp 1586364061
transform 1 0 2852 0 -1 7072
box -38 -48 1142 592
use scs8hd_buf_4  mux_left_track_17.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 4600 0 -1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 8004 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_74
timestamp 1586364061
transform 1 0 7912 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_77
timestamp 1586364061
transform 1 0 8188 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 9844 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 10212 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_81
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_85
timestamp 1586364061
transform 1 0 8924 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_91
timestamp 1586364061
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_97
timestamp 1586364061
transform 1 0 10028 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_101
timestamp 1586364061
transform 1 0 10396 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_8_113
timestamp 1586364061
transform 1 0 11500 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_119
timestamp 1586364061
transform 1 0 12052 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_131
timestamp 1586364061
transform 1 0 13156 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_143
timestamp 1586364061
transform 1 0 14260 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_151
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _092_
timestamp 1586364061
transform 1 0 24564 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_259
timestamp 1586364061
transform 1 0 24932 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_8_271
timestamp 1586364061
transform 1 0 26036 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_2  _075_
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_7
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_11
timestamp 1586364061
transform 1 0 2116 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_23
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_35
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 5888 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 6256 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_47
timestamp 1586364061
transform 1 0 5428 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_50
timestamp 1586364061
transform 1 0 5704 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_54
timestamp 1586364061
transform 1 0 6072 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_58
timestamp 1586364061
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_1.mux_l2_in_3_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 7452 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_9_68
timestamp 1586364061
transform 1 0 7360 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_71
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_75
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_buf_4  mux_left_track_3.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_88
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_92
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_95
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 11868 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 11500 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 10672 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_102
timestamp 1586364061
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_106
timestamp 1586364061
transform 1 0 10856 0 1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_9_112
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_115
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_119
timestamp 1586364061
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 13064 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 12604 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_127
timestamp 1586364061
transform 1 0 12788 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_132
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_136
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_140
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_144
timestamp 1586364061
transform 1 0 14352 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_156
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_168
timestamp 1586364061
transform 1 0 16560 0 1 7072
box -38 -48 406 592
use scs8hd_decap_8  FILLER_9_174
timestamp 1586364061
transform 1 0 17112 0 1 7072
box -38 -48 774 592
use scs8hd_buf_2  _093_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 18584 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_182
timestamp 1586364061
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_188
timestamp 1586364061
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_192
timestamp 1586364061
transform 1 0 18768 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_204
timestamp 1586364061
transform 1 0 19872 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_216
timestamp 1586364061
transform 1 0 20976 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_228
timestamp 1586364061
transform 1 0 22080 0 1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _091_
timestamp 1586364061
transform 1 0 24564 0 1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 24380 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 23828 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_240
timestamp 1586364061
transform 1 0 23184 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_249
timestamp 1586364061
transform 1 0 24012 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 25116 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_259
timestamp 1586364061
transform 1 0 24932 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_263
timestamp 1586364061
transform 1 0 25300 0 1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_9_275
timestamp 1586364061
transform 1 0 26404 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _074_
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_7
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_19
timestamp 1586364061
transform 1 0 2852 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_mux2_2  mux_left_track_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 5888 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 774 592
use scs8hd_mux2_2  mux_left_track_1.mux_l2_in_2_
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 6900 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_61
timestamp 1586364061
transform 1 0 6716 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_65
timestamp 1586364061
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_69
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 590 592
use scs8hd_mux2_2  mux_left_track_1.mux_l3_in_1_
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 590 592
use scs8hd_mux2_2  mux_left_track_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_106
timestamp 1586364061
transform 1 0 10856 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_10_114
timestamp 1586364061
transform 1 0 11592 0 -1 8160
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13432 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 13064 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_126
timestamp 1586364061
transform 1 0 12696 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_132
timestamp 1586364061
transform 1 0 13248 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_143
timestamp 1586364061
transform 1 0 14260 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_147
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_12  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use scs8hd_buf_4  mux_right_track_24.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16928 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_6  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_8  FILLER_10_178
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 18216 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_188
timestamp 1586364061
transform 1 0 18400 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_200
timestamp 1586364061
transform 1 0 19504 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_10_212
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_buf_2  _090_
timestamp 1586364061
transform 1 0 24564 0 -1 8160
box -38 -48 406 592
use scs8hd_buf_2  _104_
timestamp 1586364061
transform 1 0 23460 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 23184 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_242
timestamp 1586364061
transform 1 0 23368 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_247
timestamp 1586364061
transform 1 0 23828 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_259
timestamp 1586364061
transform 1 0 24932 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_10_271
timestamp 1586364061
transform 1 0 26036 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_buf_2  _073_
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_11
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6256 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 5888 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 5520 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_47
timestamp 1586364061
transform 1 0 5428 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_50
timestamp 1586364061
transform 1 0 5704 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_54
timestamp 1586364061
transform 1 0 6072 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_58
timestamp 1586364061
transform 1 0 6440 0 1 8160
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_5.mux_l2_in_3_
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_71
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_83
timestamp 1586364061
transform 1 0 8740 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_87
timestamp 1586364061
transform 1 0 9108 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_109
timestamp 1586364061
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_113
timestamp 1586364061
transform 1 0 11500 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_132
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_136
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_1.mux_l1_in_2_
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 866 592
use scs8hd_decap_12  FILLER_11_149
timestamp 1586364061
transform 1 0 14812 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_161
timestamp 1586364061
transform 1 0 15916 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_11_173
timestamp 1586364061
transform 1 0 17020 0 1 8160
box -38 -48 406 592
use scs8hd_buf_4  mux_right_track_32.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18216 0 1 8160
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_192
timestamp 1586364061
transform 1 0 18768 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 20976 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_11_218
timestamp 1586364061
transform 1 0 21160 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 21712 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_222
timestamp 1586364061
transform 1 0 21528 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_226
timestamp 1586364061
transform 1 0 21896 0 1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_11_234
timestamp 1586364061
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_238
timestamp 1586364061
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use scs8hd_buf_4  mux_right_track_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24380 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_242
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_251
timestamp 1586364061
transform 1 0 24196 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_255
timestamp 1586364061
transform 1 0 24564 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _089_
timestamp 1586364061
transform 1 0 24932 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 25484 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_263
timestamp 1586364061
transform 1 0 25300 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_267
timestamp 1586364061
transform 1 0 25668 0 1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_11_275
timestamp 1586364061
transform 1 0 26404 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _080_
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 1932 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_7
timestamp 1586364061
transform 1 0 1748 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_11
timestamp 1586364061
transform 1 0 2116 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 4232 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_36
timestamp 1586364061
transform 1 0 4416 0 -1 9248
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4784 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_42
timestamp 1586364061
transform 1 0 4968 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_46
timestamp 1586364061
transform 1 0 5336 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_54
timestamp 1586364061
transform 1 0 6072 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8188 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_75
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_79
timestamp 1586364061
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__S
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 10028 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_83
timestamp 1586364061
transform 1 0 8740 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_89
timestamp 1586364061
transform 1 0 9292 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_99
timestamp 1586364061
transform 1 0 10212 0 -1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 10580 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 10396 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_3.mux_l2_in_1_
timestamp 1586364061
transform 1 0 13064 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12512 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 12880 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_122
timestamp 1586364061
transform 1 0 12328 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_126
timestamp 1586364061
transform 1 0 12696 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_143
timestamp 1586364061
transform 1 0 14260 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_12_139
timestamp 1586364061
transform 1 0 13892 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_152
timestamp 1586364061
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_149
timestamp 1586364061
transform 1 0 14812 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 15456 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 14904 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_158
timestamp 1586364061
transform 1 0 15640 0 -1 9248
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 17112 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_170
timestamp 1586364061
transform 1 0 16744 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_176
timestamp 1586364061
transform 1 0 17296 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_32.mux_l1_in_2_
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_180
timestamp 1586364061
transform 1 0 17664 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_195
timestamp 1586364061
transform 1 0 19044 0 -1 9248
box -38 -48 1142 592
use scs8hd_mux2_2  mux_right_track_2.mux_l2_in_2_
timestamp 1586364061
transform 1 0 20976 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_12_207
timestamp 1586364061
transform 1 0 20148 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_213
timestamp 1586364061
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 23000 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_225
timestamp 1586364061
transform 1 0 21804 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_237
timestamp 1586364061
transform 1 0 22908 0 -1 9248
box -38 -48 130 592
use scs8hd_buf_2  _088_
timestamp 1586364061
transform 1 0 24748 0 -1 9248
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_track_8.mux_l3_in_1_
timestamp 1586364061
transform 1 0 23184 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_249
timestamp 1586364061
transform 1 0 24012 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_253
timestamp 1586364061
transform 1 0 24380 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_261
timestamp 1586364061
transform 1 0 25116 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_12_273
timestamp 1586364061
transform 1 0 26220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_buf_2  _079_
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use scs8hd_buf_2  _072_
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_7
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1932 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_11
timestamp 1586364061
transform 1 0 2116 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_11
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 2300 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 2300 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_19
timestamp 1586364061
transform 1 0 2852 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_19
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  _071_
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 406 592
use scs8hd_buf_2  _067_
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_29
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_25
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_23
timestamp 1586364061
transform 1 0 3220 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 3036 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_36
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_31
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 4600 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4784 0 -1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 406 592
use scs8hd_decap_4  FILLER_14_59
timestamp 1586364061
transform 1 0 6532 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_69
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_65
timestamp 1586364061
transform 1 0 7084 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_69
timestamp 1586364061
transform 1 0 7452 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_65
timestamp 1586364061
transform 1 0 7084 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__A1
timestamp 1586364061
transform 1 0 7268 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 6900 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_conb_1  _058_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 7544 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__A0
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_5.mux_l1_in_6_
timestamp 1586364061
transform 1 0 7728 0 -1 10336
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 1786 592
use scs8hd_decap_3  FILLER_14_81
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_86
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_90
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_92
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_97
timestamp 1586364061
transform 1 0 10028 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_96
timestamp 1586364061
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 10212 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_101
timestamp 1586364061
transform 1 0 10396 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_3  FILLER_13_109
timestamp 1586364061
transform 1 0 11132 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_3.mux_l4_in_0_
timestamp 1586364061
transform 1 0 10304 0 1 9248
box -38 -48 866 592
use scs8hd_mux2_2  mux_left_track_3.mux_l3_in_1_
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_116
timestamp 1586364061
transform 1 0 11776 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1786 592
use scs8hd_mux2_2  mux_left_track_3.mux_l2_in_3_
timestamp 1586364061
transform 1 0 12512 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12328 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_120
timestamp 1586364061
transform 1 0 12144 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_133
timestamp 1586364061
transform 1 0 13340 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_148
timestamp 1586364061
transform 1 0 14720 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_144
timestamp 1586364061
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_146
timestamp 1586364061
transform 1 0 14536 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_142
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14352 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14536 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 14720 0 1 9248
box -38 -48 222 592
use scs8hd_conb_1  _056_
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_152
timestamp 1586364061
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 14904 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_32.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use scs8hd_mux2_2  mux_left_track_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 14904 0 1 9248
box -38 -48 866 592
use scs8hd_decap_6  FILLER_13_163
timestamp 1586364061
transform 1 0 16100 0 1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_159
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 15916 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_175
timestamp 1586364061
transform 1 0 17204 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_13_169
timestamp 1586364061
transform 1 0 16652 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 16744 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 17296 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 17480 0 1 9248
box -38 -48 222 592
use scs8hd_conb_1  _064_
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_track_32.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_track_32.mux_l3_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_180
timestamp 1586364061
transform 1 0 17664 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_198
timestamp 1586364061
transform 1 0 19320 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_197
timestamp 1586364061
transform 1 0 19228 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_205
timestamp 1586364061
transform 1 0 19964 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_201
timestamp 1586364061
transform 1 0 19596 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_206
timestamp 1586364061
transform 1 0 20056 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_202
timestamp 1586364061
transform 1 0 19688 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 19504 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 19412 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 19872 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 19780 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_213
timestamp 1586364061
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_210
timestamp 1586364061
transform 1 0 20424 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 20608 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_2.mux_l3_in_1_
timestamp 1586364061
transform 1 0 20792 0 1 9248
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_13_223
timestamp 1586364061
transform 1 0 21620 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_227
timestamp 1586364061
transform 1 0 21988 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 21804 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 22172 0 1 9248
box -38 -48 222 592
use scs8hd_conb_1  _062_
timestamp 1586364061
transform 1 0 22356 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_234
timestamp 1586364061
transform 1 0 22632 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_234
timestamp 1586364061
transform 1 0 22632 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 22816 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_238
timestamp 1586364061
transform 1 0 23000 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_240
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 23184 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_8.mux_l4_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 866 592
use scs8hd_mux2_2  mux_right_track_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 23368 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_255
timestamp 1586364061
transform 1 0 24564 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_254
timestamp 1586364061
transform 1 0 24472 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 24748 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 24380 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_266
timestamp 1586364061
transform 1 0 25576 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_261
timestamp 1586364061
transform 1 0 25116 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_258
timestamp 1586364061
transform 1 0 24840 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 24932 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  _087_
timestamp 1586364061
transform 1 0 25208 0 1 9248
box -38 -48 406 592
use scs8hd_buf_2  _086_
timestamp 1586364061
transform 1 0 24932 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_276
timestamp 1586364061
transform 1 0 26496 0 1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_13_270
timestamp 1586364061
transform 1 0 25944 0 1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 25760 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_2  _070_
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 406 592
use scs8hd_buf_2  _082_
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 2300 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_11
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_19
timestamp 1586364061
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use scs8hd_buf_2  _069_
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 406 592
use scs8hd_mux2_2  mux_left_track_5.mux_l4_in_0_
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 3036 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 4140 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 4508 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_23
timestamp 1586364061
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_31
timestamp 1586364061
transform 1 0 3956 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_35
timestamp 1586364061
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 5888 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_48
timestamp 1586364061
transform 1 0 5520 0 1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_15_54
timestamp 1586364061
transform 1 0 6072 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_58
timestamp 1586364061
transform 1 0 6440 0 1 10336
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_5.mux_l1_in_2_
timestamp 1586364061
transform 1 0 6900 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_72
timestamp 1586364061
transform 1 0 7728 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_76
timestamp 1586364061
transform 1 0 8096 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9200 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_80
timestamp 1586364061
transform 1 0 8464 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_84
timestamp 1586364061
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_97
timestamp 1586364061
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_101
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_3.mux_l2_in_2_
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_136
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 14536 0 1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 14352 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_140
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_165
timestamp 1586364061
transform 1 0 16284 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_32.mux_l2_in_1_
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_track_2.mux_l2_in_3_
timestamp 1586364061
transform 1 0 19780 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 20792 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_199
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_212
timestamp 1586364061
transform 1 0 20608 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_216
timestamp 1586364061
transform 1 0 20976 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_2.mux_l4_in_0_
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 22356 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 22724 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_229
timestamp 1586364061
transform 1 0 22172 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_233
timestamp 1586364061
transform 1 0 22540 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_237
timestamp 1586364061
transform 1 0 22908 0 1 10336
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_241
timestamp 1586364061
transform 1 0 23276 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_264
timestamp 1586364061
transform 1 0 25392 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_268
timestamp 1586364061
transform 1 0 25760 0 1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_15_276
timestamp 1586364061
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use scs8hd_buf_2  _078_
timestamp 1586364061
transform 1 0 2668 0 -1 11424
box -38 -48 406 592
use scs8hd_buf_4  mux_left_track_33.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 2116 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_9
timestamp 1586364061
transform 1 0 1932 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_13
timestamp 1586364061
transform 1 0 2300 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_9.mux_l2_in_3_
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_21
timestamp 1586364061
transform 1 0 3036 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_5.mux_l3_in_1_
timestamp 1586364061
transform 1 0 5888 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 5060 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 5428 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_41
timestamp 1586364061
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_45
timestamp 1586364061
transform 1 0 5244 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_49
timestamp 1586364061
transform 1 0 5612 0 -1 11424
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_5.mux_l1_in_4_
timestamp 1586364061
transform 1 0 7728 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_5__A1
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 6900 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_61
timestamp 1586364061
transform 1 0 6716 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_65
timestamp 1586364061
transform 1 0 7084 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_69
timestamp 1586364061
transform 1 0 7452 0 -1 11424
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_5.mux_l1_in_1_
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_81
timestamp 1586364061
transform 1 0 8556 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_86
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_90
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11684 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11500 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 11132 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_102
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_107
timestamp 1586364061
transform 1 0 10948 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_111
timestamp 1586364061
transform 1 0 11316 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_134
timestamp 1586364061
transform 1 0 13432 0 -1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 15640 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14260 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_142
timestamp 1586364061
transform 1 0 14168 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_4  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_32.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16652 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 16008 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_160
timestamp 1586364061
transform 1 0 15824 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_164
timestamp 1586364061
transform 1 0 16192 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_168
timestamp 1586364061
transform 1 0 16560 0 -1 11424
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_32.mux_l2_in_0_
timestamp 1586364061
transform 1 0 19136 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 18768 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_188
timestamp 1586364061
transform 1 0 18400 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_194
timestamp 1586364061
transform 1 0 18952 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 21068 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_205
timestamp 1586364061
transform 1 0 19964 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_213
timestamp 1586364061
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 21804 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 21436 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_219
timestamp 1586364061
transform 1 0 21252 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_223
timestamp 1586364061
transform 1 0 21620 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_0.mux_l2_in_2_
timestamp 1586364061
transform 1 0 24288 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 24104 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23736 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_244
timestamp 1586364061
transform 1 0 23552 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_248
timestamp 1586364061
transform 1 0 23920 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_261
timestamp 1586364061
transform 1 0 25116 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_16_273
timestamp 1586364061
transform 1 0 26220 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_1.mux_l4_in_0_
timestamp 1586364061
transform 1 0 1656 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 2668 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_19
timestamp 1586364061
transform 1 0 2852 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_9.mux_l3_in_1_
timestamp 1586364061
transform 1 0 3220 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 3036 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_32
timestamp 1586364061
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_36
timestamp 1586364061
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_9.mux_l2_in_2_
timestamp 1586364061
transform 1 0 4784 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_49
timestamp 1586364061
transform 1 0 5612 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_5.mux_l1_in_5_
timestamp 1586364061
transform 1 0 7544 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 7360 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 6992 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_66
timestamp 1586364061
transform 1 0 7176 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_79
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_5.mux_l2_in_1_
timestamp 1586364061
transform 1 0 9108 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_5__A0
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_5__S
timestamp 1586364061
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_83
timestamp 1586364061
transform 1 0 8740 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_96
timestamp 1586364061
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_100
timestamp 1586364061
transform 1 0 10304 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 13708 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14076 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_139
timestamp 1586364061
transform 1 0 13892 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_162
timestamp 1586364061
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_166
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_17_174
timestamp 1586364061
transform 1 0 17112 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_177
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18768 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 18584 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 18216 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_181
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_188
timestamp 1586364061
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 20700 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 20516 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 20148 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 19780 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_201
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_205
timestamp 1586364061
transform 1 0 19964 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_209
timestamp 1586364061
transform 1 0 20332 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 21712 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_222
timestamp 1586364061
transform 1 0 21528 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_226
timestamp 1586364061
transform 1 0 21896 0 1 11424
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 24104 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23920 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_240
timestamp 1586364061
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use scs8hd_conb_1  _059_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_9.mux_l4_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 2116 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_6
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_10
timestamp 1586364061
transform 1 0 2024 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_13
timestamp 1586364061
transform 1 0 2300 0 -1 12512
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 6532 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 5980 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_51
timestamp 1586364061
transform 1 0 5796 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_55
timestamp 1586364061
transform 1 0 6164 0 -1 12512
box -38 -48 406 592
use scs8hd_mux2_2  mux_left_track_5.mux_l1_in_3_
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 6900 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_61
timestamp 1586364061
transform 1 0 6716 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_65
timestamp 1586364061
transform 1 0 7084 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_77
timestamp 1586364061
transform 1 0 8188 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_81
timestamp 1586364061
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_85
timestamp 1586364061
transform 1 0 8924 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_89
timestamp 1586364061
transform 1 0 9292 0 -1 12512
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 11684 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_106
timestamp 1586364061
transform 1 0 10856 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_110
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_114
timestamp 1586364061
transform 1 0 11592 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 13800 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_136
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_32.mux_l1_in_1_
timestamp 1586364061
transform 1 0 15640 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_140
timestamp 1586364061
transform 1 0 13984 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_152
timestamp 1586364061
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_32.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 17204 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 16652 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_167
timestamp 1586364061
transform 1 0 16468 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_171
timestamp 1586364061
transform 1 0 16836 0 -1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_194
timestamp 1586364061
transform 1 0 18952 0 -1 12512
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 19596 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 19964 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_199
timestamp 1586364061
transform 1 0 19412 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_203
timestamp 1586364061
transform 1 0 19780 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_207
timestamp 1586364061
transform 1 0 20148 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_213
timestamp 1586364061
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_18_234
timestamp 1586364061
transform 1 0 22632 0 -1 12512
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 23828 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 23552 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 23184 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_242
timestamp 1586364061
transform 1 0 23368 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_246
timestamp 1586364061
transform 1 0 23736 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_266
timestamp 1586364061
transform 1 0 25576 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_274
timestamp 1586364061
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 1564 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 1932 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 1932 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_11
timestamp 1586364061
transform 1 0 2116 0 -1 13600
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_17.mux_l1_in_1_
timestamp 1586364061
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 2116 0 1 12512
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_36
timestamp 1586364061
transform 1 0 4416 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_34
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_30
timestamp 1586364061
transform 1 0 3864 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 4600 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_9.mux_l2_in_1_
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 866 592
use scs8hd_buf_2  _068_
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_40
timestamp 1586364061
transform 1 0 4784 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_47
timestamp 1586364061
transform 1 0 5428 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 5336 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 4968 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 5612 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_55
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 5520 0 -1 13600
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_20_67
timestamp 1586364061
transform 1 0 7268 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 7452 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_5.mux_l2_in_2_
timestamp 1586364061
transform 1 0 6900 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_71
timestamp 1586364061
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_77
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_72
timestamp 1586364061
transform 1 0 7728 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_38.mux_l1_in_1_
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_3  FILLER_20_89
timestamp 1586364061
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_88
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_83
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 222 592
use scs8hd_conb_1  _054_
timestamp 1586364061
transform 1 0 8464 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_96
timestamp 1586364061
transform 1 0 9936 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10120 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_conb_1  _053_
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11500 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_111
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_115
timestamp 1586364061
transform 1 0 11684 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_100
timestamp 1586364061
transform 1 0 10304 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_123
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_128
timestamp 1586364061
transform 1 0 12880 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_19_121
timestamp 1586364061
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 12696 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 13064 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l1_in_3_
timestamp 1586364061
transform 1 0 13156 0 -1 13600
box -38 -48 866 592
use scs8hd_mux2_2  mux_top_track_4.mux_l1_in_2_
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_20_140
timestamp 1586364061
transform 1 0 13984 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_145
timestamp 1586364061
transform 1 0 14444 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_141
timestamp 1586364061
transform 1 0 14076 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 14260 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_148
timestamp 1586364061
transform 1 0 14720 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_156
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_153
timestamp 1586364061
transform 1 0 15180 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_149
timestamp 1586364061
transform 1 0 14812 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_20_158
timestamp 1586364061
transform 1 0 15640 0 -1 13600
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 16192 0 -1 13600
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_track_24.mux_l3_in_0_
timestamp 1586364061
transform 1 0 16192 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_160
timestamp 1586364061
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_173
timestamp 1586364061
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_177
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 590 592
use scs8hd_decap_4  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_183
timestamp 1586364061
transform 1 0 17940 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_188
timestamp 1586364061
transform 1 0 18400 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 18124 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_193
timestamp 1586364061
transform 1 0 18860 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_195
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_191
timestamp 1586364061
transform 1 0 18676 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 18492 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 18676 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 19044 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_2.mux_l1_in_1_
timestamp 1586364061
transform 1 0 19228 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_2.mux_l2_in_0_
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_210
timestamp 1586364061
transform 1 0 20424 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_212
timestamp 1586364061
transform 1 0 20608 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 21068 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 20424 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 20792 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 20976 0 1 12512
box -38 -48 866 592
use scs8hd_decap_4  FILLER_20_223
timestamp 1586364061
transform 1 0 21620 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_219
timestamp 1586364061
transform 1 0 21252 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_225
timestamp 1586364061
transform 1 0 21804 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 21436 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 21988 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_0.mux_l2_in_3_
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_236
timestamp 1586364061
transform 1 0 22816 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_237
timestamp 1586364061
transform 1 0 22908 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_233
timestamp 1586364061
transform 1 0 22540 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_229
timestamp 1586364061
transform 1 0 22172 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 22724 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 22356 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 23000 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_240
timestamp 1586364061
transform 1 0 23184 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_241
timestamp 1586364061
transform 1 0 23276 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 23368 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_0.mux_l4_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 866 592
use scs8hd_mux2_2  mux_right_track_0.mux_l3_in_1_
timestamp 1586364061
transform 1 0 23552 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_8  FILLER_20_253
timestamp 1586364061
transform 1 0 24380 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_254
timestamp 1586364061
transform 1 0 24472 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 24656 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_264
timestamp 1586364061
transform 1 0 25392 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_266
timestamp 1586364061
transform 1 0 25576 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_258
timestamp 1586364061
transform 1 0 24840 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 25024 0 1 12512
box -38 -48 222 592
use scs8hd_buf_2  _102_
timestamp 1586364061
transform 1 0 25208 0 1 12512
box -38 -48 406 592
use scs8hd_conb_1  _060_
timestamp 1586364061
transform 1 0 25116 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_272
timestamp 1586364061
transform 1 0 26128 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_6  FILLER_19_270
timestamp 1586364061
transform 1 0 25944 0 1 12512
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 25760 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_276
timestamp 1586364061
transform 1 0 26496 0 1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_0.mux_l2_in_2_
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_12
timestamp 1586364061
transform 1 0 2208 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_16
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_9.mux_l3_in_0_
timestamp 1586364061
transform 1 0 3404 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3220 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_20
timestamp 1586364061
transform 1 0 2944 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_34
timestamp 1586364061
transform 1 0 4232 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_38
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5060 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 4876 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_52
timestamp 1586364061
transform 1 0 5888 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_17.mux_l2_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use scs8hd_mux2_2  mux_left_track_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_71
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_75
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_88
timestamp 1586364061
transform 1 0 9200 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_92
timestamp 1586364061
transform 1 0 9568 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_97
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_101
timestamp 1586364061
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_24.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12880 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_127
timestamp 1586364061
transform 1 0 12788 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_130
timestamp 1586364061
transform 1 0 13064 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 14996 0 1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 14812 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 14444 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_143
timestamp 1586364061
transform 1 0 14260 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_147
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 16928 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 17296 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_170
timestamp 1586364061
transform 1 0 16744 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_174
timestamp 1586364061
transform 1 0 17112 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_178
timestamp 1586364061
transform 1 0 17480 0 1 13600
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_track_24.mux_l1_in_3_
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_193
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_197
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 19596 0 1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 21528 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_224
timestamp 1586364061
transform 1 0 21712 0 1 13600
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_21_236
timestamp 1586364061
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_240
timestamp 1586364061
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_264
timestamp 1586364061
transform 1 0 25392 0 1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_21_276
timestamp 1586364061
transform 1 0 26496 0 1 13600
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_0.mux_l2_in_3_
timestamp 1586364061
transform 1 0 1656 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 2668 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_19
timestamp 1586364061
transform 1 0 2852 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 3036 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 6440 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 5980 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_51
timestamp 1586364061
transform 1 0 5796 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_55
timestamp 1586364061
transform 1 0 6164 0 -1 14688
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_17.mux_l1_in_3_
timestamp 1586364061
transform 1 0 7176 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 8372 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 6808 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_60
timestamp 1586364061
transform 1 0 6624 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_64
timestamp 1586364061
transform 1 0 6992 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_75
timestamp 1586364061
transform 1 0 8004 0 -1 14688
box -38 -48 406 592
use scs8hd_mux2_2  mux_top_track_38.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9844 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8740 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_81
timestamp 1586364061
transform 1 0 8556 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_85
timestamp 1586364061
transform 1 0 8924 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_89
timestamp 1586364061
transform 1 0 9292 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 11408 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_104
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_108
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13432 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_131
timestamp 1586364061
transform 1 0 13156 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_136
timestamp 1586364061
transform 1 0 13616 0 -1 14688
box -38 -48 1142 592
use scs8hd_mux2_2  mux_right_track_24.mux_l1_in_1_
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_148
timestamp 1586364061
transform 1 0 14720 0 -1 14688
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_track_24.mux_l2_in_1_
timestamp 1586364061
transform 1 0 16836 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 16652 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_163
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 590 592
use scs8hd_mux2_2  mux_right_track_16.mux_l3_in_0_
timestamp 1586364061
transform 1 0 19228 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 18032 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18492 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 18860 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_180
timestamp 1586364061
transform 1 0 17664 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_3  FILLER_22_186
timestamp 1586364061
transform 1 0 18216 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_191
timestamp 1586364061
transform 1 0 18676 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_195
timestamp 1586364061
transform 1 0 19044 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 20516 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_206
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_210
timestamp 1586364061
transform 1 0 20424 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_213
timestamp 1586364061
transform 1 0 20700 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 22816 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_234
timestamp 1586364061
transform 1 0 22632 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_238
timestamp 1586364061
transform 1 0 23000 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 23368 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 23184 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 25300 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_261
timestamp 1586364061
transform 1 0 25116 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_265
timestamp 1586364061
transform 1 0 25484 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_273
timestamp 1586364061
transform 1 0 26220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_0.mux_l3_in_1_
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 2760 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_12
timestamp 1586364061
transform 1 0 2208 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_16
timestamp 1586364061
transform 1 0 2576 0 1 14688
box -38 -48 222 592
use scs8hd_buf_2  _076_
timestamp 1586364061
transform 1 0 2944 0 1 14688
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4232 0 1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 3496 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_24
timestamp 1586364061
transform 1 0 3312 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_28
timestamp 1586364061
transform 1 0 3680 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_17.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_71
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_75
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_79
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 130 592
use scs8hd_conb_1  _049_
timestamp 1586364061
transform 1 0 8464 0 1 14688
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_38.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 9292 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_38.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8924 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_83
timestamp 1586364061
transform 1 0 8740 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_87
timestamp 1586364061
transform 1 0 9108 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_91
timestamp 1586364061
transform 1 0 9476 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_136
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use scs8hd_conb_1  _050_
timestamp 1586364061
transform 1 0 13984 0 1 14688
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_track_24.mux_l2_in_0_
timestamp 1586364061
transform 1 0 14996 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 14812 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14444 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_143
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_147
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 222 592
use scs8hd_conb_1  _063_
timestamp 1586364061
transform 1 0 16928 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16744 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16376 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_160
timestamp 1586364061
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_164
timestamp 1586364061
transform 1 0 16192 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_168
timestamp 1586364061
transform 1 0 16560 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_16.mux_l2_in_1_
timestamp 1586364061
transform 1 0 20516 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 20332 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 19964 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_203
timestamp 1586364061
transform 1 0 19780 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_207
timestamp 1586364061
transform 1 0 20148 0 1 14688
box -38 -48 222 592
use scs8hd_conb_1  _061_
timestamp 1586364061
transform 1 0 22080 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 21528 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 22540 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 22908 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 21896 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_224
timestamp 1586364061
transform 1 0 21712 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_231
timestamp 1586364061
transform 1 0 22356 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_235
timestamp 1586364061
transform 1 0 22724 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_239
timestamp 1586364061
transform 1 0 23092 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_254
timestamp 1586364061
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use scs8hd_buf_2  _099_
timestamp 1586364061
transform 1 0 25208 0 1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 25760 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 25024 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_258
timestamp 1586364061
transform 1 0 24840 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_266
timestamp 1586364061
transform 1 0 25576 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_270
timestamp 1586364061
transform 1 0 25944 0 1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_23_276
timestamp 1586364061
transform 1 0 26496 0 1 14688
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 1472 0 -1 15776
box -38 -48 1786 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 130 592
use scs8hd_buf_2  _066_
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4600 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_36
timestamp 1586364061
transform 1 0 4416 0 -1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 5244 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 4968 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_40
timestamp 1586364061
transform 1 0 4784 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_17.mux_l1_in_2_
timestamp 1586364061
transform 1 0 7728 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7268 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_64
timestamp 1586364061
transform 1 0 6992 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_69
timestamp 1586364061
transform 1 0 7452 0 -1 15776
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_2.mux_l1_in_2_
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 8740 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 9108 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_81
timestamp 1586364061
transform 1 0 8556 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_85
timestamp 1586364061
transform 1 0 8924 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_89
timestamp 1586364061
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_38.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 11040 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_106
timestamp 1586364061
transform 1 0 10856 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_110
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_116
timestamp 1586364061
transform 1 0 11776 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_119
timestamp 1586364061
transform 1 0 12052 0 -1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12420 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12236 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 14812 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 15548 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_142
timestamp 1586364061
transform 1 0 14168 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_147
timestamp 1586364061
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_151
timestamp 1586364061
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use scs8hd_conb_1  _051_
timestamp 1586364061
transform 1 0 15732 0 -1 15776
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_track_16.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16744 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_162
timestamp 1586364061
transform 1 0 16008 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_168
timestamp 1586364061
transform 1 0 16560 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_16.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18492 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18032 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_179
timestamp 1586364061
transform 1 0 17572 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_183
timestamp 1586364061
transform 1 0 17940 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_24_186
timestamp 1586364061
transform 1 0 18216 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_198
timestamp 1586364061
transform 1 0 19320 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_16.mux_l1_in_3_
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 19504 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 20516 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 20148 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_202
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_206
timestamp 1586364061
transform 1 0 20056 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_209
timestamp 1586364061
transform 1 0 20332 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_213
timestamp 1586364061
transform 1 0 20700 0 -1 15776
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_16.mux_l1_in_2_
timestamp 1586364061
transform 1 0 22448 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 21896 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 22264 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_224
timestamp 1586364061
transform 1 0 21712 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_228
timestamp 1586364061
transform 1 0 22080 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_8.mux_l2_in_2_
timestamp 1586364061
transform 1 0 24012 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 23736 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_241
timestamp 1586364061
transform 1 0 23276 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_245
timestamp 1586364061
transform 1 0 23644 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_248
timestamp 1586364061
transform 1 0 23920 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 25024 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_258
timestamp 1586364061
transform 1 0 24840 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_262
timestamp 1586364061
transform 1 0 25208 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_24_274
timestamp 1586364061
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_conb_1  _034_
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2392 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 2208 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 1840 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_6
timestamp 1586364061
transform 1 0 1656 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_10
timestamp 1586364061
transform 1 0 2024 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 3404 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_23
timestamp 1586364061
transform 1 0 3220 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_31
timestamp 1586364061
transform 1 0 3956 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_34
timestamp 1586364061
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_38
timestamp 1586364061
transform 1 0 4600 0 1 15776
box -38 -48 406 592
use scs8hd_mux2_2  mux_left_track_17.mux_l3_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_17.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7268 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 8280 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7084 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_76
timestamp 1586364061
transform 1 0 8096 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_2.mux_l1_in_3_
timestamp 1586364061
transform 1 0 9108 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_80
timestamp 1586364061
transform 1 0 8464 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_84
timestamp 1586364061
transform 1 0 8832 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_96
timestamp 1586364061
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_100
timestamp 1586364061
transform 1 0 10304 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_6.mux_l1_in_3_
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 13064 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 12696 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_128
timestamp 1586364061
transform 1 0 12880 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_6.mux_l2_in_1_
timestamp 1586364061
transform 1 0 14812 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14260 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_141
timestamp 1586364061
transform 1 0 14076 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_145
timestamp 1586364061
transform 1 0 14444 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_158
timestamp 1586364061
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_162
timestamp 1586364061
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_16.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18768 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 18584 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 18216 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_179
timestamp 1586364061
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_188
timestamp 1586364061
transform 1 0 18400 0 1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 20792 0 1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20608 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 19780 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_201
timestamp 1586364061
transform 1 0 19596 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_205
timestamp 1586364061
transform 1 0 19964 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_210
timestamp 1586364061
transform 1 0 20424 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 22908 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_233
timestamp 1586364061
transform 1 0 22540 0 1 15776
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_track_8.mux_l2_in_1_
timestamp 1586364061
transform 1 0 23736 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 23276 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_239
timestamp 1586364061
transform 1 0 23092 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_243
timestamp 1586364061
transform 1 0 23460 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_255
timestamp 1586364061
transform 1 0 24564 0 1 15776
box -38 -48 222 592
use scs8hd_buf_2  _098_
timestamp 1586364061
transform 1 0 25300 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_259
timestamp 1586364061
transform 1 0 24932 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_267
timestamp 1586364061
transform 1 0 25668 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_271
timestamp 1586364061
transform 1 0 26036 0 1 15776
box -38 -48 590 592
use scs8hd_decap_4  FILLER_27_8
timestamp 1586364061
transform 1 0 1840 0 1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 1656 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 1564 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_0.mux_l4_in_0_
timestamp 1586364061
transform 1 0 1748 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_26_16
timestamp 1586364061
transform 1 0 2576 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 2760 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 2208 0 1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 2392 0 1 16864
box -38 -48 1786 592
use scs8hd_decap_3  FILLER_26_28
timestamp 1586364061
transform 1 0 3680 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_24
timestamp 1586364061
transform 1 0 3312 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_20
timestamp 1586364061
transform 1 0 2944 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 3496 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 3128 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_37
timestamp 1586364061
transform 1 0 4508 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_33
timestamp 1586364061
transform 1 0 4140 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 4324 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1786 592
use scs8hd_mux2_2  mux_top_track_36.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4876 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_36.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 5888 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_36.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 5980 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_51
timestamp 1586364061
transform 1 0 5796 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_50
timestamp 1586364061
transform 1 0 5704 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_54
timestamp 1586364061
transform 1 0 6072 0 1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_38.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 6348 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_55
timestamp 1586364061
transform 1 0 6164 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_59
timestamp 1586364061
transform 1 0 6532 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_58
timestamp 1586364061
transform 1 0 6440 0 1 16864
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_38.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1786 592
use scs8hd_mux2_2  mux_top_track_38.mux_l1_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7268 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_38.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7820 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_64
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_26_69
timestamp 1586364061
transform 1 0 7452 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_85
timestamp 1586364061
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_81
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_89
timestamp 1586364061
transform 1 0 9292 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 9108 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 9108 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 9292 0 1 16864
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_26_106
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_112
timestamp 1586364061
transform 1 0 11408 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_108
timestamp 1586364061
transform 1 0 11040 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_110
timestamp 1586364061
transform 1 0 11224 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 11040 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_116
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_119
timestamp 1586364061
transform 1 0 12052 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_116
timestamp 1586364061
transform 1 0 11776 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11868 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_123
timestamp 1586364061
transform 1 0 12420 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12236 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 12512 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_26_137
timestamp 1586364061
transform 1 0 13708 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_133
timestamp 1586364061
transform 1 0 13340 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 13524 0 -1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 12604 0 1 16864
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_27_148
timestamp 1586364061
transform 1 0 14720 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_144
timestamp 1586364061
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_141
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14628 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14260 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13892 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14536 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_149
timestamp 1586364061
transform 1 0 14812 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 14904 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_6.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_top_track_6.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15088 0 1 16864
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 17020 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 17204 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_173
timestamp 1586364061
transform 1 0 17020 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_177
timestamp 1586364061
transform 1 0 17388 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_171
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_175
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_track_24.mux_l1_in_2_
timestamp 1586364061
transform 1 0 17756 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 18768 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 19228 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_194
timestamp 1586364061
transform 1 0 18952 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_179
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_27_207
timestamp 1586364061
transform 1 0 20148 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_203
timestamp 1586364061
transform 1 0 19780 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_203
timestamp 1586364061
transform 1 0 19780 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_199
timestamp 1586364061
transform 1 0 19412 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 19596 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 19964 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_215
timestamp 1586364061
transform 1 0 20884 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 590 592
use scs8hd_decap_3  FILLER_26_211
timestamp 1586364061
transform 1 0 20516 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 21068 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_223
timestamp 1586364061
transform 1 0 21620 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_219
timestamp 1586364061
transform 1 0 21252 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_221
timestamp 1586364061
transform 1 0 21436 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 21436 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21804 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 21528 0 -1 16864
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 21712 0 -1 16864
box -38 -48 866 592
use scs8hd_mux2_2  mux_right_track_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21988 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_236
timestamp 1586364061
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_237
timestamp 1586364061
transform 1 0 22908 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_233
timestamp 1586364061
transform 1 0 22540 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 22724 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 23276 0 -1 16864
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_track_8.mux_l3_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__A0
timestamp 1586364061
transform 1 0 24656 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_240
timestamp 1586364061
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_254
timestamp 1586364061
transform 1 0 24472 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_265
timestamp 1586364061
transform 1 0 25484 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_258
timestamp 1586364061
transform 1 0 24840 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_264
timestamp 1586364061
transform 1 0 25392 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_260
timestamp 1586364061
transform 1 0 25024 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 25208 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__A1
timestamp 1586364061
transform 1 0 25024 0 1 16864
box -38 -48 222 592
use scs8hd_conb_1  _033_
timestamp 1586364061
transform 1 0 25208 0 1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_26_272
timestamp 1586364061
transform 1 0 26128 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__S
timestamp 1586364061
transform 1 0 25668 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 1656 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 2668 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_19
timestamp 1586364061
transform 1 0 2852 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 3036 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_36.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4232 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_39
timestamp 1586364061
transform 1 0 4692 0 -1 17952
box -38 -48 222 592
use scs8hd_conb_1  _048_
timestamp 1586364061
transform 1 0 4416 0 -1 17952
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_36.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 5428 0 -1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4876 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 5244 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_43
timestamp 1586364061
transform 1 0 5060 0 -1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 7636 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_66
timestamp 1586364061
transform 1 0 7176 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_70
timestamp 1586364061
transform 1 0 7544 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_73
timestamp 1586364061
transform 1 0 7820 0 -1 17952
box -38 -48 222 592
use scs8hd_conb_1  _040_
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10120 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 9292 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_84
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_88
timestamp 1586364061
transform 1 0 9200 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_91
timestamp 1586364061
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_96
timestamp 1586364061
transform 1 0 9936 0 -1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_100
timestamp 1586364061
transform 1 0 10304 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_104
timestamp 1586364061
transform 1 0 10672 0 -1 17952
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_6.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 13248 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 12696 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_124
timestamp 1586364061
transform 1 0 12512 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_128
timestamp 1586364061
transform 1 0 12880 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_134
timestamp 1586364061
transform 1 0 13432 0 -1 17952
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 14812 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_151
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_6.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 16652 0 -1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16008 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_160
timestamp 1586364061
transform 1 0 15824 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_164
timestamp 1586364061
transform 1 0 16192 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_168
timestamp 1586364061
transform 1 0 16560 0 -1 17952
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_8.mux_l2_in_3_
timestamp 1586364061
transform 1 0 19228 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_188
timestamp 1586364061
transform 1 0 18400 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_28_196
timestamp 1586364061
transform 1 0 19136 0 -1 17952
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_206
timestamp 1586364061
transform 1 0 20056 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_4  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 22172 0 -1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 21252 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_221
timestamp 1586364061
transform 1 0 21436 0 -1 17952
box -38 -48 590 592
use scs8hd_mux2_2  mux_right_track_4.mux_l1_in_5_
timestamp 1586364061
transform 1 0 24656 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A1
timestamp 1586364061
transform 1 0 24104 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 24472 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_248
timestamp 1586364061
transform 1 0 23920 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_252
timestamp 1586364061
transform 1 0 24288 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_265
timestamp 1586364061
transform 1 0 25484 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_273
timestamp 1586364061
transform 1 0 26220 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 1564 0 1 17952
box -38 -48 1786 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_36.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4232 0 1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_36.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 3496 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_24
timestamp 1586364061
transform 1 0 3312 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_28
timestamp 1586364061
transform 1 0 3680 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6256 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_58
timestamp 1586364061
transform 1 0 6440 0 1 17952
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 7452 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6992 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_66
timestamp 1586364061
transform 1 0 7176 0 1 17952
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_2.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 9936 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9568 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_90
timestamp 1586364061
transform 1 0 9384 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_94
timestamp 1586364061
transform 1 0 9752 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 11132 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 11868 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 11500 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_107
timestamp 1586364061
transform 1 0 10948 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_111
timestamp 1586364061
transform 1 0 11316 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_115
timestamp 1586364061
transform 1 0 11684 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_119
timestamp 1586364061
transform 1 0 12052 0 1 17952
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_6.mux_l1_in_1_
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13064 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12696 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_128
timestamp 1586364061
transform 1 0 12880 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_6.mux_l3_in_0_
timestamp 1586364061
transform 1 0 14812 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 14260 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_141
timestamp 1586364061
transform 1 0 14076 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_145
timestamp 1586364061
transform 1 0 14444 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_158
timestamp 1586364061
transform 1 0 15640 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_8.mux_l2_in_1_
timestamp 1586364061
transform 1 0 16376 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 16192 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 15824 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_162
timestamp 1586364061
transform 1 0 16008 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_175
timestamp 1586364061
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 19320 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 18216 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 18584 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_179
timestamp 1586364061
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_188
timestamp 1586364061
transform 1 0 18400 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_192
timestamp 1586364061
transform 1 0 18768 0 1 17952
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 19504 0 1 17952
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_track_4.mux_l2_in_3_
timestamp 1586364061
transform 1 0 21988 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 21804 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 21436 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_219
timestamp 1586364061
transform 1 0 21252 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_223
timestamp 1586364061
transform 1 0 21620 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_236
timestamp 1586364061
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_4.mux_l1_in_6_
timestamp 1586364061
transform 1 0 24012 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A0
timestamp 1586364061
transform 1 0 23828 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__S
timestamp 1586364061
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_240
timestamp 1586364061
transform 1 0 23184 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 25024 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 25392 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 25760 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_258
timestamp 1586364061
transform 1 0 24840 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_262
timestamp 1586364061
transform 1 0 25208 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_266
timestamp 1586364061
transform 1 0 25576 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_270
timestamp 1586364061
transform 1 0 25944 0 1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_29_276
timestamp 1586364061
transform 1 0 26496 0 1 17952
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_34.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2300 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 1564 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 1932 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_7
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_11
timestamp 1586364061
transform 1 0 2116 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_26
timestamp 1586364061
transform 1 0 3496 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_22
timestamp 1586364061
transform 1 0 3128 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3680 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_34.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3312 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_36
timestamp 1586364061
transform 1 0 4416 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_30
timestamp 1586364061
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_34.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 4232 0 -1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_36.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4692 0 -1 19040
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 5704 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 6072 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_48
timestamp 1586364061
transform 1 0 5520 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_52
timestamp 1586364061
transform 1 0 5888 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 8188 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_75
timestamp 1586364061
transform 1 0 8004 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_79
timestamp 1586364061
transform 1 0 8372 0 -1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 10120 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 8556 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 8924 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_83
timestamp 1586364061
transform 1 0 8740 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_87
timestamp 1586364061
transform 1 0 9108 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_97
timestamp 1586364061
transform 1 0 10028 0 -1 19040
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_4.mux_l1_in_1_
timestamp 1586364061
transform 1 0 10304 0 -1 19040
box -38 -48 866 592
use scs8hd_mux2_2  mux_top_track_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11316 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11684 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_109
timestamp 1586364061
transform 1 0 11132 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_113
timestamp 1586364061
transform 1 0 11500 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13432 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12880 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 13248 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_126
timestamp 1586364061
transform 1 0 12696 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_130
timestamp 1586364061
transform 1 0 13064 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15640 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 15456 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14812 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_143
timestamp 1586364061
transform 1 0 14260 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_147
timestamp 1586364061
transform 1 0 14628 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_151
timestamp 1586364061
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 17204 0 -1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17020 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 16652 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_167
timestamp 1586364061
transform 1 0 16468 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_171
timestamp 1586364061
transform 1 0 16836 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_194
timestamp 1586364061
transform 1 0 18952 0 -1 19040
box -38 -48 590 592
use scs8hd_conb_1  _052_
timestamp 1586364061
transform 1 0 19780 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 19504 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 21068 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_206
timestamp 1586364061
transform 1 0 20056 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 222 592
use scs8hd_buf_2  _109_
timestamp 1586364061
transform 1 0 21252 0 -1 19040
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 22356 0 -1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_223
timestamp 1586364061
transform 1 0 21620 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_30_229
timestamp 1586364061
transform 1 0 22172 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 24288 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_250
timestamp 1586364061
transform 1 0 24104 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_254
timestamp 1586364061
transform 1 0 24472 0 -1 19040
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_track_4.mux_l1_in_4_
timestamp 1586364061
transform 1 0 24840 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_267
timestamp 1586364061
transform 1 0 25668 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_34.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 2116 0 1 19040
box -38 -48 1786 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_34.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 1564 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_7
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4600 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_34.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4048 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_30
timestamp 1586364061
transform 1 0 3864 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_34
timestamp 1586364061
transform 1 0 4232 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 5612 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_47
timestamp 1586364061
transform 1 0 5428 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_25.mux_l1_in_2_
timestamp 1586364061
transform 1 0 7452 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 7268 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_66
timestamp 1586364061
transform 1 0 7176 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_78
timestamp 1586364061
transform 1 0 8280 0 1 19040
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 9108 0 1 19040
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9844 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 8464 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 8832 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_82
timestamp 1586364061
transform 1 0 8648 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_93
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_97
timestamp 1586364061
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_20.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10396 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11408 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_18.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_132
timestamp 1586364061
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_136
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_18.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 14352 0 1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_18.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14168 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_140
timestamp 1586364061
transform 1 0 13984 0 1 19040
box -38 -48 222 592
use scs8hd_conb_1  _038_
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 16284 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 16652 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17296 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_163
timestamp 1586364061
transform 1 0 16100 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_167
timestamp 1586364061
transform 1 0 16468 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_174
timestamp 1586364061
transform 1 0 17112 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_178
timestamp 1586364061
transform 1 0 17480 0 1 19040
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_track_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18492 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 18308 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_198
timestamp 1586364061
transform 1 0 19320 0 1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 20056 0 1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 19872 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 19504 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_202
timestamp 1586364061
transform 1 0 19688 0 1 19040
box -38 -48 222 592
use scs8hd_conb_1  _065_
timestamp 1586364061
transform 1 0 22540 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 22356 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23000 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_225
timestamp 1586364061
transform 1 0 21804 0 1 19040
box -38 -48 590 592
use scs8hd_fill_2  FILLER_31_236
timestamp 1586364061
transform 1 0 22816 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_4.mux_l2_in_2_
timestamp 1586364061
transform 1 0 24196 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 24012 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_240
timestamp 1586364061
transform 1 0 23184 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 25208 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 25576 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 25944 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_260
timestamp 1586364061
transform 1 0 25024 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_264
timestamp 1586364061
transform 1 0 25392 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_268
timestamp 1586364061
transform 1 0 25760 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_272
timestamp 1586364061
transform 1 0 26128 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_276
timestamp 1586364061
transform 1 0 26496 0 1 19040
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_34.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 1656 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 2024 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_8
timestamp 1586364061
transform 1 0 1840 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_12
timestamp 1586364061
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_34.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3404 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use scs8hd_buf_4  mux_left_track_25.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 6532 0 -1 20128
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 5980 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6348 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_51
timestamp 1586364061
transform 1 0 5796 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_55
timestamp 1586364061
transform 1 0 6164 0 -1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_25.mux_l1_in_1_
timestamp 1586364061
transform 1 0 7820 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 7452 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_65
timestamp 1586364061
transform 1 0 7084 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_71
timestamp 1586364061
transform 1 0 7636 0 -1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_20.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9844 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 9108 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_82
timestamp 1586364061
transform 1 0 8648 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_86
timestamp 1586364061
transform 1 0 9016 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_32_89
timestamp 1586364061
transform 1 0 9292 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_97
timestamp 1586364061
transform 1 0 10028 0 -1 20128
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_20.mux_l1_in_1_
timestamp 1586364061
transform 1 0 10304 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_20.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11316 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_109
timestamp 1586364061
transform 1 0 11132 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_113
timestamp 1586364061
transform 1 0 11500 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_119
timestamp 1586364061
transform 1 0 12052 0 -1 20128
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12328 0 -1 20128
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12144 0 -1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_6.mux_l1_in_2_
timestamp 1586364061
transform 1 0 15548 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 14628 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_141
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_32_149
timestamp 1586364061
transform 1 0 14812 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_14.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 17112 0 -1 20128
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 16928 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16560 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_170
timestamp 1586364061
transform 1 0 16744 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 19044 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_193
timestamp 1586364061
transform 1 0 18860 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_197
timestamp 1586364061
transform 1 0 19228 0 -1 20128
box -38 -48 406 592
use scs8hd_conb_1  _037_
timestamp 1586364061
transform 1 0 19596 0 -1 20128
box -38 -48 314 592
use scs8hd_buf_2  _111_
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 20056 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 20424 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_204
timestamp 1586364061
transform 1 0 19872 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_208
timestamp 1586364061
transform 1 0 20240 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_212
timestamp 1586364061
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 22356 0 -1 20128
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 21436 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 22172 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_219
timestamp 1586364061
transform 1 0 21252 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_223
timestamp 1586364061
transform 1 0 21620 0 -1 20128
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 24288 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 24656 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_250
timestamp 1586364061
transform 1 0 24104 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_254
timestamp 1586364061
transform 1 0 24472 0 -1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_4.mux_l4_in_0_
timestamp 1586364061
transform 1 0 24840 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_267
timestamp 1586364061
transform 1 0 25668 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 1656 0 1 20128
box -38 -48 1786 592
use scs8hd_mux2_2  mux_top_track_32.mux_l2_in_0_
timestamp 1586364061
transform 1 0 1564 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 2576 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_14
timestamp 1586364061
transform 1 0 2392 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_18
timestamp 1586364061
transform 1 0 2760 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_22
timestamp 1586364061
transform 1 0 3128 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 2944 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_26
timestamp 1586364061
transform 1 0 3496 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_25
timestamp 1586364061
transform 1 0 3404 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 3312 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_30
timestamp 1586364061
transform 1 0 3864 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_29
timestamp 1586364061
transform 1 0 3772 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3956 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3680 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_35
timestamp 1586364061
transform 1 0 4324 0 -1 21216
box -38 -48 222 592
use scs8hd_conb_1  _047_
timestamp 1586364061
transform 1 0 4140 0 1 20128
box -38 -48 314 592
use scs8hd_conb_1  _046_
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_39
timestamp 1586364061
transform 1 0 4692 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_36
timestamp 1586364061
transform 1 0 4416 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 4508 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 4600 0 1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 5060 0 -1 21216
box -38 -48 1786 592
use scs8hd_mux2_2  mux_left_track_25.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 4968 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 4876 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_40
timestamp 1586364061
transform 1 0 4784 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_53
timestamp 1586364061
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_57
timestamp 1586364061
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_62
timestamp 1586364061
transform 1 0 6808 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_4  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7176 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7176 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_72
timestamp 1586364061
transform 1 0 7728 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 7544 0 -1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_25.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7820 0 -1 21216
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7360 0 1 20128
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_34_82
timestamp 1586364061
transform 1 0 8648 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_87
timestamp 1586364061
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9292 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_97
timestamp 1586364061
transform 1 0 10028 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_90
timestamp 1586364061
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_91
timestamp 1586364061
transform 1 0 9476 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_20.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 10212 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 9844 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_20.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9660 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_20.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9844 0 1 20128
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_top_track_20.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10580 0 -1 21216
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_114
timestamp 1586364061
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_118
timestamp 1586364061
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_101
timestamp 1586364061
transform 1 0 10396 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_126
timestamp 1586364061
transform 1 0 12696 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_122
timestamp 1586364061
transform 1 0 12328 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12880 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12512 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_conb_1  _039_
timestamp 1586364061
transform 1 0 12696 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_133
timestamp 1586364061
transform 1 0 13340 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_129
timestamp 1586364061
transform 1 0 12972 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 13156 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_18.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_2.mux_l1_in_1_
timestamp 1586364061
transform 1 0 13064 0 -1 21216
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_top_track_18.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13708 0 1 20128
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_34_147
timestamp 1586364061
transform 1 0 14628 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_143
timestamp 1586364061
transform 1 0 14260 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_139
timestamp 1586364061
transform 1 0 13892 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14444 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_18.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_156
timestamp 1586364061
transform 1 0 15456 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 15640 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_18.mux_l1_in_1_
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_4  FILLER_34_167
timestamp 1586364061
transform 1 0 16468 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_163
timestamp 1586364061
transform 1 0 16100 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_160
timestamp 1586364061
transform 1 0 15824 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16284 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16008 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_6.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16192 0 1 20128
box -38 -48 866 592
use scs8hd_fill_1  FILLER_34_173
timestamp 1586364061
transform 1 0 17020 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_177
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_173
timestamp 1586364061
transform 1 0 17020 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 16836 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_14.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 17112 0 -1 21216
box -38 -48 1786 592
use scs8hd_mux2_2  mux_top_track_8.mux_l3_in_0_
timestamp 1586364061
transform 1 0 18216 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 19228 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 19044 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_195
timestamp 1586364061
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_193
timestamp 1586364061
transform 1 0 18860 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_197
timestamp 1586364061
transform 1 0 19228 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_205
timestamp 1586364061
transform 1 0 19964 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_199
timestamp 1586364061
transform 1 0 19412 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 19412 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 19596 0 1 20128
box -38 -48 222 592
use scs8hd_buf_2  _117_
timestamp 1586364061
transform 1 0 19596 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_212
timestamp 1586364061
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_209
timestamp 1586364061
transform 1 0 20332 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 20424 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_10.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_top_track_10.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19780 0 1 20128
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_33_222
timestamp 1586364061
transform 1 0 21528 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_226
timestamp 1586364061
transform 1 0 21896 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 21712 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_230
timestamp 1586364061
transform 1 0 22264 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 22080 0 1 20128
box -38 -48 222 592
use scs8hd_buf_2  _107_
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_234
timestamp 1586364061
transform 1 0 22632 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_236
timestamp 1586364061
transform 1 0 22816 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 22816 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_238
timestamp 1586364061
transform 1 0 23000 0 -1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 23000 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_242
timestamp 1586364061
transform 1 0 23368 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_240
timestamp 1586364061
transform 1 0 23184 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 23460 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_4.mux_l3_in_1_
timestamp 1586364061
transform 1 0 23644 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_254
timestamp 1586364061
transform 1 0 24472 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 24656 0 -1 21216
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 23920 0 1 20128
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_34_266
timestamp 1586364061
transform 1 0 25576 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_258
timestamp 1586364061
transform 1 0 24840 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 25024 0 -1 21216
box -38 -48 222 592
use scs8hd_buf_2  _108_
timestamp 1586364061
transform 1 0 25208 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_274
timestamp 1586364061
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_33_271
timestamp 1586364061
transform 1 0 26036 0 1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_267
timestamp 1586364061
transform 1 0 25668 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_32.mux_l1_in_0_
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 866 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 2392 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 2760 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_12
timestamp 1586364061
transform 1 0 2208 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_16
timestamp 1586364061
transform 1 0 2576 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2944 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3956 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 4600 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_29
timestamp 1586364061
transform 1 0 3772 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_33
timestamp 1586364061
transform 1 0 4140 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_37
timestamp 1586364061
transform 1 0 4508 0 1 21216
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_25.mux_l3_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 4968 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_40
timestamp 1586364061
transform 1 0 4784 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_53
timestamp 1586364061
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_57
timestamp 1586364061
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_33.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_conb_1  _041_
timestamp 1586364061
transform 1 0 9476 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 9936 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 8740 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 9108 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_81
timestamp 1586364061
transform 1 0 8556 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_85
timestamp 1586364061
transform 1 0 8924 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_89
timestamp 1586364061
transform 1 0 9292 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_94
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_20.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10488 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 10304 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_22.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_111
timestamp 1586364061
transform 1 0 11316 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_115
timestamp 1586364061
transform 1 0 11684 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_16.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_22.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_132
timestamp 1586364061
transform 1 0 13248 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_136
timestamp 1586364061
transform 1 0 13616 0 1 21216
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_18.mux_l2_in_0_
timestamp 1586364061
transform 1 0 14076 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 15272 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 15640 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13892 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_150
timestamp 1586364061
transform 1 0 14904 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_156
timestamp 1586364061
transform 1 0 15456 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_14.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16192 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_160
timestamp 1586364061
transform 1 0 15824 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_175
timestamp 1586364061
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_10.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18860 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 18676 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 18308 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_179
timestamp 1586364061
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_189
timestamp 1586364061
transform 1 0 18492 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 20424 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 19872 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_202
timestamp 1586364061
transform 1 0 19688 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_206
timestamp 1586364061
transform 1 0 20056 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 21988 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 23000 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 21804 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 21436 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_219
timestamp 1586364061
transform 1 0 21252 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_223
timestamp 1586364061
transform 1 0 21620 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_236
timestamp 1586364061
transform 1 0 22816 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_4.mux_l1_in_3_
timestamp 1586364061
transform 1 0 24564 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 23828 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 24380 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_240
timestamp 1586364061
transform 1 0 23184 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_249
timestamp 1586364061
transform 1 0 24012 0 1 21216
box -38 -48 406 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_264
timestamp 1586364061
transform 1 0 25392 0 1 21216
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_35_276
timestamp 1586364061
transform 1 0 26496 0 1 21216
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 1472 0 -1 22304
box -38 -48 1786 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 130 592
use scs8hd_buf_4  mux_top_track_34.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 4324 0 -1 22304
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_30.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_23
timestamp 1586364061
transform 1 0 3220 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_25.mux_l2_in_1_
timestamp 1586364061
transform 1 0 5980 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 5796 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 5060 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 5428 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_41
timestamp 1586364061
transform 1 0 4876 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_45
timestamp 1586364061
transform 1 0 5244 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_49
timestamp 1586364061
transform 1 0 5612 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_25.mux_l1_in_3_
timestamp 1586364061
transform 1 0 7544 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 6992 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_62
timestamp 1586364061
transform 1 0 6808 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_66
timestamp 1586364061
transform 1 0 7176 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_79
timestamp 1586364061
transform 1 0 8372 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_33.mux_l1_in_2_
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 8556 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 8924 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_83
timestamp 1586364061
transform 1 0 8740 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_87
timestamp 1586364061
transform 1 0 9108 0 -1 22304
box -38 -48 314 592
use scs8hd_conb_1  _042_
timestamp 1586364061
transform 1 0 11224 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10672 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12052 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11040 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11684 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_102
timestamp 1586364061
transform 1 0 10488 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_106
timestamp 1586364061
transform 1 0 10856 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_113
timestamp 1586364061
transform 1 0 11500 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_22.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12236 0 -1 22304
box -38 -48 1786 592
use scs8hd_mux2_2  mux_top_track_16.mux_l1_in_1_
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 14168 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14536 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14904 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_140
timestamp 1586364061
transform 1 0 13984 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_144
timestamp 1586364061
transform 1 0 14352 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_148
timestamp 1586364061
transform 1 0 14720 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_152
timestamp 1586364061
transform 1 0 15088 0 -1 22304
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_12.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16836 0 -1 22304
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 16652 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16284 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_163
timestamp 1586364061
transform 1 0 16100 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_167
timestamp 1586364061
transform 1 0 16468 0 -1 22304
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_10.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 19320 0 -1 22304
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18860 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_36_195
timestamp 1586364061
transform 1 0 19044 0 -1 22304
box -38 -48 314 592
use scs8hd_buf_2  _118_
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 20424 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 20056 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_204
timestamp 1586364061
transform 1 0 19872 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_208
timestamp 1586364061
transform 1 0 20240 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_212
timestamp 1586364061
transform 1 0 20608 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_4.mux_l1_in_2_
timestamp 1586364061
transform 1 0 22264 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 21436 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_219
timestamp 1586364061
transform 1 0 21252 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_223
timestamp 1586364061
transform 1 0 21620 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_229
timestamp 1586364061
transform 1 0 22172 0 -1 22304
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 23828 0 -1 22304
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 23368 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_36_244
timestamp 1586364061
transform 1 0 23552 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_266
timestamp 1586364061
transform 1 0 25576 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_1  FILLER_36_274
timestamp 1586364061
transform 1 0 26312 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_30.mux_l1_in_0_
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 866 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 2392 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_30.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 2760 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_12
timestamp 1586364061
transform 1 0 2208 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_16
timestamp 1586364061
transform 1 0 2576 0 1 22304
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 2944 0 1 22304
box -38 -48 590 592
use scs8hd_mux2_2  mux_top_track_28.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4324 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_28.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4140 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 3680 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_26
timestamp 1586364061
transform 1 0 3496 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_30
timestamp 1586364061
transform 1 0 3864 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 5336 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_28.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 5704 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 6072 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 6440 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_44
timestamp 1586364061
transform 1 0 5152 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_48
timestamp 1586364061
transform 1 0 5520 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_52
timestamp 1586364061
transform 1 0 5888 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_56
timestamp 1586364061
transform 1 0 6256 0 1 22304
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_33.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 8188 0 1 22304
box -38 -48 1786 592
use scs8hd_buf_4  mux_top_track_32.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 7636 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_60
timestamp 1586364061
transform 1 0 6624 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_37_68
timestamp 1586364061
transform 1 0 7360 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_73
timestamp 1586364061
transform 1 0 7820 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10212 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_96
timestamp 1586364061
transform 1 0 9936 0 1 22304
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_24.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 10580 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_101
timestamp 1586364061
transform 1 0 10396 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_114
timestamp 1586364061
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_118
timestamp 1586364061
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_24.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13800 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13432 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_132
timestamp 1586364061
transform 1 0 13248 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_136
timestamp 1586364061
transform 1 0 13616 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_22.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13984 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 15640 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14996 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_149
timestamp 1586364061
transform 1 0 14812 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_153
timestamp 1586364061
transform 1 0 15180 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_157
timestamp 1586364061
transform 1 0 15548 0 1 22304
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_12.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16192 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16008 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_160
timestamp 1586364061
transform 1 0 15824 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_173
timestamp 1586364061
transform 1 0 17020 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_177
timestamp 1586364061
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_10.mux_l3_in_0_
timestamp 1586364061
transform 1 0 18676 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 18492 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 17572 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_181
timestamp 1586364061
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_188
timestamp 1586364061
transform 1 0 18400 0 1 22304
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_12.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 19688 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20056 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_200
timestamp 1586364061
transform 1 0 19504 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_204
timestamp 1586364061
transform 1 0 19872 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 22172 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 23000 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_227
timestamp 1586364061
transform 1 0 21988 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_231
timestamp 1586364061
transform 1 0 22356 0 1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_37_237
timestamp 1586364061
transform 1 0 22908 0 1 22304
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 24012 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 23828 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_240
timestamp 1586364061
transform 1 0 23184 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 222 592
use scs8hd_conb_1  _035_
timestamp 1586364061
transform 1 0 25576 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 25024 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 25392 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_258
timestamp 1586364061
transform 1 0 24840 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_262
timestamp 1586364061
transform 1 0 25208 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_top_track_30.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 1472 0 -1 23392
box -38 -48 1786 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_28.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4416 0 -1 23392
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_28.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4232 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_23
timestamp 1586364061
transform 1 0 3220 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_55
timestamp 1586364061
transform 1 0 6164 0 -1 23392
box -38 -48 590 592
use scs8hd_conb_1  _057_
timestamp 1586364061
transform 1 0 6992 0 -1 23392
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_33.mux_l1_in_1_
timestamp 1586364061
transform 1 0 8004 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 7452 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 7820 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 6808 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_61
timestamp 1586364061
transform 1 0 6716 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_67
timestamp 1586364061
transform 1 0 7268 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_71
timestamp 1586364061
transform 1 0 7636 0 -1 23392
box -38 -48 222 592
use scs8hd_conb_1  _055_
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10120 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9384 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_84
timestamp 1586364061
transform 1 0 8832 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_38_96
timestamp 1586364061
transform 1 0 9936 0 -1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10856 0 -1 23392
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10488 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_100
timestamp 1586364061
transform 1 0 10304 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_104
timestamp 1586364061
transform 1 0 10672 0 -1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_22.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 13432 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_22.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 13064 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_125
timestamp 1586364061
transform 1 0 12604 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_132
timestamp 1586364061
transform 1 0 13248 0 -1 23392
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_6.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15456 0 -1 23392
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14628 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14996 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_145
timestamp 1586364061
transform 1 0 14444 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_149
timestamp 1586364061
transform 1 0 14812 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_12.mux_l1_in_1_
timestamp 1586364061
transform 1 0 16744 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16192 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16560 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_162
timestamp 1586364061
transform 1 0 16008 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_166
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_10.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19228 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 18032 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 18676 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 19044 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_179
timestamp 1586364061
transform 1 0 17572 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_183
timestamp 1586364061
transform 1 0 17940 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_186
timestamp 1586364061
transform 1 0 18216 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_193
timestamp 1586364061
transform 1 0 18860 0 -1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_10.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 20240 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_206
timestamp 1586364061
transform 1 0 20056 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_210
timestamp 1586364061
transform 1 0 20424 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_38_234
timestamp 1586364061
transform 1 0 22632 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_238
timestamp 1586364061
transform 1 0 23000 0 -1 23392
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 23368 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 24380 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 24748 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_241
timestamp 1586364061
transform 1 0 23276 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_255
timestamp 1586364061
transform 1 0 24564 0 -1 23392
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_38.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 24932 0 -1 23392
box -38 -48 590 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_265
timestamp 1586364061
transform 1 0 25484 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_38_273
timestamp 1586364061
transform 1 0 26220 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 1786 592
use scs8hd_mux2_2  mux_top_track_30.mux_l2_in_0_
timestamp 1586364061
transform 1 0 1472 0 -1 24480
box -38 -48 866 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 2852 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_40_13
timestamp 1586364061
transform 1 0 2300 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_17
timestamp 1586364061
transform 1 0 2668 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_29
timestamp 1586364061
transform 1 0 3772 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_21
timestamp 1586364061
transform 1 0 3036 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_26
timestamp 1586364061
transform 1 0 3496 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_22
timestamp 1586364061
transform 1 0 3128 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3680 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3312 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_36
timestamp 1586364061
transform 1 0 4416 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_30
timestamp 1586364061
transform 1 0 3864 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_28.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4232 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_30.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4048 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_28.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4232 0 1 23392
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_top_track_30.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4876 0 -1 24480
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_30.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_53
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_57
timestamp 1586364061
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_40
timestamp 1586364061
transform 1 0 4784 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_6  FILLER_40_60
timestamp 1586364061
transform 1 0 6624 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_39_66
timestamp 1586364061
transform 1 0 7176 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 7176 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 7268 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_33.mux_l3_in_0_
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_77
timestamp 1586364061
transform 1 0 8188 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 8372 0 -1 24480
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_33.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7452 0 1 23392
box -38 -48 1786 592
use scs8hd_decap_3  FILLER_40_89
timestamp 1586364061
transform 1 0 9292 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_81
timestamp 1586364061
transform 1 0 8556 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_88
timestamp 1586364061
transform 1 0 9200 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_92
timestamp 1586364061
transform 1 0 9568 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9752 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_mux2_2  mux_left_track_33.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9936 0 1 23392
box -38 -48 866 592
use scs8hd_conb_1  _043_
timestamp 1586364061
transform 1 0 10028 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_1  FILLER_40_107
timestamp 1586364061
transform 1 0 10948 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_104
timestamp 1586364061
transform 1 0 10672 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_100
timestamp 1586364061
transform 1 0 10304 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_3  FILLER_39_105
timestamp 1586364061
transform 1 0 10764 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11040 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_114
timestamp 1586364061
transform 1 0 11592 0 1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11408 0 1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 11040 0 -1 24480
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_40_127
timestamp 1586364061
transform 1 0 12788 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_128
timestamp 1586364061
transform 1 0 12880 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_buf_2  _125_
timestamp 1586364061
transform 1 0 12512 0 1 23392
box -38 -48 406 592
use scs8hd_decap_3  FILLER_40_131
timestamp 1586364061
transform 1 0 13156 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_132
timestamp 1586364061
transform 1 0 13248 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 13432 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_22.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13064 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 13432 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_22.mux_l1_in_1_
timestamp 1586364061
transform 1 0 13616 0 -1 24480
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_top_track_22.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 13616 0 1 23392
box -38 -48 1786 592
use scs8hd_buf_4  mux_top_track_16.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15548 0 -1 24480
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 14628 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_155
timestamp 1586364061
transform 1 0 15364 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_145
timestamp 1586364061
transform 1 0 14444 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_149
timestamp 1586364061
transform 1 0 14812 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_3  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_168
timestamp 1586364061
transform 1 0 16560 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_163
timestamp 1586364061
transform 1 0 16100 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_162
timestamp 1586364061
transform 1 0 16008 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_159
timestamp 1586364061
transform 1 0 15732 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 15824 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 16192 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_12.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_39_175
timestamp 1586364061
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 16744 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_14.mux_l1_in_1_
timestamp 1586364061
transform 1 0 16928 0 -1 24480
box -38 -48 866 592
use scs8hd_decap_3  FILLER_40_186
timestamp 1586364061
transform 1 0 18216 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_40_181
timestamp 1586364061
transform 1 0 17756 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_179
timestamp 1586364061
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 18032 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_14.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 866 592
use scs8hd_decap_4  FILLER_40_195
timestamp 1586364061
transform 1 0 19044 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_197
timestamp 1586364061
transform 1 0 19228 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_193
timestamp 1586364061
transform 1 0 18860 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 19044 0 1 23392
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18492 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_40_206
timestamp 1586364061
transform 1 0 20056 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_201
timestamp 1586364061
transform 1 0 19596 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_201
timestamp 1586364061
transform 1 0 19596 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 19412 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 20240 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 19412 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 19780 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_10.mux_l2_in_1_
timestamp 1586364061
transform 1 0 19964 0 1 23392
box -38 -48 866 592
use scs8hd_conb_1  _036_
timestamp 1586364061
transform 1 0 19780 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_4  FILLER_40_210
timestamp 1586364061
transform 1 0 20424 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_3  FILLER_39_214
timestamp 1586364061
transform 1 0 20792 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 21068 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_40_223
timestamp 1586364061
transform 1 0 21620 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_223
timestamp 1586364061
transform 1 0 21620 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_219
timestamp 1586364061
transform 1 0 21252 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 21436 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 21804 0 1 23392
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_36.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 21804 0 -1 24480
box -38 -48 590 592
use scs8hd_mux2_2  mux_right_track_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 21988 0 1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_235
timestamp 1586364061
transform 1 0 22724 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_231
timestamp 1586364061
transform 1 0 22356 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_236
timestamp 1586364061
transform 1 0 22816 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22540 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 22908 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_39_241
timestamp 1586364061
transform 1 0 23276 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 23092 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_4.mux_l1_in_1_
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 866 592
use scs8hd_decap_4  FILLER_40_252
timestamp 1586364061
transform 1 0 24288 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_248
timestamp 1586364061
transform 1 0 23920 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 24104 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23920 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _113_
timestamp 1586364061
transform 1 0 24656 0 -1 24480
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 24104 0 1 23392
box -38 -48 1786 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_269
timestamp 1586364061
transform 1 0 25852 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_260
timestamp 1586364061
transform 1 0 25024 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_40_272
timestamp 1586364061
transform 1 0 26128 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_buf_4  mux_top_track_30.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 2116 0 1 24480
box -38 -48 590 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 1564 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 1932 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2852 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_7
timestamp 1586364061
transform 1 0 1748 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_17
timestamp 1586364061
transform 1 0 2668 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_28.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4048 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 3864 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 3496 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_21
timestamp 1586364061
transform 1 0 3036 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_25
timestamp 1586364061
transform 1 0 3404 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_28
timestamp 1586364061
transform 1 0 3680 0 1 24480
box -38 -48 222 592
use scs8hd_conb_1  _044_
timestamp 1586364061
transform 1 0 5612 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 5060 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_41
timestamp 1586364061
transform 1 0 4876 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_45
timestamp 1586364061
transform 1 0 5244 0 1 24480
box -38 -48 406 592
use scs8hd_decap_8  FILLER_41_52
timestamp 1586364061
transform 1 0 5888 0 1 24480
box -38 -48 774 592
use scs8hd_mux2_2  mux_left_track_33.mux_l2_in_1_
timestamp 1586364061
transform 1 0 7636 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7452 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7084 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_60
timestamp 1586364061
transform 1 0 6624 0 1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_67
timestamp 1586364061
transform 1 0 7268 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 8648 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 10212 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_80
timestamp 1586364061
transform 1 0 8464 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_84
timestamp 1586364061
transform 1 0 8832 0 1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_41_88
timestamp 1586364061
transform 1 0 9200 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  FILLER_41_96
timestamp 1586364061
transform 1 0 9936 0 1 24480
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_24.mux_l1_in_1_
timestamp 1586364061
transform 1 0 10764 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 10580 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_101
timestamp 1586364061
transform 1 0 10396 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_114
timestamp 1586364061
transform 1 0 11592 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_118
timestamp 1586364061
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_16.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13616 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_132
timestamp 1586364061
transform 1 0 13248 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_138
timestamp 1586364061
transform 1 0 13800 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_18.mux_l1_in_0_
timestamp 1586364061
transform 1 0 14168 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13984 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 15548 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 15180 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_151
timestamp 1586364061
transform 1 0 14996 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_155
timestamp 1586364061
transform 1 0 15364 0 1 24480
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_18.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 16928 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 16468 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_165
timestamp 1586364061
transform 1 0 16284 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_169
timestamp 1586364061
transform 1 0 16652 0 1 24480
box -38 -48 314 592
use scs8hd_decap_6  FILLER_41_174
timestamp 1586364061
transform 1 0 17112 0 1 24480
box -38 -48 590 592
use scs8hd_buf_4  mux_top_track_12.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 590 592
use scs8hd_buf_4  mux_top_track_24.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 19320 0 1 24480
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 18768 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_180
timestamp 1586364061
transform 1 0 17664 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_190
timestamp 1586364061
transform 1 0 18584 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_194
timestamp 1586364061
transform 1 0 18952 0 1 24480
box -38 -48 222 592
use scs8hd_buf_2  _120_
timestamp 1586364061
transform 1 0 20608 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 21160 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20056 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_204
timestamp 1586364061
transform 1 0 19872 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_216
timestamp 1586364061
transform 1 0 20976 0 1 24480
box -38 -48 222 592
use scs8hd_buf_2  _119_
timestamp 1586364061
transform 1 0 21712 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 22264 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 21528 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 22632 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_228
timestamp 1586364061
transform 1 0 22080 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_41_236
timestamp 1586364061
transform 1 0 22816 0 1 24480
box -38 -48 590 592
use scs8hd_buf_2  _110_
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 406 592
use scs8hd_buf_2  _114_
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 24196 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 23368 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_249
timestamp 1586364061
transform 1 0 24012 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_253
timestamp 1586364061
transform 1 0 24380 0 1 24480
box -38 -48 406 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 25300 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 25668 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_261
timestamp 1586364061
transform 1 0 25116 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_265
timestamp 1586364061
transform 1 0 25484 0 1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_conb_1  _045_
timestamp 1586364061
transform 1 0 1656 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_3  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_9
timestamp 1586364061
transform 1 0 1932 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 4232 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_21
timestamp 1586364061
transform 1 0 3036 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_42_29
timestamp 1586364061
transform 1 0 3772 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_36
timestamp 1586364061
transform 1 0 4416 0 -1 25568
box -38 -48 406 592
use scs8hd_buf_4  mux_top_track_28.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 4784 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_46
timestamp 1586364061
transform 1 0 5336 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_58
timestamp 1586364061
transform 1 0 6440 0 -1 25568
box -38 -48 406 592
use scs8hd_mux2_2  mux_left_track_33.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7912 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 7636 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_1  FILLER_42_73
timestamp 1586364061
transform 1 0 7820 0 -1 25568
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_83
timestamp 1586364061
transform 1 0 8740 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_42_91
timestamp 1586364061
transform 1 0 9476 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 774 592
use scs8hd_buf_4  mux_top_track_20.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 11040 0 -1 25568
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 10764 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_102
timestamp 1586364061
transform 1 0 10488 0 -1 25568
box -38 -48 314 592
use scs8hd_fill_1  FILLER_42_107
timestamp 1586364061
transform 1 0 10948 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_114
timestamp 1586364061
transform 1 0 11592 0 -1 25568
box -38 -48 774 592
use scs8hd_buf_2  _123_
timestamp 1586364061
transform 1 0 12788 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 13340 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_122
timestamp 1586364061
transform 1 0 12328 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_131
timestamp 1586364061
transform 1 0 13156 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_135
timestamp 1586364061
transform 1 0 13524 0 -1 25568
box -38 -48 406 592
use scs8hd_buf_2  _124_
timestamp 1586364061
transform 1 0 13892 0 -1 25568
box -38 -48 406 592
use scs8hd_buf_4  mux_top_track_22.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14444 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_143
timestamp 1586364061
transform 1 0 14260 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_147
timestamp 1586364061
transform 1 0 14628 0 -1 25568
box -38 -48 774 592
use scs8hd_buf_4  mux_top_track_14.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16928 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_8  FILLER_42_162
timestamp 1586364061
transform 1 0 16008 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_42_170
timestamp 1586364061
transform 1 0 16744 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_178
timestamp 1586364061
transform 1 0 17480 0 -1 25568
box -38 -48 774 592
use scs8hd_buf_2  _122_
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_191
timestamp 1586364061
transform 1 0 18676 0 -1 25568
box -38 -48 774 592
use scs8hd_buf_2  _116_
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 406 592
use scs8hd_buf_2  _121_
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_203
timestamp 1586364061
transform 1 0 19780 0 -1 25568
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_42_215
timestamp 1586364061
transform 1 0 20884 0 -1 25568
box -38 -48 222 592
use scs8hd_buf_2  _115_
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_8  FILLER_42_222
timestamp 1586364061
transform 1 0 21528 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_12  FILLER_42_234
timestamp 1586364061
transform 1 0 22632 0 -1 25568
box -38 -48 1142 592
use scs8hd_buf_2  _112_
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_246
timestamp 1586364061
transform 1 0 23736 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_253
timestamp 1586364061
transform 1 0 24380 0 -1 25568
box -38 -48 774 592
use scs8hd_buf_2  _106_
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_265
timestamp 1586364061
transform 1 0 25484 0 -1 25568
box -38 -48 1142 592
<< labels >>
rlabel metal3 s 0 26936 480 27056 6 ccff_head
port 0 nsew default input
rlabel metal2 s 25962 27520 26018 28000 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 0 13880 480 14000 6 chanx_left_in[0]
port 2 nsew default input
rlabel metal3 s 0 20408 480 20528 6 chanx_left_in[10]
port 3 nsew default input
rlabel metal3 s 0 21088 480 21208 6 chanx_left_in[11]
port 4 nsew default input
rlabel metal3 s 0 21768 480 21888 6 chanx_left_in[12]
port 5 nsew default input
rlabel metal3 s 0 22312 480 22432 6 chanx_left_in[13]
port 6 nsew default input
rlabel metal3 s 0 22992 480 23112 6 chanx_left_in[14]
port 7 nsew default input
rlabel metal3 s 0 23672 480 23792 6 chanx_left_in[15]
port 8 nsew default input
rlabel metal3 s 0 24352 480 24472 6 chanx_left_in[16]
port 9 nsew default input
rlabel metal3 s 0 25032 480 25152 6 chanx_left_in[17]
port 10 nsew default input
rlabel metal3 s 0 25576 480 25696 6 chanx_left_in[18]
port 11 nsew default input
rlabel metal3 s 0 26256 480 26376 6 chanx_left_in[19]
port 12 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[1]
port 13 nsew default input
rlabel metal3 s 0 15240 480 15360 6 chanx_left_in[2]
port 14 nsew default input
rlabel metal3 s 0 15784 480 15904 6 chanx_left_in[3]
port 15 nsew default input
rlabel metal3 s 0 16464 480 16584 6 chanx_left_in[4]
port 16 nsew default input
rlabel metal3 s 0 17144 480 17264 6 chanx_left_in[5]
port 17 nsew default input
rlabel metal3 s 0 17824 480 17944 6 chanx_left_in[6]
port 18 nsew default input
rlabel metal3 s 0 18504 480 18624 6 chanx_left_in[7]
port 19 nsew default input
rlabel metal3 s 0 19048 480 19168 6 chanx_left_in[8]
port 20 nsew default input
rlabel metal3 s 0 19728 480 19848 6 chanx_left_in[9]
port 21 nsew default input
rlabel metal3 s 0 824 480 944 6 chanx_left_out[0]
port 22 nsew default tristate
rlabel metal3 s 0 7352 480 7472 6 chanx_left_out[10]
port 23 nsew default tristate
rlabel metal3 s 0 8032 480 8152 6 chanx_left_out[11]
port 24 nsew default tristate
rlabel metal3 s 0 8712 480 8832 6 chanx_left_out[12]
port 25 nsew default tristate
rlabel metal3 s 0 9392 480 9512 6 chanx_left_out[13]
port 26 nsew default tristate
rlabel metal3 s 0 9936 480 10056 6 chanx_left_out[14]
port 27 nsew default tristate
rlabel metal3 s 0 10616 480 10736 6 chanx_left_out[15]
port 28 nsew default tristate
rlabel metal3 s 0 11296 480 11416 6 chanx_left_out[16]
port 29 nsew default tristate
rlabel metal3 s 0 11976 480 12096 6 chanx_left_out[17]
port 30 nsew default tristate
rlabel metal3 s 0 12656 480 12776 6 chanx_left_out[18]
port 31 nsew default tristate
rlabel metal3 s 0 13200 480 13320 6 chanx_left_out[19]
port 32 nsew default tristate
rlabel metal3 s 0 1504 480 1624 6 chanx_left_out[1]
port 33 nsew default tristate
rlabel metal3 s 0 2184 480 2304 6 chanx_left_out[2]
port 34 nsew default tristate
rlabel metal3 s 0 2864 480 2984 6 chanx_left_out[3]
port 35 nsew default tristate
rlabel metal3 s 0 3408 480 3528 6 chanx_left_out[4]
port 36 nsew default tristate
rlabel metal3 s 0 4088 480 4208 6 chanx_left_out[5]
port 37 nsew default tristate
rlabel metal3 s 0 4768 480 4888 6 chanx_left_out[6]
port 38 nsew default tristate
rlabel metal3 s 0 5448 480 5568 6 chanx_left_out[7]
port 39 nsew default tristate
rlabel metal3 s 0 6128 480 6248 6 chanx_left_out[8]
port 40 nsew default tristate
rlabel metal3 s 0 6672 480 6792 6 chanx_left_out[9]
port 41 nsew default tristate
rlabel metal3 s 27520 11160 28000 11280 6 chanx_right_in[0]
port 42 nsew default input
rlabel metal3 s 27520 16464 28000 16584 6 chanx_right_in[10]
port 43 nsew default input
rlabel metal3 s 27520 17008 28000 17128 6 chanx_right_in[11]
port 44 nsew default input
rlabel metal3 s 27520 17552 28000 17672 6 chanx_right_in[12]
port 45 nsew default input
rlabel metal3 s 27520 18096 28000 18216 6 chanx_right_in[13]
port 46 nsew default input
rlabel metal3 s 27520 18640 28000 18760 6 chanx_right_in[14]
port 47 nsew default input
rlabel metal3 s 27520 19048 28000 19168 6 chanx_right_in[15]
port 48 nsew default input
rlabel metal3 s 27520 19592 28000 19712 6 chanx_right_in[16]
port 49 nsew default input
rlabel metal3 s 27520 20136 28000 20256 6 chanx_right_in[17]
port 50 nsew default input
rlabel metal3 s 27520 20680 28000 20800 6 chanx_right_in[18]
port 51 nsew default input
rlabel metal3 s 27520 21224 28000 21344 6 chanx_right_in[19]
port 52 nsew default input
rlabel metal3 s 27520 11704 28000 11824 6 chanx_right_in[1]
port 53 nsew default input
rlabel metal3 s 27520 12248 28000 12368 6 chanx_right_in[2]
port 54 nsew default input
rlabel metal3 s 27520 12792 28000 12912 6 chanx_right_in[3]
port 55 nsew default input
rlabel metal3 s 27520 13336 28000 13456 6 chanx_right_in[4]
port 56 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 chanx_right_in[5]
port 57 nsew default input
rlabel metal3 s 27520 14288 28000 14408 6 chanx_right_in[6]
port 58 nsew default input
rlabel metal3 s 27520 14832 28000 14952 6 chanx_right_in[7]
port 59 nsew default input
rlabel metal3 s 27520 15376 28000 15496 6 chanx_right_in[8]
port 60 nsew default input
rlabel metal3 s 27520 15920 28000 16040 6 chanx_right_in[9]
port 61 nsew default input
rlabel metal3 s 27520 552 28000 672 6 chanx_right_out[0]
port 62 nsew default tristate
rlabel metal3 s 27520 5856 28000 5976 6 chanx_right_out[10]
port 63 nsew default tristate
rlabel metal3 s 27520 6400 28000 6520 6 chanx_right_out[11]
port 64 nsew default tristate
rlabel metal3 s 27520 6944 28000 7064 6 chanx_right_out[12]
port 65 nsew default tristate
rlabel metal3 s 27520 7488 28000 7608 6 chanx_right_out[13]
port 66 nsew default tristate
rlabel metal3 s 27520 8032 28000 8152 6 chanx_right_out[14]
port 67 nsew default tristate
rlabel metal3 s 27520 8576 28000 8696 6 chanx_right_out[15]
port 68 nsew default tristate
rlabel metal3 s 27520 9120 28000 9240 6 chanx_right_out[16]
port 69 nsew default tristate
rlabel metal3 s 27520 9528 28000 9648 6 chanx_right_out[17]
port 70 nsew default tristate
rlabel metal3 s 27520 10072 28000 10192 6 chanx_right_out[18]
port 71 nsew default tristate
rlabel metal3 s 27520 10616 28000 10736 6 chanx_right_out[19]
port 72 nsew default tristate
rlabel metal3 s 27520 1096 28000 1216 6 chanx_right_out[1]
port 73 nsew default tristate
rlabel metal3 s 27520 1640 28000 1760 6 chanx_right_out[2]
port 74 nsew default tristate
rlabel metal3 s 27520 2184 28000 2304 6 chanx_right_out[3]
port 75 nsew default tristate
rlabel metal3 s 27520 2728 28000 2848 6 chanx_right_out[4]
port 76 nsew default tristate
rlabel metal3 s 27520 3272 28000 3392 6 chanx_right_out[5]
port 77 nsew default tristate
rlabel metal3 s 27520 3816 28000 3936 6 chanx_right_out[6]
port 78 nsew default tristate
rlabel metal3 s 27520 4360 28000 4480 6 chanx_right_out[7]
port 79 nsew default tristate
rlabel metal3 s 27520 4768 28000 4888 6 chanx_right_out[8]
port 80 nsew default tristate
rlabel metal3 s 27520 5312 28000 5432 6 chanx_right_out[9]
port 81 nsew default tristate
rlabel metal2 s 4434 27520 4490 28000 6 chany_top_in[0]
port 82 nsew default input
rlabel metal2 s 9862 27520 9918 28000 6 chany_top_in[10]
port 83 nsew default input
rlabel metal2 s 10414 27520 10470 28000 6 chany_top_in[11]
port 84 nsew default input
rlabel metal2 s 10874 27520 10930 28000 6 chany_top_in[12]
port 85 nsew default input
rlabel metal2 s 11426 27520 11482 28000 6 chany_top_in[13]
port 86 nsew default input
rlabel metal2 s 11978 27520 12034 28000 6 chany_top_in[14]
port 87 nsew default input
rlabel metal2 s 12530 27520 12586 28000 6 chany_top_in[15]
port 88 nsew default input
rlabel metal2 s 13082 27520 13138 28000 6 chany_top_in[16]
port 89 nsew default input
rlabel metal2 s 13634 27520 13690 28000 6 chany_top_in[17]
port 90 nsew default input
rlabel metal2 s 14186 27520 14242 28000 6 chany_top_in[18]
port 91 nsew default input
rlabel metal2 s 14646 27520 14702 28000 6 chany_top_in[19]
port 92 nsew default input
rlabel metal2 s 4986 27520 5042 28000 6 chany_top_in[1]
port 93 nsew default input
rlabel metal2 s 5538 27520 5594 28000 6 chany_top_in[2]
port 94 nsew default input
rlabel metal2 s 6090 27520 6146 28000 6 chany_top_in[3]
port 95 nsew default input
rlabel metal2 s 6642 27520 6698 28000 6 chany_top_in[4]
port 96 nsew default input
rlabel metal2 s 7194 27520 7250 28000 6 chany_top_in[5]
port 97 nsew default input
rlabel metal2 s 7654 27520 7710 28000 6 chany_top_in[6]
port 98 nsew default input
rlabel metal2 s 8206 27520 8262 28000 6 chany_top_in[7]
port 99 nsew default input
rlabel metal2 s 8758 27520 8814 28000 6 chany_top_in[8]
port 100 nsew default input
rlabel metal2 s 9310 27520 9366 28000 6 chany_top_in[9]
port 101 nsew default input
rlabel metal2 s 15198 27520 15254 28000 6 chany_top_out[0]
port 102 nsew default tristate
rlabel metal2 s 20626 27520 20682 28000 6 chany_top_out[10]
port 103 nsew default tristate
rlabel metal2 s 21178 27520 21234 28000 6 chany_top_out[11]
port 104 nsew default tristate
rlabel metal2 s 21638 27520 21694 28000 6 chany_top_out[12]
port 105 nsew default tristate
rlabel metal2 s 22190 27520 22246 28000 6 chany_top_out[13]
port 106 nsew default tristate
rlabel metal2 s 22742 27520 22798 28000 6 chany_top_out[14]
port 107 nsew default tristate
rlabel metal2 s 23294 27520 23350 28000 6 chany_top_out[15]
port 108 nsew default tristate
rlabel metal2 s 23846 27520 23902 28000 6 chany_top_out[16]
port 109 nsew default tristate
rlabel metal2 s 24398 27520 24454 28000 6 chany_top_out[17]
port 110 nsew default tristate
rlabel metal2 s 24858 27520 24914 28000 6 chany_top_out[18]
port 111 nsew default tristate
rlabel metal2 s 25410 27520 25466 28000 6 chany_top_out[19]
port 112 nsew default tristate
rlabel metal2 s 15750 27520 15806 28000 6 chany_top_out[1]
port 113 nsew default tristate
rlabel metal2 s 16302 27520 16358 28000 6 chany_top_out[2]
port 114 nsew default tristate
rlabel metal2 s 16854 27520 16910 28000 6 chany_top_out[3]
port 115 nsew default tristate
rlabel metal2 s 17406 27520 17462 28000 6 chany_top_out[4]
port 116 nsew default tristate
rlabel metal2 s 17866 27520 17922 28000 6 chany_top_out[5]
port 117 nsew default tristate
rlabel metal2 s 18418 27520 18474 28000 6 chany_top_out[6]
port 118 nsew default tristate
rlabel metal2 s 18970 27520 19026 28000 6 chany_top_out[7]
port 119 nsew default tristate
rlabel metal2 s 19522 27520 19578 28000 6 chany_top_out[8]
port 120 nsew default tristate
rlabel metal2 s 20074 27520 20130 28000 6 chany_top_out[9]
port 121 nsew default tristate
rlabel metal3 s 0 280 480 400 6 left_bottom_grid_pin_1_
port 122 nsew default input
rlabel metal2 s 26514 27520 26570 28000 6 left_top_grid_pin_42_
port 123 nsew default input
rlabel metal3 s 27520 25984 28000 26104 6 left_top_grid_pin_43_
port 124 nsew default input
rlabel metal3 s 27520 26528 28000 26648 6 left_top_grid_pin_44_
port 125 nsew default input
rlabel metal3 s 27520 27072 28000 27192 6 left_top_grid_pin_45_
port 126 nsew default input
rlabel metal3 s 0 27616 480 27736 6 left_top_grid_pin_46_
port 127 nsew default input
rlabel metal2 s 14002 0 14058 480 6 left_top_grid_pin_47_
port 128 nsew default input
rlabel metal3 s 27520 27616 28000 27736 6 left_top_grid_pin_48_
port 129 nsew default input
rlabel metal2 s 27066 27520 27122 28000 6 left_top_grid_pin_49_
port 130 nsew default input
rlabel metal2 s 27618 27520 27674 28000 6 prog_clk
port 131 nsew default input
rlabel metal3 s 27520 144 28000 264 6 right_bottom_grid_pin_1_
port 132 nsew default input
rlabel metal3 s 27520 21768 28000 21888 6 right_top_grid_pin_42_
port 133 nsew default input
rlabel metal3 s 27520 22312 28000 22432 6 right_top_grid_pin_43_
port 134 nsew default input
rlabel metal3 s 27520 22856 28000 22976 6 right_top_grid_pin_44_
port 135 nsew default input
rlabel metal3 s 27520 23400 28000 23520 6 right_top_grid_pin_45_
port 136 nsew default input
rlabel metal3 s 27520 23808 28000 23928 6 right_top_grid_pin_46_
port 137 nsew default input
rlabel metal3 s 27520 24352 28000 24472 6 right_top_grid_pin_47_
port 138 nsew default input
rlabel metal3 s 27520 24896 28000 25016 6 right_top_grid_pin_48_
port 139 nsew default input
rlabel metal3 s 27520 25440 28000 25560 6 right_top_grid_pin_49_
port 140 nsew default input
rlabel metal2 s 202 27520 258 28000 6 top_left_grid_pin_34_
port 141 nsew default input
rlabel metal2 s 662 27520 718 28000 6 top_left_grid_pin_35_
port 142 nsew default input
rlabel metal2 s 1214 27520 1270 28000 6 top_left_grid_pin_36_
port 143 nsew default input
rlabel metal2 s 1766 27520 1822 28000 6 top_left_grid_pin_37_
port 144 nsew default input
rlabel metal2 s 2318 27520 2374 28000 6 top_left_grid_pin_38_
port 145 nsew default input
rlabel metal2 s 2870 27520 2926 28000 6 top_left_grid_pin_39_
port 146 nsew default input
rlabel metal2 s 3422 27520 3478 28000 6 top_left_grid_pin_40_
port 147 nsew default input
rlabel metal2 s 3882 27520 3938 28000 6 top_left_grid_pin_41_
port 148 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 149 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 150 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
