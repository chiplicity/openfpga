magic
tech sky130A
magscale 1 2
timestamp 1608761684
<< checkpaint >>
rect -1260 -1260 24060 23916
<< locali >>
rect 9597 14255 9631 14425
rect 14933 14255 14967 14357
rect 16681 14255 16715 14425
rect 8125 11943 8159 12045
rect 13553 11943 13587 12249
rect 11253 7047 11287 7149
<< viali >>
rect 20177 19865 20211 19899
rect 20729 19865 20763 19899
rect 19993 19729 20027 19763
rect 20545 19729 20579 19763
rect 20453 19321 20487 19355
rect 13645 19253 13679 19287
rect 5273 19185 5307 19219
rect 8309 19185 8343 19219
rect 10241 19185 10275 19219
rect 14289 19185 14323 19219
rect 15945 19185 15979 19219
rect 16957 19185 16991 19219
rect 19717 19185 19751 19219
rect 10149 19117 10183 19151
rect 11253 19117 11287 19151
rect 17417 19117 17451 19151
rect 17969 19117 18003 19151
rect 19441 19117 19475 19151
rect 20269 19117 20303 19151
rect 8125 19049 8159 19083
rect 8769 19049 8803 19083
rect 11520 19049 11554 19083
rect 16773 19049 16807 19083
rect 18797 19049 18831 19083
rect 4721 18981 4755 19015
rect 5089 18981 5123 19015
rect 5181 18981 5215 19015
rect 7757 18981 7791 19015
rect 8217 18981 8251 19015
rect 9689 18981 9723 19015
rect 10057 18981 10091 19015
rect 12633 18981 12667 19015
rect 14013 18981 14047 19015
rect 14105 18981 14139 19015
rect 15301 18981 15335 19015
rect 15669 18981 15703 19015
rect 15761 18981 15795 19015
rect 16313 18981 16347 19015
rect 16681 18981 16715 19015
rect 17601 18981 17635 19015
rect 3525 18777 3559 18811
rect 5457 18777 5491 18811
rect 5825 18777 5859 18811
rect 11529 18777 11563 18811
rect 14013 18777 14047 18811
rect 18061 18777 18095 18811
rect 4068 18709 4102 18743
rect 8738 18709 8772 18743
rect 12878 18709 12912 18743
rect 14534 18709 14568 18743
rect 16190 18709 16224 18743
rect 19717 18709 19751 18743
rect 20453 18709 20487 18743
rect 2412 18641 2446 18675
rect 3801 18641 3835 18675
rect 6837 18641 6871 18675
rect 7104 18641 7138 18675
rect 8493 18641 8527 18675
rect 10149 18641 10183 18675
rect 10405 18641 10439 18675
rect 19441 18641 19475 18675
rect 20177 18641 20211 18675
rect 2145 18573 2179 18607
rect 5917 18573 5951 18607
rect 6009 18573 6043 18607
rect 11805 18573 11839 18607
rect 12633 18573 12667 18607
rect 14289 18573 14323 18607
rect 15945 18573 15979 18607
rect 8217 18505 8251 18539
rect 9873 18505 9907 18539
rect 5181 18437 5215 18471
rect 15669 18437 15703 18471
rect 17325 18437 17359 18471
rect 7297 18233 7331 18267
rect 7757 18233 7791 18267
rect 12357 18233 12391 18267
rect 18705 18233 18739 18267
rect 19625 18233 19659 18267
rect 20177 18233 20211 18267
rect 3341 18097 3375 18131
rect 5089 18097 5123 18131
rect 8309 18097 8343 18131
rect 11345 18097 11379 18131
rect 11529 18097 11563 18131
rect 12909 18097 12943 18131
rect 13921 18097 13955 18131
rect 17417 18097 17451 18131
rect 5917 18029 5951 18063
rect 8125 18029 8159 18063
rect 8217 18029 8251 18063
rect 11253 18029 11287 18063
rect 12817 18029 12851 18063
rect 17141 18029 17175 18063
rect 18521 18029 18555 18063
rect 19441 18029 19475 18063
rect 19993 18029 20027 18063
rect 6184 17961 6218 17995
rect 2789 17893 2823 17927
rect 3157 17893 3191 17927
rect 3249 17893 3283 17927
rect 10885 17893 10919 17927
rect 12725 17893 12759 17927
rect 2789 17689 2823 17723
rect 3433 17689 3467 17723
rect 3893 17689 3927 17723
rect 3801 17621 3835 17655
rect 18337 17621 18371 17655
rect 1409 17553 1443 17587
rect 1676 17553 1710 17587
rect 18061 17553 18095 17587
rect 19441 17553 19475 17587
rect 19717 17553 19751 17587
rect 20545 17553 20579 17587
rect 3985 17485 4019 17519
rect 20729 17349 20763 17383
rect 17785 17145 17819 17179
rect 18705 17145 18739 17179
rect 20453 17145 20487 17179
rect 6193 17077 6227 17111
rect 3157 17009 3191 17043
rect 4353 17009 4387 17043
rect 7573 17009 7607 17043
rect 8861 17009 8895 17043
rect 19349 17009 19383 17043
rect 4077 16941 4111 16975
rect 4813 16941 4847 16975
rect 7297 16941 7331 16975
rect 16405 16941 16439 16975
rect 18521 16941 18555 16975
rect 19073 16941 19107 16975
rect 20269 16941 20303 16975
rect 5080 16873 5114 16907
rect 8769 16873 8803 16907
rect 16672 16873 16706 16907
rect 8309 16805 8343 16839
rect 8677 16805 8711 16839
rect 9873 16805 9907 16839
rect 6837 16601 6871 16635
rect 10517 16601 10551 16635
rect 11345 16601 11379 16635
rect 11713 16601 11747 16635
rect 12909 16601 12943 16635
rect 14381 16601 14415 16635
rect 16865 16601 16899 16635
rect 20913 16601 20947 16635
rect 10609 16533 10643 16567
rect 19533 16533 19567 16567
rect 20269 16533 20303 16567
rect 7205 16465 7239 16499
rect 7849 16465 7883 16499
rect 8493 16465 8527 16499
rect 8760 16465 8794 16499
rect 12817 16465 12851 16499
rect 13461 16465 13495 16499
rect 14289 16465 14323 16499
rect 15752 16465 15786 16499
rect 19257 16465 19291 16499
rect 19993 16465 20027 16499
rect 20729 16465 20763 16499
rect 7297 16397 7331 16431
rect 7389 16397 7423 16431
rect 10701 16397 10735 16431
rect 11805 16397 11839 16431
rect 11897 16397 11931 16431
rect 13001 16397 13035 16431
rect 14473 16397 14507 16431
rect 15485 16397 15519 16431
rect 18061 16397 18095 16431
rect 12449 16329 12483 16363
rect 9873 16261 9907 16295
rect 10149 16261 10183 16295
rect 13921 16261 13955 16295
rect 3341 16057 3375 16091
rect 6377 16057 6411 16091
rect 7021 16057 7055 16091
rect 13001 16057 13035 16091
rect 17417 16057 17451 16091
rect 20453 16057 20487 16091
rect 16405 15989 16439 16023
rect 19901 15989 19935 16023
rect 1961 15921 1995 15955
rect 4997 15921 5031 15955
rect 7573 15921 7607 15955
rect 9965 15921 9999 15955
rect 16957 15921 16991 15955
rect 17877 15921 17911 15955
rect 17969 15921 18003 15955
rect 5264 15853 5298 15887
rect 7389 15853 7423 15887
rect 7481 15853 7515 15887
rect 10221 15853 10255 15887
rect 11621 15853 11655 15887
rect 11888 15853 11922 15887
rect 13277 15853 13311 15887
rect 13533 15853 13567 15887
rect 19717 15853 19751 15887
rect 20269 15853 20303 15887
rect 2228 15785 2262 15819
rect 16773 15785 16807 15819
rect 17785 15785 17819 15819
rect 11345 15717 11379 15751
rect 14657 15717 14691 15751
rect 15301 15717 15335 15751
rect 16865 15717 16899 15751
rect 2789 15513 2823 15547
rect 3341 15513 3375 15547
rect 3801 15513 3835 15547
rect 14749 15513 14783 15547
rect 20177 15513 20211 15547
rect 20729 15513 20763 15547
rect 3709 15445 3743 15479
rect 14841 15445 14875 15479
rect 2697 15377 2731 15411
rect 18981 15377 19015 15411
rect 19257 15377 19291 15411
rect 19993 15377 20027 15411
rect 20545 15377 20579 15411
rect 2881 15309 2915 15343
rect 3893 15309 3927 15343
rect 15025 15309 15059 15343
rect 2329 15241 2363 15275
rect 14381 15241 14415 15275
rect 2881 14969 2915 15003
rect 6377 14969 6411 15003
rect 16865 14969 16899 15003
rect 6837 14901 6871 14935
rect 13185 14901 13219 14935
rect 17141 14901 17175 14935
rect 1501 14833 1535 14867
rect 3341 14833 3375 14867
rect 4997 14833 5031 14867
rect 8493 14833 8527 14867
rect 17693 14833 17727 14867
rect 19809 14833 19843 14867
rect 7021 14765 7055 14799
rect 8217 14765 8251 14799
rect 8309 14765 8343 14799
rect 13369 14765 13403 14799
rect 15485 14765 15519 14799
rect 18889 14765 18923 14799
rect 19625 14765 19659 14799
rect 1768 14697 1802 14731
rect 5264 14697 5298 14731
rect 15752 14697 15786 14731
rect 19165 14697 19199 14731
rect 7849 14629 7883 14663
rect 9689 14629 9723 14663
rect 17509 14629 17543 14663
rect 17601 14629 17635 14663
rect 9505 14425 9539 14459
rect 9597 14425 9631 14459
rect 9781 14425 9815 14459
rect 10149 14425 10183 14459
rect 14841 14425 14875 14459
rect 16497 14425 16531 14459
rect 16681 14425 16715 14459
rect 16773 14425 16807 14459
rect 20729 14425 20763 14459
rect 3792 14357 3826 14391
rect 3525 14289 3559 14323
rect 5549 14289 5583 14323
rect 5641 14289 5675 14323
rect 8125 14289 8159 14323
rect 8392 14289 8426 14323
rect 10241 14357 10275 14391
rect 14933 14357 14967 14391
rect 15362 14357 15396 14391
rect 12817 14289 12851 14323
rect 13728 14289 13762 14323
rect 19349 14357 19383 14391
rect 17141 14289 17175 14323
rect 17233 14289 17267 14323
rect 19073 14289 19107 14323
rect 19809 14289 19843 14323
rect 20085 14289 20119 14323
rect 20545 14289 20579 14323
rect 5825 14221 5859 14255
rect 9597 14221 9631 14255
rect 10333 14221 10367 14255
rect 12909 14221 12943 14255
rect 13001 14221 13035 14255
rect 13461 14221 13495 14255
rect 14933 14221 14967 14255
rect 15117 14221 15151 14255
rect 16681 14221 16715 14255
rect 17325 14221 17359 14255
rect 4905 14085 4939 14119
rect 5181 14085 5215 14119
rect 12449 14085 12483 14119
rect 3433 13881 3467 13915
rect 4629 13881 4663 13915
rect 7021 13881 7055 13915
rect 8677 13881 8711 13915
rect 12081 13881 12115 13915
rect 12357 13881 12391 13915
rect 16681 13881 16715 13915
rect 18521 13881 18555 13915
rect 20453 13881 20487 13915
rect 2053 13745 2087 13779
rect 5089 13745 5123 13779
rect 5181 13745 5215 13779
rect 10701 13745 10735 13779
rect 13001 13745 13035 13779
rect 13369 13745 13403 13779
rect 17141 13745 17175 13779
rect 17325 13745 17359 13779
rect 2320 13677 2354 13711
rect 5641 13677 5675 13711
rect 5908 13677 5942 13711
rect 7297 13677 7331 13711
rect 9137 13677 9171 13711
rect 12817 13677 12851 13711
rect 18337 13677 18371 13711
rect 20269 13677 20303 13711
rect 7564 13609 7598 13643
rect 10968 13609 11002 13643
rect 12725 13609 12759 13643
rect 17049 13609 17083 13643
rect 17693 13609 17727 13643
rect 4997 13541 5031 13575
rect 8953 13541 8987 13575
rect 4997 13337 5031 13371
rect 11253 13337 11287 13371
rect 12817 13337 12851 13371
rect 12909 13337 12943 13371
rect 20177 13337 20211 13371
rect 20729 13337 20763 13371
rect 18889 13269 18923 13303
rect 9965 13201 9999 13235
rect 18613 13201 18647 13235
rect 19993 13201 20027 13235
rect 20545 13201 20579 13235
rect 13001 13133 13035 13167
rect 12449 12997 12483 13031
rect 11069 12793 11103 12827
rect 12449 12793 12483 12827
rect 13369 12793 13403 12827
rect 20361 12793 20395 12827
rect 19809 12725 19843 12759
rect 11437 12657 11471 12691
rect 13921 12657 13955 12691
rect 15577 12657 15611 12691
rect 9689 12589 9723 12623
rect 11161 12589 11195 12623
rect 12633 12589 12667 12623
rect 15301 12589 15335 12623
rect 16681 12589 16715 12623
rect 19625 12589 19659 12623
rect 20177 12589 20211 12623
rect 9934 12521 9968 12555
rect 13737 12521 13771 12555
rect 16948 12521 16982 12555
rect 13829 12453 13863 12487
rect 18061 12453 18095 12487
rect 7297 12249 7331 12283
rect 9965 12249 9999 12283
rect 12725 12249 12759 12283
rect 13553 12249 13587 12283
rect 14013 12249 14047 12283
rect 14473 12249 14507 12283
rect 20729 12249 20763 12283
rect 7205 12181 7239 12215
rect 10425 12181 10459 12215
rect 8033 12113 8067 12147
rect 8565 12113 8599 12147
rect 10333 12113 10367 12147
rect 13093 12113 13127 12147
rect 7481 12045 7515 12079
rect 8125 12045 8159 12079
rect 8309 12045 8343 12079
rect 10517 12045 10551 12079
rect 13185 12045 13219 12079
rect 13369 12045 13403 12079
rect 9689 11977 9723 12011
rect 6837 11909 6871 11943
rect 7849 11909 7883 11943
rect 8125 11909 8159 11943
rect 14381 12181 14415 12215
rect 15384 12181 15418 12215
rect 19533 12181 19567 12215
rect 13921 12113 13955 12147
rect 15117 12113 15151 12147
rect 18429 12113 18463 12147
rect 19257 12113 19291 12147
rect 19993 12113 20027 12147
rect 20545 12113 20579 12147
rect 14657 12045 14691 12079
rect 18521 12045 18555 12079
rect 18613 12045 18647 12079
rect 18061 11977 18095 12011
rect 20177 11977 20211 12011
rect 13553 11909 13587 11943
rect 13737 11909 13771 11943
rect 16497 11909 16531 11943
rect 10333 11705 10367 11739
rect 13645 11705 13679 11739
rect 18061 11705 18095 11739
rect 20453 11705 20487 11739
rect 7849 11637 7883 11671
rect 8677 11569 8711 11603
rect 10885 11569 10919 11603
rect 14197 11569 14231 11603
rect 18613 11569 18647 11603
rect 6469 11501 6503 11535
rect 6736 11501 6770 11535
rect 11989 11501 12023 11535
rect 12256 11501 12290 11535
rect 14105 11501 14139 11535
rect 20269 11501 20303 11535
rect 8585 11433 8619 11467
rect 10793 11433 10827 11467
rect 18429 11433 18463 11467
rect 19073 11433 19107 11467
rect 8125 11365 8159 11399
rect 8493 11365 8527 11399
rect 10701 11365 10735 11399
rect 11345 11365 11379 11399
rect 13369 11365 13403 11399
rect 14013 11365 14047 11399
rect 18521 11365 18555 11399
rect 8125 11161 8159 11195
rect 13645 11161 13679 11195
rect 15945 11161 15979 11195
rect 17417 11161 17451 11195
rect 18889 11161 18923 11195
rect 20177 11161 20211 11195
rect 20729 11161 20763 11195
rect 16405 11093 16439 11127
rect 8217 11025 8251 11059
rect 14013 11025 14047 11059
rect 14657 11025 14691 11059
rect 16313 11025 16347 11059
rect 17325 11025 17359 11059
rect 19257 11025 19291 11059
rect 19993 11025 20027 11059
rect 20545 11025 20579 11059
rect 8401 10957 8435 10991
rect 14105 10957 14139 10991
rect 14197 10957 14231 10991
rect 16497 10957 16531 10991
rect 17509 10957 17543 10991
rect 19349 10957 19383 10991
rect 19441 10957 19475 10991
rect 7757 10889 7791 10923
rect 16957 10889 16991 10923
rect 8585 10617 8619 10651
rect 16497 10617 16531 10651
rect 20453 10617 20487 10651
rect 10057 10549 10091 10583
rect 10609 10481 10643 10515
rect 11345 10481 11379 10515
rect 17141 10481 17175 10515
rect 7205 10413 7239 10447
rect 11069 10413 11103 10447
rect 20269 10413 20303 10447
rect 7472 10345 7506 10379
rect 10425 10345 10459 10379
rect 10517 10277 10551 10311
rect 16865 10277 16899 10311
rect 16957 10277 16991 10311
rect 9873 10073 9907 10107
rect 11253 10073 11287 10107
rect 11345 10073 11379 10107
rect 14197 10073 14231 10107
rect 17325 10073 17359 10107
rect 19901 10073 19935 10107
rect 20729 10073 20763 10107
rect 13084 10005 13118 10039
rect 16212 10005 16246 10039
rect 8760 9937 8794 9971
rect 12817 9937 12851 9971
rect 15945 9937 15979 9971
rect 18521 9937 18555 9971
rect 18788 9937 18822 9971
rect 20545 9937 20579 9971
rect 8493 9869 8527 9903
rect 11529 9869 11563 9903
rect 10885 9733 10919 9767
rect 9965 9529 9999 9563
rect 8953 9461 8987 9495
rect 17601 9461 17635 9495
rect 10609 9393 10643 9427
rect 11529 9393 11563 9427
rect 12725 9393 12759 9427
rect 18245 9393 18279 9427
rect 19257 9393 19291 9427
rect 7573 9325 7607 9359
rect 10333 9325 10367 9359
rect 11345 9325 11379 9359
rect 13553 9325 13587 9359
rect 13820 9325 13854 9359
rect 18981 9325 19015 9359
rect 7840 9257 7874 9291
rect 12541 9257 12575 9291
rect 17969 9257 18003 9291
rect 19625 9257 19659 9291
rect 10425 9189 10459 9223
rect 10977 9189 11011 9223
rect 11437 9189 11471 9223
rect 12081 9189 12115 9223
rect 12449 9189 12483 9223
rect 14933 9189 14967 9223
rect 18061 9189 18095 9223
rect 18613 9189 18647 9223
rect 19073 9189 19107 9223
rect 10609 8985 10643 9019
rect 11069 8985 11103 9019
rect 13369 8985 13403 9019
rect 15301 8985 15335 9019
rect 19533 8985 19567 9019
rect 20177 8985 20211 9019
rect 20729 8985 20763 9019
rect 10977 8849 11011 8883
rect 11621 8849 11655 8883
rect 13185 8849 13219 8883
rect 15117 8849 15151 8883
rect 18153 8849 18187 8883
rect 18420 8849 18454 8883
rect 19993 8849 20027 8883
rect 20545 8849 20579 8883
rect 11161 8781 11195 8815
rect 11529 8441 11563 8475
rect 20453 8441 20487 8475
rect 16221 8373 16255 8407
rect 13461 8305 13495 8339
rect 15669 8305 15703 8339
rect 16865 8305 16899 8339
rect 11345 8237 11379 8271
rect 13277 8237 13311 8271
rect 15485 8237 15519 8271
rect 16681 8237 16715 8271
rect 20269 8237 20303 8271
rect 16589 8169 16623 8203
rect 17233 8169 17267 8203
rect 13645 7897 13679 7931
rect 17417 7897 17451 7931
rect 19441 7897 19475 7931
rect 10885 7829 10919 7863
rect 18306 7829 18340 7863
rect 10609 7761 10643 7795
rect 14013 7761 14047 7795
rect 16304 7761 16338 7795
rect 19993 7761 20027 7795
rect 20545 7761 20579 7795
rect 14105 7693 14139 7727
rect 14289 7693 14323 7727
rect 16037 7693 16071 7727
rect 18061 7693 18095 7727
rect 20729 7625 20763 7659
rect 20177 7557 20211 7591
rect 10333 7353 10367 7387
rect 16681 7353 16715 7387
rect 10885 7217 10919 7251
rect 14657 7217 14691 7251
rect 15301 7217 15335 7251
rect 11253 7149 11287 7183
rect 11345 7149 11379 7183
rect 13001 7149 13035 7183
rect 13268 7149 13302 7183
rect 11590 7081 11624 7115
rect 15546 7081 15580 7115
rect 9873 7013 9907 7047
rect 10701 7013 10735 7047
rect 10793 7013 10827 7047
rect 11253 7013 11287 7047
rect 12725 7013 12759 7047
rect 14381 7013 14415 7047
rect 10609 6809 10643 6843
rect 10885 6809 10919 6843
rect 14013 6809 14047 6843
rect 17049 6809 17083 6843
rect 11253 6741 11287 6775
rect 14381 6741 14415 6775
rect 7553 6673 7587 6707
rect 9496 6673 9530 6707
rect 14473 6673 14507 6707
rect 17141 6673 17175 6707
rect 20545 6673 20579 6707
rect 7297 6605 7331 6639
rect 9229 6605 9263 6639
rect 11345 6605 11379 6639
rect 11437 6605 11471 6639
rect 14565 6605 14599 6639
rect 17233 6605 17267 6639
rect 8677 6537 8711 6571
rect 16681 6537 16715 6571
rect 20729 6469 20763 6503
rect 20729 5721 20763 5755
rect 20545 5585 20579 5619
rect 20729 4633 20763 4667
rect 20545 4497 20579 4531
<< metal1 >>
rect 1104 20010 21620 20032
rect 1104 19958 7846 20010
rect 7898 19958 7910 20010
rect 7962 19958 7974 20010
rect 8026 19958 8038 20010
rect 8090 19958 14710 20010
rect 14762 19958 14774 20010
rect 14826 19958 14838 20010
rect 14890 19958 14902 20010
rect 14954 19958 21620 20010
rect 1104 19936 21620 19958
rect 20162 19896 20168 19908
rect 20123 19868 20168 19896
rect 20162 19856 20168 19868
rect 20220 19856 20226 19908
rect 20622 19856 20628 19908
rect 20680 19896 20686 19908
rect 20717 19899 20775 19905
rect 20717 19896 20729 19899
rect 20680 19868 20729 19896
rect 20680 19856 20686 19868
rect 20717 19865 20729 19868
rect 20763 19865 20775 19899
rect 20717 19859 20775 19865
rect 19978 19760 19984 19772
rect 19939 19732 19984 19760
rect 19978 19720 19984 19732
rect 20036 19720 20042 19772
rect 20438 19720 20444 19772
rect 20496 19760 20502 19772
rect 20533 19763 20591 19769
rect 20533 19760 20545 19763
rect 20496 19732 20545 19760
rect 20496 19720 20502 19732
rect 20533 19729 20545 19732
rect 20579 19729 20591 19763
rect 20533 19723 20591 19729
rect 1104 19466 21620 19488
rect 1104 19414 4414 19466
rect 4466 19414 4478 19466
rect 4530 19414 4542 19466
rect 4594 19414 4606 19466
rect 4658 19414 11278 19466
rect 11330 19414 11342 19466
rect 11394 19414 11406 19466
rect 11458 19414 11470 19466
rect 11522 19414 18142 19466
rect 18194 19414 18206 19466
rect 18258 19414 18270 19466
rect 18322 19414 18334 19466
rect 18386 19414 21620 19466
rect 1104 19392 21620 19414
rect 20441 19355 20499 19361
rect 20441 19321 20453 19355
rect 20487 19352 20499 19355
rect 20530 19352 20536 19364
rect 20487 19324 20536 19352
rect 20487 19321 20499 19324
rect 20441 19315 20499 19321
rect 20530 19312 20536 19324
rect 20588 19312 20594 19364
rect 13633 19287 13691 19293
rect 13633 19253 13645 19287
rect 13679 19253 13691 19287
rect 13633 19247 13691 19253
rect 5166 19176 5172 19228
rect 5224 19216 5230 19228
rect 5261 19219 5319 19225
rect 5261 19216 5273 19219
rect 5224 19188 5273 19216
rect 5224 19176 5230 19188
rect 5261 19185 5273 19188
rect 5307 19185 5319 19219
rect 5261 19179 5319 19185
rect 8202 19176 8208 19228
rect 8260 19216 8266 19228
rect 8297 19219 8355 19225
rect 8297 19216 8309 19219
rect 8260 19188 8309 19216
rect 8260 19176 8266 19188
rect 8297 19185 8309 19188
rect 8343 19185 8355 19219
rect 10226 19216 10232 19228
rect 10187 19188 10232 19216
rect 8297 19179 8355 19185
rect 10226 19176 10232 19188
rect 10284 19176 10290 19228
rect 7760 19120 9076 19148
rect 4709 19015 4767 19021
rect 4709 18981 4721 19015
rect 4755 19012 4767 19015
rect 4890 19012 4896 19024
rect 4755 18984 4896 19012
rect 4755 18981 4767 18984
rect 4709 18975 4767 18981
rect 4890 18972 4896 18984
rect 4948 18972 4954 19024
rect 5074 19012 5080 19024
rect 5035 18984 5080 19012
rect 5074 18972 5080 18984
rect 5132 18972 5138 19024
rect 5169 19015 5227 19021
rect 5169 18981 5181 19015
rect 5215 19012 5227 19015
rect 5442 19012 5448 19024
rect 5215 18984 5448 19012
rect 5215 18981 5227 18984
rect 5169 18975 5227 18981
rect 5442 18972 5448 18984
rect 5500 18972 5506 19024
rect 7760 19021 7788 19120
rect 8113 19083 8171 19089
rect 8113 19049 8125 19083
rect 8159 19080 8171 19083
rect 8757 19083 8815 19089
rect 8757 19080 8769 19083
rect 8159 19052 8769 19080
rect 8159 19049 8171 19052
rect 8113 19043 8171 19049
rect 8757 19049 8769 19052
rect 8803 19049 8815 19083
rect 9048 19080 9076 19120
rect 9122 19108 9128 19160
rect 9180 19148 9186 19160
rect 10137 19151 10195 19157
rect 10137 19148 10149 19151
rect 9180 19120 10149 19148
rect 9180 19108 9186 19120
rect 10137 19117 10149 19120
rect 10183 19117 10195 19151
rect 11238 19148 11244 19160
rect 11199 19120 11244 19148
rect 10137 19111 10195 19117
rect 11238 19108 11244 19120
rect 11296 19108 11302 19160
rect 13648 19148 13676 19247
rect 14274 19216 14280 19228
rect 14235 19188 14280 19216
rect 14274 19176 14280 19188
rect 14332 19176 14338 19228
rect 15933 19219 15991 19225
rect 15933 19185 15945 19219
rect 15979 19216 15991 19219
rect 16114 19216 16120 19228
rect 15979 19188 16120 19216
rect 15979 19185 15991 19188
rect 15933 19179 15991 19185
rect 16114 19176 16120 19188
rect 16172 19176 16178 19228
rect 16945 19219 17003 19225
rect 16945 19185 16957 19219
rect 16991 19216 17003 19219
rect 17310 19216 17316 19228
rect 16991 19188 17316 19216
rect 16991 19185 17003 19188
rect 16945 19179 17003 19185
rect 17310 19176 17316 19188
rect 17368 19176 17374 19228
rect 19705 19219 19763 19225
rect 19705 19185 19717 19219
rect 19751 19216 19763 19219
rect 19978 19216 19984 19228
rect 19751 19188 19984 19216
rect 19751 19185 19763 19188
rect 19705 19179 19763 19185
rect 19978 19176 19984 19188
rect 20036 19176 20042 19228
rect 17402 19148 17408 19160
rect 11440 19120 11744 19148
rect 13648 19120 17264 19148
rect 17363 19120 17408 19148
rect 11440 19080 11468 19120
rect 11514 19089 11520 19092
rect 9048 19052 11468 19080
rect 8757 19043 8815 19049
rect 11508 19043 11520 19089
rect 11572 19080 11578 19092
rect 11716 19080 11744 19120
rect 15010 19080 15016 19092
rect 11572 19052 11608 19080
rect 11716 19052 15016 19080
rect 11514 19040 11520 19043
rect 11572 19040 11578 19052
rect 15010 19040 15016 19052
rect 15068 19040 15074 19092
rect 16761 19083 16819 19089
rect 16761 19080 16773 19083
rect 15304 19052 16773 19080
rect 7745 19015 7803 19021
rect 7745 18981 7757 19015
rect 7791 18981 7803 19015
rect 7745 18975 7803 18981
rect 8205 19015 8263 19021
rect 8205 18981 8217 19015
rect 8251 19012 8263 19015
rect 8294 19012 8300 19024
rect 8251 18984 8300 19012
rect 8251 18981 8263 18984
rect 8205 18975 8263 18981
rect 8294 18972 8300 18984
rect 8352 18972 8358 19024
rect 9674 19012 9680 19024
rect 9635 18984 9680 19012
rect 9674 18972 9680 18984
rect 9732 18972 9738 19024
rect 9950 18972 9956 19024
rect 10008 19012 10014 19024
rect 10045 19015 10103 19021
rect 10045 19012 10057 19015
rect 10008 18984 10057 19012
rect 10008 18972 10014 18984
rect 10045 18981 10057 18984
rect 10091 19012 10103 19015
rect 11146 19012 11152 19024
rect 10091 18984 11152 19012
rect 10091 18981 10103 18984
rect 10045 18975 10103 18981
rect 11146 18972 11152 18984
rect 11204 18972 11210 19024
rect 12618 19012 12624 19024
rect 12579 18984 12624 19012
rect 12618 18972 12624 18984
rect 12676 18972 12682 19024
rect 13906 18972 13912 19024
rect 13964 19012 13970 19024
rect 14001 19015 14059 19021
rect 14001 19012 14013 19015
rect 13964 18984 14013 19012
rect 13964 18972 13970 18984
rect 14001 18981 14013 18984
rect 14047 18981 14059 19015
rect 14001 18975 14059 18981
rect 14090 18972 14096 19024
rect 14148 19012 14154 19024
rect 15304 19021 15332 19052
rect 16761 19049 16773 19052
rect 16807 19049 16819 19083
rect 17236 19080 17264 19120
rect 17402 19108 17408 19120
rect 17460 19108 17466 19160
rect 17954 19148 17960 19160
rect 17915 19120 17960 19148
rect 17954 19108 17960 19120
rect 18012 19108 18018 19160
rect 19429 19151 19487 19157
rect 19429 19148 19441 19151
rect 18064 19120 19441 19148
rect 18064 19080 18092 19120
rect 19429 19117 19441 19120
rect 19475 19117 19487 19151
rect 20254 19148 20260 19160
rect 20215 19120 20260 19148
rect 19429 19111 19487 19117
rect 20254 19108 20260 19120
rect 20312 19108 20318 19160
rect 18782 19080 18788 19092
rect 17236 19052 18092 19080
rect 18743 19052 18788 19080
rect 16761 19043 16819 19049
rect 18782 19040 18788 19052
rect 18840 19040 18846 19092
rect 15289 19015 15347 19021
rect 14148 18984 14193 19012
rect 14148 18972 14154 18984
rect 15289 18981 15301 19015
rect 15335 18981 15347 19015
rect 15654 19012 15660 19024
rect 15615 18984 15660 19012
rect 15289 18975 15347 18981
rect 15654 18972 15660 18984
rect 15712 18972 15718 19024
rect 15746 18972 15752 19024
rect 15804 19012 15810 19024
rect 16298 19012 16304 19024
rect 15804 18984 15849 19012
rect 16259 18984 16304 19012
rect 15804 18972 15810 18984
rect 16298 18972 16304 18984
rect 16356 18972 16362 19024
rect 16666 19012 16672 19024
rect 16627 18984 16672 19012
rect 16666 18972 16672 18984
rect 16724 18972 16730 19024
rect 17589 19015 17647 19021
rect 17589 18981 17601 19015
rect 17635 19012 17647 19015
rect 17862 19012 17868 19024
rect 17635 18984 17868 19012
rect 17635 18981 17647 18984
rect 17589 18975 17647 18981
rect 17862 18972 17868 18984
rect 17920 18972 17926 19024
rect 1104 18922 21620 18944
rect 1104 18870 7846 18922
rect 7898 18870 7910 18922
rect 7962 18870 7974 18922
rect 8026 18870 8038 18922
rect 8090 18870 14710 18922
rect 14762 18870 14774 18922
rect 14826 18870 14838 18922
rect 14890 18870 14902 18922
rect 14954 18870 21620 18922
rect 1104 18848 21620 18870
rect 3513 18811 3571 18817
rect 3513 18777 3525 18811
rect 3559 18777 3571 18811
rect 5442 18808 5448 18820
rect 5403 18780 5448 18808
rect 3513 18771 3571 18777
rect 3528 18740 3556 18771
rect 5442 18768 5448 18780
rect 5500 18768 5506 18820
rect 5813 18811 5871 18817
rect 5813 18777 5825 18811
rect 5859 18808 5871 18811
rect 9950 18808 9956 18820
rect 5859 18780 9956 18808
rect 5859 18777 5871 18780
rect 5813 18771 5871 18777
rect 9950 18768 9956 18780
rect 10008 18768 10014 18820
rect 10134 18768 10140 18820
rect 10192 18808 10198 18820
rect 11514 18808 11520 18820
rect 10192 18780 10732 18808
rect 11475 18780 11520 18808
rect 10192 18768 10198 18780
rect 4056 18743 4114 18749
rect 4056 18740 4068 18743
rect 3528 18712 4068 18740
rect 4056 18709 4068 18712
rect 4102 18740 4114 18743
rect 4102 18712 6040 18740
rect 4102 18709 4114 18712
rect 4056 18703 4114 18709
rect 2400 18675 2458 18681
rect 2400 18641 2412 18675
rect 2446 18672 2458 18675
rect 2774 18672 2780 18684
rect 2446 18644 2780 18672
rect 2446 18641 2458 18644
rect 2400 18635 2458 18641
rect 2774 18632 2780 18644
rect 2832 18632 2838 18684
rect 3789 18675 3847 18681
rect 3789 18641 3801 18675
rect 3835 18672 3847 18675
rect 4982 18672 4988 18684
rect 3835 18644 4988 18672
rect 3835 18641 3847 18644
rect 3789 18635 3847 18641
rect 2133 18607 2191 18613
rect 2133 18573 2145 18607
rect 2179 18573 2191 18607
rect 2133 18567 2191 18573
rect 1486 18428 1492 18480
rect 1544 18468 1550 18480
rect 2148 18468 2176 18567
rect 3804 18468 3832 18635
rect 4982 18632 4988 18644
rect 5040 18632 5046 18684
rect 4798 18564 4804 18616
rect 4856 18604 4862 18616
rect 6012 18613 6040 18712
rect 6840 18712 7328 18740
rect 6546 18632 6552 18684
rect 6604 18672 6610 18684
rect 6840 18681 6868 18712
rect 7098 18681 7104 18684
rect 6825 18675 6883 18681
rect 6825 18672 6837 18675
rect 6604 18644 6837 18672
rect 6604 18632 6610 18644
rect 6825 18641 6837 18644
rect 6871 18641 6883 18675
rect 6825 18635 6883 18641
rect 7092 18635 7104 18681
rect 7156 18672 7162 18684
rect 7300 18672 7328 18712
rect 8202 18700 8208 18752
rect 8260 18740 8266 18752
rect 8726 18743 8784 18749
rect 8726 18740 8738 18743
rect 8260 18712 8738 18740
rect 8260 18700 8266 18712
rect 8726 18709 8738 18712
rect 8772 18709 8784 18743
rect 8726 18703 8784 18709
rect 8478 18672 8484 18684
rect 7156 18644 7192 18672
rect 7300 18644 8484 18672
rect 7098 18632 7104 18635
rect 7156 18632 7162 18644
rect 8478 18632 8484 18644
rect 8536 18672 8542 18684
rect 10137 18675 10195 18681
rect 10137 18672 10149 18675
rect 8536 18644 10149 18672
rect 8536 18632 8542 18644
rect 10137 18641 10149 18644
rect 10183 18641 10195 18675
rect 10137 18635 10195 18641
rect 10226 18632 10232 18684
rect 10284 18672 10290 18684
rect 10393 18675 10451 18681
rect 10393 18672 10405 18675
rect 10284 18644 10405 18672
rect 10284 18632 10290 18644
rect 10393 18641 10405 18644
rect 10439 18641 10451 18675
rect 10704 18672 10732 18780
rect 11514 18768 11520 18780
rect 11572 18768 11578 18820
rect 11606 18768 11612 18820
rect 11664 18808 11670 18820
rect 12250 18808 12256 18820
rect 11664 18780 12256 18808
rect 11664 18768 11670 18780
rect 12250 18768 12256 18780
rect 12308 18768 12314 18820
rect 14001 18811 14059 18817
rect 14001 18777 14013 18811
rect 14047 18777 14059 18811
rect 14001 18771 14059 18777
rect 12618 18700 12624 18752
rect 12676 18740 12682 18752
rect 12866 18743 12924 18749
rect 12866 18740 12878 18743
rect 12676 18712 12878 18740
rect 12676 18700 12682 18712
rect 12866 18709 12878 18712
rect 12912 18709 12924 18743
rect 14016 18740 14044 18771
rect 15010 18768 15016 18820
rect 15068 18808 15074 18820
rect 15068 18780 16344 18808
rect 15068 18768 15074 18780
rect 14274 18740 14280 18752
rect 14016 18712 14280 18740
rect 12866 18703 12924 18709
rect 14274 18700 14280 18712
rect 14332 18740 14338 18752
rect 14522 18743 14580 18749
rect 14522 18740 14534 18743
rect 14332 18712 14534 18740
rect 14332 18700 14338 18712
rect 14522 18709 14534 18712
rect 14568 18709 14580 18743
rect 14522 18703 14580 18709
rect 16114 18700 16120 18752
rect 16172 18749 16178 18752
rect 16172 18743 16236 18749
rect 16172 18709 16190 18743
rect 16224 18709 16236 18743
rect 16316 18740 16344 18780
rect 16666 18768 16672 18820
rect 16724 18808 16730 18820
rect 18049 18811 18107 18817
rect 18049 18808 18061 18811
rect 16724 18780 18061 18808
rect 16724 18768 16730 18780
rect 18049 18777 18061 18780
rect 18095 18777 18107 18811
rect 18049 18771 18107 18777
rect 19242 18768 19248 18820
rect 19300 18808 19306 18820
rect 20346 18808 20352 18820
rect 19300 18780 20352 18808
rect 19300 18768 19306 18780
rect 20346 18768 20352 18780
rect 20404 18768 20410 18820
rect 19705 18743 19763 18749
rect 16316 18712 19472 18740
rect 16172 18703 16236 18709
rect 16172 18700 16178 18703
rect 15746 18672 15752 18684
rect 10704 18644 15752 18672
rect 10393 18635 10451 18641
rect 15746 18632 15752 18644
rect 15804 18632 15810 18684
rect 15838 18632 15844 18684
rect 15896 18672 15902 18684
rect 19334 18672 19340 18684
rect 15896 18644 19340 18672
rect 15896 18632 15902 18644
rect 19334 18632 19340 18644
rect 19392 18632 19398 18684
rect 19444 18681 19472 18712
rect 19705 18709 19717 18743
rect 19751 18740 19763 18743
rect 20254 18740 20260 18752
rect 19751 18712 20260 18740
rect 19751 18709 19763 18712
rect 19705 18703 19763 18709
rect 20254 18700 20260 18712
rect 20312 18700 20318 18752
rect 20438 18740 20444 18752
rect 20399 18712 20444 18740
rect 20438 18700 20444 18712
rect 20496 18700 20502 18752
rect 19429 18675 19487 18681
rect 19429 18641 19441 18675
rect 19475 18641 19487 18675
rect 19429 18635 19487 18641
rect 19518 18632 19524 18684
rect 19576 18672 19582 18684
rect 20165 18675 20223 18681
rect 20165 18672 20177 18675
rect 19576 18644 20177 18672
rect 19576 18632 19582 18644
rect 20165 18641 20177 18644
rect 20211 18641 20223 18675
rect 20165 18635 20223 18641
rect 5905 18607 5963 18613
rect 5905 18604 5917 18607
rect 4856 18576 5917 18604
rect 4856 18564 4862 18576
rect 5905 18573 5917 18576
rect 5951 18573 5963 18607
rect 5905 18567 5963 18573
rect 5997 18607 6055 18613
rect 5997 18573 6009 18607
rect 6043 18573 6055 18607
rect 10244 18604 10272 18632
rect 11790 18604 11796 18616
rect 5997 18567 6055 18573
rect 9876 18576 10272 18604
rect 11751 18576 11796 18604
rect 8202 18536 8208 18548
rect 8163 18508 8208 18536
rect 8202 18496 8208 18508
rect 8260 18496 8266 18548
rect 9876 18545 9904 18576
rect 11790 18564 11796 18576
rect 11848 18564 11854 18616
rect 12621 18607 12679 18613
rect 12621 18573 12633 18607
rect 12667 18573 12679 18607
rect 12621 18567 12679 18573
rect 14277 18607 14335 18613
rect 14277 18573 14289 18607
rect 14323 18573 14335 18607
rect 15933 18607 15991 18613
rect 15933 18604 15945 18607
rect 14277 18567 14335 18573
rect 15304 18576 15945 18604
rect 9861 18539 9919 18545
rect 9861 18505 9873 18539
rect 9907 18505 9919 18539
rect 9861 18499 9919 18505
rect 11238 18496 11244 18548
rect 11296 18536 11302 18548
rect 12636 18536 12664 18567
rect 11296 18508 12664 18536
rect 11296 18496 11302 18508
rect 5166 18468 5172 18480
rect 1544 18440 3832 18468
rect 5127 18440 5172 18468
rect 1544 18428 1550 18440
rect 5166 18428 5172 18440
rect 5224 18428 5230 18480
rect 7006 18428 7012 18480
rect 7064 18468 7070 18480
rect 12342 18468 12348 18480
rect 7064 18440 12348 18468
rect 7064 18428 7070 18440
rect 12342 18428 12348 18440
rect 12400 18428 12406 18480
rect 12636 18468 12664 18508
rect 13262 18468 13268 18480
rect 12636 18440 13268 18468
rect 13262 18428 13268 18440
rect 13320 18468 13326 18480
rect 14292 18468 14320 18567
rect 15304 18468 15332 18576
rect 15933 18573 15945 18576
rect 15979 18573 15991 18607
rect 15933 18567 15991 18573
rect 13320 18440 15332 18468
rect 15657 18471 15715 18477
rect 13320 18428 13326 18440
rect 15657 18437 15669 18471
rect 15703 18468 15715 18471
rect 16114 18468 16120 18480
rect 15703 18440 16120 18468
rect 15703 18437 15715 18440
rect 15657 18431 15715 18437
rect 16114 18428 16120 18440
rect 16172 18428 16178 18480
rect 17310 18468 17316 18480
rect 17271 18440 17316 18468
rect 17310 18428 17316 18440
rect 17368 18428 17374 18480
rect 17494 18428 17500 18480
rect 17552 18468 17558 18480
rect 20990 18468 20996 18480
rect 17552 18440 20996 18468
rect 17552 18428 17558 18440
rect 20990 18428 20996 18440
rect 21048 18428 21054 18480
rect 1104 18378 21620 18400
rect 1104 18326 4414 18378
rect 4466 18326 4478 18378
rect 4530 18326 4542 18378
rect 4594 18326 4606 18378
rect 4658 18326 11278 18378
rect 11330 18326 11342 18378
rect 11394 18326 11406 18378
rect 11458 18326 11470 18378
rect 11522 18326 18142 18378
rect 18194 18326 18206 18378
rect 18258 18326 18270 18378
rect 18322 18326 18334 18378
rect 18386 18326 21620 18378
rect 1104 18304 21620 18326
rect 4982 18224 4988 18276
rect 5040 18264 5046 18276
rect 5040 18236 5764 18264
rect 5040 18224 5046 18236
rect 2774 18088 2780 18140
rect 2832 18128 2838 18140
rect 3329 18131 3387 18137
rect 3329 18128 3341 18131
rect 2832 18100 3341 18128
rect 2832 18088 2838 18100
rect 3329 18097 3341 18100
rect 3375 18097 3387 18131
rect 5074 18128 5080 18140
rect 5035 18100 5080 18128
rect 3329 18091 3387 18097
rect 5074 18088 5080 18100
rect 5132 18088 5138 18140
rect 290 18020 296 18072
rect 348 18060 354 18072
rect 5736 18060 5764 18236
rect 7098 18224 7104 18276
rect 7156 18264 7162 18276
rect 7285 18267 7343 18273
rect 7285 18264 7297 18267
rect 7156 18236 7297 18264
rect 7156 18224 7162 18236
rect 7285 18233 7297 18236
rect 7331 18233 7343 18267
rect 7285 18227 7343 18233
rect 7745 18267 7803 18273
rect 7745 18233 7757 18267
rect 7791 18264 7803 18267
rect 8294 18264 8300 18276
rect 7791 18236 8300 18264
rect 7791 18233 7803 18236
rect 7745 18227 7803 18233
rect 7300 18196 7328 18227
rect 8294 18224 8300 18236
rect 8352 18224 8358 18276
rect 11698 18264 11704 18276
rect 9692 18236 11704 18264
rect 7300 18168 8064 18196
rect 8036 18128 8064 18168
rect 8110 18156 8116 18208
rect 8168 18196 8174 18208
rect 9692 18196 9720 18236
rect 11698 18224 11704 18236
rect 11756 18224 11762 18276
rect 12345 18267 12403 18273
rect 12345 18233 12357 18267
rect 12391 18264 12403 18267
rect 14090 18264 14096 18276
rect 12391 18236 14096 18264
rect 12391 18233 12403 18236
rect 12345 18227 12403 18233
rect 14090 18224 14096 18236
rect 14148 18224 14154 18276
rect 18690 18264 18696 18276
rect 18651 18236 18696 18264
rect 18690 18224 18696 18236
rect 18748 18224 18754 18276
rect 19610 18264 19616 18276
rect 19571 18236 19616 18264
rect 19610 18224 19616 18236
rect 19668 18224 19674 18276
rect 20162 18264 20168 18276
rect 20123 18236 20168 18264
rect 20162 18224 20168 18236
rect 20220 18224 20226 18276
rect 8168 18168 9720 18196
rect 8168 18156 8174 18168
rect 9766 18156 9772 18208
rect 9824 18196 9830 18208
rect 9824 18168 12572 18196
rect 9824 18156 9830 18168
rect 8297 18131 8355 18137
rect 8297 18128 8309 18131
rect 8036 18100 8309 18128
rect 8297 18097 8309 18100
rect 8343 18097 8355 18131
rect 8297 18091 8355 18097
rect 9674 18088 9680 18140
rect 9732 18128 9738 18140
rect 11333 18131 11391 18137
rect 11333 18128 11345 18131
rect 9732 18100 11345 18128
rect 9732 18088 9738 18100
rect 11333 18097 11345 18100
rect 11379 18097 11391 18131
rect 11333 18091 11391 18097
rect 11517 18131 11575 18137
rect 11517 18097 11529 18131
rect 11563 18128 11575 18131
rect 11606 18128 11612 18140
rect 11563 18100 11612 18128
rect 11563 18097 11575 18100
rect 11517 18091 11575 18097
rect 11606 18088 11612 18100
rect 11664 18088 11670 18140
rect 5905 18063 5963 18069
rect 5905 18060 5917 18063
rect 348 18032 5580 18060
rect 5736 18032 5917 18060
rect 348 18020 354 18032
rect 3050 17952 3056 18004
rect 3108 17992 3114 18004
rect 3108 17964 5488 17992
rect 3108 17952 3114 17964
rect 5460 17936 5488 17964
rect 1394 17884 1400 17936
rect 1452 17924 1458 17936
rect 2682 17924 2688 17936
rect 1452 17896 2688 17924
rect 1452 17884 1458 17896
rect 2682 17884 2688 17896
rect 2740 17884 2746 17936
rect 2777 17927 2835 17933
rect 2777 17893 2789 17927
rect 2823 17924 2835 17927
rect 2958 17924 2964 17936
rect 2823 17896 2964 17924
rect 2823 17893 2835 17896
rect 2777 17887 2835 17893
rect 2958 17884 2964 17896
rect 3016 17884 3022 17936
rect 3142 17924 3148 17936
rect 3103 17896 3148 17924
rect 3142 17884 3148 17896
rect 3200 17884 3206 17936
rect 3234 17884 3240 17936
rect 3292 17924 3298 17936
rect 3292 17896 3337 17924
rect 3292 17884 3298 17896
rect 5442 17884 5448 17936
rect 5500 17884 5506 17936
rect 5552 17924 5580 18032
rect 5905 18029 5917 18032
rect 5951 18060 5963 18063
rect 6546 18060 6552 18072
rect 5951 18032 6552 18060
rect 5951 18029 5963 18032
rect 5905 18023 5963 18029
rect 6546 18020 6552 18032
rect 6604 18020 6610 18072
rect 7650 18020 7656 18072
rect 7708 18060 7714 18072
rect 8113 18063 8171 18069
rect 8113 18060 8125 18063
rect 7708 18032 8125 18060
rect 7708 18020 7714 18032
rect 8113 18029 8125 18032
rect 8159 18029 8171 18063
rect 8113 18023 8171 18029
rect 8205 18063 8263 18069
rect 8205 18029 8217 18063
rect 8251 18060 8263 18063
rect 8570 18060 8576 18072
rect 8251 18032 8576 18060
rect 8251 18029 8263 18032
rect 8205 18023 8263 18029
rect 8570 18020 8576 18032
rect 8628 18020 8634 18072
rect 11054 18060 11060 18072
rect 10796 18032 11060 18060
rect 6172 17995 6230 18001
rect 6172 17961 6184 17995
rect 6218 17992 6230 17995
rect 6362 17992 6368 18004
rect 6218 17964 6368 17992
rect 6218 17961 6230 17964
rect 6172 17955 6230 17961
rect 6362 17952 6368 17964
rect 6420 17952 6426 18004
rect 6454 17952 6460 18004
rect 6512 17992 6518 18004
rect 10796 17992 10824 18032
rect 11054 18020 11060 18032
rect 11112 18020 11118 18072
rect 11241 18063 11299 18069
rect 11241 18029 11253 18063
rect 11287 18060 11299 18063
rect 11790 18060 11796 18072
rect 11287 18032 11796 18060
rect 11287 18029 11299 18032
rect 11241 18023 11299 18029
rect 11790 18020 11796 18032
rect 11848 18020 11854 18072
rect 12544 18060 12572 18168
rect 12710 18156 12716 18208
rect 12768 18196 12774 18208
rect 17218 18196 17224 18208
rect 12768 18168 17224 18196
rect 12768 18156 12774 18168
rect 17218 18156 17224 18168
rect 17276 18156 17282 18208
rect 18506 18156 18512 18208
rect 18564 18196 18570 18208
rect 19334 18196 19340 18208
rect 18564 18168 19340 18196
rect 18564 18156 18570 18168
rect 19334 18156 19340 18168
rect 19392 18156 19398 18208
rect 12618 18088 12624 18140
rect 12676 18128 12682 18140
rect 12897 18131 12955 18137
rect 12897 18128 12909 18131
rect 12676 18100 12909 18128
rect 12676 18088 12682 18100
rect 12897 18097 12909 18100
rect 12943 18097 12955 18131
rect 13906 18128 13912 18140
rect 13867 18100 13912 18128
rect 12897 18091 12955 18097
rect 13906 18088 13912 18100
rect 13964 18088 13970 18140
rect 17402 18128 17408 18140
rect 17363 18100 17408 18128
rect 17402 18088 17408 18100
rect 17460 18088 17466 18140
rect 19610 18088 19616 18140
rect 19668 18128 19674 18140
rect 21358 18128 21364 18140
rect 19668 18100 21364 18128
rect 19668 18088 19674 18100
rect 21358 18088 21364 18100
rect 21416 18088 21422 18140
rect 12805 18063 12863 18069
rect 12805 18060 12817 18063
rect 12544 18032 12817 18060
rect 12805 18029 12817 18032
rect 12851 18029 12863 18063
rect 12805 18023 12863 18029
rect 16298 18020 16304 18072
rect 16356 18060 16362 18072
rect 17129 18063 17187 18069
rect 17129 18060 17141 18063
rect 16356 18032 17141 18060
rect 16356 18020 16362 18032
rect 17129 18029 17141 18032
rect 17175 18029 17187 18063
rect 18506 18060 18512 18072
rect 18467 18032 18512 18060
rect 17129 18023 17187 18029
rect 18506 18020 18512 18032
rect 18564 18020 18570 18072
rect 19426 18060 19432 18072
rect 19387 18032 19432 18060
rect 19426 18020 19432 18032
rect 19484 18020 19490 18072
rect 19978 18060 19984 18072
rect 19939 18032 19984 18060
rect 19978 18020 19984 18032
rect 20036 18020 20042 18072
rect 19518 17992 19524 18004
rect 6512 17964 10824 17992
rect 10888 17964 19524 17992
rect 6512 17952 6518 17964
rect 10778 17924 10784 17936
rect 5552 17896 10784 17924
rect 10778 17884 10784 17896
rect 10836 17884 10842 17936
rect 10888 17933 10916 17964
rect 19518 17952 19524 17964
rect 19576 17952 19582 18004
rect 21082 17952 21088 18004
rect 21140 17992 21146 18004
rect 22462 17992 22468 18004
rect 21140 17964 22468 17992
rect 21140 17952 21146 17964
rect 22462 17952 22468 17964
rect 22520 17952 22526 18004
rect 10873 17927 10931 17933
rect 10873 17893 10885 17927
rect 10919 17893 10931 17927
rect 10873 17887 10931 17893
rect 10962 17884 10968 17936
rect 11020 17924 11026 17936
rect 12713 17927 12771 17933
rect 12713 17924 12725 17927
rect 11020 17896 12725 17924
rect 11020 17884 11026 17896
rect 12713 17893 12725 17896
rect 12759 17893 12771 17927
rect 12713 17887 12771 17893
rect 14182 17884 14188 17936
rect 14240 17924 14246 17936
rect 15102 17924 15108 17936
rect 14240 17896 15108 17924
rect 14240 17884 14246 17896
rect 15102 17884 15108 17896
rect 15160 17884 15166 17936
rect 15286 17884 15292 17936
rect 15344 17924 15350 17936
rect 16206 17924 16212 17936
rect 15344 17896 16212 17924
rect 15344 17884 15350 17896
rect 16206 17884 16212 17896
rect 16264 17884 16270 17936
rect 16942 17884 16948 17936
rect 17000 17924 17006 17936
rect 19794 17924 19800 17936
rect 17000 17896 19800 17924
rect 17000 17884 17006 17896
rect 19794 17884 19800 17896
rect 19852 17884 19858 17936
rect 20530 17884 20536 17936
rect 20588 17924 20594 17936
rect 21910 17924 21916 17936
rect 20588 17896 21916 17924
rect 20588 17884 20594 17896
rect 21910 17884 21916 17896
rect 21968 17884 21974 17936
rect 14 17816 20 17868
rect 72 17856 78 17868
rect 842 17856 848 17868
rect 72 17828 848 17856
rect 72 17816 78 17828
rect 842 17816 848 17828
rect 900 17816 906 17868
rect 1104 17834 21620 17856
rect 1104 17782 7846 17834
rect 7898 17782 7910 17834
rect 7962 17782 7974 17834
rect 8026 17782 8038 17834
rect 8090 17782 14710 17834
rect 14762 17782 14774 17834
rect 14826 17782 14838 17834
rect 14890 17782 14902 17834
rect 14954 17782 21620 17834
rect 1104 17760 21620 17782
rect 2774 17680 2780 17732
rect 2832 17720 2838 17732
rect 2832 17692 2877 17720
rect 2832 17680 2838 17692
rect 3234 17680 3240 17732
rect 3292 17720 3298 17732
rect 3421 17723 3479 17729
rect 3421 17720 3433 17723
rect 3292 17692 3433 17720
rect 3292 17680 3298 17692
rect 3421 17689 3433 17692
rect 3467 17689 3479 17723
rect 3421 17683 3479 17689
rect 3881 17723 3939 17729
rect 3881 17689 3893 17723
rect 3927 17720 3939 17723
rect 4154 17720 4160 17732
rect 3927 17692 4160 17720
rect 3927 17689 3939 17692
rect 3881 17683 3939 17689
rect 4154 17680 4160 17692
rect 4212 17680 4218 17732
rect 4706 17680 4712 17732
rect 4764 17720 4770 17732
rect 20162 17720 20168 17732
rect 4764 17692 20168 17720
rect 4764 17680 4770 17692
rect 20162 17680 20168 17692
rect 20220 17680 20226 17732
rect 3789 17655 3847 17661
rect 3789 17621 3801 17655
rect 3835 17652 3847 17655
rect 7650 17652 7656 17664
rect 3835 17624 7656 17652
rect 3835 17621 3847 17624
rect 3789 17615 3847 17621
rect 7650 17612 7656 17624
rect 7708 17612 7714 17664
rect 18325 17655 18383 17661
rect 18325 17621 18337 17655
rect 18371 17652 18383 17655
rect 18506 17652 18512 17664
rect 18371 17624 18512 17652
rect 18371 17621 18383 17624
rect 18325 17615 18383 17621
rect 18506 17612 18512 17624
rect 18564 17612 18570 17664
rect 1397 17587 1455 17593
rect 1397 17553 1409 17587
rect 1443 17584 1455 17587
rect 1486 17584 1492 17596
rect 1443 17556 1492 17584
rect 1443 17553 1455 17556
rect 1397 17547 1455 17553
rect 1486 17544 1492 17556
rect 1544 17544 1550 17596
rect 1664 17587 1722 17593
rect 1664 17553 1676 17587
rect 1710 17584 1722 17587
rect 3418 17584 3424 17596
rect 1710 17556 3424 17584
rect 1710 17553 1722 17556
rect 1664 17547 1722 17553
rect 3418 17544 3424 17556
rect 3476 17584 3482 17596
rect 3476 17556 4016 17584
rect 3476 17544 3482 17556
rect 3988 17525 4016 17556
rect 12342 17544 12348 17596
rect 12400 17584 12406 17596
rect 12710 17584 12716 17596
rect 12400 17556 12716 17584
rect 12400 17544 12406 17556
rect 12710 17544 12716 17556
rect 12768 17544 12774 17596
rect 17954 17544 17960 17596
rect 18012 17584 18018 17596
rect 18049 17587 18107 17593
rect 18049 17584 18061 17587
rect 18012 17556 18061 17584
rect 18012 17544 18018 17556
rect 18049 17553 18061 17556
rect 18095 17553 18107 17587
rect 18049 17547 18107 17553
rect 19429 17587 19487 17593
rect 19429 17553 19441 17587
rect 19475 17553 19487 17587
rect 19429 17547 19487 17553
rect 19705 17587 19763 17593
rect 19705 17553 19717 17587
rect 19751 17584 19763 17587
rect 20533 17587 20591 17593
rect 20533 17584 20545 17587
rect 19751 17556 20545 17584
rect 19751 17553 19763 17556
rect 19705 17547 19763 17553
rect 20533 17553 20545 17556
rect 20579 17553 20591 17587
rect 20533 17547 20591 17553
rect 3973 17519 4031 17525
rect 3973 17485 3985 17519
rect 4019 17485 4031 17519
rect 3973 17479 4031 17485
rect 4890 17476 4896 17528
rect 4948 17516 4954 17528
rect 19444 17516 19472 17547
rect 4948 17488 19472 17516
rect 4948 17476 4954 17488
rect 7558 17408 7564 17460
rect 7616 17448 7622 17460
rect 19426 17448 19432 17460
rect 7616 17420 19432 17448
rect 7616 17408 7622 17420
rect 19426 17408 19432 17420
rect 19484 17408 19490 17460
rect 10870 17340 10876 17392
rect 10928 17380 10934 17392
rect 16666 17380 16672 17392
rect 10928 17352 16672 17380
rect 10928 17340 10934 17352
rect 16666 17340 16672 17352
rect 16724 17340 16730 17392
rect 20714 17380 20720 17392
rect 20675 17352 20720 17380
rect 20714 17340 20720 17352
rect 20772 17340 20778 17392
rect 1104 17290 21620 17312
rect 1104 17238 4414 17290
rect 4466 17238 4478 17290
rect 4530 17238 4542 17290
rect 4594 17238 4606 17290
rect 4658 17238 11278 17290
rect 11330 17238 11342 17290
rect 11394 17238 11406 17290
rect 11458 17238 11470 17290
rect 11522 17238 18142 17290
rect 18194 17238 18206 17290
rect 18258 17238 18270 17290
rect 18322 17238 18334 17290
rect 18386 17238 21620 17290
rect 1104 17216 21620 17238
rect 4062 17136 4068 17188
rect 4120 17176 4126 17188
rect 17678 17176 17684 17188
rect 4120 17148 17684 17176
rect 4120 17136 4126 17148
rect 17678 17136 17684 17148
rect 17736 17176 17742 17188
rect 17773 17179 17831 17185
rect 17773 17176 17785 17179
rect 17736 17148 17785 17176
rect 17736 17136 17742 17148
rect 17773 17145 17785 17148
rect 17819 17145 17831 17179
rect 18690 17176 18696 17188
rect 18651 17148 18696 17176
rect 17773 17139 17831 17145
rect 18690 17136 18696 17148
rect 18748 17136 18754 17188
rect 20438 17176 20444 17188
rect 20399 17148 20444 17176
rect 20438 17136 20444 17148
rect 20496 17136 20502 17188
rect 6181 17111 6239 17117
rect 6181 17077 6193 17111
rect 6227 17108 6239 17111
rect 6227 17080 8892 17108
rect 6227 17077 6239 17080
rect 6181 17071 6239 17077
rect 3142 17040 3148 17052
rect 3103 17012 3148 17040
rect 3142 17000 3148 17012
rect 3200 17000 3206 17052
rect 4341 17043 4399 17049
rect 4341 17009 4353 17043
rect 4387 17040 4399 17043
rect 4706 17040 4712 17052
rect 4387 17012 4712 17040
rect 4387 17009 4399 17012
rect 4341 17003 4399 17009
rect 4706 17000 4712 17012
rect 4764 17000 4770 17052
rect 7558 17040 7564 17052
rect 7519 17012 7564 17040
rect 7558 17000 7564 17012
rect 7616 17000 7622 17052
rect 8754 17000 8760 17052
rect 8812 17040 8818 17052
rect 8864 17049 8892 17080
rect 8849 17043 8907 17049
rect 8849 17040 8861 17043
rect 8812 17012 8861 17040
rect 8812 17000 8818 17012
rect 8849 17009 8861 17012
rect 8895 17009 8907 17043
rect 8849 17003 8907 17009
rect 19337 17043 19395 17049
rect 19337 17009 19349 17043
rect 19383 17040 19395 17043
rect 19978 17040 19984 17052
rect 19383 17012 19984 17040
rect 19383 17009 19395 17012
rect 19337 17003 19395 17009
rect 19978 17000 19984 17012
rect 20036 17000 20042 17052
rect 2958 16932 2964 16984
rect 3016 16972 3022 16984
rect 4065 16975 4123 16981
rect 4065 16972 4077 16975
rect 3016 16944 4077 16972
rect 3016 16932 3022 16944
rect 4065 16941 4077 16944
rect 4111 16941 4123 16975
rect 4065 16935 4123 16941
rect 4801 16975 4859 16981
rect 4801 16941 4813 16975
rect 4847 16972 4859 16975
rect 4890 16972 4896 16984
rect 4847 16944 4896 16972
rect 4847 16941 4859 16944
rect 4801 16935 4859 16941
rect 4890 16932 4896 16944
rect 4948 16932 4954 16984
rect 6822 16932 6828 16984
rect 6880 16972 6886 16984
rect 7285 16975 7343 16981
rect 7285 16972 7297 16975
rect 6880 16944 7297 16972
rect 6880 16932 6886 16944
rect 7285 16941 7297 16944
rect 7331 16941 7343 16975
rect 7285 16935 7343 16941
rect 11054 16932 11060 16984
rect 11112 16972 11118 16984
rect 13354 16972 13360 16984
rect 11112 16944 13360 16972
rect 11112 16932 11118 16944
rect 13354 16932 13360 16944
rect 13412 16932 13418 16984
rect 15470 16932 15476 16984
rect 15528 16972 15534 16984
rect 16393 16975 16451 16981
rect 16393 16972 16405 16975
rect 15528 16944 16405 16972
rect 15528 16932 15534 16944
rect 16393 16941 16405 16944
rect 16439 16941 16451 16975
rect 18506 16972 18512 16984
rect 18467 16944 18512 16972
rect 16393 16935 16451 16941
rect 18506 16932 18512 16944
rect 18564 16932 18570 16984
rect 19058 16972 19064 16984
rect 19019 16944 19064 16972
rect 19058 16932 19064 16944
rect 19116 16932 19122 16984
rect 19518 16932 19524 16984
rect 19576 16972 19582 16984
rect 20257 16975 20315 16981
rect 20257 16972 20269 16975
rect 19576 16944 20269 16972
rect 19576 16932 19582 16944
rect 20257 16941 20269 16944
rect 20303 16941 20315 16975
rect 20257 16935 20315 16941
rect 5068 16907 5126 16913
rect 5068 16873 5080 16907
rect 5114 16904 5126 16907
rect 5166 16904 5172 16916
rect 5114 16876 5172 16904
rect 5114 16873 5126 16876
rect 5068 16867 5126 16873
rect 5166 16864 5172 16876
rect 5224 16864 5230 16916
rect 5534 16864 5540 16916
rect 5592 16904 5598 16916
rect 8757 16907 8815 16913
rect 8757 16904 8769 16907
rect 5592 16876 8769 16904
rect 5592 16864 5598 16876
rect 8757 16873 8769 16876
rect 8803 16873 8815 16907
rect 10962 16904 10968 16916
rect 8757 16867 8815 16873
rect 9692 16876 10968 16904
rect 9692 16848 9720 16876
rect 10962 16864 10968 16876
rect 11020 16864 11026 16916
rect 11698 16864 11704 16916
rect 11756 16904 11762 16916
rect 15654 16904 15660 16916
rect 11756 16876 15660 16904
rect 11756 16864 11762 16876
rect 15654 16864 15660 16876
rect 15712 16864 15718 16916
rect 16660 16907 16718 16913
rect 16660 16873 16672 16907
rect 16706 16904 16718 16907
rect 16850 16904 16856 16916
rect 16706 16876 16856 16904
rect 16706 16873 16718 16876
rect 16660 16867 16718 16873
rect 16850 16864 16856 16876
rect 16908 16864 16914 16916
rect 19978 16904 19984 16916
rect 17696 16876 19984 16904
rect 8294 16836 8300 16848
rect 8255 16808 8300 16836
rect 8294 16796 8300 16808
rect 8352 16796 8358 16848
rect 8665 16839 8723 16845
rect 8665 16805 8677 16839
rect 8711 16836 8723 16839
rect 9674 16836 9680 16848
rect 8711 16808 9680 16836
rect 8711 16805 8723 16808
rect 8665 16799 8723 16805
rect 9674 16796 9680 16808
rect 9732 16836 9738 16848
rect 9861 16839 9919 16845
rect 9732 16808 9825 16836
rect 9732 16796 9738 16808
rect 9861 16805 9873 16839
rect 9907 16836 9919 16839
rect 10502 16836 10508 16848
rect 9907 16808 10508 16836
rect 9907 16805 9919 16808
rect 9861 16799 9919 16805
rect 10502 16796 10508 16808
rect 10560 16796 10566 16848
rect 12434 16796 12440 16848
rect 12492 16836 12498 16848
rect 17696 16836 17724 16876
rect 19978 16864 19984 16876
rect 20036 16864 20042 16916
rect 12492 16808 17724 16836
rect 12492 16796 12498 16808
rect 1104 16746 21620 16768
rect 1104 16694 7846 16746
rect 7898 16694 7910 16746
rect 7962 16694 7974 16746
rect 8026 16694 8038 16746
rect 8090 16694 14710 16746
rect 14762 16694 14774 16746
rect 14826 16694 14838 16746
rect 14890 16694 14902 16746
rect 14954 16694 21620 16746
rect 1104 16672 21620 16694
rect 6822 16632 6828 16644
rect 6783 16604 6828 16632
rect 6822 16592 6828 16604
rect 6880 16592 6886 16644
rect 10502 16632 10508 16644
rect 10463 16604 10508 16632
rect 10502 16592 10508 16604
rect 10560 16592 10566 16644
rect 11333 16635 11391 16641
rect 11333 16601 11345 16635
rect 11379 16601 11391 16635
rect 11698 16632 11704 16644
rect 11659 16604 11704 16632
rect 11333 16595 11391 16601
rect 8294 16524 8300 16576
rect 8352 16564 8358 16576
rect 10597 16567 10655 16573
rect 10597 16564 10609 16567
rect 8352 16536 10609 16564
rect 8352 16524 8358 16536
rect 10597 16533 10609 16536
rect 10643 16533 10655 16567
rect 11348 16564 11376 16595
rect 11698 16592 11704 16604
rect 11756 16592 11762 16644
rect 12897 16635 12955 16641
rect 12897 16632 12909 16635
rect 11808 16604 12909 16632
rect 11808 16564 11836 16604
rect 12897 16601 12909 16604
rect 12943 16601 12955 16635
rect 12897 16595 12955 16601
rect 13354 16592 13360 16644
rect 13412 16632 13418 16644
rect 14369 16635 14427 16641
rect 14369 16632 14381 16635
rect 13412 16604 14381 16632
rect 13412 16592 13418 16604
rect 14369 16601 14381 16604
rect 14415 16601 14427 16635
rect 16850 16632 16856 16644
rect 16811 16604 16856 16632
rect 14369 16595 14427 16601
rect 16850 16592 16856 16604
rect 16908 16592 16914 16644
rect 18506 16592 18512 16644
rect 18564 16632 18570 16644
rect 18564 16604 20300 16632
rect 18564 16592 18570 16604
rect 19518 16564 19524 16576
rect 11348 16536 11836 16564
rect 13740 16536 17448 16564
rect 19479 16536 19524 16564
rect 10597 16527 10655 16533
rect 7193 16499 7251 16505
rect 7193 16465 7205 16499
rect 7239 16496 7251 16499
rect 7837 16499 7895 16505
rect 7837 16496 7849 16499
rect 7239 16468 7849 16496
rect 7239 16465 7251 16468
rect 7193 16459 7251 16465
rect 7837 16465 7849 16468
rect 7883 16465 7895 16499
rect 8478 16496 8484 16508
rect 8439 16468 8484 16496
rect 7837 16459 7895 16465
rect 8478 16456 8484 16468
rect 8536 16456 8542 16508
rect 8754 16505 8760 16508
rect 8748 16496 8760 16505
rect 8715 16468 8760 16496
rect 8748 16459 8760 16468
rect 8754 16456 8760 16459
rect 8812 16456 8818 16508
rect 12805 16499 12863 16505
rect 12805 16465 12817 16499
rect 12851 16496 12863 16499
rect 13449 16499 13507 16505
rect 13449 16496 13461 16499
rect 12851 16468 13461 16496
rect 12851 16465 12863 16468
rect 12805 16459 12863 16465
rect 13449 16465 13461 16468
rect 13495 16465 13507 16499
rect 13449 16459 13507 16465
rect 7282 16428 7288 16440
rect 7243 16400 7288 16428
rect 7282 16388 7288 16400
rect 7340 16388 7346 16440
rect 7377 16431 7435 16437
rect 7377 16397 7389 16431
rect 7423 16397 7435 16431
rect 7377 16391 7435 16397
rect 10689 16431 10747 16437
rect 10689 16397 10701 16431
rect 10735 16397 10747 16431
rect 11790 16428 11796 16440
rect 11751 16400 11796 16428
rect 10689 16391 10747 16397
rect 6362 16320 6368 16372
rect 6420 16360 6426 16372
rect 7392 16360 7420 16391
rect 10704 16360 10732 16391
rect 11790 16388 11796 16400
rect 11848 16388 11854 16440
rect 11882 16388 11888 16440
rect 11940 16428 11946 16440
rect 12986 16428 12992 16440
rect 11940 16400 11985 16428
rect 12947 16400 12992 16428
rect 11940 16388 11946 16400
rect 12986 16388 12992 16400
rect 13044 16388 13050 16440
rect 6420 16332 7420 16360
rect 10060 16332 10732 16360
rect 6420 16320 6426 16332
rect 10060 16304 10088 16332
rect 12434 16320 12440 16372
rect 12492 16360 12498 16372
rect 12492 16332 12537 16360
rect 12492 16320 12498 16332
rect 2498 16252 2504 16304
rect 2556 16292 2562 16304
rect 8846 16292 8852 16304
rect 2556 16264 8852 16292
rect 2556 16252 2562 16264
rect 8846 16252 8852 16264
rect 8904 16252 8910 16304
rect 9861 16295 9919 16301
rect 9861 16261 9873 16295
rect 9907 16292 9919 16295
rect 10042 16292 10048 16304
rect 9907 16264 10048 16292
rect 9907 16261 9919 16264
rect 9861 16255 9919 16261
rect 10042 16252 10048 16264
rect 10100 16252 10106 16304
rect 10137 16295 10195 16301
rect 10137 16261 10149 16295
rect 10183 16292 10195 16295
rect 13740 16292 13768 16536
rect 14274 16496 14280 16508
rect 14235 16468 14280 16496
rect 14274 16456 14280 16468
rect 14332 16456 14338 16508
rect 15740 16499 15798 16505
rect 15740 16465 15752 16499
rect 15786 16496 15798 16499
rect 17310 16496 17316 16508
rect 15786 16468 17316 16496
rect 15786 16465 15798 16468
rect 15740 16459 15798 16465
rect 17310 16456 17316 16468
rect 17368 16456 17374 16508
rect 17420 16496 17448 16536
rect 19518 16524 19524 16536
rect 19576 16524 19582 16576
rect 20272 16573 20300 16604
rect 20622 16592 20628 16644
rect 20680 16632 20686 16644
rect 20901 16635 20959 16641
rect 20901 16632 20913 16635
rect 20680 16604 20913 16632
rect 20680 16592 20686 16604
rect 20901 16601 20913 16604
rect 20947 16601 20959 16635
rect 20901 16595 20959 16601
rect 20257 16567 20315 16573
rect 20257 16533 20269 16567
rect 20303 16533 20315 16567
rect 20257 16527 20315 16533
rect 19245 16499 19303 16505
rect 19245 16496 19257 16499
rect 17420 16468 19257 16496
rect 19245 16465 19257 16468
rect 19291 16465 19303 16499
rect 19978 16496 19984 16508
rect 19939 16468 19984 16496
rect 19245 16459 19303 16465
rect 19978 16456 19984 16468
rect 20036 16456 20042 16508
rect 20162 16456 20168 16508
rect 20220 16496 20226 16508
rect 20717 16499 20775 16505
rect 20717 16496 20729 16499
rect 20220 16468 20729 16496
rect 20220 16456 20226 16468
rect 20717 16465 20729 16468
rect 20763 16465 20775 16499
rect 20717 16459 20775 16465
rect 14458 16388 14464 16440
rect 14516 16428 14522 16440
rect 15470 16428 15476 16440
rect 14516 16400 14561 16428
rect 15431 16400 15476 16428
rect 14516 16388 14522 16400
rect 15470 16388 15476 16400
rect 15528 16388 15534 16440
rect 17954 16388 17960 16440
rect 18012 16428 18018 16440
rect 18049 16431 18107 16437
rect 18049 16428 18061 16431
rect 18012 16400 18061 16428
rect 18012 16388 18018 16400
rect 18049 16397 18061 16400
rect 18095 16397 18107 16431
rect 18049 16391 18107 16397
rect 13906 16292 13912 16304
rect 10183 16264 13768 16292
rect 13867 16264 13912 16292
rect 10183 16261 10195 16264
rect 10137 16255 10195 16261
rect 13906 16252 13912 16264
rect 13964 16252 13970 16304
rect 1104 16202 21620 16224
rect 1104 16150 4414 16202
rect 4466 16150 4478 16202
rect 4530 16150 4542 16202
rect 4594 16150 4606 16202
rect 4658 16150 11278 16202
rect 11330 16150 11342 16202
rect 11394 16150 11406 16202
rect 11458 16150 11470 16202
rect 11522 16150 18142 16202
rect 18194 16150 18206 16202
rect 18258 16150 18270 16202
rect 18322 16150 18334 16202
rect 18386 16150 21620 16202
rect 1104 16128 21620 16150
rect 3329 16091 3387 16097
rect 3329 16057 3341 16091
rect 3375 16088 3387 16091
rect 3418 16088 3424 16100
rect 3375 16060 3424 16088
rect 3375 16057 3387 16060
rect 3329 16051 3387 16057
rect 3418 16048 3424 16060
rect 3476 16048 3482 16100
rect 6362 16088 6368 16100
rect 6323 16060 6368 16088
rect 6362 16048 6368 16060
rect 6420 16048 6426 16100
rect 7009 16091 7067 16097
rect 7009 16057 7021 16091
rect 7055 16088 7067 16091
rect 7282 16088 7288 16100
rect 7055 16060 7288 16088
rect 7055 16057 7067 16060
rect 7009 16051 7067 16057
rect 7282 16048 7288 16060
rect 7340 16048 7346 16100
rect 12986 16088 12992 16100
rect 12947 16060 12992 16088
rect 12986 16048 12992 16060
rect 13044 16048 13050 16100
rect 17405 16091 17463 16097
rect 17405 16057 17417 16091
rect 17451 16088 17463 16091
rect 17862 16088 17868 16100
rect 17451 16060 17868 16088
rect 17451 16057 17463 16060
rect 17405 16051 17463 16057
rect 17862 16048 17868 16060
rect 17920 16048 17926 16100
rect 19242 16048 19248 16100
rect 19300 16088 19306 16100
rect 20441 16091 20499 16097
rect 20441 16088 20453 16091
rect 19300 16060 20453 16088
rect 19300 16048 19306 16060
rect 20441 16057 20453 16060
rect 20487 16057 20499 16091
rect 20441 16051 20499 16057
rect 1486 15912 1492 15964
rect 1544 15952 1550 15964
rect 1949 15955 2007 15961
rect 1949 15952 1961 15955
rect 1544 15924 1961 15952
rect 1544 15912 1550 15924
rect 1949 15921 1961 15924
rect 1995 15921 2007 15955
rect 4982 15952 4988 15964
rect 4943 15924 4988 15952
rect 1949 15915 2007 15921
rect 4982 15912 4988 15924
rect 5040 15912 5046 15964
rect 6362 15912 6368 15964
rect 6420 15952 6426 15964
rect 7561 15955 7619 15961
rect 7561 15952 7573 15955
rect 6420 15924 7573 15952
rect 6420 15912 6426 15924
rect 7561 15921 7573 15924
rect 7607 15921 7619 15955
rect 7561 15915 7619 15921
rect 8478 15912 8484 15964
rect 8536 15952 8542 15964
rect 9953 15955 10011 15961
rect 9953 15952 9965 15955
rect 8536 15924 9965 15952
rect 8536 15912 8542 15924
rect 9953 15921 9965 15924
rect 9999 15921 10011 15955
rect 13004 15952 13032 16048
rect 16393 16023 16451 16029
rect 16393 15989 16405 16023
rect 16439 16020 16451 16023
rect 16439 15992 17908 16020
rect 16439 15989 16451 15992
rect 16393 15983 16451 15989
rect 13004 15924 13400 15952
rect 9953 15915 10011 15921
rect 5252 15887 5310 15893
rect 5252 15853 5264 15887
rect 5298 15884 5310 15887
rect 6380 15884 6408 15912
rect 7374 15884 7380 15896
rect 5298 15856 6408 15884
rect 7335 15856 7380 15884
rect 5298 15853 5310 15856
rect 5252 15847 5310 15853
rect 7374 15844 7380 15856
rect 7432 15844 7438 15896
rect 7469 15887 7527 15893
rect 7469 15853 7481 15887
rect 7515 15884 7527 15887
rect 7742 15884 7748 15896
rect 7515 15856 7748 15884
rect 7515 15853 7527 15856
rect 7469 15847 7527 15853
rect 7742 15844 7748 15856
rect 7800 15844 7806 15896
rect 10042 15844 10048 15896
rect 10100 15884 10106 15896
rect 10209 15887 10267 15893
rect 10209 15884 10221 15887
rect 10100 15856 10221 15884
rect 10100 15844 10106 15856
rect 10209 15853 10221 15856
rect 10255 15853 10267 15887
rect 10209 15847 10267 15853
rect 10686 15844 10692 15896
rect 10744 15884 10750 15896
rect 11882 15893 11888 15896
rect 11609 15887 11667 15893
rect 11609 15884 11621 15887
rect 10744 15856 11621 15884
rect 10744 15844 10750 15856
rect 11609 15853 11621 15856
rect 11655 15853 11667 15887
rect 11876 15884 11888 15893
rect 11609 15847 11667 15853
rect 11808 15856 11888 15884
rect 2216 15819 2274 15825
rect 2216 15785 2228 15819
rect 2262 15816 2274 15819
rect 2866 15816 2872 15828
rect 2262 15788 2872 15816
rect 2262 15785 2274 15788
rect 2216 15779 2274 15785
rect 2866 15776 2872 15788
rect 2924 15776 2930 15828
rect 7558 15776 7564 15828
rect 7616 15816 7622 15828
rect 11514 15816 11520 15828
rect 7616 15788 11520 15816
rect 7616 15776 7622 15788
rect 11514 15776 11520 15788
rect 11572 15776 11578 15828
rect 11333 15751 11391 15757
rect 11333 15717 11345 15751
rect 11379 15748 11391 15751
rect 11808 15748 11836 15856
rect 11876 15847 11888 15856
rect 11882 15844 11888 15847
rect 11940 15844 11946 15896
rect 13262 15884 13268 15896
rect 13223 15856 13268 15884
rect 13262 15844 13268 15856
rect 13320 15844 13326 15896
rect 13372 15884 13400 15924
rect 16850 15912 16856 15964
rect 16908 15952 16914 15964
rect 17880 15961 17908 15992
rect 19150 15980 19156 16032
rect 19208 16020 19214 16032
rect 19889 16023 19947 16029
rect 19889 16020 19901 16023
rect 19208 15992 19901 16020
rect 19208 15980 19214 15992
rect 19889 15989 19901 15992
rect 19935 15989 19947 16023
rect 19889 15983 19947 15989
rect 16945 15955 17003 15961
rect 16945 15952 16957 15955
rect 16908 15924 16957 15952
rect 16908 15912 16914 15924
rect 16945 15921 16957 15924
rect 16991 15921 17003 15955
rect 16945 15915 17003 15921
rect 17865 15955 17923 15961
rect 17865 15921 17877 15955
rect 17911 15921 17923 15955
rect 17865 15915 17923 15921
rect 17957 15955 18015 15961
rect 17957 15921 17969 15955
rect 18003 15921 18015 15955
rect 17957 15915 18015 15921
rect 13521 15887 13579 15893
rect 13521 15884 13533 15887
rect 13372 15856 13533 15884
rect 13521 15853 13533 15856
rect 13567 15853 13579 15887
rect 13521 15847 13579 15853
rect 17678 15844 17684 15896
rect 17736 15884 17742 15896
rect 17972 15884 18000 15915
rect 19702 15884 19708 15896
rect 17736 15856 18000 15884
rect 19663 15856 19708 15884
rect 17736 15844 17742 15856
rect 19702 15844 19708 15856
rect 19760 15844 19766 15896
rect 20254 15884 20260 15896
rect 20215 15856 20260 15884
rect 20254 15844 20260 15856
rect 20312 15844 20318 15896
rect 14274 15776 14280 15828
rect 14332 15816 14338 15828
rect 16761 15819 16819 15825
rect 16761 15816 16773 15819
rect 14332 15788 16773 15816
rect 14332 15776 14338 15788
rect 16761 15785 16773 15788
rect 16807 15785 16819 15819
rect 16761 15779 16819 15785
rect 17773 15819 17831 15825
rect 17773 15785 17785 15819
rect 17819 15816 17831 15819
rect 17954 15816 17960 15828
rect 17819 15788 17960 15816
rect 17819 15785 17831 15788
rect 17773 15779 17831 15785
rect 17954 15776 17960 15788
rect 18012 15776 18018 15828
rect 11379 15720 11836 15748
rect 11379 15717 11391 15720
rect 11333 15711 11391 15717
rect 14458 15708 14464 15760
rect 14516 15748 14522 15760
rect 14645 15751 14703 15757
rect 14645 15748 14657 15751
rect 14516 15720 14657 15748
rect 14516 15708 14522 15720
rect 14645 15717 14657 15720
rect 14691 15717 14703 15751
rect 15286 15748 15292 15760
rect 15247 15720 15292 15748
rect 14645 15711 14703 15717
rect 15286 15708 15292 15720
rect 15344 15708 15350 15760
rect 16666 15708 16672 15760
rect 16724 15748 16730 15760
rect 16853 15751 16911 15757
rect 16853 15748 16865 15751
rect 16724 15720 16865 15748
rect 16724 15708 16730 15720
rect 16853 15717 16865 15720
rect 16899 15717 16911 15751
rect 16853 15711 16911 15717
rect 1104 15658 21620 15680
rect 1104 15606 7846 15658
rect 7898 15606 7910 15658
rect 7962 15606 7974 15658
rect 8026 15606 8038 15658
rect 8090 15606 14710 15658
rect 14762 15606 14774 15658
rect 14826 15606 14838 15658
rect 14890 15606 14902 15658
rect 14954 15606 21620 15658
rect 1104 15584 21620 15606
rect 2777 15547 2835 15553
rect 2777 15513 2789 15547
rect 2823 15544 2835 15547
rect 3329 15547 3387 15553
rect 3329 15544 3341 15547
rect 2823 15516 3341 15544
rect 2823 15513 2835 15516
rect 2777 15507 2835 15513
rect 3329 15513 3341 15516
rect 3375 15513 3387 15547
rect 3329 15507 3387 15513
rect 3602 15504 3608 15556
rect 3660 15544 3666 15556
rect 3789 15547 3847 15553
rect 3789 15544 3801 15547
rect 3660 15516 3801 15544
rect 3660 15504 3666 15516
rect 3789 15513 3801 15516
rect 3835 15513 3847 15547
rect 3789 15507 3847 15513
rect 14737 15547 14795 15553
rect 14737 15513 14749 15547
rect 14783 15544 14795 15547
rect 15286 15544 15292 15556
rect 14783 15516 15292 15544
rect 14783 15513 14795 15516
rect 14737 15507 14795 15513
rect 15286 15504 15292 15516
rect 15344 15504 15350 15556
rect 20162 15544 20168 15556
rect 20123 15516 20168 15544
rect 20162 15504 20168 15516
rect 20220 15504 20226 15556
rect 20714 15544 20720 15556
rect 20675 15516 20720 15544
rect 20714 15504 20720 15516
rect 20772 15504 20778 15556
rect 3697 15479 3755 15485
rect 3697 15445 3709 15479
rect 3743 15476 3755 15479
rect 7374 15476 7380 15488
rect 3743 15448 7380 15476
rect 3743 15445 3755 15448
rect 3697 15439 3755 15445
rect 7374 15436 7380 15448
rect 7432 15476 7438 15488
rect 7558 15476 7564 15488
rect 7432 15448 7564 15476
rect 7432 15436 7438 15448
rect 7558 15436 7564 15448
rect 7616 15436 7622 15488
rect 13906 15436 13912 15488
rect 13964 15476 13970 15488
rect 14829 15479 14887 15485
rect 14829 15476 14841 15479
rect 13964 15448 14841 15476
rect 13964 15436 13970 15448
rect 14829 15445 14841 15448
rect 14875 15445 14887 15479
rect 14829 15439 14887 15445
rect 2685 15411 2743 15417
rect 2685 15377 2697 15411
rect 2731 15408 2743 15411
rect 3326 15408 3332 15420
rect 2731 15380 3332 15408
rect 2731 15377 2743 15380
rect 2685 15371 2743 15377
rect 3326 15368 3332 15380
rect 3384 15368 3390 15420
rect 18969 15411 19027 15417
rect 18969 15408 18981 15411
rect 14292 15380 18981 15408
rect 2866 15340 2872 15352
rect 2827 15312 2872 15340
rect 2866 15300 2872 15312
rect 2924 15300 2930 15352
rect 3418 15300 3424 15352
rect 3476 15340 3482 15352
rect 3881 15343 3939 15349
rect 3881 15340 3893 15343
rect 3476 15312 3893 15340
rect 3476 15300 3482 15312
rect 3881 15309 3893 15312
rect 3927 15309 3939 15343
rect 3881 15303 3939 15309
rect 2317 15275 2375 15281
rect 2317 15241 2329 15275
rect 2363 15272 2375 15275
rect 14292 15272 14320 15380
rect 18969 15377 18981 15380
rect 19015 15377 19027 15411
rect 18969 15371 19027 15377
rect 19245 15411 19303 15417
rect 19245 15377 19257 15411
rect 19291 15408 19303 15411
rect 19981 15411 20039 15417
rect 19981 15408 19993 15411
rect 19291 15380 19993 15408
rect 19291 15377 19303 15380
rect 19245 15371 19303 15377
rect 19981 15377 19993 15380
rect 20027 15377 20039 15411
rect 19981 15371 20039 15377
rect 20162 15368 20168 15420
rect 20220 15408 20226 15420
rect 20533 15411 20591 15417
rect 20533 15408 20545 15411
rect 20220 15380 20545 15408
rect 20220 15368 20226 15380
rect 20533 15377 20545 15380
rect 20579 15377 20591 15411
rect 20533 15371 20591 15377
rect 15010 15340 15016 15352
rect 14971 15312 15016 15340
rect 15010 15300 15016 15312
rect 15068 15300 15074 15352
rect 2363 15244 14320 15272
rect 14369 15275 14427 15281
rect 2363 15241 2375 15244
rect 2317 15235 2375 15241
rect 14369 15241 14381 15275
rect 14415 15272 14427 15275
rect 19058 15272 19064 15284
rect 14415 15244 19064 15272
rect 14415 15241 14427 15244
rect 14369 15235 14427 15241
rect 19058 15232 19064 15244
rect 19116 15232 19122 15284
rect 1104 15114 21620 15136
rect 1104 15062 4414 15114
rect 4466 15062 4478 15114
rect 4530 15062 4542 15114
rect 4594 15062 4606 15114
rect 4658 15062 11278 15114
rect 11330 15062 11342 15114
rect 11394 15062 11406 15114
rect 11458 15062 11470 15114
rect 11522 15062 18142 15114
rect 18194 15062 18206 15114
rect 18258 15062 18270 15114
rect 18322 15062 18334 15114
rect 18386 15062 21620 15114
rect 1104 15040 21620 15062
rect 2866 15000 2872 15012
rect 2827 14972 2872 15000
rect 2866 14960 2872 14972
rect 2924 14960 2930 15012
rect 4982 14960 4988 15012
rect 5040 15000 5046 15012
rect 6362 15000 6368 15012
rect 5040 14972 6224 15000
rect 6323 14972 6368 15000
rect 5040 14960 5046 14972
rect 1486 14864 1492 14876
rect 1447 14836 1492 14864
rect 1486 14824 1492 14836
rect 1544 14824 1550 14876
rect 3326 14864 3332 14876
rect 3287 14836 3332 14864
rect 3326 14824 3332 14836
rect 3384 14824 3390 14876
rect 5000 14873 5028 14960
rect 6196 14932 6224 14972
rect 6362 14960 6368 14972
rect 6420 14960 6426 15012
rect 7466 14960 7472 15012
rect 7524 15000 7530 15012
rect 7524 14972 8340 15000
rect 7524 14960 7530 14972
rect 6825 14935 6883 14941
rect 6825 14932 6837 14935
rect 6196 14904 6837 14932
rect 6825 14901 6837 14904
rect 6871 14901 6883 14935
rect 6825 14895 6883 14901
rect 4985 14867 5043 14873
rect 4985 14833 4997 14867
rect 5031 14833 5043 14867
rect 8110 14864 8116 14876
rect 4985 14827 5043 14833
rect 7024 14836 8116 14864
rect 7024 14805 7052 14836
rect 8110 14824 8116 14836
rect 8168 14824 8174 14876
rect 7009 14799 7067 14805
rect 7009 14765 7021 14799
rect 7055 14765 7067 14799
rect 7009 14759 7067 14765
rect 7650 14756 7656 14808
rect 7708 14796 7714 14808
rect 8312 14805 8340 14972
rect 8386 14960 8392 15012
rect 8444 15000 8450 15012
rect 16853 15003 16911 15009
rect 16853 15000 16865 15003
rect 8444 14972 16865 15000
rect 8444 14960 8450 14972
rect 16853 14969 16865 14972
rect 16899 14969 16911 15003
rect 16853 14963 16911 14969
rect 10686 14892 10692 14944
rect 10744 14932 10750 14944
rect 13173 14935 13231 14941
rect 13173 14932 13185 14935
rect 10744 14904 13185 14932
rect 10744 14892 10750 14904
rect 13173 14901 13185 14904
rect 13219 14932 13231 14935
rect 13262 14932 13268 14944
rect 13219 14904 13268 14932
rect 13219 14901 13231 14904
rect 13173 14895 13231 14901
rect 13262 14892 13268 14904
rect 13320 14892 13326 14944
rect 8481 14867 8539 14873
rect 8481 14833 8493 14867
rect 8527 14864 8539 14867
rect 8662 14864 8668 14876
rect 8527 14836 8668 14864
rect 8527 14833 8539 14836
rect 8481 14827 8539 14833
rect 8662 14824 8668 14836
rect 8720 14824 8726 14876
rect 9766 14824 9772 14876
rect 9824 14864 9830 14876
rect 16868 14864 16896 14963
rect 17129 14935 17187 14941
rect 17129 14901 17141 14935
rect 17175 14932 17187 14935
rect 17175 14904 18920 14932
rect 17175 14901 17187 14904
rect 17129 14895 17187 14901
rect 17681 14867 17739 14873
rect 17681 14864 17693 14867
rect 9824 14836 15608 14864
rect 16868 14836 17693 14864
rect 9824 14824 9830 14836
rect 8205 14799 8263 14805
rect 8205 14796 8217 14799
rect 7708 14768 8217 14796
rect 7708 14756 7714 14768
rect 8205 14765 8217 14768
rect 8251 14765 8263 14799
rect 8205 14759 8263 14765
rect 8297 14799 8355 14805
rect 8297 14765 8309 14799
rect 8343 14765 8355 14799
rect 8297 14759 8355 14765
rect 12434 14756 12440 14808
rect 12492 14796 12498 14808
rect 13357 14799 13415 14805
rect 13357 14796 13369 14799
rect 12492 14768 13369 14796
rect 12492 14756 12498 14768
rect 13357 14765 13369 14768
rect 13403 14765 13415 14799
rect 13357 14759 13415 14765
rect 14550 14756 14556 14808
rect 14608 14796 14614 14808
rect 15470 14796 15476 14808
rect 14608 14768 15476 14796
rect 14608 14756 14614 14768
rect 15470 14756 15476 14768
rect 15528 14756 15534 14808
rect 15580 14796 15608 14836
rect 17681 14833 17693 14836
rect 17727 14833 17739 14867
rect 17681 14827 17739 14833
rect 18892 14805 18920 14904
rect 19702 14824 19708 14876
rect 19760 14864 19766 14876
rect 19797 14867 19855 14873
rect 19797 14864 19809 14867
rect 19760 14836 19809 14864
rect 19760 14824 19766 14836
rect 19797 14833 19809 14836
rect 19843 14833 19855 14867
rect 19797 14827 19855 14833
rect 18877 14799 18935 14805
rect 15580 14768 16068 14796
rect 1756 14731 1814 14737
rect 1756 14697 1768 14731
rect 1802 14728 1814 14731
rect 3418 14728 3424 14740
rect 1802 14700 3424 14728
rect 1802 14697 1814 14700
rect 1756 14691 1814 14697
rect 3418 14688 3424 14700
rect 3476 14688 3482 14740
rect 5252 14731 5310 14737
rect 5252 14697 5264 14731
rect 5298 14728 5310 14731
rect 9490 14728 9496 14740
rect 5298 14700 9496 14728
rect 5298 14697 5310 14700
rect 5252 14691 5310 14697
rect 9490 14688 9496 14700
rect 9548 14688 9554 14740
rect 15740 14731 15798 14737
rect 15740 14697 15752 14731
rect 15786 14697 15798 14731
rect 16040 14728 16068 14768
rect 18877 14765 18889 14799
rect 18923 14765 18935 14799
rect 19613 14799 19671 14805
rect 19613 14796 19625 14799
rect 18877 14759 18935 14765
rect 18984 14768 19625 14796
rect 18984 14728 19012 14768
rect 19613 14765 19625 14768
rect 19659 14765 19671 14799
rect 19613 14759 19671 14765
rect 16040 14700 19012 14728
rect 19153 14731 19211 14737
rect 15740 14691 15798 14697
rect 19153 14697 19165 14731
rect 19199 14728 19211 14731
rect 20254 14728 20260 14740
rect 19199 14700 20260 14728
rect 19199 14697 19211 14700
rect 19153 14691 19211 14697
rect 7837 14663 7895 14669
rect 7837 14629 7849 14663
rect 7883 14660 7895 14663
rect 9398 14660 9404 14672
rect 7883 14632 9404 14660
rect 7883 14629 7895 14632
rect 7837 14623 7895 14629
rect 9398 14620 9404 14632
rect 9456 14620 9462 14672
rect 9677 14663 9735 14669
rect 9677 14629 9689 14663
rect 9723 14660 9735 14663
rect 10134 14660 10140 14672
rect 9723 14632 10140 14660
rect 9723 14629 9735 14632
rect 9677 14623 9735 14629
rect 10134 14620 10140 14632
rect 10192 14620 10198 14672
rect 15764 14660 15792 14691
rect 20254 14688 20260 14700
rect 20312 14688 20318 14740
rect 16482 14660 16488 14672
rect 15764 14632 16488 14660
rect 16482 14620 16488 14632
rect 16540 14620 16546 14672
rect 17494 14660 17500 14672
rect 17455 14632 17500 14660
rect 17494 14620 17500 14632
rect 17552 14620 17558 14672
rect 17586 14620 17592 14672
rect 17644 14660 17650 14672
rect 17644 14632 17689 14660
rect 17644 14620 17650 14632
rect 1104 14570 21620 14592
rect 1104 14518 7846 14570
rect 7898 14518 7910 14570
rect 7962 14518 7974 14570
rect 8026 14518 8038 14570
rect 8090 14518 14710 14570
rect 14762 14518 14774 14570
rect 14826 14518 14838 14570
rect 14890 14518 14902 14570
rect 14954 14518 21620 14570
rect 1104 14496 21620 14518
rect 9490 14456 9496 14468
rect 9451 14428 9496 14456
rect 9490 14416 9496 14428
rect 9548 14456 9554 14468
rect 9585 14459 9643 14465
rect 9585 14456 9597 14459
rect 9548 14428 9597 14456
rect 9548 14416 9554 14428
rect 9585 14425 9597 14428
rect 9631 14425 9643 14459
rect 9766 14456 9772 14468
rect 9727 14428 9772 14456
rect 9585 14419 9643 14425
rect 9766 14416 9772 14428
rect 9824 14416 9830 14468
rect 10134 14456 10140 14468
rect 10095 14428 10140 14456
rect 10134 14416 10140 14428
rect 10192 14416 10198 14468
rect 13262 14416 13268 14468
rect 13320 14456 13326 14468
rect 14550 14456 14556 14468
rect 13320 14428 14556 14456
rect 13320 14416 13326 14428
rect 14550 14416 14556 14428
rect 14608 14456 14614 14468
rect 14829 14459 14887 14465
rect 14608 14428 14780 14456
rect 14608 14416 14614 14428
rect 3780 14391 3838 14397
rect 3780 14357 3792 14391
rect 3826 14388 3838 14391
rect 8294 14388 8300 14400
rect 3826 14360 5856 14388
rect 3826 14357 3838 14360
rect 3780 14351 3838 14357
rect 3513 14323 3571 14329
rect 3513 14289 3525 14323
rect 3559 14320 3571 14323
rect 4982 14320 4988 14332
rect 3559 14292 4988 14320
rect 3559 14289 3571 14292
rect 3513 14283 3571 14289
rect 4982 14280 4988 14292
rect 5040 14280 5046 14332
rect 5537 14323 5595 14329
rect 5537 14289 5549 14323
rect 5583 14289 5595 14323
rect 5537 14283 5595 14289
rect 5552 14184 5580 14283
rect 5626 14280 5632 14332
rect 5684 14320 5690 14332
rect 5684 14292 5729 14320
rect 5684 14280 5690 14292
rect 5828 14261 5856 14360
rect 8128 14360 8300 14388
rect 8128 14329 8156 14360
rect 8294 14348 8300 14360
rect 8352 14348 8358 14400
rect 9398 14348 9404 14400
rect 9456 14388 9462 14400
rect 10229 14391 10287 14397
rect 10229 14388 10241 14391
rect 9456 14360 10241 14388
rect 9456 14348 9462 14360
rect 10229 14357 10241 14360
rect 10275 14357 10287 14391
rect 14752 14388 14780 14428
rect 14829 14425 14841 14459
rect 14875 14456 14887 14459
rect 15010 14456 15016 14468
rect 14875 14428 15016 14456
rect 14875 14425 14887 14428
rect 14829 14419 14887 14425
rect 15010 14416 15016 14428
rect 15068 14416 15074 14468
rect 16482 14456 16488 14468
rect 16443 14428 16488 14456
rect 16482 14416 16488 14428
rect 16540 14456 16546 14468
rect 16669 14459 16727 14465
rect 16669 14456 16681 14459
rect 16540 14428 16681 14456
rect 16540 14416 16546 14428
rect 16669 14425 16681 14428
rect 16715 14425 16727 14459
rect 16669 14419 16727 14425
rect 16761 14459 16819 14465
rect 16761 14425 16773 14459
rect 16807 14456 16819 14459
rect 17586 14456 17592 14468
rect 16807 14428 17592 14456
rect 16807 14425 16819 14428
rect 16761 14419 16819 14425
rect 17586 14416 17592 14428
rect 17644 14416 17650 14468
rect 20714 14456 20720 14468
rect 20675 14428 20720 14456
rect 20714 14416 20720 14428
rect 20772 14416 20778 14468
rect 14921 14391 14979 14397
rect 14921 14388 14933 14391
rect 10229 14351 10287 14357
rect 12360 14360 14596 14388
rect 14752 14360 14933 14388
rect 8113 14323 8171 14329
rect 8113 14289 8125 14323
rect 8159 14289 8171 14323
rect 8113 14283 8171 14289
rect 8380 14323 8438 14329
rect 8380 14289 8392 14323
rect 8426 14320 8438 14323
rect 8662 14320 8668 14332
rect 8426 14292 8668 14320
rect 8426 14289 8438 14292
rect 8380 14283 8438 14289
rect 8662 14280 8668 14292
rect 8720 14280 8726 14332
rect 8846 14280 8852 14332
rect 8904 14320 8910 14332
rect 11882 14320 11888 14332
rect 8904 14292 11888 14320
rect 8904 14280 8910 14292
rect 11882 14280 11888 14292
rect 11940 14280 11946 14332
rect 5813 14255 5871 14261
rect 5813 14221 5825 14255
rect 5859 14252 5871 14255
rect 7006 14252 7012 14264
rect 5859 14224 7012 14252
rect 5859 14221 5871 14224
rect 5813 14215 5871 14221
rect 7006 14212 7012 14224
rect 7064 14212 7070 14264
rect 9585 14255 9643 14261
rect 9585 14221 9597 14255
rect 9631 14252 9643 14255
rect 10321 14255 10379 14261
rect 10321 14252 10333 14255
rect 9631 14224 10333 14252
rect 9631 14221 9643 14224
rect 9585 14215 9643 14221
rect 10321 14221 10333 14224
rect 10367 14221 10379 14255
rect 10321 14215 10379 14221
rect 7650 14184 7656 14196
rect 5552 14156 7656 14184
rect 7650 14144 7656 14156
rect 7708 14144 7714 14196
rect 4890 14116 4896 14128
rect 4851 14088 4896 14116
rect 4890 14076 4896 14088
rect 4948 14076 4954 14128
rect 5074 14076 5080 14128
rect 5132 14116 5138 14128
rect 5169 14119 5227 14125
rect 5169 14116 5181 14119
rect 5132 14088 5181 14116
rect 5132 14076 5138 14088
rect 5169 14085 5181 14088
rect 5215 14085 5227 14119
rect 5169 14079 5227 14085
rect 5258 14076 5264 14128
rect 5316 14116 5322 14128
rect 12360 14116 12388 14360
rect 12805 14323 12863 14329
rect 12805 14289 12817 14323
rect 12851 14320 12863 14323
rect 13354 14320 13360 14332
rect 12851 14292 13360 14320
rect 12851 14289 12863 14292
rect 12805 14283 12863 14289
rect 13354 14280 13360 14292
rect 13412 14280 13418 14332
rect 13716 14323 13774 14329
rect 13716 14289 13728 14323
rect 13762 14320 13774 14323
rect 14458 14320 14464 14332
rect 13762 14292 14464 14320
rect 13762 14289 13774 14292
rect 13716 14283 13774 14289
rect 14458 14280 14464 14292
rect 14516 14280 14522 14332
rect 14568 14320 14596 14360
rect 14921 14357 14933 14360
rect 14967 14357 14979 14391
rect 15028 14388 15056 14416
rect 15350 14391 15408 14397
rect 15350 14388 15362 14391
rect 15028 14360 15362 14388
rect 14921 14351 14979 14357
rect 15350 14357 15362 14360
rect 15396 14357 15408 14391
rect 19337 14391 19395 14397
rect 15350 14351 15408 14357
rect 15488 14360 19104 14388
rect 15488 14320 15516 14360
rect 14568 14292 15516 14320
rect 16942 14280 16948 14332
rect 17000 14320 17006 14332
rect 17129 14323 17187 14329
rect 17129 14320 17141 14323
rect 17000 14292 17141 14320
rect 17000 14280 17006 14292
rect 17129 14289 17141 14292
rect 17175 14289 17187 14323
rect 17129 14283 17187 14289
rect 17218 14280 17224 14332
rect 17276 14320 17282 14332
rect 19076 14329 19104 14360
rect 19337 14357 19349 14391
rect 19383 14388 19395 14391
rect 20162 14388 20168 14400
rect 19383 14360 20168 14388
rect 19383 14357 19395 14360
rect 19337 14351 19395 14357
rect 20162 14348 20168 14360
rect 20220 14348 20226 14400
rect 19061 14323 19119 14329
rect 17276 14292 17321 14320
rect 17276 14280 17282 14292
rect 19061 14289 19073 14323
rect 19107 14289 19119 14323
rect 19061 14283 19119 14289
rect 19797 14323 19855 14329
rect 19797 14289 19809 14323
rect 19843 14289 19855 14323
rect 19797 14283 19855 14289
rect 20073 14323 20131 14329
rect 20073 14289 20085 14323
rect 20119 14320 20131 14323
rect 20533 14323 20591 14329
rect 20533 14320 20545 14323
rect 20119 14292 20545 14320
rect 20119 14289 20131 14292
rect 20073 14283 20131 14289
rect 20533 14289 20545 14292
rect 20579 14289 20591 14323
rect 20533 14283 20591 14289
rect 12897 14255 12955 14261
rect 12897 14221 12909 14255
rect 12943 14221 12955 14255
rect 12897 14215 12955 14221
rect 5316 14088 12388 14116
rect 12437 14119 12495 14125
rect 5316 14076 5322 14088
rect 12437 14085 12449 14119
rect 12483 14116 12495 14119
rect 12802 14116 12808 14128
rect 12483 14088 12808 14116
rect 12483 14085 12495 14088
rect 12437 14079 12495 14085
rect 12802 14076 12808 14088
rect 12860 14076 12866 14128
rect 12912 14116 12940 14215
rect 12986 14212 12992 14264
rect 13044 14252 13050 14264
rect 13044 14224 13089 14252
rect 13044 14212 13050 14224
rect 13262 14212 13268 14264
rect 13320 14252 13326 14264
rect 13449 14255 13507 14261
rect 13449 14252 13461 14255
rect 13320 14224 13461 14252
rect 13320 14212 13326 14224
rect 13449 14221 13461 14224
rect 13495 14221 13507 14255
rect 13449 14215 13507 14221
rect 14921 14255 14979 14261
rect 14921 14221 14933 14255
rect 14967 14252 14979 14255
rect 15105 14255 15163 14261
rect 15105 14252 15117 14255
rect 14967 14224 15117 14252
rect 14967 14221 14979 14224
rect 14921 14215 14979 14221
rect 15105 14221 15117 14224
rect 15151 14221 15163 14255
rect 15105 14215 15163 14221
rect 16669 14255 16727 14261
rect 16669 14221 16681 14255
rect 16715 14252 16727 14255
rect 17310 14252 17316 14264
rect 16715 14224 17316 14252
rect 16715 14221 16727 14224
rect 16669 14215 16727 14221
rect 17310 14212 17316 14224
rect 17368 14212 17374 14264
rect 17402 14212 17408 14264
rect 17460 14252 17466 14264
rect 19812 14252 19840 14283
rect 17460 14224 19840 14252
rect 17460 14212 17466 14224
rect 17126 14116 17132 14128
rect 12912 14088 17132 14116
rect 17126 14076 17132 14088
rect 17184 14076 17190 14128
rect 1104 14026 21620 14048
rect 1104 13974 4414 14026
rect 4466 13974 4478 14026
rect 4530 13974 4542 14026
rect 4594 13974 4606 14026
rect 4658 13974 11278 14026
rect 11330 13974 11342 14026
rect 11394 13974 11406 14026
rect 11458 13974 11470 14026
rect 11522 13974 18142 14026
rect 18194 13974 18206 14026
rect 18258 13974 18270 14026
rect 18322 13974 18334 14026
rect 18386 13974 21620 14026
rect 1104 13952 21620 13974
rect 3418 13912 3424 13924
rect 3379 13884 3424 13912
rect 3418 13872 3424 13884
rect 3476 13872 3482 13924
rect 4617 13915 4675 13921
rect 4617 13881 4629 13915
rect 4663 13912 4675 13915
rect 5258 13912 5264 13924
rect 4663 13884 5264 13912
rect 4663 13881 4675 13884
rect 4617 13875 4675 13881
rect 5258 13872 5264 13884
rect 5316 13872 5322 13924
rect 7006 13912 7012 13924
rect 6967 13884 7012 13912
rect 7006 13872 7012 13884
rect 7064 13872 7070 13924
rect 8662 13912 8668 13924
rect 7208 13884 8524 13912
rect 8623 13884 8668 13912
rect 1486 13736 1492 13788
rect 1544 13776 1550 13788
rect 2041 13779 2099 13785
rect 2041 13776 2053 13779
rect 1544 13748 2053 13776
rect 1544 13736 1550 13748
rect 2041 13745 2053 13748
rect 2087 13745 2099 13779
rect 5074 13776 5080 13788
rect 5035 13748 5080 13776
rect 2041 13739 2099 13745
rect 5074 13736 5080 13748
rect 5132 13736 5138 13788
rect 5169 13779 5227 13785
rect 5169 13745 5181 13779
rect 5215 13745 5227 13779
rect 5169 13739 5227 13745
rect 2308 13711 2366 13717
rect 2308 13677 2320 13711
rect 2354 13708 2366 13711
rect 4890 13708 4896 13720
rect 2354 13680 4896 13708
rect 2354 13677 2366 13680
rect 2308 13671 2366 13677
rect 4890 13668 4896 13680
rect 4948 13708 4954 13720
rect 5184 13708 5212 13739
rect 4948 13680 5212 13708
rect 5629 13711 5687 13717
rect 4948 13668 4954 13680
rect 5629 13677 5641 13711
rect 5675 13708 5687 13711
rect 5896 13711 5954 13717
rect 5675 13680 5856 13708
rect 5675 13677 5687 13680
rect 5629 13671 5687 13677
rect 5828 13640 5856 13680
rect 5896 13677 5908 13711
rect 5942 13708 5954 13711
rect 7208 13708 7236 13884
rect 8496 13844 8524 13884
rect 8662 13872 8668 13884
rect 8720 13872 8726 13924
rect 12066 13912 12072 13924
rect 10152 13884 12072 13912
rect 10152 13844 10180 13884
rect 12066 13872 12072 13884
rect 12124 13872 12130 13924
rect 12345 13915 12403 13921
rect 12345 13881 12357 13915
rect 12391 13912 12403 13915
rect 12894 13912 12900 13924
rect 12391 13884 12900 13912
rect 12391 13881 12403 13884
rect 12345 13875 12403 13881
rect 12894 13872 12900 13884
rect 12952 13872 12958 13924
rect 16669 13915 16727 13921
rect 16669 13881 16681 13915
rect 16715 13912 16727 13915
rect 17494 13912 17500 13924
rect 16715 13884 17500 13912
rect 16715 13881 16727 13884
rect 16669 13875 16727 13881
rect 17494 13872 17500 13884
rect 17552 13872 17558 13924
rect 18509 13915 18567 13921
rect 18509 13881 18521 13915
rect 18555 13912 18567 13915
rect 18598 13912 18604 13924
rect 18555 13884 18604 13912
rect 18555 13881 18567 13884
rect 18509 13875 18567 13881
rect 18598 13872 18604 13884
rect 18656 13872 18662 13924
rect 20441 13915 20499 13921
rect 20441 13881 20453 13915
rect 20487 13912 20499 13915
rect 20530 13912 20536 13924
rect 20487 13884 20536 13912
rect 20487 13881 20499 13884
rect 20441 13875 20499 13881
rect 20530 13872 20536 13884
rect 20588 13872 20594 13924
rect 8496 13816 10180 13844
rect 10686 13776 10692 13788
rect 10647 13748 10692 13776
rect 10686 13736 10692 13748
rect 10744 13736 10750 13788
rect 12986 13776 12992 13788
rect 11808 13748 12992 13776
rect 5942 13680 7236 13708
rect 7285 13711 7343 13717
rect 5942 13677 5954 13680
rect 5896 13671 5954 13677
rect 7285 13677 7297 13711
rect 7331 13708 7343 13711
rect 8294 13708 8300 13720
rect 7331 13680 8300 13708
rect 7331 13677 7343 13680
rect 7285 13671 7343 13677
rect 7190 13640 7196 13652
rect 5828 13612 7196 13640
rect 7190 13600 7196 13612
rect 7248 13640 7254 13652
rect 7300 13640 7328 13671
rect 8294 13668 8300 13680
rect 8352 13668 8358 13720
rect 9125 13711 9183 13717
rect 9125 13677 9137 13711
rect 9171 13708 9183 13711
rect 10594 13708 10600 13720
rect 9171 13680 10600 13708
rect 9171 13677 9183 13680
rect 9125 13671 9183 13677
rect 10594 13668 10600 13680
rect 10652 13668 10658 13720
rect 7248 13612 7328 13640
rect 7552 13643 7610 13649
rect 7248 13600 7254 13612
rect 7552 13609 7564 13643
rect 7598 13640 7610 13643
rect 8386 13640 8392 13652
rect 7598 13612 8392 13640
rect 7598 13609 7610 13612
rect 7552 13603 7610 13609
rect 8386 13600 8392 13612
rect 8444 13600 8450 13652
rect 10956 13643 11014 13649
rect 10956 13609 10968 13643
rect 11002 13640 11014 13643
rect 11054 13640 11060 13652
rect 11002 13612 11060 13640
rect 11002 13609 11014 13612
rect 10956 13603 11014 13609
rect 11054 13600 11060 13612
rect 11112 13640 11118 13652
rect 11808 13640 11836 13748
rect 12986 13736 12992 13748
rect 13044 13736 13050 13788
rect 13354 13776 13360 13788
rect 13315 13748 13360 13776
rect 13354 13736 13360 13748
rect 13412 13736 13418 13788
rect 17126 13776 17132 13788
rect 17087 13748 17132 13776
rect 17126 13736 17132 13748
rect 17184 13736 17190 13788
rect 17310 13776 17316 13788
rect 17271 13748 17316 13776
rect 17310 13736 17316 13748
rect 17368 13736 17374 13788
rect 11882 13668 11888 13720
rect 11940 13708 11946 13720
rect 12805 13711 12863 13717
rect 12805 13708 12817 13711
rect 11940 13680 12817 13708
rect 11940 13668 11946 13680
rect 12805 13677 12817 13680
rect 12851 13677 12863 13711
rect 18322 13708 18328 13720
rect 18283 13680 18328 13708
rect 12805 13671 12863 13677
rect 18322 13668 18328 13680
rect 18380 13668 18386 13720
rect 20254 13708 20260 13720
rect 20215 13680 20260 13708
rect 20254 13668 20260 13680
rect 20312 13668 20318 13720
rect 11112 13612 11836 13640
rect 12713 13643 12771 13649
rect 11112 13600 11118 13612
rect 12713 13609 12725 13643
rect 12759 13640 12771 13643
rect 16114 13640 16120 13652
rect 12759 13612 16120 13640
rect 12759 13609 12771 13612
rect 12713 13603 12771 13609
rect 16114 13600 16120 13612
rect 16172 13640 16178 13652
rect 16942 13640 16948 13652
rect 16172 13612 16948 13640
rect 16172 13600 16178 13612
rect 16942 13600 16948 13612
rect 17000 13600 17006 13652
rect 17037 13643 17095 13649
rect 17037 13609 17049 13643
rect 17083 13640 17095 13643
rect 17681 13643 17739 13649
rect 17681 13640 17693 13643
rect 17083 13612 17693 13640
rect 17083 13609 17095 13612
rect 17037 13603 17095 13609
rect 17681 13609 17693 13612
rect 17727 13609 17739 13643
rect 17681 13603 17739 13609
rect 4982 13572 4988 13584
rect 4943 13544 4988 13572
rect 4982 13532 4988 13544
rect 5040 13532 5046 13584
rect 8202 13532 8208 13584
rect 8260 13572 8266 13584
rect 8941 13575 8999 13581
rect 8941 13572 8953 13575
rect 8260 13544 8953 13572
rect 8260 13532 8266 13544
rect 8941 13541 8953 13544
rect 8987 13541 8999 13575
rect 8941 13535 8999 13541
rect 11146 13532 11152 13584
rect 11204 13572 11210 13584
rect 11698 13572 11704 13584
rect 11204 13544 11704 13572
rect 11204 13532 11210 13544
rect 11698 13532 11704 13544
rect 11756 13532 11762 13584
rect 1104 13482 21620 13504
rect 1104 13430 7846 13482
rect 7898 13430 7910 13482
rect 7962 13430 7974 13482
rect 8026 13430 8038 13482
rect 8090 13430 14710 13482
rect 14762 13430 14774 13482
rect 14826 13430 14838 13482
rect 14890 13430 14902 13482
rect 14954 13430 21620 13482
rect 1104 13408 21620 13430
rect 4982 13368 4988 13380
rect 4943 13340 4988 13368
rect 4982 13328 4988 13340
rect 5040 13328 5046 13380
rect 10594 13328 10600 13380
rect 10652 13368 10658 13380
rect 10962 13368 10968 13380
rect 10652 13340 10968 13368
rect 10652 13328 10658 13340
rect 10962 13328 10968 13340
rect 11020 13368 11026 13380
rect 11241 13371 11299 13377
rect 11241 13368 11253 13371
rect 11020 13340 11253 13368
rect 11020 13328 11026 13340
rect 11241 13337 11253 13340
rect 11287 13337 11299 13371
rect 12802 13368 12808 13380
rect 12763 13340 12808 13368
rect 11241 13331 11299 13337
rect 12802 13328 12808 13340
rect 12860 13328 12866 13380
rect 12894 13328 12900 13380
rect 12952 13368 12958 13380
rect 18782 13368 18788 13380
rect 12952 13340 12997 13368
rect 14384 13340 18788 13368
rect 12952 13328 12958 13340
rect 9953 13235 10011 13241
rect 9953 13201 9965 13235
rect 9999 13232 10011 13235
rect 14384 13232 14412 13340
rect 18782 13328 18788 13340
rect 18840 13328 18846 13380
rect 20165 13371 20223 13377
rect 20165 13337 20177 13371
rect 20211 13368 20223 13371
rect 20346 13368 20352 13380
rect 20211 13340 20352 13368
rect 20211 13337 20223 13340
rect 20165 13331 20223 13337
rect 20346 13328 20352 13340
rect 20404 13328 20410 13380
rect 20714 13368 20720 13380
rect 20675 13340 20720 13368
rect 20714 13328 20720 13340
rect 20772 13328 20778 13380
rect 18322 13260 18328 13312
rect 18380 13300 18386 13312
rect 18877 13303 18935 13309
rect 18877 13300 18889 13303
rect 18380 13272 18889 13300
rect 18380 13260 18386 13272
rect 18877 13269 18889 13272
rect 18923 13269 18935 13303
rect 18877 13263 18935 13269
rect 9999 13204 14412 13232
rect 9999 13201 10011 13204
rect 9953 13195 10011 13201
rect 17586 13192 17592 13244
rect 17644 13232 17650 13244
rect 18601 13235 18659 13241
rect 18601 13232 18613 13235
rect 17644 13204 18613 13232
rect 17644 13192 17650 13204
rect 18601 13201 18613 13204
rect 18647 13201 18659 13235
rect 19978 13232 19984 13244
rect 19939 13204 19984 13232
rect 18601 13195 18659 13201
rect 19978 13192 19984 13204
rect 20036 13192 20042 13244
rect 20533 13235 20591 13241
rect 20533 13201 20545 13235
rect 20579 13201 20591 13235
rect 20533 13195 20591 13201
rect 12066 13124 12072 13176
rect 12124 13164 12130 13176
rect 12989 13167 13047 13173
rect 12989 13164 13001 13167
rect 12124 13136 13001 13164
rect 12124 13124 12130 13136
rect 12989 13133 13001 13136
rect 13035 13133 13047 13167
rect 12989 13127 13047 13133
rect 15562 13124 15568 13176
rect 15620 13164 15626 13176
rect 20548 13164 20576 13195
rect 15620 13136 20576 13164
rect 15620 13124 15626 13136
rect 12437 13031 12495 13037
rect 12437 12997 12449 13031
rect 12483 13028 12495 13031
rect 17402 13028 17408 13040
rect 12483 13000 17408 13028
rect 12483 12997 12495 13000
rect 12437 12991 12495 12997
rect 17402 12988 17408 13000
rect 17460 12988 17466 13040
rect 1104 12938 21620 12960
rect 1104 12886 4414 12938
rect 4466 12886 4478 12938
rect 4530 12886 4542 12938
rect 4594 12886 4606 12938
rect 4658 12886 11278 12938
rect 11330 12886 11342 12938
rect 11394 12886 11406 12938
rect 11458 12886 11470 12938
rect 11522 12886 18142 12938
rect 18194 12886 18206 12938
rect 18258 12886 18270 12938
rect 18322 12886 18334 12938
rect 18386 12886 21620 12938
rect 1104 12864 21620 12886
rect 11054 12824 11060 12836
rect 11015 12796 11060 12824
rect 11054 12784 11060 12796
rect 11112 12784 11118 12836
rect 12434 12824 12440 12836
rect 12395 12796 12440 12824
rect 12434 12784 12440 12796
rect 12492 12784 12498 12836
rect 13357 12827 13415 12833
rect 13357 12793 13369 12827
rect 13403 12824 13415 12827
rect 14090 12824 14096 12836
rect 13403 12796 14096 12824
rect 13403 12793 13415 12796
rect 13357 12787 13415 12793
rect 14090 12784 14096 12796
rect 14148 12784 14154 12836
rect 19978 12824 19984 12836
rect 16224 12796 19984 12824
rect 16224 12756 16252 12796
rect 19978 12784 19984 12796
rect 20036 12784 20042 12836
rect 20346 12824 20352 12836
rect 20307 12796 20352 12824
rect 20346 12784 20352 12796
rect 20404 12784 20410 12836
rect 11440 12728 16252 12756
rect 10962 12648 10968 12700
rect 11020 12688 11026 12700
rect 11440 12697 11468 12728
rect 19610 12716 19616 12768
rect 19668 12756 19674 12768
rect 19797 12759 19855 12765
rect 19797 12756 19809 12759
rect 19668 12728 19809 12756
rect 19668 12716 19674 12728
rect 19797 12725 19809 12728
rect 19843 12725 19855 12759
rect 19797 12719 19855 12725
rect 11425 12691 11483 12697
rect 11020 12660 11284 12688
rect 11020 12648 11026 12660
rect 8294 12580 8300 12632
rect 8352 12620 8358 12632
rect 9677 12623 9735 12629
rect 9677 12620 9689 12623
rect 8352 12592 9689 12620
rect 8352 12580 8358 12592
rect 9677 12589 9689 12592
rect 9723 12589 9735 12623
rect 11146 12620 11152 12632
rect 11107 12592 11152 12620
rect 9677 12583 9735 12589
rect 11146 12580 11152 12592
rect 11204 12580 11210 12632
rect 11256 12620 11284 12660
rect 11425 12657 11437 12691
rect 11471 12657 11483 12691
rect 11425 12651 11483 12657
rect 12434 12648 12440 12700
rect 12492 12688 12498 12700
rect 12492 12660 13308 12688
rect 12492 12648 12498 12660
rect 12621 12623 12679 12629
rect 12621 12620 12633 12623
rect 11256 12592 12633 12620
rect 12621 12589 12633 12592
rect 12667 12589 12679 12623
rect 13280 12620 13308 12660
rect 13354 12648 13360 12700
rect 13412 12688 13418 12700
rect 13909 12691 13967 12697
rect 13909 12688 13921 12691
rect 13412 12660 13921 12688
rect 13412 12648 13418 12660
rect 13909 12657 13921 12660
rect 13955 12657 13967 12691
rect 15562 12688 15568 12700
rect 15523 12660 15568 12688
rect 13909 12651 13967 12657
rect 15562 12648 15568 12660
rect 15620 12648 15626 12700
rect 14182 12620 14188 12632
rect 13280 12592 14188 12620
rect 12621 12583 12679 12589
rect 14182 12580 14188 12592
rect 14240 12580 14246 12632
rect 14458 12580 14464 12632
rect 14516 12620 14522 12632
rect 15289 12623 15347 12629
rect 15289 12620 15301 12623
rect 14516 12592 15301 12620
rect 14516 12580 14522 12592
rect 15289 12589 15301 12592
rect 15335 12589 15347 12623
rect 16666 12620 16672 12632
rect 16627 12592 16672 12620
rect 15289 12583 15347 12589
rect 16666 12580 16672 12592
rect 16724 12580 16730 12632
rect 19242 12580 19248 12632
rect 19300 12620 19306 12632
rect 19613 12623 19671 12629
rect 19613 12620 19625 12623
rect 19300 12592 19625 12620
rect 19300 12580 19306 12592
rect 19613 12589 19625 12592
rect 19659 12589 19671 12623
rect 20162 12620 20168 12632
rect 20123 12592 20168 12620
rect 19613 12583 19671 12589
rect 20162 12580 20168 12592
rect 20220 12580 20226 12632
rect 9858 12512 9864 12564
rect 9916 12561 9922 12564
rect 9916 12555 9980 12561
rect 9916 12521 9934 12555
rect 9968 12521 9980 12555
rect 9916 12515 9980 12521
rect 13725 12555 13783 12561
rect 13725 12521 13737 12555
rect 13771 12552 13783 12555
rect 13998 12552 14004 12564
rect 13771 12524 14004 12552
rect 13771 12521 13783 12524
rect 13725 12515 13783 12521
rect 9916 12512 9922 12515
rect 13998 12512 14004 12524
rect 14056 12512 14062 12564
rect 16936 12555 16994 12561
rect 16936 12521 16948 12555
rect 16982 12552 16994 12555
rect 17494 12552 17500 12564
rect 16982 12524 17500 12552
rect 16982 12521 16994 12524
rect 16936 12515 16994 12521
rect 17494 12512 17500 12524
rect 17552 12512 17558 12564
rect 19794 12512 19800 12564
rect 19852 12552 19858 12564
rect 20070 12552 20076 12564
rect 19852 12524 20076 12552
rect 19852 12512 19858 12524
rect 20070 12512 20076 12524
rect 20128 12512 20134 12564
rect 8478 12444 8484 12496
rect 8536 12484 8542 12496
rect 9674 12484 9680 12496
rect 8536 12456 9680 12484
rect 8536 12444 8542 12456
rect 9674 12444 9680 12456
rect 9732 12444 9738 12496
rect 13446 12444 13452 12496
rect 13504 12484 13510 12496
rect 13817 12487 13875 12493
rect 13817 12484 13829 12487
rect 13504 12456 13829 12484
rect 13504 12444 13510 12456
rect 13817 12453 13829 12456
rect 13863 12453 13875 12487
rect 18046 12484 18052 12496
rect 18007 12456 18052 12484
rect 13817 12447 13875 12453
rect 18046 12444 18052 12456
rect 18104 12444 18110 12496
rect 1104 12394 21620 12416
rect 1104 12342 7846 12394
rect 7898 12342 7910 12394
rect 7962 12342 7974 12394
rect 8026 12342 8038 12394
rect 8090 12342 14710 12394
rect 14762 12342 14774 12394
rect 14826 12342 14838 12394
rect 14890 12342 14902 12394
rect 14954 12342 21620 12394
rect 1104 12320 21620 12342
rect 1946 12240 1952 12292
rect 2004 12280 2010 12292
rect 7285 12283 7343 12289
rect 7285 12280 7297 12283
rect 2004 12252 7297 12280
rect 2004 12240 2010 12252
rect 7285 12249 7297 12252
rect 7331 12249 7343 12283
rect 7285 12243 7343 12249
rect 7650 12240 7656 12292
rect 7708 12280 7714 12292
rect 9953 12283 10011 12289
rect 7708 12252 9352 12280
rect 7708 12240 7714 12252
rect 7193 12215 7251 12221
rect 7193 12181 7205 12215
rect 7239 12212 7251 12215
rect 7668 12212 7696 12240
rect 7239 12184 7696 12212
rect 7239 12181 7251 12184
rect 7193 12175 7251 12181
rect 8021 12147 8079 12153
rect 8021 12113 8033 12147
rect 8067 12144 8079 12147
rect 8202 12144 8208 12156
rect 8067 12116 8208 12144
rect 8067 12113 8079 12116
rect 8021 12107 8079 12113
rect 8202 12104 8208 12116
rect 8260 12104 8266 12156
rect 8386 12104 8392 12156
rect 8444 12144 8450 12156
rect 8553 12147 8611 12153
rect 8553 12144 8565 12147
rect 8444 12116 8565 12144
rect 8444 12104 8450 12116
rect 8553 12113 8565 12116
rect 8599 12113 8611 12147
rect 8553 12107 8611 12113
rect 7469 12079 7527 12085
rect 7469 12045 7481 12079
rect 7515 12076 7527 12079
rect 8113 12079 8171 12085
rect 8113 12076 8125 12079
rect 7515 12048 8125 12076
rect 7515 12045 7527 12048
rect 7469 12039 7527 12045
rect 8113 12045 8125 12048
rect 8159 12045 8171 12079
rect 8294 12076 8300 12088
rect 8207 12048 8300 12076
rect 8113 12039 8171 12045
rect 8294 12036 8300 12048
rect 8352 12036 8358 12088
rect 9324 12076 9352 12252
rect 9953 12249 9965 12283
rect 9999 12280 10011 12283
rect 11146 12280 11152 12292
rect 9999 12252 11152 12280
rect 9999 12249 10011 12252
rect 9953 12243 10011 12249
rect 11146 12240 11152 12252
rect 11204 12240 11210 12292
rect 12713 12283 12771 12289
rect 12713 12249 12725 12283
rect 12759 12280 12771 12283
rect 13446 12280 13452 12292
rect 12759 12252 13452 12280
rect 12759 12249 12771 12252
rect 12713 12243 12771 12249
rect 13446 12240 13452 12252
rect 13504 12240 13510 12292
rect 13541 12283 13599 12289
rect 13541 12249 13553 12283
rect 13587 12280 13599 12283
rect 13998 12280 14004 12292
rect 13587 12252 13851 12280
rect 13959 12252 14004 12280
rect 13587 12249 13599 12252
rect 13541 12243 13599 12249
rect 10410 12212 10416 12224
rect 10371 12184 10416 12212
rect 10410 12172 10416 12184
rect 10468 12172 10474 12224
rect 13823 12212 13851 12252
rect 13998 12240 14004 12252
rect 14056 12240 14062 12292
rect 14461 12283 14519 12289
rect 14461 12280 14473 12283
rect 14108 12252 14473 12280
rect 14108 12212 14136 12252
rect 14461 12249 14473 12252
rect 14507 12280 14519 12283
rect 18782 12280 18788 12292
rect 14507 12252 18788 12280
rect 14507 12249 14519 12252
rect 14461 12243 14519 12249
rect 18782 12240 18788 12252
rect 18840 12240 18846 12292
rect 20254 12240 20260 12292
rect 20312 12280 20318 12292
rect 20717 12283 20775 12289
rect 20717 12280 20729 12283
rect 20312 12252 20729 12280
rect 20312 12240 20318 12252
rect 20717 12249 20729 12252
rect 20763 12249 20775 12283
rect 20717 12243 20775 12249
rect 13823 12184 14136 12212
rect 14369 12215 14427 12221
rect 14369 12181 14381 12215
rect 14415 12212 14427 12215
rect 14550 12212 14556 12224
rect 14415 12184 14556 12212
rect 14415 12181 14427 12184
rect 14369 12175 14427 12181
rect 14550 12172 14556 12184
rect 14608 12212 14614 12224
rect 15372 12215 15430 12221
rect 14608 12184 15240 12212
rect 14608 12172 14614 12184
rect 10318 12144 10324 12156
rect 10279 12116 10324 12144
rect 10318 12104 10324 12116
rect 10376 12104 10382 12156
rect 12986 12144 12992 12156
rect 10428 12116 12992 12144
rect 10428 12076 10456 12116
rect 12986 12104 12992 12116
rect 13044 12144 13050 12156
rect 13081 12147 13139 12153
rect 13081 12144 13093 12147
rect 13044 12116 13093 12144
rect 13044 12104 13050 12116
rect 13081 12113 13093 12116
rect 13127 12113 13139 12147
rect 13081 12107 13139 12113
rect 13909 12147 13967 12153
rect 13909 12113 13921 12147
rect 13955 12144 13967 12147
rect 14182 12144 14188 12156
rect 13955 12116 14188 12144
rect 13955 12113 13967 12116
rect 13909 12107 13967 12113
rect 14182 12104 14188 12116
rect 14240 12104 14246 12156
rect 15105 12147 15163 12153
rect 15105 12144 15117 12147
rect 14476 12116 15117 12144
rect 9324 12048 10456 12076
rect 10505 12079 10563 12085
rect 10505 12045 10517 12079
rect 10551 12045 10563 12079
rect 13170 12076 13176 12088
rect 13131 12048 13176 12076
rect 10505 12039 10563 12045
rect 8312 12008 8340 12036
rect 7852 11980 8340 12008
rect 9677 12011 9735 12017
rect 6822 11940 6828 11952
rect 6783 11912 6828 11940
rect 6822 11900 6828 11912
rect 6880 11900 6886 11952
rect 7190 11900 7196 11952
rect 7248 11940 7254 11952
rect 7558 11940 7564 11952
rect 7248 11912 7564 11940
rect 7248 11900 7254 11912
rect 7558 11900 7564 11912
rect 7616 11940 7622 11952
rect 7852 11949 7880 11980
rect 9677 11977 9689 12011
rect 9723 12008 9735 12011
rect 9858 12008 9864 12020
rect 9723 11980 9864 12008
rect 9723 11977 9735 11980
rect 9677 11971 9735 11977
rect 9858 11968 9864 11980
rect 9916 12008 9922 12020
rect 10520 12008 10548 12039
rect 13170 12036 13176 12048
rect 13228 12036 13234 12088
rect 13357 12079 13415 12085
rect 13357 12045 13369 12079
rect 13403 12045 13415 12079
rect 13357 12039 13415 12045
rect 9916 11980 10548 12008
rect 9916 11968 9922 11980
rect 12618 11968 12624 12020
rect 12676 12008 12682 12020
rect 13372 12008 13400 12039
rect 13722 12036 13728 12088
rect 13780 12076 13786 12088
rect 14476 12076 14504 12116
rect 15105 12113 15117 12116
rect 15151 12113 15163 12147
rect 15212 12144 15240 12184
rect 15372 12181 15384 12215
rect 15418 12212 15430 12215
rect 18046 12212 18052 12224
rect 15418 12184 18052 12212
rect 15418 12181 15430 12184
rect 15372 12175 15430 12181
rect 18046 12172 18052 12184
rect 18104 12212 18110 12224
rect 19521 12215 19579 12221
rect 18104 12184 18644 12212
rect 18104 12172 18110 12184
rect 15212 12116 16620 12144
rect 15105 12107 15163 12113
rect 13780 12048 14504 12076
rect 14645 12079 14703 12085
rect 13780 12036 13786 12048
rect 14645 12045 14657 12079
rect 14691 12076 14703 12079
rect 14691 12048 14780 12076
rect 14691 12045 14703 12048
rect 14645 12039 14703 12045
rect 12676 11980 13851 12008
rect 12676 11968 12682 11980
rect 7837 11943 7895 11949
rect 7837 11940 7849 11943
rect 7616 11912 7849 11940
rect 7616 11900 7622 11912
rect 7837 11909 7849 11912
rect 7883 11909 7895 11943
rect 7837 11903 7895 11909
rect 8113 11943 8171 11949
rect 8113 11909 8125 11943
rect 8159 11940 8171 11943
rect 8570 11940 8576 11952
rect 8159 11912 8576 11940
rect 8159 11909 8171 11912
rect 8113 11903 8171 11909
rect 8570 11900 8576 11912
rect 8628 11900 8634 11952
rect 8938 11900 8944 11952
rect 8996 11940 9002 11952
rect 13541 11943 13599 11949
rect 13541 11940 13553 11943
rect 8996 11912 13553 11940
rect 8996 11900 9002 11912
rect 13541 11909 13553 11912
rect 13587 11909 13599 11943
rect 13722 11940 13728 11952
rect 13683 11912 13728 11940
rect 13541 11903 13599 11909
rect 13722 11900 13728 11912
rect 13780 11900 13786 11952
rect 13823 11940 13851 11980
rect 14752 11940 14780 12048
rect 16485 11943 16543 11949
rect 16485 11940 16497 11943
rect 13823 11912 16497 11940
rect 16485 11909 16497 11912
rect 16531 11909 16543 11943
rect 16592 11940 16620 12116
rect 17954 12104 17960 12156
rect 18012 12144 18018 12156
rect 18417 12147 18475 12153
rect 18417 12144 18429 12147
rect 18012 12116 18429 12144
rect 18012 12104 18018 12116
rect 18417 12113 18429 12116
rect 18463 12113 18475 12147
rect 18417 12107 18475 12113
rect 16942 12036 16948 12088
rect 17000 12076 17006 12088
rect 18616 12085 18644 12184
rect 19521 12181 19533 12215
rect 19567 12212 19579 12215
rect 20162 12212 20168 12224
rect 19567 12184 20168 12212
rect 19567 12181 19579 12184
rect 19521 12175 19579 12181
rect 20162 12172 20168 12184
rect 20220 12172 20226 12224
rect 19245 12147 19303 12153
rect 19245 12144 19257 12147
rect 18708 12116 19257 12144
rect 18509 12079 18567 12085
rect 18509 12076 18521 12079
rect 17000 12048 18521 12076
rect 17000 12036 17006 12048
rect 18509 12045 18521 12048
rect 18555 12045 18567 12079
rect 18509 12039 18567 12045
rect 18601 12079 18659 12085
rect 18601 12045 18613 12079
rect 18647 12045 18659 12079
rect 18601 12039 18659 12045
rect 18049 12011 18107 12017
rect 18049 11977 18061 12011
rect 18095 12008 18107 12011
rect 18708 12008 18736 12116
rect 19245 12113 19257 12116
rect 19291 12113 19303 12147
rect 19978 12144 19984 12156
rect 19939 12116 19984 12144
rect 19245 12107 19303 12113
rect 19978 12104 19984 12116
rect 20036 12104 20042 12156
rect 20530 12144 20536 12156
rect 20491 12116 20536 12144
rect 20530 12104 20536 12116
rect 20588 12104 20594 12156
rect 18095 11980 18736 12008
rect 20165 12011 20223 12017
rect 18095 11977 18107 11980
rect 18049 11971 18107 11977
rect 20165 11977 20177 12011
rect 20211 12008 20223 12011
rect 20898 12008 20904 12020
rect 20211 11980 20904 12008
rect 20211 11977 20223 11980
rect 20165 11971 20223 11977
rect 20898 11968 20904 11980
rect 20956 11968 20962 12020
rect 18598 11940 18604 11952
rect 16592 11912 18604 11940
rect 16485 11903 16543 11909
rect 18598 11900 18604 11912
rect 18656 11900 18662 11952
rect 1104 11850 21620 11872
rect 1104 11798 4414 11850
rect 4466 11798 4478 11850
rect 4530 11798 4542 11850
rect 4594 11798 4606 11850
rect 4658 11798 11278 11850
rect 11330 11798 11342 11850
rect 11394 11798 11406 11850
rect 11458 11798 11470 11850
rect 11522 11798 18142 11850
rect 18194 11798 18206 11850
rect 18258 11798 18270 11850
rect 18322 11798 18334 11850
rect 18386 11798 21620 11850
rect 1104 11776 21620 11798
rect 10318 11736 10324 11748
rect 10279 11708 10324 11736
rect 10318 11696 10324 11708
rect 10376 11696 10382 11748
rect 13633 11739 13691 11745
rect 13633 11705 13645 11739
rect 13679 11736 13691 11739
rect 14458 11736 14464 11748
rect 13679 11708 14464 11736
rect 13679 11705 13691 11708
rect 13633 11699 13691 11705
rect 14458 11696 14464 11708
rect 14516 11696 14522 11748
rect 17954 11696 17960 11748
rect 18012 11736 18018 11748
rect 18049 11739 18107 11745
rect 18049 11736 18061 11739
rect 18012 11708 18061 11736
rect 18012 11696 18018 11708
rect 18049 11705 18061 11708
rect 18095 11705 18107 11739
rect 18049 11699 18107 11705
rect 19886 11696 19892 11748
rect 19944 11736 19950 11748
rect 20441 11739 20499 11745
rect 20441 11736 20453 11739
rect 19944 11708 20453 11736
rect 19944 11696 19950 11708
rect 20441 11705 20453 11708
rect 20487 11705 20499 11739
rect 20441 11699 20499 11705
rect 7837 11671 7895 11677
rect 7837 11637 7849 11671
rect 7883 11668 7895 11671
rect 8386 11668 8392 11680
rect 7883 11640 8392 11668
rect 7883 11637 7895 11640
rect 7837 11631 7895 11637
rect 8386 11628 8392 11640
rect 8444 11668 8450 11680
rect 8444 11640 10916 11668
rect 8444 11628 8450 11640
rect 8570 11560 8576 11612
rect 8628 11600 8634 11612
rect 10888 11609 10916 11640
rect 12986 11628 12992 11680
rect 13044 11668 13050 11680
rect 18506 11668 18512 11680
rect 13044 11640 18512 11668
rect 13044 11628 13050 11640
rect 18506 11628 18512 11640
rect 18564 11628 18570 11680
rect 8665 11603 8723 11609
rect 8665 11600 8677 11603
rect 8628 11572 8677 11600
rect 8628 11560 8634 11572
rect 8665 11569 8677 11572
rect 8711 11569 8723 11603
rect 8665 11563 8723 11569
rect 10873 11603 10931 11609
rect 10873 11569 10885 11603
rect 10919 11569 10931 11603
rect 14182 11600 14188 11612
rect 14143 11572 14188 11600
rect 10873 11563 10931 11569
rect 14182 11560 14188 11572
rect 14240 11560 14246 11612
rect 17494 11560 17500 11612
rect 17552 11600 17558 11612
rect 18601 11603 18659 11609
rect 18601 11600 18613 11603
rect 17552 11572 18613 11600
rect 17552 11560 17558 11572
rect 18601 11569 18613 11572
rect 18647 11569 18659 11603
rect 18601 11563 18659 11569
rect 6457 11535 6515 11541
rect 6457 11501 6469 11535
rect 6503 11501 6515 11535
rect 6457 11495 6515 11501
rect 6724 11535 6782 11541
rect 6724 11501 6736 11535
rect 6770 11532 6782 11535
rect 8588 11532 8616 11560
rect 6770 11504 8616 11532
rect 11977 11535 12035 11541
rect 6770 11501 6782 11504
rect 6724 11495 6782 11501
rect 11977 11501 11989 11535
rect 12023 11501 12035 11535
rect 11977 11495 12035 11501
rect 12244 11535 12302 11541
rect 12244 11501 12256 11535
rect 12290 11532 12302 11535
rect 12618 11532 12624 11544
rect 12290 11504 12624 11532
rect 12290 11501 12302 11504
rect 12244 11495 12302 11501
rect 6472 11464 6500 11495
rect 7558 11464 7564 11476
rect 6472 11436 7564 11464
rect 7558 11424 7564 11436
rect 7616 11424 7622 11476
rect 7742 11424 7748 11476
rect 7800 11464 7806 11476
rect 8573 11467 8631 11473
rect 8573 11464 8585 11467
rect 7800 11436 8585 11464
rect 7800 11424 7806 11436
rect 8573 11433 8585 11436
rect 8619 11464 8631 11467
rect 8938 11464 8944 11476
rect 8619 11436 8944 11464
rect 8619 11433 8631 11436
rect 8573 11427 8631 11433
rect 8938 11424 8944 11436
rect 8996 11424 9002 11476
rect 10781 11467 10839 11473
rect 10781 11433 10793 11467
rect 10827 11464 10839 11467
rect 11992 11464 12020 11495
rect 12618 11492 12624 11504
rect 12676 11492 12682 11544
rect 14090 11532 14096 11544
rect 14051 11504 14096 11532
rect 14090 11492 14096 11504
rect 14148 11492 14154 11544
rect 20254 11532 20260 11544
rect 20215 11504 20260 11532
rect 20254 11492 20260 11504
rect 20312 11492 20318 11544
rect 12802 11464 12808 11476
rect 10827 11436 11652 11464
rect 11992 11436 12808 11464
rect 10827 11433 10839 11436
rect 10781 11427 10839 11433
rect 8113 11399 8171 11405
rect 8113 11365 8125 11399
rect 8159 11396 8171 11399
rect 8202 11396 8208 11408
rect 8159 11368 8208 11396
rect 8159 11365 8171 11368
rect 8113 11359 8171 11365
rect 8202 11356 8208 11368
rect 8260 11356 8266 11408
rect 8478 11396 8484 11408
rect 8391 11368 8484 11396
rect 8478 11356 8484 11368
rect 8536 11396 8542 11408
rect 10594 11396 10600 11408
rect 8536 11368 10600 11396
rect 8536 11356 8542 11368
rect 10594 11356 10600 11368
rect 10652 11356 10658 11408
rect 10689 11399 10747 11405
rect 10689 11365 10701 11399
rect 10735 11396 10747 11399
rect 11333 11399 11391 11405
rect 11333 11396 11345 11399
rect 10735 11368 11345 11396
rect 10735 11365 10747 11368
rect 10689 11359 10747 11365
rect 11333 11365 11345 11368
rect 11379 11365 11391 11399
rect 11624 11396 11652 11436
rect 12802 11424 12808 11436
rect 12860 11464 12866 11476
rect 13722 11464 13728 11476
rect 12860 11436 13728 11464
rect 12860 11424 12866 11436
rect 13722 11424 13728 11436
rect 13780 11424 13786 11476
rect 18417 11467 18475 11473
rect 18417 11433 18429 11467
rect 18463 11464 18475 11467
rect 19061 11467 19119 11473
rect 19061 11464 19073 11467
rect 18463 11436 19073 11464
rect 18463 11433 18475 11436
rect 18417 11427 18475 11433
rect 19061 11433 19073 11436
rect 19107 11433 19119 11467
rect 19061 11427 19119 11433
rect 12986 11396 12992 11408
rect 11624 11368 12992 11396
rect 11333 11359 11391 11365
rect 12986 11356 12992 11368
rect 13044 11356 13050 11408
rect 13354 11396 13360 11408
rect 13315 11368 13360 11396
rect 13354 11356 13360 11368
rect 13412 11356 13418 11408
rect 13998 11396 14004 11408
rect 13959 11368 14004 11396
rect 13998 11356 14004 11368
rect 14056 11356 14062 11408
rect 18509 11399 18567 11405
rect 18509 11365 18521 11399
rect 18555 11396 18567 11399
rect 18874 11396 18880 11408
rect 18555 11368 18880 11396
rect 18555 11365 18567 11368
rect 18509 11359 18567 11365
rect 18874 11356 18880 11368
rect 18932 11356 18938 11408
rect 1104 11306 21620 11328
rect 1104 11254 7846 11306
rect 7898 11254 7910 11306
rect 7962 11254 7974 11306
rect 8026 11254 8038 11306
rect 8090 11254 14710 11306
rect 14762 11254 14774 11306
rect 14826 11254 14838 11306
rect 14890 11254 14902 11306
rect 14954 11254 21620 11306
rect 1104 11232 21620 11254
rect 8113 11195 8171 11201
rect 8113 11161 8125 11195
rect 8159 11192 8171 11195
rect 8202 11192 8208 11204
rect 8159 11164 8208 11192
rect 8159 11161 8171 11164
rect 8113 11155 8171 11161
rect 8202 11152 8208 11164
rect 8260 11152 8266 11204
rect 12250 11152 12256 11204
rect 12308 11192 12314 11204
rect 13633 11195 13691 11201
rect 12308 11164 13584 11192
rect 12308 11152 12314 11164
rect 14 11084 20 11136
rect 72 11124 78 11136
rect 13170 11124 13176 11136
rect 72 11096 13176 11124
rect 72 11084 78 11096
rect 13170 11084 13176 11096
rect 13228 11084 13234 11136
rect 13556 11124 13584 11164
rect 13633 11161 13645 11195
rect 13679 11192 13691 11195
rect 13998 11192 14004 11204
rect 13679 11164 14004 11192
rect 13679 11161 13691 11164
rect 13633 11155 13691 11161
rect 13998 11152 14004 11164
rect 14056 11152 14062 11204
rect 14090 11152 14096 11204
rect 14148 11192 14154 11204
rect 14274 11192 14280 11204
rect 14148 11164 14280 11192
rect 14148 11152 14154 11164
rect 14274 11152 14280 11164
rect 14332 11152 14338 11204
rect 15933 11195 15991 11201
rect 15933 11161 15945 11195
rect 15979 11192 15991 11195
rect 17405 11195 17463 11201
rect 17405 11192 17417 11195
rect 15979 11164 17417 11192
rect 15979 11161 15991 11164
rect 15933 11155 15991 11161
rect 17405 11161 17417 11164
rect 17451 11161 17463 11195
rect 18874 11192 18880 11204
rect 18835 11164 18880 11192
rect 17405 11155 17463 11161
rect 18874 11152 18880 11164
rect 18932 11152 18938 11204
rect 20165 11195 20223 11201
rect 20165 11161 20177 11195
rect 20211 11192 20223 11195
rect 20622 11192 20628 11204
rect 20211 11164 20628 11192
rect 20211 11161 20223 11164
rect 20165 11155 20223 11161
rect 20622 11152 20628 11164
rect 20680 11152 20686 11204
rect 20717 11195 20775 11201
rect 20717 11161 20729 11195
rect 20763 11192 20775 11195
rect 20806 11192 20812 11204
rect 20763 11164 20812 11192
rect 20763 11161 20775 11164
rect 20717 11155 20775 11161
rect 20806 11152 20812 11164
rect 20864 11152 20870 11204
rect 16393 11127 16451 11133
rect 16393 11124 16405 11127
rect 13556 11096 16405 11124
rect 16393 11093 16405 11096
rect 16439 11093 16451 11127
rect 16393 11087 16451 11093
rect 16482 11084 16488 11136
rect 16540 11124 16546 11136
rect 16540 11096 20576 11124
rect 16540 11084 16546 11096
rect 6822 11016 6828 11068
rect 6880 11056 6886 11068
rect 8205 11059 8263 11065
rect 8205 11056 8217 11059
rect 6880 11028 8217 11056
rect 6880 11016 6886 11028
rect 8205 11025 8217 11028
rect 8251 11025 8263 11059
rect 8205 11019 8263 11025
rect 14001 11059 14059 11065
rect 14001 11025 14013 11059
rect 14047 11056 14059 11059
rect 14645 11059 14703 11065
rect 14645 11056 14657 11059
rect 14047 11028 14657 11056
rect 14047 11025 14059 11028
rect 14001 11019 14059 11025
rect 14645 11025 14657 11028
rect 14691 11025 14703 11059
rect 14645 11019 14703 11025
rect 16114 11016 16120 11068
rect 16172 11056 16178 11068
rect 16301 11059 16359 11065
rect 16301 11056 16313 11059
rect 16172 11028 16313 11056
rect 16172 11016 16178 11028
rect 16301 11025 16313 11028
rect 16347 11025 16359 11059
rect 17310 11056 17316 11068
rect 17271 11028 17316 11056
rect 16301 11019 16359 11025
rect 17310 11016 17316 11028
rect 17368 11016 17374 11068
rect 17402 11016 17408 11068
rect 17460 11056 17466 11068
rect 17862 11056 17868 11068
rect 17460 11028 17868 11056
rect 17460 11016 17466 11028
rect 17862 11016 17868 11028
rect 17920 11056 17926 11068
rect 19245 11059 19303 11065
rect 19245 11056 19257 11059
rect 17920 11028 19257 11056
rect 17920 11016 17926 11028
rect 19245 11025 19257 11028
rect 19291 11025 19303 11059
rect 19978 11056 19984 11068
rect 19939 11028 19984 11056
rect 19245 11019 19303 11025
rect 19978 11016 19984 11028
rect 20036 11016 20042 11068
rect 20548 11065 20576 11096
rect 20533 11059 20591 11065
rect 20533 11025 20545 11059
rect 20579 11025 20591 11059
rect 20533 11019 20591 11025
rect 8386 10988 8392 11000
rect 8347 10960 8392 10988
rect 8386 10948 8392 10960
rect 8444 10948 8450 11000
rect 12986 10948 12992 11000
rect 13044 10988 13050 11000
rect 14090 10988 14096 11000
rect 13044 10960 14096 10988
rect 13044 10948 13050 10960
rect 14090 10948 14096 10960
rect 14148 10948 14154 11000
rect 14185 10991 14243 10997
rect 14185 10957 14197 10991
rect 14231 10957 14243 10991
rect 16482 10988 16488 11000
rect 16443 10960 16488 10988
rect 14185 10951 14243 10957
rect 7745 10923 7803 10929
rect 7745 10889 7757 10923
rect 7791 10920 7803 10923
rect 10410 10920 10416 10932
rect 7791 10892 10416 10920
rect 7791 10889 7803 10892
rect 7745 10883 7803 10889
rect 10410 10880 10416 10892
rect 10468 10880 10474 10932
rect 13354 10880 13360 10932
rect 13412 10920 13418 10932
rect 14200 10920 14228 10951
rect 16482 10948 16488 10960
rect 16540 10948 16546 11000
rect 17494 10988 17500 11000
rect 16776 10960 17356 10988
rect 17455 10960 17500 10988
rect 13412 10892 14228 10920
rect 13412 10880 13418 10892
rect 15654 10880 15660 10932
rect 15712 10920 15718 10932
rect 15930 10920 15936 10932
rect 15712 10892 15936 10920
rect 15712 10880 15718 10892
rect 15930 10880 15936 10892
rect 15988 10920 15994 10932
rect 16776 10920 16804 10960
rect 16942 10920 16948 10932
rect 15988 10892 16804 10920
rect 16903 10892 16948 10920
rect 15988 10880 15994 10892
rect 16942 10880 16948 10892
rect 17000 10880 17006 10932
rect 17328 10920 17356 10960
rect 17494 10948 17500 10960
rect 17552 10948 17558 11000
rect 19337 10991 19395 10997
rect 19337 10988 19349 10991
rect 17604 10960 19349 10988
rect 17604 10920 17632 10960
rect 19337 10957 19349 10960
rect 19383 10957 19395 10991
rect 19337 10951 19395 10957
rect 19429 10991 19487 10997
rect 19429 10957 19441 10991
rect 19475 10957 19487 10991
rect 19429 10951 19487 10957
rect 17328 10892 17632 10920
rect 19242 10880 19248 10932
rect 19300 10920 19306 10932
rect 19444 10920 19472 10951
rect 19300 10892 19472 10920
rect 19300 10880 19306 10892
rect 1104 10762 21620 10784
rect 1104 10710 4414 10762
rect 4466 10710 4478 10762
rect 4530 10710 4542 10762
rect 4594 10710 4606 10762
rect 4658 10710 11278 10762
rect 11330 10710 11342 10762
rect 11394 10710 11406 10762
rect 11458 10710 11470 10762
rect 11522 10710 18142 10762
rect 18194 10710 18206 10762
rect 18258 10710 18270 10762
rect 18322 10710 18334 10762
rect 18386 10710 21620 10762
rect 1104 10688 21620 10710
rect 8570 10648 8576 10660
rect 8531 10620 8576 10648
rect 8570 10608 8576 10620
rect 8628 10608 8634 10660
rect 16485 10651 16543 10657
rect 16485 10617 16497 10651
rect 16531 10648 16543 10651
rect 17310 10648 17316 10660
rect 16531 10620 17316 10648
rect 16531 10617 16543 10620
rect 16485 10611 16543 10617
rect 17310 10608 17316 10620
rect 17368 10608 17374 10660
rect 19334 10608 19340 10660
rect 19392 10648 19398 10660
rect 20441 10651 20499 10657
rect 20441 10648 20453 10651
rect 19392 10620 20453 10648
rect 19392 10608 19398 10620
rect 20441 10617 20453 10620
rect 20487 10617 20499 10651
rect 20441 10611 20499 10617
rect 10045 10583 10103 10589
rect 10045 10549 10057 10583
rect 10091 10580 10103 10583
rect 16390 10580 16396 10592
rect 10091 10552 11100 10580
rect 10091 10549 10103 10552
rect 10045 10543 10103 10549
rect 10597 10515 10655 10521
rect 10597 10512 10609 10515
rect 10152 10484 10609 10512
rect 7193 10447 7251 10453
rect 7193 10413 7205 10447
rect 7239 10413 7251 10447
rect 7193 10407 7251 10413
rect 7208 10308 7236 10407
rect 7460 10379 7518 10385
rect 7460 10345 7472 10379
rect 7506 10376 7518 10379
rect 9858 10376 9864 10388
rect 7506 10348 9864 10376
rect 7506 10345 7518 10348
rect 7460 10339 7518 10345
rect 9858 10336 9864 10348
rect 9916 10376 9922 10388
rect 10152 10376 10180 10484
rect 10597 10481 10609 10484
rect 10643 10481 10655 10515
rect 10597 10475 10655 10481
rect 11072 10453 11100 10552
rect 11348 10552 16396 10580
rect 11348 10521 11376 10552
rect 16390 10540 16396 10552
rect 16448 10540 16454 10592
rect 11333 10515 11391 10521
rect 11333 10481 11345 10515
rect 11379 10481 11391 10515
rect 11333 10475 11391 10481
rect 16482 10472 16488 10524
rect 16540 10512 16546 10524
rect 17129 10515 17187 10521
rect 17129 10512 17141 10515
rect 16540 10484 17141 10512
rect 16540 10472 16546 10484
rect 17129 10481 17141 10484
rect 17175 10512 17187 10515
rect 19242 10512 19248 10524
rect 17175 10484 19248 10512
rect 17175 10481 17187 10484
rect 17129 10475 17187 10481
rect 19242 10472 19248 10484
rect 19300 10472 19306 10524
rect 11057 10447 11115 10453
rect 11057 10413 11069 10447
rect 11103 10413 11115 10447
rect 11057 10407 11115 10413
rect 11606 10404 11612 10456
rect 11664 10444 11670 10456
rect 20254 10444 20260 10456
rect 11664 10416 16988 10444
rect 20215 10416 20260 10444
rect 11664 10404 11670 10416
rect 10410 10376 10416 10388
rect 9916 10348 10180 10376
rect 10371 10348 10416 10376
rect 9916 10336 9922 10348
rect 10410 10336 10416 10348
rect 10468 10336 10474 10388
rect 11238 10336 11244 10388
rect 11296 10376 11302 10388
rect 11790 10376 11796 10388
rect 11296 10348 11796 10376
rect 11296 10336 11302 10348
rect 11790 10336 11796 10348
rect 11848 10376 11854 10388
rect 11848 10348 16804 10376
rect 11848 10336 11854 10348
rect 16776 10320 16804 10348
rect 7558 10308 7564 10320
rect 7208 10280 7564 10308
rect 7558 10268 7564 10280
rect 7616 10268 7622 10320
rect 10502 10308 10508 10320
rect 10463 10280 10508 10308
rect 10502 10268 10508 10280
rect 10560 10268 10566 10320
rect 16758 10268 16764 10320
rect 16816 10308 16822 10320
rect 16960 10317 16988 10416
rect 20254 10404 20260 10416
rect 20312 10404 20318 10456
rect 16853 10311 16911 10317
rect 16853 10308 16865 10311
rect 16816 10280 16865 10308
rect 16816 10268 16822 10280
rect 16853 10277 16865 10280
rect 16899 10277 16911 10311
rect 16853 10271 16911 10277
rect 16945 10311 17003 10317
rect 16945 10277 16957 10311
rect 16991 10308 17003 10311
rect 18690 10308 18696 10320
rect 16991 10280 18696 10308
rect 16991 10277 17003 10280
rect 16945 10271 17003 10277
rect 18690 10268 18696 10280
rect 18748 10268 18754 10320
rect 1104 10218 21620 10240
rect 1104 10166 7846 10218
rect 7898 10166 7910 10218
rect 7962 10166 7974 10218
rect 8026 10166 8038 10218
rect 8090 10166 14710 10218
rect 14762 10166 14774 10218
rect 14826 10166 14838 10218
rect 14890 10166 14902 10218
rect 14954 10166 21620 10218
rect 1104 10144 21620 10166
rect 9858 10104 9864 10116
rect 9819 10076 9864 10104
rect 9858 10064 9864 10076
rect 9916 10064 9922 10116
rect 11238 10104 11244 10116
rect 11199 10076 11244 10104
rect 11238 10064 11244 10076
rect 11296 10064 11302 10116
rect 11333 10107 11391 10113
rect 11333 10073 11345 10107
rect 11379 10104 11391 10107
rect 11606 10104 11612 10116
rect 11379 10076 11612 10104
rect 11379 10073 11391 10076
rect 11333 10067 11391 10073
rect 11606 10064 11612 10076
rect 11664 10064 11670 10116
rect 14182 10104 14188 10116
rect 14143 10076 14188 10104
rect 14182 10064 14188 10076
rect 14240 10064 14246 10116
rect 17313 10107 17371 10113
rect 17313 10073 17325 10107
rect 17359 10104 17371 10107
rect 17494 10104 17500 10116
rect 17359 10076 17500 10104
rect 17359 10073 17371 10076
rect 17313 10067 17371 10073
rect 17494 10064 17500 10076
rect 17552 10064 17558 10116
rect 19242 10064 19248 10116
rect 19300 10104 19306 10116
rect 19889 10107 19947 10113
rect 19889 10104 19901 10107
rect 19300 10076 19901 10104
rect 19300 10064 19306 10076
rect 19889 10073 19901 10076
rect 19935 10073 19947 10107
rect 19889 10067 19947 10073
rect 20717 10107 20775 10113
rect 20717 10073 20729 10107
rect 20763 10104 20775 10107
rect 20990 10104 20996 10116
rect 20763 10076 20996 10104
rect 20763 10073 20775 10076
rect 20717 10067 20775 10073
rect 20990 10064 20996 10076
rect 21048 10064 21054 10116
rect 13072 10039 13130 10045
rect 13072 10005 13084 10039
rect 13118 10036 13130 10039
rect 13354 10036 13360 10048
rect 13118 10008 13360 10036
rect 13118 10005 13130 10008
rect 13072 9999 13130 10005
rect 13354 9996 13360 10008
rect 13412 9996 13418 10048
rect 16200 10039 16258 10045
rect 16200 10005 16212 10039
rect 16246 10036 16258 10039
rect 16482 10036 16488 10048
rect 16246 10008 16488 10036
rect 16246 10005 16258 10008
rect 16200 9999 16258 10005
rect 16482 9996 16488 10008
rect 16540 9996 16546 10048
rect 8754 9977 8760 9980
rect 8748 9968 8760 9977
rect 8715 9940 8760 9968
rect 8748 9931 8760 9940
rect 8754 9928 8760 9931
rect 8812 9928 8818 9980
rect 12802 9968 12808 9980
rect 12715 9940 12808 9968
rect 12802 9928 12808 9940
rect 12860 9968 12866 9980
rect 13630 9968 13636 9980
rect 12860 9940 13636 9968
rect 12860 9928 12866 9940
rect 13630 9928 13636 9940
rect 13688 9968 13694 9980
rect 15933 9971 15991 9977
rect 15933 9968 15945 9971
rect 13688 9940 15945 9968
rect 13688 9928 13694 9940
rect 15933 9937 15945 9940
rect 15979 9968 15991 9971
rect 16666 9968 16672 9980
rect 15979 9940 16672 9968
rect 15979 9937 15991 9940
rect 15933 9931 15991 9937
rect 16666 9928 16672 9940
rect 16724 9968 16730 9980
rect 17954 9968 17960 9980
rect 16724 9940 17960 9968
rect 16724 9928 16730 9940
rect 17954 9928 17960 9940
rect 18012 9968 18018 9980
rect 18782 9977 18788 9980
rect 18509 9971 18567 9977
rect 18509 9968 18521 9971
rect 18012 9940 18521 9968
rect 18012 9928 18018 9940
rect 18509 9937 18521 9940
rect 18555 9937 18567 9971
rect 18776 9968 18788 9977
rect 18743 9940 18788 9968
rect 18509 9931 18567 9937
rect 18776 9931 18788 9940
rect 18782 9928 18788 9931
rect 18840 9928 18846 9980
rect 20530 9968 20536 9980
rect 20491 9940 20536 9968
rect 20530 9928 20536 9940
rect 20588 9928 20594 9980
rect 7558 9860 7564 9912
rect 7616 9900 7622 9912
rect 8481 9903 8539 9909
rect 8481 9900 8493 9903
rect 7616 9872 8493 9900
rect 7616 9860 7622 9872
rect 8481 9869 8493 9872
rect 8527 9869 8539 9903
rect 8481 9863 8539 9869
rect 11517 9903 11575 9909
rect 11517 9869 11529 9903
rect 11563 9900 11575 9903
rect 11606 9900 11612 9912
rect 11563 9872 11612 9900
rect 11563 9869 11575 9872
rect 11517 9863 11575 9869
rect 11606 9860 11612 9872
rect 11664 9860 11670 9912
rect 10870 9764 10876 9776
rect 10831 9736 10876 9764
rect 10870 9724 10876 9736
rect 10928 9724 10934 9776
rect 1104 9674 21620 9696
rect 1104 9622 4414 9674
rect 4466 9622 4478 9674
rect 4530 9622 4542 9674
rect 4594 9622 4606 9674
rect 4658 9622 11278 9674
rect 11330 9622 11342 9674
rect 11394 9622 11406 9674
rect 11458 9622 11470 9674
rect 11522 9622 18142 9674
rect 18194 9622 18206 9674
rect 18258 9622 18270 9674
rect 18322 9622 18334 9674
rect 18386 9622 21620 9674
rect 1104 9600 21620 9622
rect 9953 9563 10011 9569
rect 9953 9529 9965 9563
rect 9999 9560 10011 9563
rect 10502 9560 10508 9572
rect 9999 9532 10508 9560
rect 9999 9529 10011 9532
rect 9953 9523 10011 9529
rect 10502 9520 10508 9532
rect 10560 9520 10566 9572
rect 8754 9452 8760 9504
rect 8812 9492 8818 9504
rect 8941 9495 8999 9501
rect 8941 9492 8953 9495
rect 8812 9464 8953 9492
rect 8812 9452 8818 9464
rect 8941 9461 8953 9464
rect 8987 9461 8999 9495
rect 8941 9455 8999 9461
rect 11256 9464 13492 9492
rect 8956 9424 8984 9455
rect 10594 9424 10600 9436
rect 8956 9396 10600 9424
rect 10594 9384 10600 9396
rect 10652 9384 10658 9436
rect 7558 9356 7564 9368
rect 7519 9328 7564 9356
rect 7558 9316 7564 9328
rect 7616 9316 7622 9368
rect 10321 9359 10379 9365
rect 10321 9325 10333 9359
rect 10367 9356 10379 9359
rect 10870 9356 10876 9368
rect 10367 9328 10876 9356
rect 10367 9325 10379 9328
rect 10321 9319 10379 9325
rect 10870 9316 10876 9328
rect 10928 9316 10934 9368
rect 11256 9356 11284 9464
rect 11517 9427 11575 9433
rect 11517 9424 11529 9427
rect 11440 9396 11529 9424
rect 11333 9359 11391 9365
rect 11333 9356 11345 9359
rect 11256 9328 11345 9356
rect 11333 9325 11345 9328
rect 11379 9325 11391 9359
rect 11333 9319 11391 9325
rect 7828 9291 7886 9297
rect 7828 9257 7840 9291
rect 7874 9288 7886 9291
rect 11440 9288 11468 9396
rect 11517 9393 11529 9396
rect 11563 9424 11575 9427
rect 11606 9424 11612 9436
rect 11563 9396 11612 9424
rect 11563 9393 11575 9396
rect 11517 9387 11575 9393
rect 11606 9384 11612 9396
rect 11664 9424 11670 9436
rect 12713 9427 12771 9433
rect 12713 9424 12725 9427
rect 11664 9396 12725 9424
rect 11664 9384 11670 9396
rect 12713 9393 12725 9396
rect 12759 9393 12771 9427
rect 12713 9387 12771 9393
rect 7874 9260 11468 9288
rect 7874 9257 7886 9260
rect 7828 9251 7886 9257
rect 12342 9248 12348 9300
rect 12400 9288 12406 9300
rect 12529 9291 12587 9297
rect 12529 9288 12541 9291
rect 12400 9260 12541 9288
rect 12400 9248 12406 9260
rect 12529 9257 12541 9260
rect 12575 9257 12587 9291
rect 12529 9251 12587 9257
rect 10413 9223 10471 9229
rect 10413 9189 10425 9223
rect 10459 9220 10471 9223
rect 10965 9223 11023 9229
rect 10965 9220 10977 9223
rect 10459 9192 10977 9220
rect 10459 9189 10471 9192
rect 10413 9183 10471 9189
rect 10965 9189 10977 9192
rect 11011 9189 11023 9223
rect 11422 9220 11428 9232
rect 11383 9192 11428 9220
rect 10965 9183 11023 9189
rect 11422 9180 11428 9192
rect 11480 9180 11486 9232
rect 12066 9220 12072 9232
rect 12027 9192 12072 9220
rect 12066 9180 12072 9192
rect 12124 9180 12130 9232
rect 12434 9180 12440 9232
rect 12492 9220 12498 9232
rect 12728 9220 12756 9387
rect 13464 9288 13492 9464
rect 16114 9452 16120 9504
rect 16172 9492 16178 9504
rect 16390 9492 16396 9504
rect 16172 9464 16396 9492
rect 16172 9452 16178 9464
rect 16390 9452 16396 9464
rect 16448 9452 16454 9504
rect 17586 9492 17592 9504
rect 17547 9464 17592 9492
rect 17586 9452 17592 9464
rect 17644 9452 17650 9504
rect 13541 9359 13599 9365
rect 13541 9325 13553 9359
rect 13587 9356 13599 9359
rect 13630 9356 13636 9368
rect 13587 9328 13636 9356
rect 13587 9325 13599 9328
rect 13541 9319 13599 9325
rect 13630 9316 13636 9328
rect 13688 9316 13694 9368
rect 13808 9359 13866 9365
rect 13808 9325 13820 9359
rect 13854 9356 13866 9359
rect 14182 9356 14188 9368
rect 13854 9328 14188 9356
rect 13854 9325 13866 9328
rect 13808 9319 13866 9325
rect 14182 9316 14188 9328
rect 14240 9316 14246 9368
rect 16132 9288 16160 9452
rect 18230 9424 18236 9436
rect 18191 9396 18236 9424
rect 18230 9384 18236 9396
rect 18288 9384 18294 9436
rect 19245 9427 19303 9433
rect 19245 9393 19257 9427
rect 19291 9424 19303 9427
rect 19426 9424 19432 9436
rect 19291 9396 19432 9424
rect 19291 9393 19303 9396
rect 19245 9387 19303 9393
rect 19426 9384 19432 9396
rect 19484 9384 19490 9436
rect 18966 9356 18972 9368
rect 18927 9328 18972 9356
rect 18966 9316 18972 9328
rect 19024 9316 19030 9368
rect 13464 9260 16160 9288
rect 17957 9291 18015 9297
rect 17957 9257 17969 9291
rect 18003 9288 18015 9291
rect 19613 9291 19671 9297
rect 19613 9288 19625 9291
rect 18003 9260 19625 9288
rect 18003 9257 18015 9260
rect 17957 9251 18015 9257
rect 19613 9257 19625 9260
rect 19659 9257 19671 9291
rect 19613 9251 19671 9257
rect 14921 9223 14979 9229
rect 14921 9220 14933 9223
rect 12492 9192 12537 9220
rect 12728 9192 14933 9220
rect 12492 9180 12498 9192
rect 14921 9189 14933 9192
rect 14967 9189 14979 9223
rect 14921 9183 14979 9189
rect 18049 9223 18107 9229
rect 18049 9189 18061 9223
rect 18095 9220 18107 9223
rect 18601 9223 18659 9229
rect 18601 9220 18613 9223
rect 18095 9192 18613 9220
rect 18095 9189 18107 9192
rect 18049 9183 18107 9189
rect 18601 9189 18613 9192
rect 18647 9189 18659 9223
rect 19058 9220 19064 9232
rect 19019 9192 19064 9220
rect 18601 9183 18659 9189
rect 19058 9180 19064 9192
rect 19116 9180 19122 9232
rect 1104 9130 21620 9152
rect 1104 9078 7846 9130
rect 7898 9078 7910 9130
rect 7962 9078 7974 9130
rect 8026 9078 8038 9130
rect 8090 9078 14710 9130
rect 14762 9078 14774 9130
rect 14826 9078 14838 9130
rect 14890 9078 14902 9130
rect 14954 9078 21620 9130
rect 1104 9056 21620 9078
rect 10410 8976 10416 9028
rect 10468 9016 10474 9028
rect 10597 9019 10655 9025
rect 10597 9016 10609 9019
rect 10468 8988 10609 9016
rect 10468 8976 10474 8988
rect 10597 8985 10609 8988
rect 10643 8985 10655 9019
rect 10597 8979 10655 8985
rect 11057 9019 11115 9025
rect 11057 8985 11069 9019
rect 11103 9016 11115 9019
rect 12066 9016 12072 9028
rect 11103 8988 12072 9016
rect 11103 8985 11115 8988
rect 11057 8979 11115 8985
rect 12066 8976 12072 8988
rect 12124 8976 12130 9028
rect 13078 8976 13084 9028
rect 13136 9016 13142 9028
rect 13357 9019 13415 9025
rect 13357 9016 13369 9019
rect 13136 8988 13369 9016
rect 13136 8976 13142 8988
rect 13357 8985 13369 8988
rect 13403 8985 13415 9019
rect 13357 8979 13415 8985
rect 15102 8976 15108 9028
rect 15160 9016 15166 9028
rect 15289 9019 15347 9025
rect 15289 9016 15301 9019
rect 15160 8988 15301 9016
rect 15160 8976 15166 8988
rect 15289 8985 15301 8988
rect 15335 8985 15347 9019
rect 17862 9016 17868 9028
rect 15289 8979 15347 8985
rect 15396 8988 17868 9016
rect 2682 8908 2688 8960
rect 2740 8948 2746 8960
rect 11422 8948 11428 8960
rect 2740 8920 11428 8948
rect 2740 8908 2746 8920
rect 11422 8908 11428 8920
rect 11480 8908 11486 8960
rect 12434 8908 12440 8960
rect 12492 8948 12498 8960
rect 15396 8948 15424 8988
rect 17862 8976 17868 8988
rect 17920 8976 17926 9028
rect 18230 8976 18236 9028
rect 18288 9016 18294 9028
rect 18782 9016 18788 9028
rect 18288 8988 18788 9016
rect 18288 8976 18294 8988
rect 18782 8976 18788 8988
rect 18840 9016 18846 9028
rect 19521 9019 19579 9025
rect 19521 9016 19533 9019
rect 18840 8988 19533 9016
rect 18840 8976 18846 8988
rect 19521 8985 19533 8988
rect 19567 8985 19579 9019
rect 19521 8979 19579 8985
rect 20070 8976 20076 9028
rect 20128 9016 20134 9028
rect 20165 9019 20223 9025
rect 20165 9016 20177 9019
rect 20128 8988 20177 9016
rect 20128 8976 20134 8988
rect 20165 8985 20177 8988
rect 20211 8985 20223 9019
rect 20165 8979 20223 8985
rect 20717 9019 20775 9025
rect 20717 8985 20729 9019
rect 20763 8985 20775 9019
rect 20717 8979 20775 8985
rect 12492 8920 15424 8948
rect 12492 8908 12498 8920
rect 16298 8908 16304 8960
rect 16356 8948 16362 8960
rect 20732 8948 20760 8979
rect 16356 8920 20760 8948
rect 16356 8908 16362 8920
rect 10965 8883 11023 8889
rect 10965 8849 10977 8883
rect 11011 8880 11023 8883
rect 11609 8883 11667 8889
rect 11609 8880 11621 8883
rect 11011 8852 11621 8880
rect 11011 8849 11023 8852
rect 10965 8843 11023 8849
rect 11609 8849 11621 8852
rect 11655 8849 11667 8883
rect 11609 8843 11667 8849
rect 13173 8883 13231 8889
rect 13173 8849 13185 8883
rect 13219 8880 13231 8883
rect 13446 8880 13452 8892
rect 13219 8852 13452 8880
rect 13219 8849 13231 8852
rect 13173 8843 13231 8849
rect 13446 8840 13452 8852
rect 13504 8840 13510 8892
rect 15105 8883 15163 8889
rect 15105 8849 15117 8883
rect 15151 8880 15163 8883
rect 15654 8880 15660 8892
rect 15151 8852 15660 8880
rect 15151 8849 15163 8852
rect 15105 8843 15163 8849
rect 15654 8840 15660 8852
rect 15712 8840 15718 8892
rect 17954 8840 17960 8892
rect 18012 8880 18018 8892
rect 18141 8883 18199 8889
rect 18141 8880 18153 8883
rect 18012 8852 18153 8880
rect 18012 8840 18018 8852
rect 18141 8849 18153 8852
rect 18187 8849 18199 8883
rect 18141 8843 18199 8849
rect 18408 8883 18466 8889
rect 18408 8849 18420 8883
rect 18454 8880 18466 8883
rect 19426 8880 19432 8892
rect 18454 8852 19432 8880
rect 18454 8849 18466 8852
rect 18408 8843 18466 8849
rect 19426 8840 19432 8852
rect 19484 8840 19490 8892
rect 19978 8880 19984 8892
rect 19939 8852 19984 8880
rect 19978 8840 19984 8852
rect 20036 8840 20042 8892
rect 20530 8880 20536 8892
rect 20491 8852 20536 8880
rect 20530 8840 20536 8852
rect 20588 8840 20594 8892
rect 10594 8772 10600 8824
rect 10652 8812 10658 8824
rect 11149 8815 11207 8821
rect 11149 8812 11161 8815
rect 10652 8784 11161 8812
rect 10652 8772 10658 8784
rect 11149 8781 11161 8784
rect 11195 8781 11207 8815
rect 11149 8775 11207 8781
rect 12342 8772 12348 8824
rect 12400 8812 12406 8824
rect 15930 8812 15936 8824
rect 12400 8784 15936 8812
rect 12400 8772 12406 8784
rect 15930 8772 15936 8784
rect 15988 8772 15994 8824
rect 18506 8636 18512 8688
rect 18564 8676 18570 8688
rect 18782 8676 18788 8688
rect 18564 8648 18788 8676
rect 18564 8636 18570 8648
rect 18782 8636 18788 8648
rect 18840 8636 18846 8688
rect 1104 8586 21620 8608
rect 1104 8534 4414 8586
rect 4466 8534 4478 8586
rect 4530 8534 4542 8586
rect 4594 8534 4606 8586
rect 4658 8534 11278 8586
rect 11330 8534 11342 8586
rect 11394 8534 11406 8586
rect 11458 8534 11470 8586
rect 11522 8534 18142 8586
rect 18194 8534 18206 8586
rect 18258 8534 18270 8586
rect 18322 8534 18334 8586
rect 18386 8534 21620 8586
rect 1104 8512 21620 8534
rect 11517 8475 11575 8481
rect 11517 8441 11529 8475
rect 11563 8472 11575 8475
rect 11974 8472 11980 8484
rect 11563 8444 11980 8472
rect 11563 8441 11575 8444
rect 11517 8435 11575 8441
rect 11974 8432 11980 8444
rect 12032 8432 12038 8484
rect 20438 8472 20444 8484
rect 20399 8444 20444 8472
rect 20438 8432 20444 8444
rect 20496 8432 20502 8484
rect 16209 8407 16267 8413
rect 16209 8373 16221 8407
rect 16255 8373 16267 8407
rect 16209 8367 16267 8373
rect 13446 8336 13452 8348
rect 13407 8308 13452 8336
rect 13446 8296 13452 8308
rect 13504 8296 13510 8348
rect 15654 8336 15660 8348
rect 15615 8308 15660 8336
rect 15654 8296 15660 8308
rect 15712 8296 15718 8348
rect 11330 8268 11336 8280
rect 11291 8240 11336 8268
rect 11330 8228 11336 8240
rect 11388 8228 11394 8280
rect 13262 8268 13268 8280
rect 13223 8240 13268 8268
rect 13262 8228 13268 8240
rect 13320 8228 13326 8280
rect 15473 8271 15531 8277
rect 15473 8237 15485 8271
rect 15519 8268 15531 8271
rect 16224 8268 16252 8367
rect 16853 8339 16911 8345
rect 16853 8305 16865 8339
rect 16899 8336 16911 8339
rect 17402 8336 17408 8348
rect 16899 8308 17408 8336
rect 16899 8305 16911 8308
rect 16853 8299 16911 8305
rect 17402 8296 17408 8308
rect 17460 8296 17466 8348
rect 16666 8268 16672 8280
rect 15519 8240 16252 8268
rect 16627 8240 16672 8268
rect 15519 8237 15531 8240
rect 15473 8231 15531 8237
rect 16666 8228 16672 8240
rect 16724 8228 16730 8280
rect 20254 8268 20260 8280
rect 20215 8240 20260 8268
rect 20254 8228 20260 8240
rect 20312 8228 20318 8280
rect 16577 8203 16635 8209
rect 16577 8169 16589 8203
rect 16623 8200 16635 8203
rect 17221 8203 17279 8209
rect 17221 8200 17233 8203
rect 16623 8172 17233 8200
rect 16623 8169 16635 8172
rect 16577 8163 16635 8169
rect 17221 8169 17233 8172
rect 17267 8169 17279 8203
rect 17221 8163 17279 8169
rect 1104 8042 21620 8064
rect 1104 7990 7846 8042
rect 7898 7990 7910 8042
rect 7962 7990 7974 8042
rect 8026 7990 8038 8042
rect 8090 7990 14710 8042
rect 14762 7990 14774 8042
rect 14826 7990 14838 8042
rect 14890 7990 14902 8042
rect 14954 7990 21620 8042
rect 1104 7968 21620 7990
rect 13262 7888 13268 7940
rect 13320 7928 13326 7940
rect 13633 7931 13691 7937
rect 13633 7928 13645 7931
rect 13320 7900 13645 7928
rect 13320 7888 13326 7900
rect 13633 7897 13645 7900
rect 13679 7897 13691 7931
rect 17402 7928 17408 7940
rect 17363 7900 17408 7928
rect 13633 7891 13691 7897
rect 17402 7888 17408 7900
rect 17460 7888 17466 7940
rect 19426 7928 19432 7940
rect 19387 7900 19432 7928
rect 19426 7888 19432 7900
rect 19484 7888 19490 7940
rect 10873 7863 10931 7869
rect 10873 7829 10885 7863
rect 10919 7860 10931 7863
rect 11330 7860 11336 7872
rect 10919 7832 11336 7860
rect 10919 7829 10931 7832
rect 10873 7823 10931 7829
rect 11330 7820 11336 7832
rect 11388 7820 11394 7872
rect 14366 7820 14372 7872
rect 14424 7860 14430 7872
rect 17420 7860 17448 7888
rect 18294 7863 18352 7869
rect 18294 7860 18306 7863
rect 14424 7832 17356 7860
rect 17420 7832 18306 7860
rect 14424 7820 14430 7832
rect 10318 7752 10324 7804
rect 10376 7792 10382 7804
rect 10597 7795 10655 7801
rect 10597 7792 10609 7795
rect 10376 7764 10609 7792
rect 10376 7752 10382 7764
rect 10597 7761 10609 7764
rect 10643 7761 10655 7795
rect 10597 7755 10655 7761
rect 14001 7795 14059 7801
rect 14001 7761 14013 7795
rect 14047 7792 14059 7795
rect 14642 7792 14648 7804
rect 14047 7764 14648 7792
rect 14047 7761 14059 7764
rect 14001 7755 14059 7761
rect 14642 7752 14648 7764
rect 14700 7752 14706 7804
rect 16292 7795 16350 7801
rect 16292 7761 16304 7795
rect 16338 7792 16350 7795
rect 16574 7792 16580 7804
rect 16338 7764 16580 7792
rect 16338 7761 16350 7764
rect 16292 7755 16350 7761
rect 16574 7752 16580 7764
rect 16632 7752 16638 7804
rect 17328 7792 17356 7832
rect 18294 7829 18306 7832
rect 18340 7829 18352 7863
rect 18294 7823 18352 7829
rect 19978 7792 19984 7804
rect 17328 7764 19104 7792
rect 19939 7764 19984 7792
rect 14090 7724 14096 7736
rect 14051 7696 14096 7724
rect 14090 7684 14096 7696
rect 14148 7684 14154 7736
rect 14274 7724 14280 7736
rect 14235 7696 14280 7724
rect 14274 7684 14280 7696
rect 14332 7684 14338 7736
rect 16022 7724 16028 7736
rect 15983 7696 16028 7724
rect 16022 7684 16028 7696
rect 16080 7684 16086 7736
rect 17954 7684 17960 7736
rect 18012 7724 18018 7736
rect 18049 7727 18107 7733
rect 18049 7724 18061 7727
rect 18012 7696 18061 7724
rect 18012 7684 18018 7696
rect 18049 7693 18061 7696
rect 18095 7693 18107 7727
rect 18049 7687 18107 7693
rect 19076 7656 19104 7764
rect 19978 7752 19984 7764
rect 20036 7752 20042 7804
rect 20530 7792 20536 7804
rect 20491 7764 20536 7792
rect 20530 7752 20536 7764
rect 20588 7752 20594 7804
rect 20717 7659 20775 7665
rect 20717 7656 20729 7659
rect 19076 7628 20729 7656
rect 20717 7625 20729 7628
rect 20763 7625 20775 7659
rect 20717 7619 20775 7625
rect 16206 7548 16212 7600
rect 16264 7588 16270 7600
rect 20165 7591 20223 7597
rect 20165 7588 20177 7591
rect 16264 7560 20177 7588
rect 16264 7548 16270 7560
rect 20165 7557 20177 7560
rect 20211 7557 20223 7591
rect 20165 7551 20223 7557
rect 1104 7498 21620 7520
rect 1104 7446 4414 7498
rect 4466 7446 4478 7498
rect 4530 7446 4542 7498
rect 4594 7446 4606 7498
rect 4658 7446 11278 7498
rect 11330 7446 11342 7498
rect 11394 7446 11406 7498
rect 11458 7446 11470 7498
rect 11522 7446 18142 7498
rect 18194 7446 18206 7498
rect 18258 7446 18270 7498
rect 18322 7446 18334 7498
rect 18386 7446 21620 7498
rect 1104 7424 21620 7446
rect 10318 7384 10324 7396
rect 10279 7356 10324 7384
rect 10318 7344 10324 7356
rect 10376 7344 10382 7396
rect 13630 7384 13636 7396
rect 13004 7356 13636 7384
rect 10594 7208 10600 7260
rect 10652 7248 10658 7260
rect 10873 7251 10931 7257
rect 10873 7248 10885 7251
rect 10652 7220 10885 7248
rect 10652 7208 10658 7220
rect 10873 7217 10885 7220
rect 10919 7217 10931 7251
rect 10873 7211 10931 7217
rect 10888 7112 10916 7211
rect 13004 7189 13032 7356
rect 13630 7344 13636 7356
rect 13688 7384 13694 7396
rect 16022 7384 16028 7396
rect 13688 7356 16028 7384
rect 13688 7344 13694 7356
rect 14642 7248 14648 7260
rect 14603 7220 14648 7248
rect 14642 7208 14648 7220
rect 14700 7208 14706 7260
rect 15120 7248 15148 7356
rect 16022 7344 16028 7356
rect 16080 7344 16086 7396
rect 16574 7344 16580 7396
rect 16632 7384 16638 7396
rect 16669 7387 16727 7393
rect 16669 7384 16681 7387
rect 16632 7356 16681 7384
rect 16632 7344 16638 7356
rect 16669 7353 16681 7356
rect 16715 7384 16727 7387
rect 17218 7384 17224 7396
rect 16715 7356 17224 7384
rect 16715 7353 16727 7356
rect 16669 7347 16727 7353
rect 17218 7344 17224 7356
rect 17276 7344 17282 7396
rect 15289 7251 15347 7257
rect 15289 7248 15301 7251
rect 15120 7220 15301 7248
rect 15289 7217 15301 7220
rect 15335 7217 15347 7251
rect 15289 7211 15347 7217
rect 11241 7183 11299 7189
rect 11241 7149 11253 7183
rect 11287 7180 11299 7183
rect 11333 7183 11391 7189
rect 11333 7180 11345 7183
rect 11287 7152 11345 7180
rect 11287 7149 11299 7152
rect 11241 7143 11299 7149
rect 11333 7149 11345 7152
rect 11379 7149 11391 7183
rect 11333 7143 11391 7149
rect 12989 7183 13047 7189
rect 12989 7149 13001 7183
rect 13035 7149 13047 7183
rect 13256 7183 13314 7189
rect 13256 7180 13268 7183
rect 12989 7143 13047 7149
rect 13188 7152 13268 7180
rect 11578 7115 11636 7121
rect 11578 7112 11590 7115
rect 10888 7084 11590 7112
rect 11578 7081 11590 7084
rect 11624 7081 11636 7115
rect 13004 7112 13032 7143
rect 11578 7075 11636 7081
rect 12360 7084 13032 7112
rect 9861 7047 9919 7053
rect 9861 7013 9873 7047
rect 9907 7044 9919 7047
rect 10689 7047 10747 7053
rect 10689 7044 10701 7047
rect 9907 7016 10701 7044
rect 9907 7013 9919 7016
rect 9861 7007 9919 7013
rect 10689 7013 10701 7016
rect 10735 7013 10747 7047
rect 10689 7007 10747 7013
rect 10778 7004 10784 7056
rect 10836 7044 10842 7056
rect 11241 7047 11299 7053
rect 10836 7016 10881 7044
rect 10836 7004 10842 7016
rect 11241 7013 11253 7047
rect 11287 7044 11299 7047
rect 12360 7044 12388 7084
rect 11287 7016 12388 7044
rect 12713 7047 12771 7053
rect 11287 7013 11299 7016
rect 11241 7007 11299 7013
rect 12713 7013 12725 7047
rect 12759 7044 12771 7047
rect 13188 7044 13216 7152
rect 13256 7149 13268 7152
rect 13302 7180 13314 7183
rect 14550 7180 14556 7192
rect 13302 7152 14556 7180
rect 13302 7149 13314 7152
rect 13256 7143 13314 7149
rect 14550 7140 14556 7152
rect 14608 7140 14614 7192
rect 14274 7072 14280 7124
rect 14332 7112 14338 7124
rect 15534 7115 15592 7121
rect 15534 7112 15546 7115
rect 14332 7084 15546 7112
rect 14332 7072 14338 7084
rect 14384 7053 14412 7084
rect 15534 7081 15546 7084
rect 15580 7081 15592 7115
rect 15534 7075 15592 7081
rect 12759 7016 13216 7044
rect 14369 7047 14427 7053
rect 12759 7013 12771 7016
rect 12713 7007 12771 7013
rect 14369 7013 14381 7047
rect 14415 7013 14427 7047
rect 14369 7007 14427 7013
rect 1104 6954 21620 6976
rect 1104 6902 7846 6954
rect 7898 6902 7910 6954
rect 7962 6902 7974 6954
rect 8026 6902 8038 6954
rect 8090 6902 14710 6954
rect 14762 6902 14774 6954
rect 14826 6902 14838 6954
rect 14890 6902 14902 6954
rect 14954 6902 21620 6954
rect 1104 6880 21620 6902
rect 10594 6840 10600 6852
rect 10555 6812 10600 6840
rect 10594 6800 10600 6812
rect 10652 6800 10658 6852
rect 10778 6800 10784 6852
rect 10836 6840 10842 6852
rect 10873 6843 10931 6849
rect 10873 6840 10885 6843
rect 10836 6812 10885 6840
rect 10836 6800 10842 6812
rect 10873 6809 10885 6812
rect 10919 6809 10931 6843
rect 10873 6803 10931 6809
rect 14001 6843 14059 6849
rect 14001 6809 14013 6843
rect 14047 6840 14059 6843
rect 14090 6840 14096 6852
rect 14047 6812 14096 6840
rect 14047 6809 14059 6812
rect 14001 6803 14059 6809
rect 14090 6800 14096 6812
rect 14148 6800 14154 6852
rect 16942 6840 16948 6852
rect 14292 6812 16948 6840
rect 11241 6775 11299 6781
rect 11241 6741 11253 6775
rect 11287 6772 11299 6775
rect 14292 6772 14320 6812
rect 16942 6800 16948 6812
rect 17000 6800 17006 6852
rect 17037 6843 17095 6849
rect 17037 6809 17049 6843
rect 17083 6840 17095 6843
rect 18506 6840 18512 6852
rect 17083 6812 18512 6840
rect 17083 6809 17095 6812
rect 17037 6803 17095 6809
rect 18506 6800 18512 6812
rect 18564 6800 18570 6852
rect 11287 6744 14320 6772
rect 14369 6775 14427 6781
rect 11287 6741 11299 6744
rect 11241 6735 11299 6741
rect 14369 6741 14381 6775
rect 14415 6772 14427 6775
rect 15194 6772 15200 6784
rect 14415 6744 15200 6772
rect 14415 6741 14427 6744
rect 14369 6735 14427 6741
rect 15194 6732 15200 6744
rect 15252 6732 15258 6784
rect 2958 6664 2964 6716
rect 3016 6704 3022 6716
rect 7541 6707 7599 6713
rect 7541 6704 7553 6707
rect 3016 6676 7553 6704
rect 3016 6664 3022 6676
rect 7541 6673 7553 6676
rect 7587 6673 7599 6707
rect 9484 6707 9542 6713
rect 9484 6704 9496 6707
rect 7541 6667 7599 6673
rect 8680 6676 9496 6704
rect 7285 6639 7343 6645
rect 7285 6605 7297 6639
rect 7331 6605 7343 6639
rect 7285 6599 7343 6605
rect 7300 6500 7328 6599
rect 8680 6577 8708 6676
rect 9484 6673 9496 6676
rect 9530 6704 9542 6707
rect 9530 6676 11468 6704
rect 9530 6673 9542 6676
rect 9484 6667 9542 6673
rect 11440 6645 11468 6676
rect 11698 6664 11704 6716
rect 11756 6704 11762 6716
rect 14461 6707 14519 6713
rect 14461 6704 14473 6707
rect 11756 6676 14473 6704
rect 11756 6664 11762 6676
rect 14461 6673 14473 6676
rect 14507 6704 14519 6707
rect 17129 6707 17187 6713
rect 14507 6676 15792 6704
rect 14507 6673 14519 6676
rect 14461 6667 14519 6673
rect 9217 6639 9275 6645
rect 9217 6605 9229 6639
rect 9263 6605 9275 6639
rect 9217 6599 9275 6605
rect 11333 6639 11391 6645
rect 11333 6605 11345 6639
rect 11379 6605 11391 6639
rect 11333 6599 11391 6605
rect 11425 6639 11483 6645
rect 11425 6605 11437 6639
rect 11471 6605 11483 6639
rect 14550 6636 14556 6648
rect 14511 6608 14556 6636
rect 11425 6599 11483 6605
rect 8665 6571 8723 6577
rect 8665 6537 8677 6571
rect 8711 6537 8723 6571
rect 8665 6531 8723 6537
rect 7558 6500 7564 6512
rect 7300 6472 7564 6500
rect 7558 6460 7564 6472
rect 7616 6500 7622 6512
rect 9232 6500 9260 6599
rect 11348 6568 11376 6599
rect 14550 6596 14556 6608
rect 14608 6596 14614 6648
rect 15764 6636 15792 6676
rect 17129 6673 17141 6707
rect 17175 6704 17187 6707
rect 19058 6704 19064 6716
rect 17175 6676 19064 6704
rect 17175 6673 17187 6676
rect 17129 6667 17187 6673
rect 17144 6636 17172 6667
rect 19058 6664 19064 6676
rect 19116 6664 19122 6716
rect 20530 6704 20536 6716
rect 20491 6676 20536 6704
rect 20530 6664 20536 6676
rect 20588 6664 20594 6716
rect 15764 6608 17172 6636
rect 17218 6596 17224 6648
rect 17276 6636 17282 6648
rect 17276 6608 17321 6636
rect 17276 6596 17282 6608
rect 11698 6568 11704 6580
rect 11348 6540 11704 6568
rect 11698 6528 11704 6540
rect 11756 6528 11762 6580
rect 16666 6568 16672 6580
rect 16627 6540 16672 6568
rect 16666 6528 16672 6540
rect 16724 6528 16730 6580
rect 18598 6528 18604 6580
rect 18656 6568 18662 6580
rect 19058 6568 19064 6580
rect 18656 6540 19064 6568
rect 18656 6528 18662 6540
rect 19058 6528 19064 6540
rect 19116 6528 19122 6580
rect 7616 6472 9260 6500
rect 7616 6460 7622 6472
rect 13722 6460 13728 6512
rect 13780 6500 13786 6512
rect 20717 6503 20775 6509
rect 20717 6500 20729 6503
rect 13780 6472 20729 6500
rect 13780 6460 13786 6472
rect 20717 6469 20729 6472
rect 20763 6469 20775 6503
rect 20717 6463 20775 6469
rect 1104 6410 21620 6432
rect 1104 6358 4414 6410
rect 4466 6358 4478 6410
rect 4530 6358 4542 6410
rect 4594 6358 4606 6410
rect 4658 6358 11278 6410
rect 11330 6358 11342 6410
rect 11394 6358 11406 6410
rect 11458 6358 11470 6410
rect 11522 6358 18142 6410
rect 18194 6358 18206 6410
rect 18258 6358 18270 6410
rect 18322 6358 18334 6410
rect 18386 6358 21620 6410
rect 1104 6336 21620 6358
rect 15194 6256 15200 6308
rect 15252 6296 15258 6308
rect 17954 6296 17960 6308
rect 15252 6268 17960 6296
rect 15252 6256 15258 6268
rect 17954 6256 17960 6268
rect 18012 6256 18018 6308
rect 1104 5866 21620 5888
rect 1104 5814 7846 5866
rect 7898 5814 7910 5866
rect 7962 5814 7974 5866
rect 8026 5814 8038 5866
rect 8090 5814 14710 5866
rect 14762 5814 14774 5866
rect 14826 5814 14838 5866
rect 14890 5814 14902 5866
rect 14954 5814 21620 5866
rect 1104 5792 21620 5814
rect 12526 5712 12532 5764
rect 12584 5752 12590 5764
rect 20717 5755 20775 5761
rect 20717 5752 20729 5755
rect 12584 5724 20729 5752
rect 12584 5712 12590 5724
rect 20717 5721 20729 5724
rect 20763 5721 20775 5755
rect 20717 5715 20775 5721
rect 20530 5616 20536 5628
rect 20491 5588 20536 5616
rect 20530 5576 20536 5588
rect 20588 5576 20594 5628
rect 1104 5322 21620 5344
rect 1104 5270 4414 5322
rect 4466 5270 4478 5322
rect 4530 5270 4542 5322
rect 4594 5270 4606 5322
rect 4658 5270 11278 5322
rect 11330 5270 11342 5322
rect 11394 5270 11406 5322
rect 11458 5270 11470 5322
rect 11522 5270 18142 5322
rect 18194 5270 18206 5322
rect 18258 5270 18270 5322
rect 18322 5270 18334 5322
rect 18386 5270 21620 5322
rect 1104 5248 21620 5270
rect 16942 5168 16948 5220
rect 17000 5208 17006 5220
rect 17954 5208 17960 5220
rect 17000 5180 17960 5208
rect 17000 5168 17006 5180
rect 17954 5168 17960 5180
rect 18012 5168 18018 5220
rect 1104 4778 21620 4800
rect 1104 4726 7846 4778
rect 7898 4726 7910 4778
rect 7962 4726 7974 4778
rect 8026 4726 8038 4778
rect 8090 4726 14710 4778
rect 14762 4726 14774 4778
rect 14826 4726 14838 4778
rect 14890 4726 14902 4778
rect 14954 4726 21620 4778
rect 1104 4704 21620 4726
rect 20717 4667 20775 4673
rect 20717 4633 20729 4667
rect 20763 4664 20775 4667
rect 21082 4664 21088 4676
rect 20763 4636 21088 4664
rect 20763 4633 20775 4636
rect 20717 4627 20775 4633
rect 21082 4624 21088 4636
rect 21140 4624 21146 4676
rect 20530 4528 20536 4540
rect 20491 4500 20536 4528
rect 20530 4488 20536 4500
rect 20588 4488 20594 4540
rect 1104 4234 21620 4256
rect 1104 4182 4414 4234
rect 4466 4182 4478 4234
rect 4530 4182 4542 4234
rect 4594 4182 4606 4234
rect 4658 4182 11278 4234
rect 11330 4182 11342 4234
rect 11394 4182 11406 4234
rect 11458 4182 11470 4234
rect 11522 4182 18142 4234
rect 18194 4182 18206 4234
rect 18258 4182 18270 4234
rect 18322 4182 18334 4234
rect 18386 4182 21620 4234
rect 1104 4160 21620 4182
rect 14182 3944 14188 3996
rect 14240 3984 14246 3996
rect 18506 3984 18512 3996
rect 14240 3956 18512 3984
rect 14240 3944 14246 3956
rect 18506 3944 18512 3956
rect 18564 3944 18570 3996
rect 15930 3876 15936 3928
rect 15988 3916 15994 3928
rect 19242 3916 19248 3928
rect 15988 3888 19248 3916
rect 15988 3876 15994 3888
rect 19242 3876 19248 3888
rect 19300 3876 19306 3928
rect 1104 3690 21620 3712
rect 1104 3638 7846 3690
rect 7898 3638 7910 3690
rect 7962 3638 7974 3690
rect 8026 3638 8038 3690
rect 8090 3638 14710 3690
rect 14762 3638 14774 3690
rect 14826 3638 14838 3690
rect 14890 3638 14902 3690
rect 14954 3638 21620 3690
rect 1104 3616 21620 3638
rect 1104 3146 21620 3168
rect 1104 3094 4414 3146
rect 4466 3094 4478 3146
rect 4530 3094 4542 3146
rect 4594 3094 4606 3146
rect 4658 3094 11278 3146
rect 11330 3094 11342 3146
rect 11394 3094 11406 3146
rect 11458 3094 11470 3146
rect 11522 3094 18142 3146
rect 18194 3094 18206 3146
rect 18258 3094 18270 3146
rect 18322 3094 18334 3146
rect 18386 3094 21620 3146
rect 1104 3072 21620 3094
rect 1104 2602 21620 2624
rect 1104 2550 7846 2602
rect 7898 2550 7910 2602
rect 7962 2550 7974 2602
rect 8026 2550 8038 2602
rect 8090 2550 14710 2602
rect 14762 2550 14774 2602
rect 14826 2550 14838 2602
rect 14890 2550 14902 2602
rect 14954 2550 21620 2602
rect 1104 2528 21620 2550
rect 16850 2244 16856 2296
rect 16908 2284 16914 2296
rect 19242 2284 19248 2296
rect 16908 2256 19248 2284
rect 16908 2244 16914 2256
rect 19242 2244 19248 2256
rect 19300 2244 19306 2296
rect 1104 2058 21620 2080
rect 1104 2006 4414 2058
rect 4466 2006 4478 2058
rect 4530 2006 4542 2058
rect 4594 2006 4606 2058
rect 4658 2006 11278 2058
rect 11330 2006 11342 2058
rect 11394 2006 11406 2058
rect 11458 2006 11470 2058
rect 11522 2006 18142 2058
rect 18194 2006 18206 2058
rect 18258 2006 18270 2058
rect 18322 2006 18334 2058
rect 18386 2006 21620 2058
rect 1104 1984 21620 2006
rect 16390 1156 16396 1208
rect 16448 1196 16454 1208
rect 17954 1196 17960 1208
rect 16448 1168 17960 1196
rect 16448 1156 16454 1168
rect 17954 1156 17960 1168
rect 18012 1156 18018 1208
<< via1 >>
rect 7846 19958 7898 20010
rect 7910 19958 7962 20010
rect 7974 19958 8026 20010
rect 8038 19958 8090 20010
rect 14710 19958 14762 20010
rect 14774 19958 14826 20010
rect 14838 19958 14890 20010
rect 14902 19958 14954 20010
rect 20168 19899 20220 19908
rect 20168 19865 20177 19899
rect 20177 19865 20211 19899
rect 20211 19865 20220 19899
rect 20168 19856 20220 19865
rect 20628 19856 20680 19908
rect 19984 19763 20036 19772
rect 19984 19729 19993 19763
rect 19993 19729 20027 19763
rect 20027 19729 20036 19763
rect 19984 19720 20036 19729
rect 20444 19720 20496 19772
rect 4414 19414 4466 19466
rect 4478 19414 4530 19466
rect 4542 19414 4594 19466
rect 4606 19414 4658 19466
rect 11278 19414 11330 19466
rect 11342 19414 11394 19466
rect 11406 19414 11458 19466
rect 11470 19414 11522 19466
rect 18142 19414 18194 19466
rect 18206 19414 18258 19466
rect 18270 19414 18322 19466
rect 18334 19414 18386 19466
rect 20536 19312 20588 19364
rect 5172 19176 5224 19228
rect 8208 19176 8260 19228
rect 10232 19219 10284 19228
rect 10232 19185 10241 19219
rect 10241 19185 10275 19219
rect 10275 19185 10284 19219
rect 10232 19176 10284 19185
rect 4896 18972 4948 19024
rect 5080 19015 5132 19024
rect 5080 18981 5089 19015
rect 5089 18981 5123 19015
rect 5123 18981 5132 19015
rect 5080 18972 5132 18981
rect 5448 18972 5500 19024
rect 9128 19108 9180 19160
rect 11244 19151 11296 19160
rect 11244 19117 11253 19151
rect 11253 19117 11287 19151
rect 11287 19117 11296 19151
rect 11244 19108 11296 19117
rect 14280 19219 14332 19228
rect 14280 19185 14289 19219
rect 14289 19185 14323 19219
rect 14323 19185 14332 19219
rect 14280 19176 14332 19185
rect 16120 19176 16172 19228
rect 17316 19176 17368 19228
rect 19984 19176 20036 19228
rect 17408 19151 17460 19160
rect 11520 19083 11572 19092
rect 11520 19049 11554 19083
rect 11554 19049 11572 19083
rect 11520 19040 11572 19049
rect 15016 19040 15068 19092
rect 8300 18972 8352 19024
rect 9680 19015 9732 19024
rect 9680 18981 9689 19015
rect 9689 18981 9723 19015
rect 9723 18981 9732 19015
rect 9680 18972 9732 18981
rect 9956 18972 10008 19024
rect 11152 18972 11204 19024
rect 12624 19015 12676 19024
rect 12624 18981 12633 19015
rect 12633 18981 12667 19015
rect 12667 18981 12676 19015
rect 12624 18972 12676 18981
rect 13912 18972 13964 19024
rect 14096 19015 14148 19024
rect 14096 18981 14105 19015
rect 14105 18981 14139 19015
rect 14139 18981 14148 19015
rect 17408 19117 17417 19151
rect 17417 19117 17451 19151
rect 17451 19117 17460 19151
rect 17408 19108 17460 19117
rect 17960 19151 18012 19160
rect 17960 19117 17969 19151
rect 17969 19117 18003 19151
rect 18003 19117 18012 19151
rect 17960 19108 18012 19117
rect 20260 19151 20312 19160
rect 20260 19117 20269 19151
rect 20269 19117 20303 19151
rect 20303 19117 20312 19151
rect 20260 19108 20312 19117
rect 18788 19083 18840 19092
rect 18788 19049 18797 19083
rect 18797 19049 18831 19083
rect 18831 19049 18840 19083
rect 18788 19040 18840 19049
rect 14096 18972 14148 18981
rect 15660 19015 15712 19024
rect 15660 18981 15669 19015
rect 15669 18981 15703 19015
rect 15703 18981 15712 19015
rect 15660 18972 15712 18981
rect 15752 19015 15804 19024
rect 15752 18981 15761 19015
rect 15761 18981 15795 19015
rect 15795 18981 15804 19015
rect 16304 19015 16356 19024
rect 15752 18972 15804 18981
rect 16304 18981 16313 19015
rect 16313 18981 16347 19015
rect 16347 18981 16356 19015
rect 16304 18972 16356 18981
rect 16672 19015 16724 19024
rect 16672 18981 16681 19015
rect 16681 18981 16715 19015
rect 16715 18981 16724 19015
rect 16672 18972 16724 18981
rect 17868 18972 17920 19024
rect 7846 18870 7898 18922
rect 7910 18870 7962 18922
rect 7974 18870 8026 18922
rect 8038 18870 8090 18922
rect 14710 18870 14762 18922
rect 14774 18870 14826 18922
rect 14838 18870 14890 18922
rect 14902 18870 14954 18922
rect 5448 18811 5500 18820
rect 5448 18777 5457 18811
rect 5457 18777 5491 18811
rect 5491 18777 5500 18811
rect 5448 18768 5500 18777
rect 9956 18768 10008 18820
rect 10140 18768 10192 18820
rect 11520 18811 11572 18820
rect 2780 18632 2832 18684
rect 1492 18428 1544 18480
rect 4988 18632 5040 18684
rect 4804 18564 4856 18616
rect 6552 18632 6604 18684
rect 7104 18675 7156 18684
rect 7104 18641 7138 18675
rect 7138 18641 7156 18675
rect 8208 18700 8260 18752
rect 8484 18675 8536 18684
rect 7104 18632 7156 18641
rect 8484 18641 8493 18675
rect 8493 18641 8527 18675
rect 8527 18641 8536 18675
rect 8484 18632 8536 18641
rect 10232 18632 10284 18684
rect 11520 18777 11529 18811
rect 11529 18777 11563 18811
rect 11563 18777 11572 18811
rect 11520 18768 11572 18777
rect 11612 18768 11664 18820
rect 12256 18768 12308 18820
rect 12624 18700 12676 18752
rect 15016 18768 15068 18820
rect 14280 18700 14332 18752
rect 16120 18700 16172 18752
rect 16672 18768 16724 18820
rect 19248 18768 19300 18820
rect 20352 18768 20404 18820
rect 15752 18632 15804 18684
rect 15844 18632 15896 18684
rect 19340 18632 19392 18684
rect 20260 18700 20312 18752
rect 20444 18743 20496 18752
rect 20444 18709 20453 18743
rect 20453 18709 20487 18743
rect 20487 18709 20496 18743
rect 20444 18700 20496 18709
rect 19524 18632 19576 18684
rect 11796 18607 11848 18616
rect 8208 18539 8260 18548
rect 8208 18505 8217 18539
rect 8217 18505 8251 18539
rect 8251 18505 8260 18539
rect 8208 18496 8260 18505
rect 11796 18573 11805 18607
rect 11805 18573 11839 18607
rect 11839 18573 11848 18607
rect 11796 18564 11848 18573
rect 11244 18496 11296 18548
rect 5172 18471 5224 18480
rect 5172 18437 5181 18471
rect 5181 18437 5215 18471
rect 5215 18437 5224 18471
rect 5172 18428 5224 18437
rect 7012 18428 7064 18480
rect 12348 18428 12400 18480
rect 13268 18428 13320 18480
rect 16120 18428 16172 18480
rect 17316 18471 17368 18480
rect 17316 18437 17325 18471
rect 17325 18437 17359 18471
rect 17359 18437 17368 18471
rect 17316 18428 17368 18437
rect 17500 18428 17552 18480
rect 20996 18428 21048 18480
rect 4414 18326 4466 18378
rect 4478 18326 4530 18378
rect 4542 18326 4594 18378
rect 4606 18326 4658 18378
rect 11278 18326 11330 18378
rect 11342 18326 11394 18378
rect 11406 18326 11458 18378
rect 11470 18326 11522 18378
rect 18142 18326 18194 18378
rect 18206 18326 18258 18378
rect 18270 18326 18322 18378
rect 18334 18326 18386 18378
rect 4988 18224 5040 18276
rect 2780 18088 2832 18140
rect 5080 18131 5132 18140
rect 5080 18097 5089 18131
rect 5089 18097 5123 18131
rect 5123 18097 5132 18131
rect 5080 18088 5132 18097
rect 296 18020 348 18072
rect 7104 18224 7156 18276
rect 8300 18224 8352 18276
rect 8116 18156 8168 18208
rect 11704 18224 11756 18276
rect 14096 18224 14148 18276
rect 18696 18267 18748 18276
rect 18696 18233 18705 18267
rect 18705 18233 18739 18267
rect 18739 18233 18748 18267
rect 18696 18224 18748 18233
rect 19616 18267 19668 18276
rect 19616 18233 19625 18267
rect 19625 18233 19659 18267
rect 19659 18233 19668 18267
rect 19616 18224 19668 18233
rect 20168 18267 20220 18276
rect 20168 18233 20177 18267
rect 20177 18233 20211 18267
rect 20211 18233 20220 18267
rect 20168 18224 20220 18233
rect 9772 18156 9824 18208
rect 9680 18088 9732 18140
rect 11612 18088 11664 18140
rect 3056 17952 3108 18004
rect 1400 17884 1452 17936
rect 2688 17884 2740 17936
rect 2964 17884 3016 17936
rect 3148 17927 3200 17936
rect 3148 17893 3157 17927
rect 3157 17893 3191 17927
rect 3191 17893 3200 17927
rect 3148 17884 3200 17893
rect 3240 17927 3292 17936
rect 3240 17893 3249 17927
rect 3249 17893 3283 17927
rect 3283 17893 3292 17927
rect 3240 17884 3292 17893
rect 5448 17884 5500 17936
rect 6552 18020 6604 18072
rect 7656 18020 7708 18072
rect 8576 18020 8628 18072
rect 6368 17952 6420 18004
rect 6460 17952 6512 18004
rect 11060 18020 11112 18072
rect 11796 18020 11848 18072
rect 12716 18156 12768 18208
rect 17224 18156 17276 18208
rect 18512 18156 18564 18208
rect 19340 18156 19392 18208
rect 12624 18088 12676 18140
rect 13912 18131 13964 18140
rect 13912 18097 13921 18131
rect 13921 18097 13955 18131
rect 13955 18097 13964 18131
rect 13912 18088 13964 18097
rect 17408 18131 17460 18140
rect 17408 18097 17417 18131
rect 17417 18097 17451 18131
rect 17451 18097 17460 18131
rect 17408 18088 17460 18097
rect 19616 18088 19668 18140
rect 21364 18088 21416 18140
rect 16304 18020 16356 18072
rect 18512 18063 18564 18072
rect 18512 18029 18521 18063
rect 18521 18029 18555 18063
rect 18555 18029 18564 18063
rect 18512 18020 18564 18029
rect 19432 18063 19484 18072
rect 19432 18029 19441 18063
rect 19441 18029 19475 18063
rect 19475 18029 19484 18063
rect 19432 18020 19484 18029
rect 19984 18063 20036 18072
rect 19984 18029 19993 18063
rect 19993 18029 20027 18063
rect 20027 18029 20036 18063
rect 19984 18020 20036 18029
rect 10784 17884 10836 17936
rect 19524 17952 19576 18004
rect 21088 17952 21140 18004
rect 22468 17952 22520 18004
rect 10968 17884 11020 17936
rect 14188 17884 14240 17936
rect 15108 17884 15160 17936
rect 15292 17884 15344 17936
rect 16212 17884 16264 17936
rect 16948 17884 17000 17936
rect 19800 17884 19852 17936
rect 20536 17884 20588 17936
rect 21916 17884 21968 17936
rect 20 17816 72 17868
rect 848 17816 900 17868
rect 7846 17782 7898 17834
rect 7910 17782 7962 17834
rect 7974 17782 8026 17834
rect 8038 17782 8090 17834
rect 14710 17782 14762 17834
rect 14774 17782 14826 17834
rect 14838 17782 14890 17834
rect 14902 17782 14954 17834
rect 2780 17723 2832 17732
rect 2780 17689 2789 17723
rect 2789 17689 2823 17723
rect 2823 17689 2832 17723
rect 2780 17680 2832 17689
rect 3240 17680 3292 17732
rect 4160 17680 4212 17732
rect 4712 17680 4764 17732
rect 20168 17680 20220 17732
rect 7656 17612 7708 17664
rect 18512 17612 18564 17664
rect 1492 17544 1544 17596
rect 3424 17544 3476 17596
rect 12348 17544 12400 17596
rect 12716 17544 12768 17596
rect 17960 17544 18012 17596
rect 4896 17476 4948 17528
rect 7564 17408 7616 17460
rect 19432 17408 19484 17460
rect 10876 17340 10928 17392
rect 16672 17340 16724 17392
rect 20720 17383 20772 17392
rect 20720 17349 20729 17383
rect 20729 17349 20763 17383
rect 20763 17349 20772 17383
rect 20720 17340 20772 17349
rect 4414 17238 4466 17290
rect 4478 17238 4530 17290
rect 4542 17238 4594 17290
rect 4606 17238 4658 17290
rect 11278 17238 11330 17290
rect 11342 17238 11394 17290
rect 11406 17238 11458 17290
rect 11470 17238 11522 17290
rect 18142 17238 18194 17290
rect 18206 17238 18258 17290
rect 18270 17238 18322 17290
rect 18334 17238 18386 17290
rect 4068 17136 4120 17188
rect 17684 17136 17736 17188
rect 18696 17179 18748 17188
rect 18696 17145 18705 17179
rect 18705 17145 18739 17179
rect 18739 17145 18748 17179
rect 18696 17136 18748 17145
rect 20444 17179 20496 17188
rect 20444 17145 20453 17179
rect 20453 17145 20487 17179
rect 20487 17145 20496 17179
rect 20444 17136 20496 17145
rect 3148 17043 3200 17052
rect 3148 17009 3157 17043
rect 3157 17009 3191 17043
rect 3191 17009 3200 17043
rect 3148 17000 3200 17009
rect 4712 17000 4764 17052
rect 7564 17043 7616 17052
rect 7564 17009 7573 17043
rect 7573 17009 7607 17043
rect 7607 17009 7616 17043
rect 7564 17000 7616 17009
rect 8760 17000 8812 17052
rect 19984 17000 20036 17052
rect 2964 16932 3016 16984
rect 4896 16932 4948 16984
rect 6828 16932 6880 16984
rect 11060 16932 11112 16984
rect 13360 16932 13412 16984
rect 15476 16932 15528 16984
rect 18512 16975 18564 16984
rect 18512 16941 18521 16975
rect 18521 16941 18555 16975
rect 18555 16941 18564 16975
rect 18512 16932 18564 16941
rect 19064 16975 19116 16984
rect 19064 16941 19073 16975
rect 19073 16941 19107 16975
rect 19107 16941 19116 16975
rect 19064 16932 19116 16941
rect 19524 16932 19576 16984
rect 5172 16864 5224 16916
rect 5540 16864 5592 16916
rect 10968 16864 11020 16916
rect 11704 16864 11756 16916
rect 15660 16864 15712 16916
rect 16856 16864 16908 16916
rect 8300 16839 8352 16848
rect 8300 16805 8309 16839
rect 8309 16805 8343 16839
rect 8343 16805 8352 16839
rect 8300 16796 8352 16805
rect 9680 16796 9732 16848
rect 10508 16796 10560 16848
rect 12440 16796 12492 16848
rect 19984 16864 20036 16916
rect 7846 16694 7898 16746
rect 7910 16694 7962 16746
rect 7974 16694 8026 16746
rect 8038 16694 8090 16746
rect 14710 16694 14762 16746
rect 14774 16694 14826 16746
rect 14838 16694 14890 16746
rect 14902 16694 14954 16746
rect 6828 16635 6880 16644
rect 6828 16601 6837 16635
rect 6837 16601 6871 16635
rect 6871 16601 6880 16635
rect 6828 16592 6880 16601
rect 10508 16635 10560 16644
rect 10508 16601 10517 16635
rect 10517 16601 10551 16635
rect 10551 16601 10560 16635
rect 10508 16592 10560 16601
rect 11704 16635 11756 16644
rect 8300 16524 8352 16576
rect 11704 16601 11713 16635
rect 11713 16601 11747 16635
rect 11747 16601 11756 16635
rect 11704 16592 11756 16601
rect 13360 16592 13412 16644
rect 16856 16635 16908 16644
rect 16856 16601 16865 16635
rect 16865 16601 16899 16635
rect 16899 16601 16908 16635
rect 16856 16592 16908 16601
rect 18512 16592 18564 16644
rect 19524 16567 19576 16576
rect 8484 16499 8536 16508
rect 8484 16465 8493 16499
rect 8493 16465 8527 16499
rect 8527 16465 8536 16499
rect 8484 16456 8536 16465
rect 8760 16499 8812 16508
rect 8760 16465 8794 16499
rect 8794 16465 8812 16499
rect 8760 16456 8812 16465
rect 7288 16431 7340 16440
rect 7288 16397 7297 16431
rect 7297 16397 7331 16431
rect 7331 16397 7340 16431
rect 7288 16388 7340 16397
rect 11796 16431 11848 16440
rect 6368 16320 6420 16372
rect 11796 16397 11805 16431
rect 11805 16397 11839 16431
rect 11839 16397 11848 16431
rect 11796 16388 11848 16397
rect 11888 16431 11940 16440
rect 11888 16397 11897 16431
rect 11897 16397 11931 16431
rect 11931 16397 11940 16431
rect 12992 16431 13044 16440
rect 11888 16388 11940 16397
rect 12992 16397 13001 16431
rect 13001 16397 13035 16431
rect 13035 16397 13044 16431
rect 12992 16388 13044 16397
rect 12440 16363 12492 16372
rect 12440 16329 12449 16363
rect 12449 16329 12483 16363
rect 12483 16329 12492 16363
rect 12440 16320 12492 16329
rect 2504 16252 2556 16304
rect 8852 16252 8904 16304
rect 10048 16252 10100 16304
rect 14280 16499 14332 16508
rect 14280 16465 14289 16499
rect 14289 16465 14323 16499
rect 14323 16465 14332 16499
rect 14280 16456 14332 16465
rect 17316 16456 17368 16508
rect 19524 16533 19533 16567
rect 19533 16533 19567 16567
rect 19567 16533 19576 16567
rect 19524 16524 19576 16533
rect 20628 16592 20680 16644
rect 19984 16499 20036 16508
rect 19984 16465 19993 16499
rect 19993 16465 20027 16499
rect 20027 16465 20036 16499
rect 19984 16456 20036 16465
rect 20168 16456 20220 16508
rect 14464 16431 14516 16440
rect 14464 16397 14473 16431
rect 14473 16397 14507 16431
rect 14507 16397 14516 16431
rect 15476 16431 15528 16440
rect 14464 16388 14516 16397
rect 15476 16397 15485 16431
rect 15485 16397 15519 16431
rect 15519 16397 15528 16431
rect 15476 16388 15528 16397
rect 17960 16388 18012 16440
rect 13912 16295 13964 16304
rect 13912 16261 13921 16295
rect 13921 16261 13955 16295
rect 13955 16261 13964 16295
rect 13912 16252 13964 16261
rect 4414 16150 4466 16202
rect 4478 16150 4530 16202
rect 4542 16150 4594 16202
rect 4606 16150 4658 16202
rect 11278 16150 11330 16202
rect 11342 16150 11394 16202
rect 11406 16150 11458 16202
rect 11470 16150 11522 16202
rect 18142 16150 18194 16202
rect 18206 16150 18258 16202
rect 18270 16150 18322 16202
rect 18334 16150 18386 16202
rect 3424 16048 3476 16100
rect 6368 16091 6420 16100
rect 6368 16057 6377 16091
rect 6377 16057 6411 16091
rect 6411 16057 6420 16091
rect 6368 16048 6420 16057
rect 7288 16048 7340 16100
rect 12992 16091 13044 16100
rect 12992 16057 13001 16091
rect 13001 16057 13035 16091
rect 13035 16057 13044 16091
rect 12992 16048 13044 16057
rect 17868 16048 17920 16100
rect 19248 16048 19300 16100
rect 1492 15912 1544 15964
rect 4988 15955 5040 15964
rect 4988 15921 4997 15955
rect 4997 15921 5031 15955
rect 5031 15921 5040 15955
rect 4988 15912 5040 15921
rect 6368 15912 6420 15964
rect 8484 15912 8536 15964
rect 7380 15887 7432 15896
rect 7380 15853 7389 15887
rect 7389 15853 7423 15887
rect 7423 15853 7432 15887
rect 7380 15844 7432 15853
rect 7748 15844 7800 15896
rect 10048 15844 10100 15896
rect 10692 15844 10744 15896
rect 11888 15887 11940 15896
rect 2872 15776 2924 15828
rect 7564 15776 7616 15828
rect 11520 15776 11572 15828
rect 11888 15853 11922 15887
rect 11922 15853 11940 15887
rect 11888 15844 11940 15853
rect 13268 15887 13320 15896
rect 13268 15853 13277 15887
rect 13277 15853 13311 15887
rect 13311 15853 13320 15887
rect 13268 15844 13320 15853
rect 16856 15912 16908 15964
rect 19156 15980 19208 16032
rect 17684 15844 17736 15896
rect 19708 15887 19760 15896
rect 19708 15853 19717 15887
rect 19717 15853 19751 15887
rect 19751 15853 19760 15887
rect 19708 15844 19760 15853
rect 20260 15887 20312 15896
rect 20260 15853 20269 15887
rect 20269 15853 20303 15887
rect 20303 15853 20312 15887
rect 20260 15844 20312 15853
rect 14280 15776 14332 15828
rect 17960 15776 18012 15828
rect 14464 15708 14516 15760
rect 15292 15751 15344 15760
rect 15292 15717 15301 15751
rect 15301 15717 15335 15751
rect 15335 15717 15344 15751
rect 15292 15708 15344 15717
rect 16672 15708 16724 15760
rect 7846 15606 7898 15658
rect 7910 15606 7962 15658
rect 7974 15606 8026 15658
rect 8038 15606 8090 15658
rect 14710 15606 14762 15658
rect 14774 15606 14826 15658
rect 14838 15606 14890 15658
rect 14902 15606 14954 15658
rect 3608 15504 3660 15556
rect 15292 15504 15344 15556
rect 20168 15547 20220 15556
rect 20168 15513 20177 15547
rect 20177 15513 20211 15547
rect 20211 15513 20220 15547
rect 20168 15504 20220 15513
rect 20720 15547 20772 15556
rect 20720 15513 20729 15547
rect 20729 15513 20763 15547
rect 20763 15513 20772 15547
rect 20720 15504 20772 15513
rect 7380 15436 7432 15488
rect 7564 15436 7616 15488
rect 13912 15436 13964 15488
rect 3332 15368 3384 15420
rect 2872 15343 2924 15352
rect 2872 15309 2881 15343
rect 2881 15309 2915 15343
rect 2915 15309 2924 15343
rect 2872 15300 2924 15309
rect 3424 15300 3476 15352
rect 20168 15368 20220 15420
rect 15016 15343 15068 15352
rect 15016 15309 15025 15343
rect 15025 15309 15059 15343
rect 15059 15309 15068 15343
rect 15016 15300 15068 15309
rect 19064 15232 19116 15284
rect 4414 15062 4466 15114
rect 4478 15062 4530 15114
rect 4542 15062 4594 15114
rect 4606 15062 4658 15114
rect 11278 15062 11330 15114
rect 11342 15062 11394 15114
rect 11406 15062 11458 15114
rect 11470 15062 11522 15114
rect 18142 15062 18194 15114
rect 18206 15062 18258 15114
rect 18270 15062 18322 15114
rect 18334 15062 18386 15114
rect 2872 15003 2924 15012
rect 2872 14969 2881 15003
rect 2881 14969 2915 15003
rect 2915 14969 2924 15003
rect 2872 14960 2924 14969
rect 4988 14960 5040 15012
rect 6368 15003 6420 15012
rect 1492 14867 1544 14876
rect 1492 14833 1501 14867
rect 1501 14833 1535 14867
rect 1535 14833 1544 14867
rect 1492 14824 1544 14833
rect 3332 14867 3384 14876
rect 3332 14833 3341 14867
rect 3341 14833 3375 14867
rect 3375 14833 3384 14867
rect 3332 14824 3384 14833
rect 6368 14969 6377 15003
rect 6377 14969 6411 15003
rect 6411 14969 6420 15003
rect 6368 14960 6420 14969
rect 7472 14960 7524 15012
rect 8116 14824 8168 14876
rect 7656 14756 7708 14808
rect 8392 14960 8444 15012
rect 10692 14892 10744 14944
rect 13268 14892 13320 14944
rect 8668 14824 8720 14876
rect 9772 14824 9824 14876
rect 12440 14756 12492 14808
rect 14556 14756 14608 14808
rect 15476 14799 15528 14808
rect 15476 14765 15485 14799
rect 15485 14765 15519 14799
rect 15519 14765 15528 14799
rect 15476 14756 15528 14765
rect 19708 14824 19760 14876
rect 3424 14688 3476 14740
rect 9496 14688 9548 14740
rect 9404 14620 9456 14672
rect 10140 14620 10192 14672
rect 20260 14688 20312 14740
rect 16488 14620 16540 14672
rect 17500 14663 17552 14672
rect 17500 14629 17509 14663
rect 17509 14629 17543 14663
rect 17543 14629 17552 14663
rect 17500 14620 17552 14629
rect 17592 14663 17644 14672
rect 17592 14629 17601 14663
rect 17601 14629 17635 14663
rect 17635 14629 17644 14663
rect 17592 14620 17644 14629
rect 7846 14518 7898 14570
rect 7910 14518 7962 14570
rect 7974 14518 8026 14570
rect 8038 14518 8090 14570
rect 14710 14518 14762 14570
rect 14774 14518 14826 14570
rect 14838 14518 14890 14570
rect 14902 14518 14954 14570
rect 9496 14459 9548 14468
rect 9496 14425 9505 14459
rect 9505 14425 9539 14459
rect 9539 14425 9548 14459
rect 9496 14416 9548 14425
rect 9772 14459 9824 14468
rect 9772 14425 9781 14459
rect 9781 14425 9815 14459
rect 9815 14425 9824 14459
rect 9772 14416 9824 14425
rect 10140 14459 10192 14468
rect 10140 14425 10149 14459
rect 10149 14425 10183 14459
rect 10183 14425 10192 14459
rect 10140 14416 10192 14425
rect 13268 14416 13320 14468
rect 14556 14416 14608 14468
rect 4988 14280 5040 14332
rect 5632 14323 5684 14332
rect 5632 14289 5641 14323
rect 5641 14289 5675 14323
rect 5675 14289 5684 14323
rect 5632 14280 5684 14289
rect 8300 14348 8352 14400
rect 9404 14348 9456 14400
rect 15016 14416 15068 14468
rect 16488 14459 16540 14468
rect 16488 14425 16497 14459
rect 16497 14425 16531 14459
rect 16531 14425 16540 14459
rect 16488 14416 16540 14425
rect 17592 14416 17644 14468
rect 20720 14459 20772 14468
rect 20720 14425 20729 14459
rect 20729 14425 20763 14459
rect 20763 14425 20772 14459
rect 20720 14416 20772 14425
rect 8668 14280 8720 14332
rect 8852 14280 8904 14332
rect 11888 14280 11940 14332
rect 7012 14212 7064 14264
rect 7656 14144 7708 14196
rect 4896 14119 4948 14128
rect 4896 14085 4905 14119
rect 4905 14085 4939 14119
rect 4939 14085 4948 14119
rect 4896 14076 4948 14085
rect 5080 14076 5132 14128
rect 5264 14076 5316 14128
rect 13360 14280 13412 14332
rect 14464 14280 14516 14332
rect 16948 14280 17000 14332
rect 17224 14323 17276 14332
rect 17224 14289 17233 14323
rect 17233 14289 17267 14323
rect 17267 14289 17276 14323
rect 20168 14348 20220 14400
rect 17224 14280 17276 14289
rect 12808 14076 12860 14128
rect 12992 14255 13044 14264
rect 12992 14221 13001 14255
rect 13001 14221 13035 14255
rect 13035 14221 13044 14255
rect 12992 14212 13044 14221
rect 13268 14212 13320 14264
rect 17316 14255 17368 14264
rect 17316 14221 17325 14255
rect 17325 14221 17359 14255
rect 17359 14221 17368 14255
rect 17316 14212 17368 14221
rect 17408 14212 17460 14264
rect 17132 14076 17184 14128
rect 4414 13974 4466 14026
rect 4478 13974 4530 14026
rect 4542 13974 4594 14026
rect 4606 13974 4658 14026
rect 11278 13974 11330 14026
rect 11342 13974 11394 14026
rect 11406 13974 11458 14026
rect 11470 13974 11522 14026
rect 18142 13974 18194 14026
rect 18206 13974 18258 14026
rect 18270 13974 18322 14026
rect 18334 13974 18386 14026
rect 3424 13915 3476 13924
rect 3424 13881 3433 13915
rect 3433 13881 3467 13915
rect 3467 13881 3476 13915
rect 3424 13872 3476 13881
rect 5264 13872 5316 13924
rect 7012 13915 7064 13924
rect 7012 13881 7021 13915
rect 7021 13881 7055 13915
rect 7055 13881 7064 13915
rect 7012 13872 7064 13881
rect 8668 13915 8720 13924
rect 1492 13736 1544 13788
rect 5080 13779 5132 13788
rect 5080 13745 5089 13779
rect 5089 13745 5123 13779
rect 5123 13745 5132 13779
rect 5080 13736 5132 13745
rect 4896 13668 4948 13720
rect 8668 13881 8677 13915
rect 8677 13881 8711 13915
rect 8711 13881 8720 13915
rect 8668 13872 8720 13881
rect 12072 13915 12124 13924
rect 12072 13881 12081 13915
rect 12081 13881 12115 13915
rect 12115 13881 12124 13915
rect 12072 13872 12124 13881
rect 12900 13872 12952 13924
rect 17500 13872 17552 13924
rect 18604 13872 18656 13924
rect 20536 13872 20588 13924
rect 10692 13779 10744 13788
rect 10692 13745 10701 13779
rect 10701 13745 10735 13779
rect 10735 13745 10744 13779
rect 10692 13736 10744 13745
rect 12992 13779 13044 13788
rect 7196 13600 7248 13652
rect 8300 13668 8352 13720
rect 10600 13668 10652 13720
rect 8392 13600 8444 13652
rect 11060 13600 11112 13652
rect 12992 13745 13001 13779
rect 13001 13745 13035 13779
rect 13035 13745 13044 13779
rect 12992 13736 13044 13745
rect 13360 13779 13412 13788
rect 13360 13745 13369 13779
rect 13369 13745 13403 13779
rect 13403 13745 13412 13779
rect 13360 13736 13412 13745
rect 17132 13779 17184 13788
rect 17132 13745 17141 13779
rect 17141 13745 17175 13779
rect 17175 13745 17184 13779
rect 17132 13736 17184 13745
rect 17316 13779 17368 13788
rect 17316 13745 17325 13779
rect 17325 13745 17359 13779
rect 17359 13745 17368 13779
rect 17316 13736 17368 13745
rect 11888 13668 11940 13720
rect 18328 13711 18380 13720
rect 18328 13677 18337 13711
rect 18337 13677 18371 13711
rect 18371 13677 18380 13711
rect 18328 13668 18380 13677
rect 20260 13711 20312 13720
rect 20260 13677 20269 13711
rect 20269 13677 20303 13711
rect 20303 13677 20312 13711
rect 20260 13668 20312 13677
rect 16120 13600 16172 13652
rect 16948 13600 17000 13652
rect 4988 13575 5040 13584
rect 4988 13541 4997 13575
rect 4997 13541 5031 13575
rect 5031 13541 5040 13575
rect 4988 13532 5040 13541
rect 8208 13532 8260 13584
rect 11152 13532 11204 13584
rect 11704 13532 11756 13584
rect 7846 13430 7898 13482
rect 7910 13430 7962 13482
rect 7974 13430 8026 13482
rect 8038 13430 8090 13482
rect 14710 13430 14762 13482
rect 14774 13430 14826 13482
rect 14838 13430 14890 13482
rect 14902 13430 14954 13482
rect 4988 13371 5040 13380
rect 4988 13337 4997 13371
rect 4997 13337 5031 13371
rect 5031 13337 5040 13371
rect 4988 13328 5040 13337
rect 10600 13328 10652 13380
rect 10968 13328 11020 13380
rect 12808 13371 12860 13380
rect 12808 13337 12817 13371
rect 12817 13337 12851 13371
rect 12851 13337 12860 13371
rect 12808 13328 12860 13337
rect 12900 13371 12952 13380
rect 12900 13337 12909 13371
rect 12909 13337 12943 13371
rect 12943 13337 12952 13371
rect 12900 13328 12952 13337
rect 18788 13328 18840 13380
rect 20352 13328 20404 13380
rect 20720 13371 20772 13380
rect 20720 13337 20729 13371
rect 20729 13337 20763 13371
rect 20763 13337 20772 13371
rect 20720 13328 20772 13337
rect 18328 13260 18380 13312
rect 17592 13192 17644 13244
rect 19984 13235 20036 13244
rect 19984 13201 19993 13235
rect 19993 13201 20027 13235
rect 20027 13201 20036 13235
rect 19984 13192 20036 13201
rect 12072 13124 12124 13176
rect 15568 13124 15620 13176
rect 17408 12988 17460 13040
rect 4414 12886 4466 12938
rect 4478 12886 4530 12938
rect 4542 12886 4594 12938
rect 4606 12886 4658 12938
rect 11278 12886 11330 12938
rect 11342 12886 11394 12938
rect 11406 12886 11458 12938
rect 11470 12886 11522 12938
rect 18142 12886 18194 12938
rect 18206 12886 18258 12938
rect 18270 12886 18322 12938
rect 18334 12886 18386 12938
rect 11060 12827 11112 12836
rect 11060 12793 11069 12827
rect 11069 12793 11103 12827
rect 11103 12793 11112 12827
rect 11060 12784 11112 12793
rect 12440 12827 12492 12836
rect 12440 12793 12449 12827
rect 12449 12793 12483 12827
rect 12483 12793 12492 12827
rect 12440 12784 12492 12793
rect 14096 12784 14148 12836
rect 19984 12784 20036 12836
rect 20352 12827 20404 12836
rect 20352 12793 20361 12827
rect 20361 12793 20395 12827
rect 20395 12793 20404 12827
rect 20352 12784 20404 12793
rect 10968 12648 11020 12700
rect 19616 12716 19668 12768
rect 8300 12580 8352 12632
rect 11152 12623 11204 12632
rect 11152 12589 11161 12623
rect 11161 12589 11195 12623
rect 11195 12589 11204 12623
rect 11152 12580 11204 12589
rect 12440 12648 12492 12700
rect 13360 12648 13412 12700
rect 15568 12691 15620 12700
rect 15568 12657 15577 12691
rect 15577 12657 15611 12691
rect 15611 12657 15620 12691
rect 15568 12648 15620 12657
rect 14188 12580 14240 12632
rect 14464 12580 14516 12632
rect 16672 12623 16724 12632
rect 16672 12589 16681 12623
rect 16681 12589 16715 12623
rect 16715 12589 16724 12623
rect 16672 12580 16724 12589
rect 19248 12580 19300 12632
rect 20168 12623 20220 12632
rect 20168 12589 20177 12623
rect 20177 12589 20211 12623
rect 20211 12589 20220 12623
rect 20168 12580 20220 12589
rect 9864 12512 9916 12564
rect 14004 12512 14056 12564
rect 17500 12512 17552 12564
rect 19800 12512 19852 12564
rect 20076 12512 20128 12564
rect 8484 12444 8536 12496
rect 9680 12444 9732 12496
rect 13452 12444 13504 12496
rect 18052 12487 18104 12496
rect 18052 12453 18061 12487
rect 18061 12453 18095 12487
rect 18095 12453 18104 12487
rect 18052 12444 18104 12453
rect 7846 12342 7898 12394
rect 7910 12342 7962 12394
rect 7974 12342 8026 12394
rect 8038 12342 8090 12394
rect 14710 12342 14762 12394
rect 14774 12342 14826 12394
rect 14838 12342 14890 12394
rect 14902 12342 14954 12394
rect 1952 12240 2004 12292
rect 7656 12240 7708 12292
rect 8208 12104 8260 12156
rect 8392 12104 8444 12156
rect 8300 12079 8352 12088
rect 8300 12045 8309 12079
rect 8309 12045 8343 12079
rect 8343 12045 8352 12079
rect 8300 12036 8352 12045
rect 11152 12240 11204 12292
rect 13452 12240 13504 12292
rect 14004 12283 14056 12292
rect 10416 12215 10468 12224
rect 10416 12181 10425 12215
rect 10425 12181 10459 12215
rect 10459 12181 10468 12215
rect 10416 12172 10468 12181
rect 14004 12249 14013 12283
rect 14013 12249 14047 12283
rect 14047 12249 14056 12283
rect 14004 12240 14056 12249
rect 18788 12240 18840 12292
rect 20260 12240 20312 12292
rect 14556 12172 14608 12224
rect 10324 12147 10376 12156
rect 10324 12113 10333 12147
rect 10333 12113 10367 12147
rect 10367 12113 10376 12147
rect 10324 12104 10376 12113
rect 12992 12104 13044 12156
rect 14188 12104 14240 12156
rect 13176 12079 13228 12088
rect 6828 11943 6880 11952
rect 6828 11909 6837 11943
rect 6837 11909 6871 11943
rect 6871 11909 6880 11943
rect 6828 11900 6880 11909
rect 7196 11900 7248 11952
rect 7564 11900 7616 11952
rect 9864 11968 9916 12020
rect 13176 12045 13185 12079
rect 13185 12045 13219 12079
rect 13219 12045 13228 12079
rect 13176 12036 13228 12045
rect 12624 11968 12676 12020
rect 13728 12036 13780 12088
rect 18052 12172 18104 12224
rect 8576 11900 8628 11952
rect 8944 11900 8996 11952
rect 13728 11943 13780 11952
rect 13728 11909 13737 11943
rect 13737 11909 13771 11943
rect 13771 11909 13780 11943
rect 13728 11900 13780 11909
rect 17960 12104 18012 12156
rect 16948 12036 17000 12088
rect 20168 12172 20220 12224
rect 19984 12147 20036 12156
rect 19984 12113 19993 12147
rect 19993 12113 20027 12147
rect 20027 12113 20036 12147
rect 19984 12104 20036 12113
rect 20536 12147 20588 12156
rect 20536 12113 20545 12147
rect 20545 12113 20579 12147
rect 20579 12113 20588 12147
rect 20536 12104 20588 12113
rect 20904 11968 20956 12020
rect 18604 11900 18656 11952
rect 4414 11798 4466 11850
rect 4478 11798 4530 11850
rect 4542 11798 4594 11850
rect 4606 11798 4658 11850
rect 11278 11798 11330 11850
rect 11342 11798 11394 11850
rect 11406 11798 11458 11850
rect 11470 11798 11522 11850
rect 18142 11798 18194 11850
rect 18206 11798 18258 11850
rect 18270 11798 18322 11850
rect 18334 11798 18386 11850
rect 10324 11739 10376 11748
rect 10324 11705 10333 11739
rect 10333 11705 10367 11739
rect 10367 11705 10376 11739
rect 10324 11696 10376 11705
rect 14464 11696 14516 11748
rect 17960 11696 18012 11748
rect 19892 11696 19944 11748
rect 8392 11628 8444 11680
rect 8576 11560 8628 11612
rect 12992 11628 13044 11680
rect 18512 11628 18564 11680
rect 14188 11603 14240 11612
rect 14188 11569 14197 11603
rect 14197 11569 14231 11603
rect 14231 11569 14240 11603
rect 14188 11560 14240 11569
rect 17500 11560 17552 11612
rect 7564 11424 7616 11476
rect 7748 11424 7800 11476
rect 8944 11424 8996 11476
rect 12624 11492 12676 11544
rect 14096 11535 14148 11544
rect 14096 11501 14105 11535
rect 14105 11501 14139 11535
rect 14139 11501 14148 11535
rect 14096 11492 14148 11501
rect 20260 11535 20312 11544
rect 20260 11501 20269 11535
rect 20269 11501 20303 11535
rect 20303 11501 20312 11535
rect 20260 11492 20312 11501
rect 8208 11356 8260 11408
rect 8484 11399 8536 11408
rect 8484 11365 8493 11399
rect 8493 11365 8527 11399
rect 8527 11365 8536 11399
rect 8484 11356 8536 11365
rect 10600 11356 10652 11408
rect 12808 11424 12860 11476
rect 13728 11424 13780 11476
rect 12992 11356 13044 11408
rect 13360 11399 13412 11408
rect 13360 11365 13369 11399
rect 13369 11365 13403 11399
rect 13403 11365 13412 11399
rect 13360 11356 13412 11365
rect 14004 11399 14056 11408
rect 14004 11365 14013 11399
rect 14013 11365 14047 11399
rect 14047 11365 14056 11399
rect 14004 11356 14056 11365
rect 18880 11356 18932 11408
rect 7846 11254 7898 11306
rect 7910 11254 7962 11306
rect 7974 11254 8026 11306
rect 8038 11254 8090 11306
rect 14710 11254 14762 11306
rect 14774 11254 14826 11306
rect 14838 11254 14890 11306
rect 14902 11254 14954 11306
rect 8208 11152 8260 11204
rect 12256 11152 12308 11204
rect 20 11084 72 11136
rect 13176 11084 13228 11136
rect 14004 11152 14056 11204
rect 14096 11152 14148 11204
rect 14280 11152 14332 11204
rect 18880 11195 18932 11204
rect 18880 11161 18889 11195
rect 18889 11161 18923 11195
rect 18923 11161 18932 11195
rect 18880 11152 18932 11161
rect 20628 11152 20680 11204
rect 20812 11152 20864 11204
rect 16488 11084 16540 11136
rect 6828 11016 6880 11068
rect 16120 11016 16172 11068
rect 17316 11059 17368 11068
rect 17316 11025 17325 11059
rect 17325 11025 17359 11059
rect 17359 11025 17368 11059
rect 17316 11016 17368 11025
rect 17408 11016 17460 11068
rect 17868 11016 17920 11068
rect 19984 11059 20036 11068
rect 19984 11025 19993 11059
rect 19993 11025 20027 11059
rect 20027 11025 20036 11059
rect 19984 11016 20036 11025
rect 8392 10991 8444 11000
rect 8392 10957 8401 10991
rect 8401 10957 8435 10991
rect 8435 10957 8444 10991
rect 8392 10948 8444 10957
rect 12992 10948 13044 11000
rect 14096 10991 14148 11000
rect 14096 10957 14105 10991
rect 14105 10957 14139 10991
rect 14139 10957 14148 10991
rect 14096 10948 14148 10957
rect 16488 10991 16540 11000
rect 10416 10880 10468 10932
rect 13360 10880 13412 10932
rect 16488 10957 16497 10991
rect 16497 10957 16531 10991
rect 16531 10957 16540 10991
rect 16488 10948 16540 10957
rect 17500 10991 17552 11000
rect 15660 10880 15712 10932
rect 15936 10880 15988 10932
rect 16948 10923 17000 10932
rect 16948 10889 16957 10923
rect 16957 10889 16991 10923
rect 16991 10889 17000 10923
rect 16948 10880 17000 10889
rect 17500 10957 17509 10991
rect 17509 10957 17543 10991
rect 17543 10957 17552 10991
rect 17500 10948 17552 10957
rect 19248 10880 19300 10932
rect 4414 10710 4466 10762
rect 4478 10710 4530 10762
rect 4542 10710 4594 10762
rect 4606 10710 4658 10762
rect 11278 10710 11330 10762
rect 11342 10710 11394 10762
rect 11406 10710 11458 10762
rect 11470 10710 11522 10762
rect 18142 10710 18194 10762
rect 18206 10710 18258 10762
rect 18270 10710 18322 10762
rect 18334 10710 18386 10762
rect 8576 10651 8628 10660
rect 8576 10617 8585 10651
rect 8585 10617 8619 10651
rect 8619 10617 8628 10651
rect 8576 10608 8628 10617
rect 17316 10608 17368 10660
rect 19340 10608 19392 10660
rect 9864 10336 9916 10388
rect 16396 10540 16448 10592
rect 16488 10472 16540 10524
rect 19248 10472 19300 10524
rect 11612 10404 11664 10456
rect 20260 10447 20312 10456
rect 10416 10379 10468 10388
rect 10416 10345 10425 10379
rect 10425 10345 10459 10379
rect 10459 10345 10468 10379
rect 10416 10336 10468 10345
rect 11244 10336 11296 10388
rect 11796 10336 11848 10388
rect 7564 10268 7616 10320
rect 10508 10311 10560 10320
rect 10508 10277 10517 10311
rect 10517 10277 10551 10311
rect 10551 10277 10560 10311
rect 10508 10268 10560 10277
rect 16764 10268 16816 10320
rect 20260 10413 20269 10447
rect 20269 10413 20303 10447
rect 20303 10413 20312 10447
rect 20260 10404 20312 10413
rect 18696 10268 18748 10320
rect 7846 10166 7898 10218
rect 7910 10166 7962 10218
rect 7974 10166 8026 10218
rect 8038 10166 8090 10218
rect 14710 10166 14762 10218
rect 14774 10166 14826 10218
rect 14838 10166 14890 10218
rect 14902 10166 14954 10218
rect 9864 10107 9916 10116
rect 9864 10073 9873 10107
rect 9873 10073 9907 10107
rect 9907 10073 9916 10107
rect 9864 10064 9916 10073
rect 11244 10107 11296 10116
rect 11244 10073 11253 10107
rect 11253 10073 11287 10107
rect 11287 10073 11296 10107
rect 11244 10064 11296 10073
rect 11612 10064 11664 10116
rect 14188 10107 14240 10116
rect 14188 10073 14197 10107
rect 14197 10073 14231 10107
rect 14231 10073 14240 10107
rect 14188 10064 14240 10073
rect 17500 10064 17552 10116
rect 19248 10064 19300 10116
rect 20996 10064 21048 10116
rect 13360 9996 13412 10048
rect 16488 9996 16540 10048
rect 8760 9971 8812 9980
rect 8760 9937 8794 9971
rect 8794 9937 8812 9971
rect 8760 9928 8812 9937
rect 12808 9971 12860 9980
rect 12808 9937 12817 9971
rect 12817 9937 12851 9971
rect 12851 9937 12860 9971
rect 12808 9928 12860 9937
rect 13636 9928 13688 9980
rect 16672 9928 16724 9980
rect 17960 9928 18012 9980
rect 18788 9971 18840 9980
rect 18788 9937 18822 9971
rect 18822 9937 18840 9971
rect 18788 9928 18840 9937
rect 20536 9971 20588 9980
rect 20536 9937 20545 9971
rect 20545 9937 20579 9971
rect 20579 9937 20588 9971
rect 20536 9928 20588 9937
rect 7564 9860 7616 9912
rect 11612 9860 11664 9912
rect 10876 9767 10928 9776
rect 10876 9733 10885 9767
rect 10885 9733 10919 9767
rect 10919 9733 10928 9767
rect 10876 9724 10928 9733
rect 4414 9622 4466 9674
rect 4478 9622 4530 9674
rect 4542 9622 4594 9674
rect 4606 9622 4658 9674
rect 11278 9622 11330 9674
rect 11342 9622 11394 9674
rect 11406 9622 11458 9674
rect 11470 9622 11522 9674
rect 18142 9622 18194 9674
rect 18206 9622 18258 9674
rect 18270 9622 18322 9674
rect 18334 9622 18386 9674
rect 10508 9520 10560 9572
rect 8760 9452 8812 9504
rect 10600 9427 10652 9436
rect 10600 9393 10609 9427
rect 10609 9393 10643 9427
rect 10643 9393 10652 9427
rect 10600 9384 10652 9393
rect 7564 9359 7616 9368
rect 7564 9325 7573 9359
rect 7573 9325 7607 9359
rect 7607 9325 7616 9359
rect 7564 9316 7616 9325
rect 10876 9316 10928 9368
rect 11612 9384 11664 9436
rect 12348 9248 12400 9300
rect 11428 9223 11480 9232
rect 11428 9189 11437 9223
rect 11437 9189 11471 9223
rect 11471 9189 11480 9223
rect 11428 9180 11480 9189
rect 12072 9223 12124 9232
rect 12072 9189 12081 9223
rect 12081 9189 12115 9223
rect 12115 9189 12124 9223
rect 12072 9180 12124 9189
rect 12440 9223 12492 9232
rect 12440 9189 12449 9223
rect 12449 9189 12483 9223
rect 12483 9189 12492 9223
rect 16120 9452 16172 9504
rect 16396 9452 16448 9504
rect 17592 9495 17644 9504
rect 17592 9461 17601 9495
rect 17601 9461 17635 9495
rect 17635 9461 17644 9495
rect 17592 9452 17644 9461
rect 13636 9316 13688 9368
rect 14188 9316 14240 9368
rect 18236 9427 18288 9436
rect 18236 9393 18245 9427
rect 18245 9393 18279 9427
rect 18279 9393 18288 9427
rect 18236 9384 18288 9393
rect 19432 9384 19484 9436
rect 18972 9359 19024 9368
rect 18972 9325 18981 9359
rect 18981 9325 19015 9359
rect 19015 9325 19024 9359
rect 18972 9316 19024 9325
rect 12440 9180 12492 9189
rect 19064 9223 19116 9232
rect 19064 9189 19073 9223
rect 19073 9189 19107 9223
rect 19107 9189 19116 9223
rect 19064 9180 19116 9189
rect 7846 9078 7898 9130
rect 7910 9078 7962 9130
rect 7974 9078 8026 9130
rect 8038 9078 8090 9130
rect 14710 9078 14762 9130
rect 14774 9078 14826 9130
rect 14838 9078 14890 9130
rect 14902 9078 14954 9130
rect 10416 8976 10468 9028
rect 12072 8976 12124 9028
rect 13084 8976 13136 9028
rect 15108 8976 15160 9028
rect 2688 8908 2740 8960
rect 11428 8908 11480 8960
rect 12440 8908 12492 8960
rect 17868 8976 17920 9028
rect 18236 8976 18288 9028
rect 18788 8976 18840 9028
rect 20076 8976 20128 9028
rect 16304 8908 16356 8960
rect 13452 8840 13504 8892
rect 15660 8840 15712 8892
rect 17960 8840 18012 8892
rect 19432 8840 19484 8892
rect 19984 8883 20036 8892
rect 19984 8849 19993 8883
rect 19993 8849 20027 8883
rect 20027 8849 20036 8883
rect 19984 8840 20036 8849
rect 20536 8883 20588 8892
rect 20536 8849 20545 8883
rect 20545 8849 20579 8883
rect 20579 8849 20588 8883
rect 20536 8840 20588 8849
rect 10600 8772 10652 8824
rect 12348 8772 12400 8824
rect 15936 8772 15988 8824
rect 18512 8636 18564 8688
rect 18788 8636 18840 8688
rect 4414 8534 4466 8586
rect 4478 8534 4530 8586
rect 4542 8534 4594 8586
rect 4606 8534 4658 8586
rect 11278 8534 11330 8586
rect 11342 8534 11394 8586
rect 11406 8534 11458 8586
rect 11470 8534 11522 8586
rect 18142 8534 18194 8586
rect 18206 8534 18258 8586
rect 18270 8534 18322 8586
rect 18334 8534 18386 8586
rect 11980 8432 12032 8484
rect 20444 8475 20496 8484
rect 20444 8441 20453 8475
rect 20453 8441 20487 8475
rect 20487 8441 20496 8475
rect 20444 8432 20496 8441
rect 13452 8339 13504 8348
rect 13452 8305 13461 8339
rect 13461 8305 13495 8339
rect 13495 8305 13504 8339
rect 13452 8296 13504 8305
rect 15660 8339 15712 8348
rect 15660 8305 15669 8339
rect 15669 8305 15703 8339
rect 15703 8305 15712 8339
rect 15660 8296 15712 8305
rect 11336 8271 11388 8280
rect 11336 8237 11345 8271
rect 11345 8237 11379 8271
rect 11379 8237 11388 8271
rect 11336 8228 11388 8237
rect 13268 8271 13320 8280
rect 13268 8237 13277 8271
rect 13277 8237 13311 8271
rect 13311 8237 13320 8271
rect 13268 8228 13320 8237
rect 17408 8296 17460 8348
rect 16672 8271 16724 8280
rect 16672 8237 16681 8271
rect 16681 8237 16715 8271
rect 16715 8237 16724 8271
rect 16672 8228 16724 8237
rect 20260 8271 20312 8280
rect 20260 8237 20269 8271
rect 20269 8237 20303 8271
rect 20303 8237 20312 8271
rect 20260 8228 20312 8237
rect 7846 7990 7898 8042
rect 7910 7990 7962 8042
rect 7974 7990 8026 8042
rect 8038 7990 8090 8042
rect 14710 7990 14762 8042
rect 14774 7990 14826 8042
rect 14838 7990 14890 8042
rect 14902 7990 14954 8042
rect 13268 7888 13320 7940
rect 17408 7931 17460 7940
rect 17408 7897 17417 7931
rect 17417 7897 17451 7931
rect 17451 7897 17460 7931
rect 17408 7888 17460 7897
rect 19432 7931 19484 7940
rect 19432 7897 19441 7931
rect 19441 7897 19475 7931
rect 19475 7897 19484 7931
rect 19432 7888 19484 7897
rect 11336 7820 11388 7872
rect 14372 7820 14424 7872
rect 10324 7752 10376 7804
rect 14648 7752 14700 7804
rect 16580 7752 16632 7804
rect 19984 7795 20036 7804
rect 14096 7727 14148 7736
rect 14096 7693 14105 7727
rect 14105 7693 14139 7727
rect 14139 7693 14148 7727
rect 14096 7684 14148 7693
rect 14280 7727 14332 7736
rect 14280 7693 14289 7727
rect 14289 7693 14323 7727
rect 14323 7693 14332 7727
rect 14280 7684 14332 7693
rect 16028 7727 16080 7736
rect 16028 7693 16037 7727
rect 16037 7693 16071 7727
rect 16071 7693 16080 7727
rect 16028 7684 16080 7693
rect 17960 7684 18012 7736
rect 19984 7761 19993 7795
rect 19993 7761 20027 7795
rect 20027 7761 20036 7795
rect 19984 7752 20036 7761
rect 20536 7795 20588 7804
rect 20536 7761 20545 7795
rect 20545 7761 20579 7795
rect 20579 7761 20588 7795
rect 20536 7752 20588 7761
rect 16212 7548 16264 7600
rect 4414 7446 4466 7498
rect 4478 7446 4530 7498
rect 4542 7446 4594 7498
rect 4606 7446 4658 7498
rect 11278 7446 11330 7498
rect 11342 7446 11394 7498
rect 11406 7446 11458 7498
rect 11470 7446 11522 7498
rect 18142 7446 18194 7498
rect 18206 7446 18258 7498
rect 18270 7446 18322 7498
rect 18334 7446 18386 7498
rect 10324 7387 10376 7396
rect 10324 7353 10333 7387
rect 10333 7353 10367 7387
rect 10367 7353 10376 7387
rect 10324 7344 10376 7353
rect 10600 7208 10652 7260
rect 13636 7344 13688 7396
rect 14648 7251 14700 7260
rect 14648 7217 14657 7251
rect 14657 7217 14691 7251
rect 14691 7217 14700 7251
rect 14648 7208 14700 7217
rect 16028 7344 16080 7396
rect 16580 7344 16632 7396
rect 17224 7344 17276 7396
rect 10784 7047 10836 7056
rect 10784 7013 10793 7047
rect 10793 7013 10827 7047
rect 10827 7013 10836 7047
rect 10784 7004 10836 7013
rect 14556 7140 14608 7192
rect 14280 7072 14332 7124
rect 7846 6902 7898 6954
rect 7910 6902 7962 6954
rect 7974 6902 8026 6954
rect 8038 6902 8090 6954
rect 14710 6902 14762 6954
rect 14774 6902 14826 6954
rect 14838 6902 14890 6954
rect 14902 6902 14954 6954
rect 10600 6843 10652 6852
rect 10600 6809 10609 6843
rect 10609 6809 10643 6843
rect 10643 6809 10652 6843
rect 10600 6800 10652 6809
rect 10784 6800 10836 6852
rect 14096 6800 14148 6852
rect 16948 6800 17000 6852
rect 18512 6800 18564 6852
rect 15200 6732 15252 6784
rect 2964 6664 3016 6716
rect 11704 6664 11756 6716
rect 14556 6639 14608 6648
rect 7564 6460 7616 6512
rect 14556 6605 14565 6639
rect 14565 6605 14599 6639
rect 14599 6605 14608 6639
rect 14556 6596 14608 6605
rect 19064 6664 19116 6716
rect 20536 6707 20588 6716
rect 20536 6673 20545 6707
rect 20545 6673 20579 6707
rect 20579 6673 20588 6707
rect 20536 6664 20588 6673
rect 17224 6639 17276 6648
rect 17224 6605 17233 6639
rect 17233 6605 17267 6639
rect 17267 6605 17276 6639
rect 17224 6596 17276 6605
rect 11704 6528 11756 6580
rect 16672 6571 16724 6580
rect 16672 6537 16681 6571
rect 16681 6537 16715 6571
rect 16715 6537 16724 6571
rect 16672 6528 16724 6537
rect 18604 6528 18656 6580
rect 19064 6528 19116 6580
rect 13728 6460 13780 6512
rect 4414 6358 4466 6410
rect 4478 6358 4530 6410
rect 4542 6358 4594 6410
rect 4606 6358 4658 6410
rect 11278 6358 11330 6410
rect 11342 6358 11394 6410
rect 11406 6358 11458 6410
rect 11470 6358 11522 6410
rect 18142 6358 18194 6410
rect 18206 6358 18258 6410
rect 18270 6358 18322 6410
rect 18334 6358 18386 6410
rect 15200 6256 15252 6308
rect 17960 6256 18012 6308
rect 7846 5814 7898 5866
rect 7910 5814 7962 5866
rect 7974 5814 8026 5866
rect 8038 5814 8090 5866
rect 14710 5814 14762 5866
rect 14774 5814 14826 5866
rect 14838 5814 14890 5866
rect 14902 5814 14954 5866
rect 12532 5712 12584 5764
rect 20536 5619 20588 5628
rect 20536 5585 20545 5619
rect 20545 5585 20579 5619
rect 20579 5585 20588 5619
rect 20536 5576 20588 5585
rect 4414 5270 4466 5322
rect 4478 5270 4530 5322
rect 4542 5270 4594 5322
rect 4606 5270 4658 5322
rect 11278 5270 11330 5322
rect 11342 5270 11394 5322
rect 11406 5270 11458 5322
rect 11470 5270 11522 5322
rect 18142 5270 18194 5322
rect 18206 5270 18258 5322
rect 18270 5270 18322 5322
rect 18334 5270 18386 5322
rect 16948 5168 17000 5220
rect 17960 5168 18012 5220
rect 7846 4726 7898 4778
rect 7910 4726 7962 4778
rect 7974 4726 8026 4778
rect 8038 4726 8090 4778
rect 14710 4726 14762 4778
rect 14774 4726 14826 4778
rect 14838 4726 14890 4778
rect 14902 4726 14954 4778
rect 21088 4624 21140 4676
rect 20536 4531 20588 4540
rect 20536 4497 20545 4531
rect 20545 4497 20579 4531
rect 20579 4497 20588 4531
rect 20536 4488 20588 4497
rect 4414 4182 4466 4234
rect 4478 4182 4530 4234
rect 4542 4182 4594 4234
rect 4606 4182 4658 4234
rect 11278 4182 11330 4234
rect 11342 4182 11394 4234
rect 11406 4182 11458 4234
rect 11470 4182 11522 4234
rect 18142 4182 18194 4234
rect 18206 4182 18258 4234
rect 18270 4182 18322 4234
rect 18334 4182 18386 4234
rect 14188 3944 14240 3996
rect 18512 3944 18564 3996
rect 15936 3876 15988 3928
rect 19248 3876 19300 3928
rect 7846 3638 7898 3690
rect 7910 3638 7962 3690
rect 7974 3638 8026 3690
rect 8038 3638 8090 3690
rect 14710 3638 14762 3690
rect 14774 3638 14826 3690
rect 14838 3638 14890 3690
rect 14902 3638 14954 3690
rect 4414 3094 4466 3146
rect 4478 3094 4530 3146
rect 4542 3094 4594 3146
rect 4606 3094 4658 3146
rect 11278 3094 11330 3146
rect 11342 3094 11394 3146
rect 11406 3094 11458 3146
rect 11470 3094 11522 3146
rect 18142 3094 18194 3146
rect 18206 3094 18258 3146
rect 18270 3094 18322 3146
rect 18334 3094 18386 3146
rect 7846 2550 7898 2602
rect 7910 2550 7962 2602
rect 7974 2550 8026 2602
rect 8038 2550 8090 2602
rect 14710 2550 14762 2602
rect 14774 2550 14826 2602
rect 14838 2550 14890 2602
rect 14902 2550 14954 2602
rect 16856 2244 16908 2296
rect 19248 2244 19300 2296
rect 4414 2006 4466 2058
rect 4478 2006 4530 2058
rect 4542 2006 4594 2058
rect 4606 2006 4658 2058
rect 11278 2006 11330 2058
rect 11342 2006 11394 2058
rect 11406 2006 11458 2058
rect 11470 2006 11522 2058
rect 18142 2006 18194 2058
rect 18206 2006 18258 2058
rect 18270 2006 18322 2058
rect 18334 2006 18386 2058
rect 16396 1156 16448 1208
rect 17960 1156 18012 1208
<< metal2 >>
rect 294 21856 350 22656
rect 846 21856 902 22656
rect 1398 21856 1454 22656
rect 1950 21856 2006 22656
rect 2502 21856 2558 22656
rect 3054 21856 3110 22656
rect 3606 21856 3662 22656
rect 4158 21856 4214 22656
rect 4710 21856 4766 22656
rect 5262 21856 5318 22656
rect 5814 21856 5870 22656
rect 6366 21856 6422 22656
rect 6918 21856 6974 22656
rect 7470 21856 7526 22656
rect 8022 21856 8078 22656
rect 8574 21856 8630 22656
rect 9126 21856 9182 22656
rect 9678 21856 9734 22656
rect 10230 21856 10286 22656
rect 10782 21856 10838 22656
rect 11334 21856 11390 22656
rect 11978 21856 12034 22656
rect 12530 21856 12586 22656
rect 13082 21856 13138 22656
rect 13634 21856 13690 22656
rect 14186 21856 14242 22656
rect 14738 21856 14794 22656
rect 15290 21856 15346 22656
rect 15842 21856 15898 22656
rect 16394 21856 16450 22656
rect 16946 21856 17002 22656
rect 17498 21856 17554 22656
rect 17958 22392 18014 22401
rect 17958 22327 18014 22336
rect 308 18078 336 21856
rect 296 18072 348 18078
rect 296 18014 348 18020
rect 860 17874 888 21856
rect 1412 17942 1440 21856
rect 1492 18480 1544 18486
rect 1492 18422 1544 18428
rect 1400 17936 1452 17942
rect 1400 17878 1452 17884
rect 20 17868 72 17874
rect 20 17810 72 17816
rect 848 17868 900 17874
rect 848 17810 900 17816
rect 32 11142 60 17810
rect 1504 17602 1532 18422
rect 1492 17596 1544 17602
rect 1492 17538 1544 17544
rect 1504 15970 1532 17538
rect 1492 15964 1544 15970
rect 1492 15906 1544 15912
rect 1504 14882 1532 15906
rect 1492 14876 1544 14882
rect 1492 14818 1544 14824
rect 1504 13794 1532 14818
rect 1492 13788 1544 13794
rect 1492 13730 1544 13736
rect 1964 12298 1992 21856
rect 2516 16310 2544 21856
rect 2780 18684 2832 18690
rect 2780 18626 2832 18632
rect 2792 18146 2820 18626
rect 2780 18140 2832 18146
rect 2780 18082 2832 18088
rect 2688 17936 2740 17942
rect 2688 17878 2740 17884
rect 2504 16304 2556 16310
rect 2504 16246 2556 16252
rect 1952 12292 2004 12298
rect 1952 12234 2004 12240
rect 20 11136 72 11142
rect 20 11078 72 11084
rect 2700 8966 2728 17878
rect 2792 17738 2820 18082
rect 3068 18010 3096 21856
rect 3056 18004 3108 18010
rect 3056 17946 3108 17952
rect 2964 17936 3016 17942
rect 2964 17878 3016 17884
rect 3148 17936 3200 17942
rect 3148 17878 3200 17884
rect 3240 17936 3292 17942
rect 3240 17878 3292 17884
rect 2780 17732 2832 17738
rect 2780 17674 2832 17680
rect 2976 16990 3004 17878
rect 3160 17058 3188 17878
rect 3252 17738 3280 17878
rect 3240 17732 3292 17738
rect 3240 17674 3292 17680
rect 3424 17596 3476 17602
rect 3424 17538 3476 17544
rect 3148 17052 3200 17058
rect 3148 16994 3200 17000
rect 2964 16984 3016 16990
rect 2964 16926 3016 16932
rect 3436 16106 3464 17538
rect 3424 16100 3476 16106
rect 3424 16042 3476 16048
rect 2872 15828 2924 15834
rect 2872 15770 2924 15776
rect 2884 15358 2912 15770
rect 3620 15562 3648 21856
rect 4172 17738 4200 21856
rect 4388 19468 4684 19488
rect 4444 19466 4468 19468
rect 4524 19466 4548 19468
rect 4604 19466 4628 19468
rect 4466 19414 4468 19466
rect 4530 19414 4542 19466
rect 4604 19414 4606 19466
rect 4444 19412 4468 19414
rect 4524 19412 4548 19414
rect 4604 19412 4628 19414
rect 4388 19392 4684 19412
rect 4724 18706 4752 21856
rect 5172 19228 5224 19234
rect 5172 19170 5224 19176
rect 4896 19024 4948 19030
rect 4896 18966 4948 18972
rect 5080 19024 5132 19030
rect 5080 18966 5132 18972
rect 4724 18678 4844 18706
rect 4816 18622 4844 18678
rect 4804 18616 4856 18622
rect 4804 18558 4856 18564
rect 4388 18380 4684 18400
rect 4444 18378 4468 18380
rect 4524 18378 4548 18380
rect 4604 18378 4628 18380
rect 4466 18326 4468 18378
rect 4530 18326 4542 18378
rect 4604 18326 4606 18378
rect 4444 18324 4468 18326
rect 4524 18324 4548 18326
rect 4604 18324 4628 18326
rect 4388 18304 4684 18324
rect 4160 17732 4212 17738
rect 4160 17674 4212 17680
rect 4712 17732 4764 17738
rect 4712 17674 4764 17680
rect 4388 17292 4684 17312
rect 4444 17290 4468 17292
rect 4524 17290 4548 17292
rect 4604 17290 4628 17292
rect 4466 17238 4468 17290
rect 4530 17238 4542 17290
rect 4604 17238 4606 17290
rect 4444 17236 4468 17238
rect 4524 17236 4548 17238
rect 4604 17236 4628 17238
rect 4388 17216 4684 17236
rect 4068 17188 4120 17194
rect 4068 17130 4120 17136
rect 4080 17097 4108 17130
rect 4066 17088 4122 17097
rect 4724 17058 4752 17674
rect 4908 17534 4936 18966
rect 4988 18684 5040 18690
rect 4988 18626 5040 18632
rect 5000 18282 5028 18626
rect 4988 18276 5040 18282
rect 4988 18218 5040 18224
rect 4896 17528 4948 17534
rect 4896 17470 4948 17476
rect 4066 17023 4122 17032
rect 4712 17052 4764 17058
rect 4712 16994 4764 17000
rect 4896 16984 4948 16990
rect 5000 16938 5028 18218
rect 5092 18146 5120 18966
rect 5184 18486 5212 19170
rect 5172 18480 5224 18486
rect 5172 18422 5224 18428
rect 5080 18140 5132 18146
rect 5080 18082 5132 18088
rect 4948 16932 5028 16938
rect 4896 16926 5028 16932
rect 4908 16910 5028 16926
rect 5184 16922 5212 18422
rect 5276 18026 5304 21856
rect 5448 19024 5500 19030
rect 5448 18966 5500 18972
rect 5460 18826 5488 18966
rect 5448 18820 5500 18826
rect 5448 18762 5500 18768
rect 5828 18729 5856 21856
rect 5814 18720 5870 18729
rect 5814 18655 5870 18664
rect 6380 18162 6408 21856
rect 6552 18684 6604 18690
rect 6552 18626 6604 18632
rect 6380 18134 6500 18162
rect 5276 17998 5580 18026
rect 6472 18010 6500 18134
rect 6564 18078 6592 18626
rect 6932 18570 6960 21856
rect 7104 18684 7156 18690
rect 7104 18626 7156 18632
rect 6932 18542 7052 18570
rect 7024 18486 7052 18542
rect 7012 18480 7064 18486
rect 7012 18422 7064 18428
rect 7116 18282 7144 18626
rect 7104 18276 7156 18282
rect 7104 18218 7156 18224
rect 6552 18072 6604 18078
rect 6552 18014 6604 18020
rect 5448 17936 5500 17942
rect 5448 17878 5500 17884
rect 4388 16204 4684 16224
rect 4444 16202 4468 16204
rect 4524 16202 4548 16204
rect 4604 16202 4628 16204
rect 4466 16150 4468 16202
rect 4530 16150 4542 16202
rect 4604 16150 4606 16202
rect 4444 16148 4468 16150
rect 4524 16148 4548 16150
rect 4604 16148 4628 16150
rect 4388 16128 4684 16148
rect 5000 15970 5028 16910
rect 5172 16916 5224 16922
rect 5172 16858 5224 16864
rect 4988 15964 5040 15970
rect 4988 15906 5040 15912
rect 3608 15556 3660 15562
rect 3608 15498 3660 15504
rect 3332 15420 3384 15426
rect 3332 15362 3384 15368
rect 2872 15352 2924 15358
rect 2872 15294 2924 15300
rect 2884 15018 2912 15294
rect 2872 15012 2924 15018
rect 2872 14954 2924 14960
rect 3344 14882 3372 15362
rect 3424 15352 3476 15358
rect 3424 15294 3476 15300
rect 3332 14876 3384 14882
rect 3332 14818 3384 14824
rect 3436 14746 3464 15294
rect 4388 15116 4684 15136
rect 4444 15114 4468 15116
rect 4524 15114 4548 15116
rect 4604 15114 4628 15116
rect 4466 15062 4468 15114
rect 4530 15062 4542 15114
rect 4604 15062 4606 15114
rect 4444 15060 4468 15062
rect 4524 15060 4548 15062
rect 4604 15060 4628 15062
rect 4388 15040 4684 15060
rect 5000 15018 5028 15906
rect 4988 15012 5040 15018
rect 4988 14954 5040 14960
rect 3424 14740 3476 14746
rect 3424 14682 3476 14688
rect 3436 13930 3464 14682
rect 5000 14338 5028 14954
rect 5460 14354 5488 17878
rect 5552 16922 5580 17998
rect 6368 18004 6420 18010
rect 6368 17946 6420 17952
rect 6460 18004 6512 18010
rect 6460 17946 6512 17952
rect 5540 16916 5592 16922
rect 5540 16858 5592 16864
rect 6380 16378 6408 17946
rect 6828 16984 6880 16990
rect 6828 16926 6880 16932
rect 6840 16650 6868 16926
rect 6828 16644 6880 16650
rect 6828 16586 6880 16592
rect 7288 16440 7340 16446
rect 7288 16382 7340 16388
rect 6368 16372 6420 16378
rect 6368 16314 6420 16320
rect 6380 16106 6408 16314
rect 7300 16106 7328 16382
rect 6368 16100 6420 16106
rect 6368 16042 6420 16048
rect 7288 16100 7340 16106
rect 7288 16042 7340 16048
rect 6368 15964 6420 15970
rect 6368 15906 6420 15912
rect 6380 15018 6408 15906
rect 7380 15896 7432 15902
rect 7380 15838 7432 15844
rect 7392 15494 7420 15838
rect 7380 15488 7432 15494
rect 7380 15430 7432 15436
rect 7484 15018 7512 21856
rect 8036 20202 8064 21856
rect 7760 20174 8064 20202
rect 7656 18072 7708 18078
rect 7656 18014 7708 18020
rect 7668 17670 7696 18014
rect 7656 17664 7708 17670
rect 7656 17606 7708 17612
rect 7564 17460 7616 17466
rect 7564 17402 7616 17408
rect 7576 17058 7604 17402
rect 7564 17052 7616 17058
rect 7564 16994 7616 17000
rect 7564 15828 7616 15834
rect 7564 15770 7616 15776
rect 7576 15494 7604 15770
rect 7564 15488 7616 15494
rect 7564 15430 7616 15436
rect 6368 15012 6420 15018
rect 6368 14954 6420 14960
rect 7472 15012 7524 15018
rect 7472 14954 7524 14960
rect 7668 14898 7696 17606
rect 7760 15902 7788 20174
rect 7820 20012 8116 20032
rect 7876 20010 7900 20012
rect 7956 20010 7980 20012
rect 8036 20010 8060 20012
rect 7898 19958 7900 20010
rect 7962 19958 7974 20010
rect 8036 19958 8038 20010
rect 7876 19956 7900 19958
rect 7956 19956 7980 19958
rect 8036 19956 8060 19958
rect 7820 19936 8116 19956
rect 8208 19228 8260 19234
rect 8208 19170 8260 19176
rect 7820 18924 8116 18944
rect 7876 18922 7900 18924
rect 7956 18922 7980 18924
rect 8036 18922 8060 18924
rect 7898 18870 7900 18922
rect 7962 18870 7974 18922
rect 8036 18870 8038 18922
rect 7876 18868 7900 18870
rect 7956 18868 7980 18870
rect 8036 18868 8060 18870
rect 7820 18848 8116 18868
rect 8220 18758 8248 19170
rect 8300 19024 8352 19030
rect 8300 18966 8352 18972
rect 8208 18752 8260 18758
rect 8114 18720 8170 18729
rect 8208 18694 8260 18700
rect 8114 18655 8170 18664
rect 8128 18214 8156 18655
rect 8220 18554 8248 18694
rect 8208 18548 8260 18554
rect 8208 18490 8260 18496
rect 8312 18282 8340 18966
rect 8484 18684 8536 18690
rect 8484 18626 8536 18632
rect 8300 18276 8352 18282
rect 8300 18218 8352 18224
rect 8116 18208 8168 18214
rect 8116 18150 8168 18156
rect 7820 17836 8116 17856
rect 7876 17834 7900 17836
rect 7956 17834 7980 17836
rect 8036 17834 8060 17836
rect 7898 17782 7900 17834
rect 7962 17782 7974 17834
rect 8036 17782 8038 17834
rect 7876 17780 7900 17782
rect 7956 17780 7980 17782
rect 8036 17780 8060 17782
rect 7820 17760 8116 17780
rect 8300 16848 8352 16854
rect 8300 16790 8352 16796
rect 7820 16748 8116 16768
rect 7876 16746 7900 16748
rect 7956 16746 7980 16748
rect 8036 16746 8060 16748
rect 7898 16694 7900 16746
rect 7962 16694 7974 16746
rect 8036 16694 8038 16746
rect 7876 16692 7900 16694
rect 7956 16692 7980 16694
rect 8036 16692 8060 16694
rect 7820 16672 8116 16692
rect 8312 16582 8340 16790
rect 8300 16576 8352 16582
rect 8300 16518 8352 16524
rect 8496 16514 8524 18626
rect 8588 18078 8616 21856
rect 9140 19166 9168 21856
rect 9128 19160 9180 19166
rect 9128 19102 9180 19108
rect 9692 19114 9720 21856
rect 10244 19794 10272 21856
rect 10152 19766 10272 19794
rect 9692 19086 9812 19114
rect 9680 19024 9732 19030
rect 9680 18966 9732 18972
rect 9692 18146 9720 18966
rect 9784 18214 9812 19086
rect 9956 19024 10008 19030
rect 9956 18966 10008 18972
rect 9968 18826 9996 18966
rect 10152 18826 10180 19766
rect 10232 19228 10284 19234
rect 10232 19170 10284 19176
rect 9956 18820 10008 18826
rect 9956 18762 10008 18768
rect 10140 18820 10192 18826
rect 10140 18762 10192 18768
rect 10244 18690 10272 19170
rect 10232 18684 10284 18690
rect 10232 18626 10284 18632
rect 9772 18208 9824 18214
rect 9772 18150 9824 18156
rect 9680 18140 9732 18146
rect 9680 18082 9732 18088
rect 8576 18072 8628 18078
rect 8576 18014 8628 18020
rect 10796 18026 10824 21856
rect 11348 19658 11376 21856
rect 11348 19630 11652 19658
rect 11252 19468 11548 19488
rect 11308 19466 11332 19468
rect 11388 19466 11412 19468
rect 11468 19466 11492 19468
rect 11330 19414 11332 19466
rect 11394 19414 11406 19466
rect 11468 19414 11470 19466
rect 11308 19412 11332 19414
rect 11388 19412 11412 19414
rect 11468 19412 11492 19414
rect 11252 19392 11548 19412
rect 11244 19160 11296 19166
rect 11244 19102 11296 19108
rect 11152 19024 11204 19030
rect 11152 18966 11204 18972
rect 11060 18072 11112 18078
rect 10796 17998 10916 18026
rect 11060 18014 11112 18020
rect 10784 17936 10836 17942
rect 10784 17878 10836 17884
rect 8760 17052 8812 17058
rect 8760 16994 8812 17000
rect 8772 16514 8800 16994
rect 9680 16848 9732 16854
rect 9680 16790 9732 16796
rect 10508 16848 10560 16854
rect 10508 16790 10560 16796
rect 10796 16802 10824 17878
rect 10888 17398 10916 17998
rect 10968 17936 11020 17942
rect 10968 17878 11020 17884
rect 10876 17392 10928 17398
rect 10876 17334 10928 17340
rect 10980 16922 11008 17878
rect 11072 16990 11100 18014
rect 11060 16984 11112 16990
rect 11060 16926 11112 16932
rect 10968 16916 11020 16922
rect 10968 16858 11020 16864
rect 8484 16508 8536 16514
rect 8484 16450 8536 16456
rect 8760 16508 8812 16514
rect 8760 16450 8812 16456
rect 8496 15970 8524 16450
rect 8852 16304 8904 16310
rect 8852 16246 8904 16252
rect 8484 15964 8536 15970
rect 8484 15906 8536 15912
rect 7748 15896 7800 15902
rect 7748 15838 7800 15844
rect 7820 15660 8116 15680
rect 7876 15658 7900 15660
rect 7956 15658 7980 15660
rect 8036 15658 8060 15660
rect 7898 15606 7900 15658
rect 7962 15606 7974 15658
rect 8036 15606 8038 15658
rect 7876 15604 7900 15606
rect 7956 15604 7980 15606
rect 8036 15604 8060 15606
rect 7820 15584 8116 15604
rect 8392 15012 8444 15018
rect 8392 14954 8444 14960
rect 7668 14870 7788 14898
rect 7656 14808 7708 14814
rect 7656 14750 7708 14756
rect 5460 14338 5672 14354
rect 4988 14332 5040 14338
rect 5460 14332 5684 14338
rect 5460 14326 5632 14332
rect 4988 14274 5040 14280
rect 5632 14274 5684 14280
rect 7012 14264 7064 14270
rect 7012 14206 7064 14212
rect 4896 14128 4948 14134
rect 4896 14070 4948 14076
rect 5080 14128 5132 14134
rect 5080 14070 5132 14076
rect 5264 14128 5316 14134
rect 5264 14070 5316 14076
rect 4388 14028 4684 14048
rect 4444 14026 4468 14028
rect 4524 14026 4548 14028
rect 4604 14026 4628 14028
rect 4466 13974 4468 14026
rect 4530 13974 4542 14026
rect 4604 13974 4606 14026
rect 4444 13972 4468 13974
rect 4524 13972 4548 13974
rect 4604 13972 4628 13974
rect 4388 13952 4684 13972
rect 3424 13924 3476 13930
rect 3424 13866 3476 13872
rect 4908 13726 4936 14070
rect 5092 13794 5120 14070
rect 5276 13930 5304 14070
rect 7024 13930 7052 14206
rect 7668 14202 7696 14750
rect 7656 14196 7708 14202
rect 7656 14138 7708 14144
rect 5264 13924 5316 13930
rect 5264 13866 5316 13872
rect 7012 13924 7064 13930
rect 7012 13866 7064 13872
rect 5080 13788 5132 13794
rect 5080 13730 5132 13736
rect 4896 13720 4948 13726
rect 4896 13662 4948 13668
rect 7196 13652 7248 13658
rect 7196 13594 7248 13600
rect 4988 13584 5040 13590
rect 4988 13526 5040 13532
rect 5000 13386 5028 13526
rect 4988 13380 5040 13386
rect 4988 13322 5040 13328
rect 4388 12940 4684 12960
rect 4444 12938 4468 12940
rect 4524 12938 4548 12940
rect 4604 12938 4628 12940
rect 4466 12886 4468 12938
rect 4530 12886 4542 12938
rect 4604 12886 4606 12938
rect 4444 12884 4468 12886
rect 4524 12884 4548 12886
rect 4604 12884 4628 12886
rect 4388 12864 4684 12884
rect 7208 11958 7236 13594
rect 7668 12298 7696 14138
rect 7656 12292 7708 12298
rect 7656 12234 7708 12240
rect 6828 11952 6880 11958
rect 6828 11894 6880 11900
rect 7196 11952 7248 11958
rect 7196 11894 7248 11900
rect 7564 11952 7616 11958
rect 7564 11894 7616 11900
rect 4388 11852 4684 11872
rect 4444 11850 4468 11852
rect 4524 11850 4548 11852
rect 4604 11850 4628 11852
rect 4466 11798 4468 11850
rect 4530 11798 4542 11850
rect 4604 11798 4606 11850
rect 4444 11796 4468 11798
rect 4524 11796 4548 11798
rect 4604 11796 4628 11798
rect 4388 11776 4684 11796
rect 6840 11074 6868 11894
rect 7576 11482 7604 11894
rect 7760 11482 7788 14870
rect 8116 14876 8168 14882
rect 8116 14818 8168 14824
rect 8128 14762 8156 14818
rect 8128 14734 8248 14762
rect 7820 14572 8116 14592
rect 7876 14570 7900 14572
rect 7956 14570 7980 14572
rect 8036 14570 8060 14572
rect 7898 14518 7900 14570
rect 7962 14518 7974 14570
rect 8036 14518 8038 14570
rect 7876 14516 7900 14518
rect 7956 14516 7980 14518
rect 8036 14516 8060 14518
rect 7820 14496 8116 14516
rect 8220 13590 8248 14734
rect 8300 14400 8352 14406
rect 8300 14342 8352 14348
rect 8312 13726 8340 14342
rect 8300 13720 8352 13726
rect 8300 13662 8352 13668
rect 8404 13658 8432 14954
rect 8668 14876 8720 14882
rect 8668 14818 8720 14824
rect 8680 14338 8708 14818
rect 8864 14338 8892 16246
rect 9496 14740 9548 14746
rect 9496 14682 9548 14688
rect 9404 14672 9456 14678
rect 9404 14614 9456 14620
rect 9416 14406 9444 14614
rect 9508 14474 9536 14682
rect 9496 14468 9548 14474
rect 9496 14410 9548 14416
rect 9404 14400 9456 14406
rect 9404 14342 9456 14348
rect 8668 14332 8720 14338
rect 8668 14274 8720 14280
rect 8852 14332 8904 14338
rect 8852 14274 8904 14280
rect 8680 13930 8708 14274
rect 8668 13924 8720 13930
rect 8668 13866 8720 13872
rect 8392 13652 8444 13658
rect 8392 13594 8444 13600
rect 8208 13584 8260 13590
rect 8208 13526 8260 13532
rect 7820 13484 8116 13504
rect 7876 13482 7900 13484
rect 7956 13482 7980 13484
rect 8036 13482 8060 13484
rect 7898 13430 7900 13482
rect 7962 13430 7974 13482
rect 8036 13430 8038 13482
rect 7876 13428 7900 13430
rect 7956 13428 7980 13430
rect 8036 13428 8060 13430
rect 7820 13408 8116 13428
rect 7820 12396 8116 12416
rect 7876 12394 7900 12396
rect 7956 12394 7980 12396
rect 8036 12394 8060 12396
rect 7898 12342 7900 12394
rect 7962 12342 7974 12394
rect 8036 12342 8038 12394
rect 7876 12340 7900 12342
rect 7956 12340 7980 12342
rect 8036 12340 8060 12342
rect 7820 12320 8116 12340
rect 8220 12162 8248 13526
rect 8300 12632 8352 12638
rect 8300 12574 8352 12580
rect 8208 12156 8260 12162
rect 8208 12098 8260 12104
rect 8312 12094 8340 12574
rect 9692 12502 9720 16790
rect 10520 16650 10548 16790
rect 10796 16774 11100 16802
rect 10508 16644 10560 16650
rect 10508 16586 10560 16592
rect 10048 16304 10100 16310
rect 10048 16246 10100 16252
rect 10060 15902 10088 16246
rect 10048 15896 10100 15902
rect 10048 15838 10100 15844
rect 10692 15896 10744 15902
rect 10692 15838 10744 15844
rect 11072 15850 11100 16774
rect 11164 15986 11192 18966
rect 11256 18554 11284 19102
rect 11520 19092 11572 19098
rect 11520 19034 11572 19040
rect 11532 18826 11560 19034
rect 11624 18826 11652 19630
rect 11520 18820 11572 18826
rect 11520 18762 11572 18768
rect 11612 18820 11664 18826
rect 11612 18762 11664 18768
rect 11532 18570 11560 18762
rect 11796 18616 11848 18622
rect 11244 18548 11296 18554
rect 11532 18542 11652 18570
rect 11796 18558 11848 18564
rect 11244 18490 11296 18496
rect 11252 18380 11548 18400
rect 11308 18378 11332 18380
rect 11388 18378 11412 18380
rect 11468 18378 11492 18380
rect 11330 18326 11332 18378
rect 11394 18326 11406 18378
rect 11468 18326 11470 18378
rect 11308 18324 11332 18326
rect 11388 18324 11412 18326
rect 11468 18324 11492 18326
rect 11252 18304 11548 18324
rect 11624 18146 11652 18542
rect 11704 18276 11756 18282
rect 11704 18218 11756 18224
rect 11612 18140 11664 18146
rect 11612 18082 11664 18088
rect 11716 17924 11744 18218
rect 11808 18078 11836 18558
rect 11796 18072 11848 18078
rect 11796 18014 11848 18020
rect 11716 17896 11836 17924
rect 11252 17292 11548 17312
rect 11308 17290 11332 17292
rect 11388 17290 11412 17292
rect 11468 17290 11492 17292
rect 11330 17238 11332 17290
rect 11394 17238 11406 17290
rect 11468 17238 11470 17290
rect 11308 17236 11332 17238
rect 11388 17236 11412 17238
rect 11468 17236 11492 17238
rect 11252 17216 11548 17236
rect 11704 16916 11756 16922
rect 11704 16858 11756 16864
rect 11716 16650 11744 16858
rect 11704 16644 11756 16650
rect 11704 16586 11756 16592
rect 11808 16446 11836 17896
rect 11796 16440 11848 16446
rect 11796 16382 11848 16388
rect 11888 16440 11940 16446
rect 11888 16382 11940 16388
rect 11252 16204 11548 16224
rect 11308 16202 11332 16204
rect 11388 16202 11412 16204
rect 11468 16202 11492 16204
rect 11330 16150 11332 16202
rect 11394 16150 11406 16202
rect 11468 16150 11470 16202
rect 11308 16148 11332 16150
rect 11388 16148 11412 16150
rect 11468 16148 11492 16150
rect 11252 16128 11548 16148
rect 11164 15958 11836 15986
rect 10704 14950 10732 15838
rect 11072 15822 11192 15850
rect 10692 14944 10744 14950
rect 10692 14886 10744 14892
rect 9772 14876 9824 14882
rect 9772 14818 9824 14824
rect 9784 14474 9812 14818
rect 10140 14672 10192 14678
rect 10140 14614 10192 14620
rect 10152 14474 10180 14614
rect 9772 14468 9824 14474
rect 9772 14410 9824 14416
rect 10140 14468 10192 14474
rect 10140 14410 10192 14416
rect 10704 13794 10732 14886
rect 10692 13788 10744 13794
rect 10692 13730 10744 13736
rect 10600 13720 10652 13726
rect 10600 13662 10652 13668
rect 10612 13386 10640 13662
rect 11060 13652 11112 13658
rect 11060 13594 11112 13600
rect 10600 13380 10652 13386
rect 10600 13322 10652 13328
rect 10968 13380 11020 13386
rect 10968 13322 11020 13328
rect 10980 12706 11008 13322
rect 11072 12842 11100 13594
rect 11164 13590 11192 15822
rect 11520 15828 11572 15834
rect 11520 15770 11572 15776
rect 11532 15714 11560 15770
rect 11532 15686 11652 15714
rect 11252 15116 11548 15136
rect 11308 15114 11332 15116
rect 11388 15114 11412 15116
rect 11468 15114 11492 15116
rect 11330 15062 11332 15114
rect 11394 15062 11406 15114
rect 11468 15062 11470 15114
rect 11308 15060 11332 15062
rect 11388 15060 11412 15062
rect 11468 15060 11492 15062
rect 11252 15040 11548 15060
rect 11252 14028 11548 14048
rect 11308 14026 11332 14028
rect 11388 14026 11412 14028
rect 11468 14026 11492 14028
rect 11330 13974 11332 14026
rect 11394 13974 11406 14026
rect 11468 13974 11470 14026
rect 11308 13972 11332 13974
rect 11388 13972 11412 13974
rect 11468 13972 11492 13974
rect 11252 13952 11548 13972
rect 11152 13584 11204 13590
rect 11152 13526 11204 13532
rect 11252 12940 11548 12960
rect 11308 12938 11332 12940
rect 11388 12938 11412 12940
rect 11468 12938 11492 12940
rect 11330 12886 11332 12938
rect 11394 12886 11406 12938
rect 11468 12886 11470 12938
rect 11308 12884 11332 12886
rect 11388 12884 11412 12886
rect 11468 12884 11492 12886
rect 11252 12864 11548 12884
rect 11060 12836 11112 12842
rect 11060 12778 11112 12784
rect 10968 12700 11020 12706
rect 10968 12642 11020 12648
rect 11152 12632 11204 12638
rect 11152 12574 11204 12580
rect 9864 12564 9916 12570
rect 9864 12506 9916 12512
rect 8484 12496 8536 12502
rect 8484 12438 8536 12444
rect 9680 12496 9732 12502
rect 9680 12438 9732 12444
rect 8392 12156 8444 12162
rect 8392 12098 8444 12104
rect 8300 12088 8352 12094
rect 8300 12030 8352 12036
rect 8404 11686 8432 12098
rect 8392 11680 8444 11686
rect 8392 11622 8444 11628
rect 7564 11476 7616 11482
rect 7564 11418 7616 11424
rect 7748 11476 7800 11482
rect 7748 11418 7800 11424
rect 6828 11068 6880 11074
rect 6828 11010 6880 11016
rect 4388 10764 4684 10784
rect 4444 10762 4468 10764
rect 4524 10762 4548 10764
rect 4604 10762 4628 10764
rect 4466 10710 4468 10762
rect 4530 10710 4542 10762
rect 4604 10710 4606 10762
rect 4444 10708 4468 10710
rect 4524 10708 4548 10710
rect 4604 10708 4628 10710
rect 4388 10688 4684 10708
rect 7576 10326 7604 11418
rect 8208 11408 8260 11414
rect 8208 11350 8260 11356
rect 7820 11308 8116 11328
rect 7876 11306 7900 11308
rect 7956 11306 7980 11308
rect 8036 11306 8060 11308
rect 7898 11254 7900 11306
rect 7962 11254 7974 11306
rect 8036 11254 8038 11306
rect 7876 11252 7900 11254
rect 7956 11252 7980 11254
rect 8036 11252 8060 11254
rect 7820 11232 8116 11252
rect 8220 11210 8248 11350
rect 8208 11204 8260 11210
rect 8208 11146 8260 11152
rect 8404 11006 8432 11622
rect 8496 11414 8524 12438
rect 9876 12026 9904 12506
rect 11164 12298 11192 12574
rect 11152 12292 11204 12298
rect 11152 12234 11204 12240
rect 10416 12224 10468 12230
rect 10416 12166 10468 12172
rect 10324 12156 10376 12162
rect 10324 12098 10376 12104
rect 9864 12020 9916 12026
rect 9864 11962 9916 11968
rect 8576 11952 8628 11958
rect 8576 11894 8628 11900
rect 8944 11952 8996 11958
rect 8944 11894 8996 11900
rect 8588 11618 8616 11894
rect 8576 11612 8628 11618
rect 8576 11554 8628 11560
rect 8484 11408 8536 11414
rect 8484 11350 8536 11356
rect 8392 11000 8444 11006
rect 8392 10942 8444 10948
rect 8588 10666 8616 11554
rect 8956 11482 8984 11894
rect 10336 11754 10364 12098
rect 10324 11748 10376 11754
rect 10324 11690 10376 11696
rect 8944 11476 8996 11482
rect 8944 11418 8996 11424
rect 10428 10938 10456 12166
rect 11252 11852 11548 11872
rect 11308 11850 11332 11852
rect 11388 11850 11412 11852
rect 11468 11850 11492 11852
rect 11330 11798 11332 11850
rect 11394 11798 11406 11850
rect 11468 11798 11470 11850
rect 11308 11796 11332 11798
rect 11388 11796 11412 11798
rect 11468 11796 11492 11798
rect 11252 11776 11548 11796
rect 10598 11512 10654 11521
rect 10598 11447 10654 11456
rect 10612 11414 10640 11447
rect 10600 11408 10652 11414
rect 10600 11350 10652 11356
rect 10416 10932 10468 10938
rect 10416 10874 10468 10880
rect 11252 10764 11548 10784
rect 11308 10762 11332 10764
rect 11388 10762 11412 10764
rect 11468 10762 11492 10764
rect 11330 10710 11332 10762
rect 11394 10710 11406 10762
rect 11468 10710 11470 10762
rect 11308 10708 11332 10710
rect 11388 10708 11412 10710
rect 11468 10708 11492 10710
rect 11252 10688 11548 10708
rect 8576 10660 8628 10666
rect 8576 10602 8628 10608
rect 11624 10462 11652 15686
rect 11704 13584 11756 13590
rect 11704 13526 11756 13532
rect 11612 10456 11664 10462
rect 11612 10398 11664 10404
rect 9864 10388 9916 10394
rect 9864 10330 9916 10336
rect 10416 10388 10468 10394
rect 10416 10330 10468 10336
rect 11244 10388 11296 10394
rect 11244 10330 11296 10336
rect 7564 10320 7616 10326
rect 7564 10262 7616 10268
rect 7576 9918 7604 10262
rect 7820 10220 8116 10240
rect 7876 10218 7900 10220
rect 7956 10218 7980 10220
rect 8036 10218 8060 10220
rect 7898 10166 7900 10218
rect 7962 10166 7974 10218
rect 8036 10166 8038 10218
rect 7876 10164 7900 10166
rect 7956 10164 7980 10166
rect 8036 10164 8060 10166
rect 7820 10144 8116 10164
rect 9876 10122 9904 10330
rect 9864 10116 9916 10122
rect 9864 10058 9916 10064
rect 8760 9980 8812 9986
rect 8760 9922 8812 9928
rect 7564 9912 7616 9918
rect 7564 9854 7616 9860
rect 4388 9676 4684 9696
rect 4444 9674 4468 9676
rect 4524 9674 4548 9676
rect 4604 9674 4628 9676
rect 4466 9622 4468 9674
rect 4530 9622 4542 9674
rect 4604 9622 4606 9674
rect 4444 9620 4468 9622
rect 4524 9620 4548 9622
rect 4604 9620 4628 9622
rect 4388 9600 4684 9620
rect 7576 9374 7604 9854
rect 8772 9510 8800 9922
rect 8760 9504 8812 9510
rect 8760 9446 8812 9452
rect 7564 9368 7616 9374
rect 7564 9310 7616 9316
rect 2688 8960 2740 8966
rect 2688 8902 2740 8908
rect 4388 8588 4684 8608
rect 4444 8586 4468 8588
rect 4524 8586 4548 8588
rect 4604 8586 4628 8588
rect 4466 8534 4468 8586
rect 4530 8534 4542 8586
rect 4604 8534 4606 8586
rect 4444 8532 4468 8534
rect 4524 8532 4548 8534
rect 4604 8532 4628 8534
rect 4388 8512 4684 8532
rect 4388 7500 4684 7520
rect 4444 7498 4468 7500
rect 4524 7498 4548 7500
rect 4604 7498 4628 7500
rect 4466 7446 4468 7498
rect 4530 7446 4542 7498
rect 4604 7446 4606 7498
rect 4444 7444 4468 7446
rect 4524 7444 4548 7446
rect 4604 7444 4628 7446
rect 4388 7424 4684 7444
rect 2964 6716 3016 6722
rect 2964 6658 3016 6664
rect 2976 5673 3004 6658
rect 7576 6518 7604 9310
rect 7820 9132 8116 9152
rect 7876 9130 7900 9132
rect 7956 9130 7980 9132
rect 8036 9130 8060 9132
rect 7898 9078 7900 9130
rect 7962 9078 7974 9130
rect 8036 9078 8038 9130
rect 7876 9076 7900 9078
rect 7956 9076 7980 9078
rect 8036 9076 8060 9078
rect 7820 9056 8116 9076
rect 10428 9034 10456 10330
rect 10508 10320 10560 10326
rect 10508 10262 10560 10268
rect 10520 9578 10548 10262
rect 11256 10122 11284 10330
rect 11624 10122 11652 10398
rect 11244 10116 11296 10122
rect 11244 10058 11296 10064
rect 11612 10116 11664 10122
rect 11612 10058 11664 10064
rect 11612 9912 11664 9918
rect 11612 9854 11664 9860
rect 10876 9776 10928 9782
rect 10876 9718 10928 9724
rect 10508 9572 10560 9578
rect 10508 9514 10560 9520
rect 10600 9436 10652 9442
rect 10600 9378 10652 9384
rect 10416 9028 10468 9034
rect 10416 8970 10468 8976
rect 10612 8830 10640 9378
rect 10888 9374 10916 9718
rect 11252 9676 11548 9696
rect 11308 9674 11332 9676
rect 11388 9674 11412 9676
rect 11468 9674 11492 9676
rect 11330 9622 11332 9674
rect 11394 9622 11406 9674
rect 11468 9622 11470 9674
rect 11308 9620 11332 9622
rect 11388 9620 11412 9622
rect 11468 9620 11492 9622
rect 11252 9600 11548 9620
rect 11624 9442 11652 9854
rect 11612 9436 11664 9442
rect 11612 9378 11664 9384
rect 10876 9368 10928 9374
rect 10876 9310 10928 9316
rect 11428 9232 11480 9238
rect 11428 9174 11480 9180
rect 11440 8966 11468 9174
rect 11428 8960 11480 8966
rect 11428 8902 11480 8908
rect 10600 8824 10652 8830
rect 10600 8766 10652 8772
rect 11252 8588 11548 8608
rect 11308 8586 11332 8588
rect 11388 8586 11412 8588
rect 11468 8586 11492 8588
rect 11330 8534 11332 8586
rect 11394 8534 11406 8586
rect 11468 8534 11470 8586
rect 11308 8532 11332 8534
rect 11388 8532 11412 8534
rect 11468 8532 11492 8534
rect 11252 8512 11548 8532
rect 11336 8280 11388 8286
rect 11336 8222 11388 8228
rect 7820 8044 8116 8064
rect 7876 8042 7900 8044
rect 7956 8042 7980 8044
rect 8036 8042 8060 8044
rect 7898 7990 7900 8042
rect 7962 7990 7974 8042
rect 8036 7990 8038 8042
rect 7876 7988 7900 7990
rect 7956 7988 7980 7990
rect 8036 7988 8060 7990
rect 7820 7968 8116 7988
rect 11348 7878 11376 8222
rect 11336 7872 11388 7878
rect 11336 7814 11388 7820
rect 10324 7804 10376 7810
rect 10324 7746 10376 7752
rect 10336 7402 10364 7746
rect 11252 7500 11548 7520
rect 11308 7498 11332 7500
rect 11388 7498 11412 7500
rect 11468 7498 11492 7500
rect 11330 7446 11332 7498
rect 11394 7446 11406 7498
rect 11468 7446 11470 7498
rect 11308 7444 11332 7446
rect 11388 7444 11412 7446
rect 11468 7444 11492 7446
rect 11252 7424 11548 7444
rect 10324 7396 10376 7402
rect 10324 7338 10376 7344
rect 10600 7260 10652 7266
rect 10600 7202 10652 7208
rect 7820 6956 8116 6976
rect 7876 6954 7900 6956
rect 7956 6954 7980 6956
rect 8036 6954 8060 6956
rect 7898 6902 7900 6954
rect 7962 6902 7974 6954
rect 8036 6902 8038 6954
rect 7876 6900 7900 6902
rect 7956 6900 7980 6902
rect 8036 6900 8060 6902
rect 7820 6880 8116 6900
rect 10612 6858 10640 7202
rect 10784 7056 10836 7062
rect 10784 6998 10836 7004
rect 10796 6858 10824 6998
rect 10600 6852 10652 6858
rect 10600 6794 10652 6800
rect 10784 6852 10836 6858
rect 10784 6794 10836 6800
rect 11716 6722 11744 13526
rect 11808 10394 11836 15958
rect 11900 15902 11928 16382
rect 11888 15896 11940 15902
rect 11888 15838 11940 15844
rect 11888 14332 11940 14338
rect 11888 14274 11940 14280
rect 11900 13726 11928 14274
rect 11888 13720 11940 13726
rect 11888 13662 11940 13668
rect 11796 10388 11848 10394
rect 11796 10330 11848 10336
rect 11992 8490 12020 21856
rect 12256 18820 12308 18826
rect 12256 18762 12308 18768
rect 12072 13924 12124 13930
rect 12072 13866 12124 13872
rect 12084 13182 12112 13866
rect 12072 13176 12124 13182
rect 12072 13118 12124 13124
rect 12268 11210 12296 18762
rect 12348 18480 12400 18486
rect 12348 18422 12400 18428
rect 12360 17602 12388 18422
rect 12348 17596 12400 17602
rect 12348 17538 12400 17544
rect 12440 16848 12492 16854
rect 12440 16790 12492 16796
rect 12452 16378 12480 16790
rect 12440 16372 12492 16378
rect 12440 16314 12492 16320
rect 12440 14808 12492 14814
rect 12440 14750 12492 14756
rect 12452 12842 12480 14750
rect 12440 12836 12492 12842
rect 12440 12778 12492 12784
rect 12452 12706 12480 12778
rect 12440 12700 12492 12706
rect 12440 12642 12492 12648
rect 12256 11204 12308 11210
rect 12256 11146 12308 11152
rect 12348 9300 12400 9306
rect 12348 9242 12400 9248
rect 12072 9232 12124 9238
rect 12072 9174 12124 9180
rect 12084 9034 12112 9174
rect 12072 9028 12124 9034
rect 12072 8970 12124 8976
rect 12360 8830 12388 9242
rect 12440 9232 12492 9238
rect 12440 9174 12492 9180
rect 12452 8966 12480 9174
rect 12440 8960 12492 8966
rect 12440 8902 12492 8908
rect 12348 8824 12400 8830
rect 12348 8766 12400 8772
rect 11980 8484 12032 8490
rect 11980 8426 12032 8432
rect 11704 6716 11756 6722
rect 11704 6658 11756 6664
rect 11716 6586 11744 6658
rect 11704 6580 11756 6586
rect 11704 6522 11756 6528
rect 7564 6512 7616 6518
rect 7564 6454 7616 6460
rect 4388 6412 4684 6432
rect 4444 6410 4468 6412
rect 4524 6410 4548 6412
rect 4604 6410 4628 6412
rect 4466 6358 4468 6410
rect 4530 6358 4542 6410
rect 4604 6358 4606 6410
rect 4444 6356 4468 6358
rect 4524 6356 4548 6358
rect 4604 6356 4628 6358
rect 4388 6336 4684 6356
rect 11252 6412 11548 6432
rect 11308 6410 11332 6412
rect 11388 6410 11412 6412
rect 11468 6410 11492 6412
rect 11330 6358 11332 6410
rect 11394 6358 11406 6410
rect 11468 6358 11470 6410
rect 11308 6356 11332 6358
rect 11388 6356 11412 6358
rect 11468 6356 11492 6358
rect 11252 6336 11548 6356
rect 7820 5868 8116 5888
rect 7876 5866 7900 5868
rect 7956 5866 7980 5868
rect 8036 5866 8060 5868
rect 7898 5814 7900 5866
rect 7962 5814 7974 5866
rect 8036 5814 8038 5866
rect 7876 5812 7900 5814
rect 7956 5812 7980 5814
rect 8036 5812 8060 5814
rect 7820 5792 8116 5812
rect 12544 5770 12572 21856
rect 12624 19024 12676 19030
rect 12624 18966 12676 18972
rect 12636 18758 12664 18966
rect 12624 18752 12676 18758
rect 12624 18694 12676 18700
rect 12636 18146 12664 18694
rect 12716 18208 12768 18214
rect 12716 18150 12768 18156
rect 12624 18140 12676 18146
rect 12624 18082 12676 18088
rect 12728 17602 12756 18150
rect 12716 17596 12768 17602
rect 12716 17538 12768 17544
rect 12992 16440 13044 16446
rect 12992 16382 13044 16388
rect 13004 16106 13032 16382
rect 12992 16100 13044 16106
rect 12992 16042 13044 16048
rect 12992 14264 13044 14270
rect 12992 14206 13044 14212
rect 12808 14128 12860 14134
rect 12808 14070 12860 14076
rect 12820 13386 12848 14070
rect 12900 13924 12952 13930
rect 12900 13866 12952 13872
rect 12912 13386 12940 13866
rect 13004 13794 13032 14206
rect 12992 13788 13044 13794
rect 12992 13730 13044 13736
rect 12808 13380 12860 13386
rect 12808 13322 12860 13328
rect 12900 13380 12952 13386
rect 12900 13322 12952 13328
rect 12992 12156 13044 12162
rect 12992 12098 13044 12104
rect 12624 12020 12676 12026
rect 12624 11962 12676 11968
rect 12636 11550 12664 11962
rect 13004 11686 13032 12098
rect 12992 11680 13044 11686
rect 12992 11622 13044 11628
rect 12624 11544 12676 11550
rect 12624 11486 12676 11492
rect 12808 11476 12860 11482
rect 12808 11418 12860 11424
rect 12820 9986 12848 11418
rect 12992 11408 13044 11414
rect 12992 11350 13044 11356
rect 13004 11006 13032 11350
rect 12992 11000 13044 11006
rect 12992 10942 13044 10948
rect 12808 9980 12860 9986
rect 12808 9922 12860 9928
rect 13096 9034 13124 21856
rect 13268 18480 13320 18486
rect 13268 18422 13320 18428
rect 13280 15902 13308 18422
rect 13360 16984 13412 16990
rect 13360 16926 13412 16932
rect 13372 16650 13400 16926
rect 13360 16644 13412 16650
rect 13360 16586 13412 16592
rect 13268 15896 13320 15902
rect 13268 15838 13320 15844
rect 13280 14950 13308 15838
rect 13268 14944 13320 14950
rect 13268 14886 13320 14892
rect 13280 14474 13308 14886
rect 13268 14468 13320 14474
rect 13268 14410 13320 14416
rect 13280 14270 13308 14410
rect 13360 14332 13412 14338
rect 13360 14274 13412 14280
rect 13268 14264 13320 14270
rect 13268 14206 13320 14212
rect 13372 13794 13400 14274
rect 13360 13788 13412 13794
rect 13360 13730 13412 13736
rect 13360 12700 13412 12706
rect 13360 12642 13412 12648
rect 13176 12088 13228 12094
rect 13176 12030 13228 12036
rect 13188 11142 13216 12030
rect 13372 11414 13400 12642
rect 13452 12496 13504 12502
rect 13452 12438 13504 12444
rect 13464 12298 13492 12438
rect 13452 12292 13504 12298
rect 13452 12234 13504 12240
rect 13360 11408 13412 11414
rect 13360 11350 13412 11356
rect 13176 11136 13228 11142
rect 13176 11078 13228 11084
rect 13372 10938 13400 11350
rect 13360 10932 13412 10938
rect 13360 10874 13412 10880
rect 13372 10054 13400 10874
rect 13648 10138 13676 21856
rect 13912 19024 13964 19030
rect 13912 18966 13964 18972
rect 14096 19024 14148 19030
rect 14096 18966 14148 18972
rect 13924 18146 13952 18966
rect 14108 18282 14136 18966
rect 14096 18276 14148 18282
rect 14096 18218 14148 18224
rect 13912 18140 13964 18146
rect 13912 18082 13964 18088
rect 14200 17942 14228 21856
rect 14752 20202 14780 21856
rect 14384 20174 14780 20202
rect 14280 19228 14332 19234
rect 14280 19170 14332 19176
rect 14292 18758 14320 19170
rect 14280 18752 14332 18758
rect 14280 18694 14332 18700
rect 14188 17936 14240 17942
rect 14188 17878 14240 17884
rect 14280 16508 14332 16514
rect 14280 16450 14332 16456
rect 13912 16304 13964 16310
rect 13912 16246 13964 16252
rect 13924 15494 13952 16246
rect 14292 15834 14320 16450
rect 14280 15828 14332 15834
rect 14280 15770 14332 15776
rect 13912 15488 13964 15494
rect 13912 15430 13964 15436
rect 14096 12836 14148 12842
rect 14096 12778 14148 12784
rect 14004 12564 14056 12570
rect 14004 12506 14056 12512
rect 14016 12298 14044 12506
rect 14004 12292 14056 12298
rect 14004 12234 14056 12240
rect 13728 12088 13780 12094
rect 13728 12030 13780 12036
rect 13740 11958 13768 12030
rect 13728 11952 13780 11958
rect 13728 11894 13780 11900
rect 13740 11482 13768 11894
rect 14108 11550 14136 12778
rect 14188 12632 14240 12638
rect 14188 12574 14240 12580
rect 14200 12162 14228 12574
rect 14188 12156 14240 12162
rect 14188 12098 14240 12104
rect 14188 11612 14240 11618
rect 14188 11554 14240 11560
rect 14096 11544 14148 11550
rect 14096 11486 14148 11492
rect 13728 11476 13780 11482
rect 13728 11418 13780 11424
rect 14004 11408 14056 11414
rect 14004 11350 14056 11356
rect 14016 11210 14044 11350
rect 14004 11204 14056 11210
rect 14004 11146 14056 11152
rect 14096 11204 14148 11210
rect 14096 11146 14148 11152
rect 14108 11006 14136 11146
rect 14096 11000 14148 11006
rect 14096 10942 14148 10948
rect 13648 10110 13768 10138
rect 13360 10048 13412 10054
rect 13360 9990 13412 9996
rect 13636 9980 13688 9986
rect 13636 9922 13688 9928
rect 13648 9374 13676 9922
rect 13636 9368 13688 9374
rect 13636 9310 13688 9316
rect 13084 9028 13136 9034
rect 13084 8970 13136 8976
rect 13452 8892 13504 8898
rect 13452 8834 13504 8840
rect 13464 8354 13492 8834
rect 13452 8348 13504 8354
rect 13452 8290 13504 8296
rect 13268 8280 13320 8286
rect 13268 8222 13320 8228
rect 13280 7946 13308 8222
rect 13268 7940 13320 7946
rect 13268 7882 13320 7888
rect 13648 7402 13676 9310
rect 13636 7396 13688 7402
rect 13636 7338 13688 7344
rect 13740 6518 13768 10110
rect 14108 9220 14136 10942
rect 14200 10122 14228 11554
rect 14292 11210 14320 15770
rect 14280 11204 14332 11210
rect 14280 11146 14332 11152
rect 14188 10116 14240 10122
rect 14188 10058 14240 10064
rect 14200 9374 14228 10058
rect 14188 9368 14240 9374
rect 14188 9310 14240 9316
rect 14108 9192 14228 9220
rect 14096 7736 14148 7742
rect 14096 7678 14148 7684
rect 14108 6858 14136 7678
rect 14096 6852 14148 6858
rect 14096 6794 14148 6800
rect 13728 6512 13780 6518
rect 13728 6454 13780 6460
rect 12532 5764 12584 5770
rect 12532 5706 12584 5712
rect 2962 5664 3018 5673
rect 2962 5599 3018 5608
rect 4388 5324 4684 5344
rect 4444 5322 4468 5324
rect 4524 5322 4548 5324
rect 4604 5322 4628 5324
rect 4466 5270 4468 5322
rect 4530 5270 4542 5322
rect 4604 5270 4606 5322
rect 4444 5268 4468 5270
rect 4524 5268 4548 5270
rect 4604 5268 4628 5270
rect 4388 5248 4684 5268
rect 11252 5324 11548 5344
rect 11308 5322 11332 5324
rect 11388 5322 11412 5324
rect 11468 5322 11492 5324
rect 11330 5270 11332 5322
rect 11394 5270 11406 5322
rect 11468 5270 11470 5322
rect 11308 5268 11332 5270
rect 11388 5268 11412 5270
rect 11468 5268 11492 5270
rect 11252 5248 11548 5268
rect 7820 4780 8116 4800
rect 7876 4778 7900 4780
rect 7956 4778 7980 4780
rect 8036 4778 8060 4780
rect 7898 4726 7900 4778
rect 7962 4726 7974 4778
rect 8036 4726 8038 4778
rect 7876 4724 7900 4726
rect 7956 4724 7980 4726
rect 8036 4724 8060 4726
rect 7820 4704 8116 4724
rect 4388 4236 4684 4256
rect 4444 4234 4468 4236
rect 4524 4234 4548 4236
rect 4604 4234 4628 4236
rect 4466 4182 4468 4234
rect 4530 4182 4542 4234
rect 4604 4182 4606 4234
rect 4444 4180 4468 4182
rect 4524 4180 4548 4182
rect 4604 4180 4628 4182
rect 4388 4160 4684 4180
rect 11252 4236 11548 4256
rect 11308 4234 11332 4236
rect 11388 4234 11412 4236
rect 11468 4234 11492 4236
rect 11330 4182 11332 4234
rect 11394 4182 11406 4234
rect 11468 4182 11470 4234
rect 11308 4180 11332 4182
rect 11388 4180 11412 4182
rect 11468 4180 11492 4182
rect 11252 4160 11548 4180
rect 14200 4002 14228 9192
rect 14384 7878 14412 20174
rect 14684 20012 14980 20032
rect 14740 20010 14764 20012
rect 14820 20010 14844 20012
rect 14900 20010 14924 20012
rect 14762 19958 14764 20010
rect 14826 19958 14838 20010
rect 14900 19958 14902 20010
rect 14740 19956 14764 19958
rect 14820 19956 14844 19958
rect 14900 19956 14924 19958
rect 14684 19936 14980 19956
rect 15016 19092 15068 19098
rect 15016 19034 15068 19040
rect 14684 18924 14980 18944
rect 14740 18922 14764 18924
rect 14820 18922 14844 18924
rect 14900 18922 14924 18924
rect 14762 18870 14764 18922
rect 14826 18870 14838 18922
rect 14900 18870 14902 18922
rect 14740 18868 14764 18870
rect 14820 18868 14844 18870
rect 14900 18868 14924 18870
rect 14684 18848 14980 18868
rect 15028 18826 15056 19034
rect 15016 18820 15068 18826
rect 15016 18762 15068 18768
rect 15304 17942 15332 21856
rect 15660 19024 15712 19030
rect 15660 18966 15712 18972
rect 15752 19024 15804 19030
rect 15752 18966 15804 18972
rect 15108 17936 15160 17942
rect 15108 17878 15160 17884
rect 15292 17936 15344 17942
rect 15292 17878 15344 17884
rect 14684 17836 14980 17856
rect 14740 17834 14764 17836
rect 14820 17834 14844 17836
rect 14900 17834 14924 17836
rect 14762 17782 14764 17834
rect 14826 17782 14838 17834
rect 14900 17782 14902 17834
rect 14740 17780 14764 17782
rect 14820 17780 14844 17782
rect 14900 17780 14924 17782
rect 14684 17760 14980 17780
rect 14684 16748 14980 16768
rect 14740 16746 14764 16748
rect 14820 16746 14844 16748
rect 14900 16746 14924 16748
rect 14762 16694 14764 16746
rect 14826 16694 14838 16746
rect 14900 16694 14902 16746
rect 14740 16692 14764 16694
rect 14820 16692 14844 16694
rect 14900 16692 14924 16694
rect 14684 16672 14980 16692
rect 14464 16440 14516 16446
rect 14464 16382 14516 16388
rect 14476 15766 14504 16382
rect 14464 15760 14516 15766
rect 14464 15702 14516 15708
rect 14476 14338 14504 15702
rect 14684 15660 14980 15680
rect 14740 15658 14764 15660
rect 14820 15658 14844 15660
rect 14900 15658 14924 15660
rect 14762 15606 14764 15658
rect 14826 15606 14838 15658
rect 14900 15606 14902 15658
rect 14740 15604 14764 15606
rect 14820 15604 14844 15606
rect 14900 15604 14924 15606
rect 14684 15584 14980 15604
rect 15016 15352 15068 15358
rect 15016 15294 15068 15300
rect 14556 14808 14608 14814
rect 14556 14750 14608 14756
rect 14568 14474 14596 14750
rect 14684 14572 14980 14592
rect 14740 14570 14764 14572
rect 14820 14570 14844 14572
rect 14900 14570 14924 14572
rect 14762 14518 14764 14570
rect 14826 14518 14838 14570
rect 14900 14518 14902 14570
rect 14740 14516 14764 14518
rect 14820 14516 14844 14518
rect 14900 14516 14924 14518
rect 14684 14496 14980 14516
rect 15028 14474 15056 15294
rect 14556 14468 14608 14474
rect 14556 14410 14608 14416
rect 15016 14468 15068 14474
rect 15016 14410 15068 14416
rect 14464 14332 14516 14338
rect 14464 14274 14516 14280
rect 14684 13484 14980 13504
rect 14740 13482 14764 13484
rect 14820 13482 14844 13484
rect 14900 13482 14924 13484
rect 14762 13430 14764 13482
rect 14826 13430 14838 13482
rect 14900 13430 14902 13482
rect 14740 13428 14764 13430
rect 14820 13428 14844 13430
rect 14900 13428 14924 13430
rect 14684 13408 14980 13428
rect 14464 12632 14516 12638
rect 14464 12574 14516 12580
rect 14476 11754 14504 12574
rect 14684 12396 14980 12416
rect 14740 12394 14764 12396
rect 14820 12394 14844 12396
rect 14900 12394 14924 12396
rect 14762 12342 14764 12394
rect 14826 12342 14838 12394
rect 14900 12342 14902 12394
rect 14740 12340 14764 12342
rect 14820 12340 14844 12342
rect 14900 12340 14924 12342
rect 14684 12320 14980 12340
rect 14556 12224 14608 12230
rect 14556 12166 14608 12172
rect 14464 11748 14516 11754
rect 14464 11690 14516 11696
rect 14568 11521 14596 12166
rect 14554 11512 14610 11521
rect 14554 11447 14610 11456
rect 14684 11308 14980 11328
rect 14740 11306 14764 11308
rect 14820 11306 14844 11308
rect 14900 11306 14924 11308
rect 14762 11254 14764 11306
rect 14826 11254 14838 11306
rect 14900 11254 14902 11306
rect 14740 11252 14764 11254
rect 14820 11252 14844 11254
rect 14900 11252 14924 11254
rect 14684 11232 14980 11252
rect 14684 10220 14980 10240
rect 14740 10218 14764 10220
rect 14820 10218 14844 10220
rect 14900 10218 14924 10220
rect 14762 10166 14764 10218
rect 14826 10166 14838 10218
rect 14900 10166 14902 10218
rect 14740 10164 14764 10166
rect 14820 10164 14844 10166
rect 14900 10164 14924 10166
rect 14684 10144 14980 10164
rect 14684 9132 14980 9152
rect 14740 9130 14764 9132
rect 14820 9130 14844 9132
rect 14900 9130 14924 9132
rect 14762 9078 14764 9130
rect 14826 9078 14838 9130
rect 14900 9078 14902 9130
rect 14740 9076 14764 9078
rect 14820 9076 14844 9078
rect 14900 9076 14924 9078
rect 14684 9056 14980 9076
rect 15120 9034 15148 17878
rect 15476 16984 15528 16990
rect 15476 16926 15528 16932
rect 15488 16446 15516 16926
rect 15672 16922 15700 18966
rect 15764 18690 15792 18966
rect 15856 18690 15884 21856
rect 16120 19228 16172 19234
rect 16120 19170 16172 19176
rect 16132 18758 16160 19170
rect 16304 19024 16356 19030
rect 16304 18966 16356 18972
rect 16120 18752 16172 18758
rect 16120 18694 16172 18700
rect 15752 18684 15804 18690
rect 15752 18626 15804 18632
rect 15844 18684 15896 18690
rect 15844 18626 15896 18632
rect 16132 18486 16160 18694
rect 16120 18480 16172 18486
rect 16120 18422 16172 18428
rect 16316 18078 16344 18966
rect 16304 18072 16356 18078
rect 16304 18014 16356 18020
rect 16212 17936 16264 17942
rect 16212 17878 16264 17884
rect 15660 16916 15712 16922
rect 15660 16858 15712 16864
rect 15476 16440 15528 16446
rect 15476 16382 15528 16388
rect 15292 15760 15344 15766
rect 15292 15702 15344 15708
rect 15304 15562 15332 15702
rect 15292 15556 15344 15562
rect 15292 15498 15344 15504
rect 15488 14814 15516 16382
rect 15476 14808 15528 14814
rect 15476 14750 15528 14756
rect 15568 13176 15620 13182
rect 15568 13118 15620 13124
rect 15580 12706 15608 13118
rect 15568 12700 15620 12706
rect 15568 12642 15620 12648
rect 15672 10938 15700 16858
rect 16120 13652 16172 13658
rect 16120 13594 16172 13600
rect 16132 11074 16160 13594
rect 16120 11068 16172 11074
rect 16120 11010 16172 11016
rect 15660 10932 15712 10938
rect 15660 10874 15712 10880
rect 15936 10932 15988 10938
rect 15936 10874 15988 10880
rect 15108 9028 15160 9034
rect 15108 8970 15160 8976
rect 15660 8892 15712 8898
rect 15660 8834 15712 8840
rect 15672 8354 15700 8834
rect 15948 8830 15976 10874
rect 16132 9510 16160 11010
rect 16120 9504 16172 9510
rect 16120 9446 16172 9452
rect 15936 8824 15988 8830
rect 15936 8766 15988 8772
rect 15660 8348 15712 8354
rect 15660 8290 15712 8296
rect 14684 8044 14980 8064
rect 14740 8042 14764 8044
rect 14820 8042 14844 8044
rect 14900 8042 14924 8044
rect 14762 7990 14764 8042
rect 14826 7990 14838 8042
rect 14900 7990 14902 8042
rect 14740 7988 14764 7990
rect 14820 7988 14844 7990
rect 14900 7988 14924 7990
rect 14684 7968 14980 7988
rect 14372 7872 14424 7878
rect 14372 7814 14424 7820
rect 14648 7804 14700 7810
rect 14648 7746 14700 7752
rect 14280 7736 14332 7742
rect 14280 7678 14332 7684
rect 14292 7130 14320 7678
rect 14660 7266 14688 7746
rect 14648 7260 14700 7266
rect 14648 7202 14700 7208
rect 14556 7192 14608 7198
rect 14556 7134 14608 7140
rect 14280 7124 14332 7130
rect 14280 7066 14332 7072
rect 14568 6654 14596 7134
rect 14684 6956 14980 6976
rect 14740 6954 14764 6956
rect 14820 6954 14844 6956
rect 14900 6954 14924 6956
rect 14762 6902 14764 6954
rect 14826 6902 14838 6954
rect 14900 6902 14902 6954
rect 14740 6900 14764 6902
rect 14820 6900 14844 6902
rect 14900 6900 14924 6902
rect 14684 6880 14980 6900
rect 15200 6784 15252 6790
rect 15200 6726 15252 6732
rect 14556 6648 14608 6654
rect 14556 6590 14608 6596
rect 15212 6314 15240 6726
rect 15200 6308 15252 6314
rect 15200 6250 15252 6256
rect 14684 5868 14980 5888
rect 14740 5866 14764 5868
rect 14820 5866 14844 5868
rect 14900 5866 14924 5868
rect 14762 5814 14764 5866
rect 14826 5814 14838 5866
rect 14900 5814 14902 5866
rect 14740 5812 14764 5814
rect 14820 5812 14844 5814
rect 14900 5812 14924 5814
rect 14684 5792 14980 5812
rect 14684 4780 14980 4800
rect 14740 4778 14764 4780
rect 14820 4778 14844 4780
rect 14900 4778 14924 4780
rect 14762 4726 14764 4778
rect 14826 4726 14838 4778
rect 14900 4726 14902 4778
rect 14740 4724 14764 4726
rect 14820 4724 14844 4726
rect 14900 4724 14924 4726
rect 14684 4704 14980 4724
rect 14188 3996 14240 4002
rect 14188 3938 14240 3944
rect 15948 3934 15976 8766
rect 16028 7736 16080 7742
rect 16028 7678 16080 7684
rect 16040 7402 16068 7678
rect 16224 7606 16252 17878
rect 16408 11192 16436 21856
rect 16672 19024 16724 19030
rect 16672 18966 16724 18972
rect 16684 18826 16712 18966
rect 16672 18820 16724 18826
rect 16672 18762 16724 18768
rect 16960 17942 16988 21856
rect 17316 19228 17368 19234
rect 17316 19170 17368 19176
rect 17328 18486 17356 19170
rect 17408 19160 17460 19166
rect 17408 19102 17460 19108
rect 17316 18480 17368 18486
rect 17316 18422 17368 18428
rect 17224 18208 17276 18214
rect 17224 18150 17276 18156
rect 16948 17936 17000 17942
rect 16948 17878 17000 17884
rect 16672 17392 16724 17398
rect 16672 17334 16724 17340
rect 16684 15766 16712 17334
rect 16856 16916 16908 16922
rect 16856 16858 16908 16864
rect 16868 16650 16896 16858
rect 16856 16644 16908 16650
rect 16856 16586 16908 16592
rect 16868 15970 16896 16586
rect 16856 15964 16908 15970
rect 16856 15906 16908 15912
rect 16672 15760 16724 15766
rect 16672 15702 16724 15708
rect 16488 14672 16540 14678
rect 16488 14614 16540 14620
rect 16500 14474 16528 14614
rect 16488 14468 16540 14474
rect 16488 14410 16540 14416
rect 17236 14338 17264 18150
rect 17328 16514 17356 18422
rect 17420 18146 17448 19102
rect 17512 18486 17540 21856
rect 17866 21440 17922 21449
rect 17866 21375 17922 21384
rect 17880 19030 17908 21375
rect 17972 19166 18000 22327
rect 18050 21856 18106 22656
rect 18602 21856 18658 22656
rect 18694 21984 18750 21993
rect 18694 21919 18750 21928
rect 18064 19658 18092 21856
rect 18064 19630 18552 19658
rect 18116 19468 18412 19488
rect 18172 19466 18196 19468
rect 18252 19466 18276 19468
rect 18332 19466 18356 19468
rect 18194 19414 18196 19466
rect 18258 19414 18270 19466
rect 18332 19414 18334 19466
rect 18172 19412 18196 19414
rect 18252 19412 18276 19414
rect 18332 19412 18356 19414
rect 18116 19392 18412 19412
rect 17960 19160 18012 19166
rect 17960 19102 18012 19108
rect 17868 19024 17920 19030
rect 17868 18966 17920 18972
rect 17500 18480 17552 18486
rect 17500 18422 17552 18428
rect 18116 18380 18412 18400
rect 18172 18378 18196 18380
rect 18252 18378 18276 18380
rect 18332 18378 18356 18380
rect 18194 18326 18196 18378
rect 18258 18326 18270 18378
rect 18332 18326 18334 18378
rect 18172 18324 18196 18326
rect 18252 18324 18276 18326
rect 18332 18324 18356 18326
rect 18116 18304 18412 18324
rect 18524 18214 18552 19630
rect 18512 18208 18564 18214
rect 18512 18150 18564 18156
rect 17408 18140 17460 18146
rect 17408 18082 17460 18088
rect 18512 18072 18564 18078
rect 18512 18014 18564 18020
rect 18524 17670 18552 18014
rect 18512 17664 18564 17670
rect 18512 17606 18564 17612
rect 17960 17596 18012 17602
rect 17960 17538 18012 17544
rect 17684 17188 17736 17194
rect 17684 17130 17736 17136
rect 17316 16508 17368 16514
rect 17316 16450 17368 16456
rect 17696 15902 17724 17130
rect 17972 16530 18000 17538
rect 18116 17292 18412 17312
rect 18172 17290 18196 17292
rect 18252 17290 18276 17292
rect 18332 17290 18356 17292
rect 18194 17238 18196 17290
rect 18258 17238 18270 17290
rect 18332 17238 18334 17290
rect 18172 17236 18196 17238
rect 18252 17236 18276 17238
rect 18332 17236 18356 17238
rect 18116 17216 18412 17236
rect 18512 16984 18564 16990
rect 18512 16926 18564 16932
rect 18524 16650 18552 16926
rect 18512 16644 18564 16650
rect 18512 16586 18564 16592
rect 17880 16502 18000 16530
rect 17880 16106 17908 16502
rect 17960 16440 18012 16446
rect 17960 16382 18012 16388
rect 17868 16100 17920 16106
rect 17868 16042 17920 16048
rect 17684 15896 17736 15902
rect 17684 15838 17736 15844
rect 17972 15834 18000 16382
rect 18116 16204 18412 16224
rect 18172 16202 18196 16204
rect 18252 16202 18276 16204
rect 18332 16202 18356 16204
rect 18194 16150 18196 16202
rect 18258 16150 18270 16202
rect 18332 16150 18334 16202
rect 18172 16148 18196 16150
rect 18252 16148 18276 16150
rect 18332 16148 18356 16150
rect 18116 16128 18412 16148
rect 17960 15828 18012 15834
rect 17960 15770 18012 15776
rect 18116 15116 18412 15136
rect 18172 15114 18196 15116
rect 18252 15114 18276 15116
rect 18332 15114 18356 15116
rect 18194 15062 18196 15114
rect 18258 15062 18270 15114
rect 18332 15062 18334 15114
rect 18172 15060 18196 15062
rect 18252 15060 18276 15062
rect 18332 15060 18356 15062
rect 18116 15040 18412 15060
rect 17500 14672 17552 14678
rect 17500 14614 17552 14620
rect 17592 14672 17644 14678
rect 17592 14614 17644 14620
rect 16948 14332 17000 14338
rect 16948 14274 17000 14280
rect 17224 14332 17276 14338
rect 17224 14274 17276 14280
rect 16960 13658 16988 14274
rect 17316 14264 17368 14270
rect 17316 14206 17368 14212
rect 17408 14264 17460 14270
rect 17408 14206 17460 14212
rect 17132 14128 17184 14134
rect 17132 14070 17184 14076
rect 17144 13794 17172 14070
rect 17328 13794 17356 14206
rect 17132 13788 17184 13794
rect 17132 13730 17184 13736
rect 17316 13788 17368 13794
rect 17316 13730 17368 13736
rect 16948 13652 17000 13658
rect 16948 13594 17000 13600
rect 16672 12632 16724 12638
rect 16672 12574 16724 12580
rect 17144 12586 17172 13730
rect 17420 13046 17448 14206
rect 17512 13930 17540 14614
rect 17604 14474 17632 14614
rect 17592 14468 17644 14474
rect 17592 14410 17644 14416
rect 18116 14028 18412 14048
rect 18172 14026 18196 14028
rect 18252 14026 18276 14028
rect 18332 14026 18356 14028
rect 18194 13974 18196 14026
rect 18258 13974 18270 14026
rect 18332 13974 18334 14026
rect 18172 13972 18196 13974
rect 18252 13972 18276 13974
rect 18332 13972 18356 13974
rect 18116 13952 18412 13972
rect 18616 13930 18644 21856
rect 18708 18282 18736 21919
rect 19154 21856 19210 22656
rect 19706 21856 19762 22656
rect 20258 21856 20314 22656
rect 20810 21856 20866 22656
rect 21362 21856 21418 22656
rect 21914 21856 21970 22656
rect 22466 21856 22522 22656
rect 19168 19386 19196 21856
rect 19614 19672 19670 19681
rect 19614 19607 19670 19616
rect 19168 19358 19288 19386
rect 19154 19264 19210 19273
rect 19154 19199 19210 19208
rect 18788 19092 18840 19098
rect 18788 19034 18840 19040
rect 18696 18276 18748 18282
rect 18696 18218 18748 18224
rect 18694 17904 18750 17913
rect 18694 17839 18750 17848
rect 18708 17194 18736 17839
rect 18696 17188 18748 17194
rect 18696 17130 18748 17136
rect 17500 13924 17552 13930
rect 17500 13866 17552 13872
rect 18604 13924 18656 13930
rect 18604 13866 18656 13872
rect 18328 13720 18380 13726
rect 18328 13662 18380 13668
rect 18340 13318 18368 13662
rect 18800 13386 18828 19034
rect 19064 16984 19116 16990
rect 19064 16926 19116 16932
rect 19076 15290 19104 16926
rect 19168 16038 19196 19199
rect 19260 18826 19288 19358
rect 19248 18820 19300 18826
rect 19248 18762 19300 18768
rect 19246 18720 19302 18729
rect 19246 18655 19302 18664
rect 19340 18684 19392 18690
rect 19260 16106 19288 18655
rect 19340 18626 19392 18632
rect 19524 18684 19576 18690
rect 19524 18626 19576 18632
rect 19352 18593 19380 18626
rect 19338 18584 19394 18593
rect 19338 18519 19394 18528
rect 19340 18208 19392 18214
rect 19340 18150 19392 18156
rect 19248 16100 19300 16106
rect 19248 16042 19300 16048
rect 19156 16032 19208 16038
rect 19156 15974 19208 15980
rect 19064 15284 19116 15290
rect 19064 15226 19116 15232
rect 18788 13380 18840 13386
rect 18788 13322 18840 13328
rect 18328 13312 18380 13318
rect 18328 13254 18380 13260
rect 17592 13244 17644 13250
rect 17592 13186 17644 13192
rect 17408 13040 17460 13046
rect 17408 12982 17460 12988
rect 16316 11164 16436 11192
rect 16316 8966 16344 11164
rect 16488 11136 16540 11142
rect 16408 11084 16488 11090
rect 16408 11078 16540 11084
rect 16408 11062 16528 11078
rect 16408 10598 16436 11062
rect 16488 11000 16540 11006
rect 16488 10942 16540 10948
rect 16396 10592 16448 10598
rect 16396 10534 16448 10540
rect 16500 10530 16528 10942
rect 16488 10524 16540 10530
rect 16488 10466 16540 10472
rect 16500 10054 16528 10466
rect 16488 10048 16540 10054
rect 16488 9990 16540 9996
rect 16684 9986 16712 12574
rect 17144 12558 17448 12586
rect 16948 12088 17000 12094
rect 16948 12030 17000 12036
rect 16960 10938 16988 12030
rect 17420 11074 17448 12558
rect 17500 12564 17552 12570
rect 17500 12506 17552 12512
rect 17512 11618 17540 12506
rect 17500 11612 17552 11618
rect 17500 11554 17552 11560
rect 17316 11068 17368 11074
rect 17316 11010 17368 11016
rect 17408 11068 17460 11074
rect 17408 11010 17460 11016
rect 16948 10932 17000 10938
rect 16948 10874 17000 10880
rect 17328 10666 17356 11010
rect 17512 11006 17540 11554
rect 17500 11000 17552 11006
rect 17500 10942 17552 10948
rect 17316 10660 17368 10666
rect 17316 10602 17368 10608
rect 16764 10320 16816 10326
rect 16816 10268 16896 10274
rect 16764 10262 16896 10268
rect 16776 10246 16896 10262
rect 16672 9980 16724 9986
rect 16672 9922 16724 9928
rect 16396 9504 16448 9510
rect 16396 9446 16448 9452
rect 16304 8960 16356 8966
rect 16304 8902 16356 8908
rect 16212 7600 16264 7606
rect 16212 7542 16264 7548
rect 16028 7396 16080 7402
rect 16028 7338 16080 7344
rect 15936 3928 15988 3934
rect 15936 3870 15988 3876
rect 7820 3692 8116 3712
rect 7876 3690 7900 3692
rect 7956 3690 7980 3692
rect 8036 3690 8060 3692
rect 7898 3638 7900 3690
rect 7962 3638 7974 3690
rect 8036 3638 8038 3690
rect 7876 3636 7900 3638
rect 7956 3636 7980 3638
rect 8036 3636 8060 3638
rect 7820 3616 8116 3636
rect 14684 3692 14980 3712
rect 14740 3690 14764 3692
rect 14820 3690 14844 3692
rect 14900 3690 14924 3692
rect 14762 3638 14764 3690
rect 14826 3638 14838 3690
rect 14900 3638 14902 3690
rect 14740 3636 14764 3638
rect 14820 3636 14844 3638
rect 14900 3636 14924 3638
rect 14684 3616 14980 3636
rect 4388 3148 4684 3168
rect 4444 3146 4468 3148
rect 4524 3146 4548 3148
rect 4604 3146 4628 3148
rect 4466 3094 4468 3146
rect 4530 3094 4542 3146
rect 4604 3094 4606 3146
rect 4444 3092 4468 3094
rect 4524 3092 4548 3094
rect 4604 3092 4628 3094
rect 4388 3072 4684 3092
rect 11252 3148 11548 3168
rect 11308 3146 11332 3148
rect 11388 3146 11412 3148
rect 11468 3146 11492 3148
rect 11330 3094 11332 3146
rect 11394 3094 11406 3146
rect 11468 3094 11470 3146
rect 11308 3092 11332 3094
rect 11388 3092 11412 3094
rect 11468 3092 11492 3094
rect 11252 3072 11548 3092
rect 7820 2604 8116 2624
rect 7876 2602 7900 2604
rect 7956 2602 7980 2604
rect 8036 2602 8060 2604
rect 7898 2550 7900 2602
rect 7962 2550 7974 2602
rect 8036 2550 8038 2602
rect 7876 2548 7900 2550
rect 7956 2548 7980 2550
rect 8036 2548 8060 2550
rect 7820 2528 8116 2548
rect 14684 2604 14980 2624
rect 14740 2602 14764 2604
rect 14820 2602 14844 2604
rect 14900 2602 14924 2604
rect 14762 2550 14764 2602
rect 14826 2550 14838 2602
rect 14900 2550 14902 2602
rect 14740 2548 14764 2550
rect 14820 2548 14844 2550
rect 14900 2548 14924 2550
rect 14684 2528 14980 2548
rect 4388 2060 4684 2080
rect 4444 2058 4468 2060
rect 4524 2058 4548 2060
rect 4604 2058 4628 2060
rect 4466 2006 4468 2058
rect 4530 2006 4542 2058
rect 4604 2006 4606 2058
rect 4444 2004 4468 2006
rect 4524 2004 4548 2006
rect 4604 2004 4628 2006
rect 4388 1984 4684 2004
rect 11252 2060 11548 2080
rect 11308 2058 11332 2060
rect 11388 2058 11412 2060
rect 11468 2058 11492 2060
rect 11330 2006 11332 2058
rect 11394 2006 11406 2058
rect 11468 2006 11470 2058
rect 11308 2004 11332 2006
rect 11388 2004 11412 2006
rect 11468 2004 11492 2006
rect 11252 1984 11548 2004
rect 16408 1214 16436 9446
rect 16672 8280 16724 8286
rect 16672 8222 16724 8228
rect 16580 7804 16632 7810
rect 16580 7746 16632 7752
rect 16592 7402 16620 7746
rect 16580 7396 16632 7402
rect 16580 7338 16632 7344
rect 16684 6586 16712 8222
rect 16672 6580 16724 6586
rect 16672 6522 16724 6528
rect 16868 2302 16896 10246
rect 17512 10122 17540 10942
rect 17500 10116 17552 10122
rect 17500 10058 17552 10064
rect 17604 9510 17632 13186
rect 18116 12940 18412 12960
rect 18172 12938 18196 12940
rect 18252 12938 18276 12940
rect 18332 12938 18356 12940
rect 18194 12886 18196 12938
rect 18258 12886 18270 12938
rect 18332 12886 18334 12938
rect 18172 12884 18196 12886
rect 18252 12884 18276 12886
rect 18332 12884 18356 12886
rect 18116 12864 18412 12884
rect 19248 12632 19300 12638
rect 19248 12574 19300 12580
rect 18052 12496 18104 12502
rect 18052 12438 18104 12444
rect 18064 12230 18092 12438
rect 19260 12337 19288 12574
rect 19246 12328 19302 12337
rect 18788 12292 18840 12298
rect 19246 12263 19302 12272
rect 18788 12234 18840 12240
rect 18052 12224 18104 12230
rect 18052 12166 18104 12172
rect 17960 12156 18012 12162
rect 17960 12098 18012 12104
rect 17972 11754 18000 12098
rect 18604 11952 18656 11958
rect 18604 11894 18656 11900
rect 18116 11852 18412 11872
rect 18172 11850 18196 11852
rect 18252 11850 18276 11852
rect 18332 11850 18356 11852
rect 18194 11798 18196 11850
rect 18258 11798 18270 11850
rect 18332 11798 18334 11850
rect 18172 11796 18196 11798
rect 18252 11796 18276 11798
rect 18332 11796 18356 11798
rect 18116 11776 18412 11796
rect 17960 11748 18012 11754
rect 17960 11690 18012 11696
rect 18512 11680 18564 11686
rect 18512 11622 18564 11628
rect 17868 11068 17920 11074
rect 17868 11010 17920 11016
rect 17592 9504 17644 9510
rect 17592 9446 17644 9452
rect 17880 9034 17908 11010
rect 18116 10764 18412 10784
rect 18172 10762 18196 10764
rect 18252 10762 18276 10764
rect 18332 10762 18356 10764
rect 18194 10710 18196 10762
rect 18258 10710 18270 10762
rect 18332 10710 18334 10762
rect 18172 10708 18196 10710
rect 18252 10708 18276 10710
rect 18332 10708 18356 10710
rect 18116 10688 18412 10708
rect 17960 9980 18012 9986
rect 17960 9922 18012 9928
rect 17868 9028 17920 9034
rect 17868 8970 17920 8976
rect 17408 8348 17460 8354
rect 17408 8290 17460 8296
rect 17420 7946 17448 8290
rect 17408 7940 17460 7946
rect 17408 7882 17460 7888
rect 17224 7396 17276 7402
rect 17224 7338 17276 7344
rect 16948 6852 17000 6858
rect 16948 6794 17000 6800
rect 16960 5226 16988 6794
rect 17236 6654 17264 7338
rect 17224 6648 17276 6654
rect 17224 6590 17276 6596
rect 16948 5220 17000 5226
rect 16948 5162 17000 5168
rect 17880 3633 17908 8970
rect 17972 8898 18000 9922
rect 18116 9676 18412 9696
rect 18172 9674 18196 9676
rect 18252 9674 18276 9676
rect 18332 9674 18356 9676
rect 18194 9622 18196 9674
rect 18258 9622 18270 9674
rect 18332 9622 18334 9674
rect 18172 9620 18196 9622
rect 18252 9620 18276 9622
rect 18332 9620 18356 9622
rect 18116 9600 18412 9620
rect 18236 9436 18288 9442
rect 18236 9378 18288 9384
rect 18248 9034 18276 9378
rect 18236 9028 18288 9034
rect 18236 8970 18288 8976
rect 17960 8892 18012 8898
rect 17960 8834 18012 8840
rect 17972 7742 18000 8834
rect 18524 8694 18552 11622
rect 18512 8688 18564 8694
rect 18512 8630 18564 8636
rect 18116 8588 18412 8608
rect 18172 8586 18196 8588
rect 18252 8586 18276 8588
rect 18332 8586 18356 8588
rect 18194 8534 18196 8586
rect 18258 8534 18270 8586
rect 18332 8534 18334 8586
rect 18172 8532 18196 8534
rect 18252 8532 18276 8534
rect 18332 8532 18356 8534
rect 18116 8512 18412 8532
rect 17960 7736 18012 7742
rect 17960 7678 18012 7684
rect 18116 7500 18412 7520
rect 18172 7498 18196 7500
rect 18252 7498 18276 7500
rect 18332 7498 18356 7500
rect 18194 7446 18196 7498
rect 18258 7446 18270 7498
rect 18332 7446 18334 7498
rect 18172 7444 18196 7446
rect 18252 7444 18276 7446
rect 18332 7444 18356 7446
rect 18116 7424 18412 7444
rect 18512 6852 18564 6858
rect 18512 6794 18564 6800
rect 18524 6489 18552 6794
rect 18616 6586 18644 11894
rect 18800 11090 18828 12234
rect 18880 11408 18932 11414
rect 18880 11350 18932 11356
rect 18892 11210 18920 11350
rect 18880 11204 18932 11210
rect 18880 11146 18932 11152
rect 18800 11062 18920 11090
rect 18696 10320 18748 10326
rect 18696 10262 18748 10268
rect 18604 6580 18656 6586
rect 18604 6522 18656 6528
rect 18510 6480 18566 6489
rect 18116 6412 18412 6432
rect 18510 6415 18566 6424
rect 18172 6410 18196 6412
rect 18252 6410 18276 6412
rect 18332 6410 18356 6412
rect 18194 6358 18196 6410
rect 18258 6358 18270 6410
rect 18332 6358 18334 6410
rect 18172 6356 18196 6358
rect 18252 6356 18276 6358
rect 18332 6356 18356 6358
rect 18116 6336 18412 6356
rect 17960 6308 18012 6314
rect 17960 6250 18012 6256
rect 17972 5537 18000 6250
rect 17958 5528 18014 5537
rect 17958 5463 18014 5472
rect 18116 5324 18412 5344
rect 18172 5322 18196 5324
rect 18252 5322 18276 5324
rect 18332 5322 18356 5324
rect 18194 5270 18196 5322
rect 18258 5270 18270 5322
rect 18332 5270 18334 5322
rect 18172 5268 18196 5270
rect 18252 5268 18276 5270
rect 18332 5268 18356 5270
rect 18116 5248 18412 5268
rect 17960 5220 18012 5226
rect 17960 5162 18012 5168
rect 17972 4585 18000 5162
rect 17958 4576 18014 4585
rect 17958 4511 18014 4520
rect 18116 4236 18412 4256
rect 18172 4234 18196 4236
rect 18252 4234 18276 4236
rect 18332 4234 18356 4236
rect 18194 4182 18196 4234
rect 18258 4182 18270 4234
rect 18332 4182 18334 4234
rect 18172 4180 18196 4182
rect 18252 4180 18276 4182
rect 18332 4180 18356 4182
rect 18116 4160 18412 4180
rect 18512 3996 18564 4002
rect 18512 3938 18564 3944
rect 17866 3624 17922 3633
rect 17866 3559 17922 3568
rect 18524 3225 18552 3938
rect 18510 3216 18566 3225
rect 18116 3148 18412 3168
rect 18510 3151 18566 3160
rect 18172 3146 18196 3148
rect 18252 3146 18276 3148
rect 18332 3146 18356 3148
rect 18194 3094 18196 3146
rect 18258 3094 18270 3146
rect 18332 3094 18334 3146
rect 18172 3092 18196 3094
rect 18252 3092 18276 3094
rect 18332 3092 18356 3094
rect 18116 3072 18412 3092
rect 16856 2296 16908 2302
rect 16856 2238 16908 2244
rect 18116 2060 18412 2080
rect 18172 2058 18196 2060
rect 18252 2058 18276 2060
rect 18332 2058 18356 2060
rect 18194 2006 18196 2058
rect 18258 2006 18270 2058
rect 18332 2006 18334 2058
rect 18172 2004 18196 2006
rect 18252 2004 18276 2006
rect 18332 2004 18356 2006
rect 18116 1984 18412 2004
rect 16396 1208 16448 1214
rect 16396 1150 16448 1156
rect 17960 1208 18012 1214
rect 17960 1150 18012 1156
rect 17972 97 18000 1150
rect 18708 913 18736 10262
rect 18788 9980 18840 9986
rect 18788 9922 18840 9928
rect 18800 9034 18828 9922
rect 18788 9028 18840 9034
rect 18788 8970 18840 8976
rect 18788 8688 18840 8694
rect 18788 8630 18840 8636
rect 18694 904 18750 913
rect 18694 839 18750 848
rect 18800 505 18828 8630
rect 18892 1457 18920 11062
rect 19248 10932 19300 10938
rect 19248 10874 19300 10880
rect 19260 10530 19288 10874
rect 19352 10666 19380 18150
rect 19432 18072 19484 18078
rect 19432 18014 19484 18020
rect 19444 17466 19472 18014
rect 19536 18010 19564 18626
rect 19628 18282 19656 19607
rect 19616 18276 19668 18282
rect 19616 18218 19668 18224
rect 19616 18140 19668 18146
rect 19616 18082 19668 18088
rect 19524 18004 19576 18010
rect 19524 17946 19576 17952
rect 19432 17460 19484 17466
rect 19432 17402 19484 17408
rect 19524 16984 19576 16990
rect 19524 16926 19576 16932
rect 19536 16582 19564 16926
rect 19524 16576 19576 16582
rect 19524 16518 19576 16524
rect 19628 12774 19656 18082
rect 19720 18026 19748 21856
rect 20166 21032 20222 21041
rect 20166 20967 20222 20976
rect 20180 19914 20208 20967
rect 20168 19908 20220 19914
rect 20168 19850 20220 19856
rect 19984 19772 20036 19778
rect 19984 19714 20036 19720
rect 19996 19234 20024 19714
rect 20272 19250 20300 21856
rect 20626 20624 20682 20633
rect 20626 20559 20682 20568
rect 20534 20080 20590 20089
rect 20534 20015 20590 20024
rect 20444 19772 20496 19778
rect 20444 19714 20496 19720
rect 19984 19228 20036 19234
rect 19984 19170 20036 19176
rect 20088 19222 20300 19250
rect 19984 18072 20036 18078
rect 19720 17998 19932 18026
rect 19984 18014 20036 18020
rect 19800 17936 19852 17942
rect 19800 17878 19852 17884
rect 19708 15896 19760 15902
rect 19708 15838 19760 15844
rect 19720 14882 19748 15838
rect 19708 14876 19760 14882
rect 19708 14818 19760 14824
rect 19616 12768 19668 12774
rect 19616 12710 19668 12716
rect 19812 12570 19840 17878
rect 19800 12564 19852 12570
rect 19800 12506 19852 12512
rect 19904 11754 19932 17998
rect 19996 17058 20024 18014
rect 19984 17052 20036 17058
rect 19984 16994 20036 17000
rect 19984 16916 20036 16922
rect 19984 16858 20036 16864
rect 19996 16514 20024 16858
rect 19984 16508 20036 16514
rect 19984 16450 20036 16456
rect 20088 16394 20116 19222
rect 20260 19160 20312 19166
rect 20260 19102 20312 19108
rect 20272 18758 20300 19102
rect 20352 18820 20404 18826
rect 20352 18762 20404 18768
rect 20260 18752 20312 18758
rect 20260 18694 20312 18700
rect 20166 18312 20222 18321
rect 20166 18247 20168 18256
rect 20220 18247 20222 18256
rect 20168 18218 20220 18224
rect 20168 17732 20220 17738
rect 20168 17674 20220 17680
rect 20180 16514 20208 17674
rect 20168 16508 20220 16514
rect 20168 16450 20220 16456
rect 20088 16366 20208 16394
rect 20180 16088 20208 16366
rect 20088 16060 20208 16088
rect 19984 13244 20036 13250
rect 19984 13186 20036 13192
rect 19996 12842 20024 13186
rect 19984 12836 20036 12842
rect 19984 12778 20036 12784
rect 20088 12722 20116 16060
rect 20166 16000 20222 16009
rect 20166 15935 20222 15944
rect 20180 15562 20208 15935
rect 20260 15896 20312 15902
rect 20260 15838 20312 15844
rect 20168 15556 20220 15562
rect 20168 15498 20220 15504
rect 20168 15420 20220 15426
rect 20168 15362 20220 15368
rect 20180 14406 20208 15362
rect 20272 14746 20300 15838
rect 20364 14762 20392 18762
rect 20456 18758 20484 19714
rect 20548 19370 20576 20015
rect 20640 19914 20668 20559
rect 20628 19908 20680 19914
rect 20628 19850 20680 19856
rect 20536 19364 20588 19370
rect 20536 19306 20588 19312
rect 20444 18752 20496 18758
rect 20444 18694 20496 18700
rect 20536 17936 20588 17942
rect 20536 17878 20588 17884
rect 20442 17360 20498 17369
rect 20442 17295 20498 17304
rect 20456 17194 20484 17295
rect 20444 17188 20496 17194
rect 20444 17130 20496 17136
rect 20260 14740 20312 14746
rect 20364 14734 20484 14762
rect 20260 14682 20312 14688
rect 20350 14640 20406 14649
rect 20350 14575 20406 14584
rect 20168 14400 20220 14406
rect 20168 14342 20220 14348
rect 20260 13720 20312 13726
rect 20260 13662 20312 13668
rect 20272 12881 20300 13662
rect 20364 13386 20392 14575
rect 20456 13810 20484 14734
rect 20548 13930 20576 17878
rect 20720 17392 20772 17398
rect 20720 17334 20772 17340
rect 20732 16961 20760 17334
rect 20824 17074 20852 21856
rect 20996 18480 21048 18486
rect 20996 18422 21048 18428
rect 20824 17046 20944 17074
rect 20718 16952 20774 16961
rect 20718 16887 20774 16896
rect 20628 16644 20680 16650
rect 20628 16586 20680 16592
rect 20640 16417 20668 16586
rect 20626 16408 20682 16417
rect 20626 16343 20682 16352
rect 20718 15592 20774 15601
rect 20718 15527 20720 15536
rect 20772 15527 20774 15536
rect 20720 15498 20772 15504
rect 20718 15048 20774 15057
rect 20718 14983 20774 14992
rect 20732 14474 20760 14983
rect 20720 14468 20772 14474
rect 20720 14410 20772 14416
rect 20810 14232 20866 14241
rect 20810 14167 20866 14176
rect 20536 13924 20588 13930
rect 20536 13866 20588 13872
rect 20456 13782 20668 13810
rect 20442 13688 20498 13697
rect 20442 13623 20498 13632
rect 20352 13380 20404 13386
rect 20352 13322 20404 13328
rect 20350 13280 20406 13289
rect 20350 13215 20406 13224
rect 20258 12872 20314 12881
rect 20364 12842 20392 13215
rect 20258 12807 20314 12816
rect 20352 12836 20404 12842
rect 20352 12778 20404 12784
rect 20088 12694 20300 12722
rect 20168 12632 20220 12638
rect 20168 12574 20220 12580
rect 20076 12564 20128 12570
rect 20076 12506 20128 12512
rect 19984 12156 20036 12162
rect 19984 12098 20036 12104
rect 19996 11929 20024 12098
rect 19982 11920 20038 11929
rect 19982 11855 20038 11864
rect 19892 11748 19944 11754
rect 19892 11690 19944 11696
rect 19984 11068 20036 11074
rect 19984 11010 20036 11016
rect 19340 10660 19392 10666
rect 19340 10602 19392 10608
rect 19996 10569 20024 11010
rect 19982 10560 20038 10569
rect 19248 10524 19300 10530
rect 19982 10495 20038 10504
rect 19248 10466 19300 10472
rect 19260 10122 19288 10466
rect 19248 10116 19300 10122
rect 19248 10058 19300 10064
rect 18970 10016 19026 10025
rect 18970 9951 19026 9960
rect 18984 9374 19012 9951
rect 19432 9436 19484 9442
rect 19432 9378 19484 9384
rect 18972 9368 19024 9374
rect 18972 9310 19024 9316
rect 19064 9232 19116 9238
rect 19064 9174 19116 9180
rect 19076 6722 19104 9174
rect 19444 8898 19472 9378
rect 20088 9034 20116 12506
rect 20180 12230 20208 12574
rect 20272 12298 20300 12694
rect 20260 12292 20312 12298
rect 20260 12234 20312 12240
rect 20168 12224 20220 12230
rect 20168 12166 20220 12172
rect 20260 11544 20312 11550
rect 20260 11486 20312 11492
rect 20272 10977 20300 11486
rect 20258 10968 20314 10977
rect 20258 10903 20314 10912
rect 20260 10456 20312 10462
rect 20260 10398 20312 10404
rect 20272 9617 20300 10398
rect 20258 9608 20314 9617
rect 20258 9543 20314 9552
rect 20076 9028 20128 9034
rect 20076 8970 20128 8976
rect 19432 8892 19484 8898
rect 19432 8834 19484 8840
rect 19984 8892 20036 8898
rect 19984 8834 20036 8840
rect 19444 7946 19472 8834
rect 19996 8665 20024 8834
rect 19982 8656 20038 8665
rect 19982 8591 20038 8600
rect 20456 8490 20484 13623
rect 20536 12156 20588 12162
rect 20536 12098 20588 12104
rect 20548 11521 20576 12098
rect 20534 11512 20590 11521
rect 20534 11447 20590 11456
rect 20640 11210 20668 13782
rect 20718 13688 20774 13697
rect 20718 13623 20774 13632
rect 20732 13386 20760 13623
rect 20720 13380 20772 13386
rect 20720 13322 20772 13328
rect 20824 11210 20852 14167
rect 20916 12026 20944 17046
rect 20904 12020 20956 12026
rect 20904 11962 20956 11968
rect 20628 11204 20680 11210
rect 20628 11146 20680 11152
rect 20812 11204 20864 11210
rect 20812 11146 20864 11152
rect 21008 10122 21036 18422
rect 21376 18146 21404 21856
rect 21364 18140 21416 18146
rect 21364 18082 21416 18088
rect 21088 18004 21140 18010
rect 21088 17946 21140 17952
rect 20996 10116 21048 10122
rect 20996 10058 21048 10064
rect 20536 9980 20588 9986
rect 20536 9922 20588 9928
rect 20548 9209 20576 9922
rect 20534 9200 20590 9209
rect 20534 9135 20590 9144
rect 20536 8892 20588 8898
rect 20536 8834 20588 8840
rect 20444 8484 20496 8490
rect 20444 8426 20496 8432
rect 20260 8280 20312 8286
rect 20548 8257 20576 8834
rect 20260 8222 20312 8228
rect 20534 8248 20590 8257
rect 19432 7940 19484 7946
rect 19432 7882 19484 7888
rect 20272 7849 20300 8222
rect 20534 8183 20590 8192
rect 20258 7840 20314 7849
rect 19984 7804 20036 7810
rect 20258 7775 20314 7784
rect 20536 7804 20588 7810
rect 19984 7746 20036 7752
rect 20536 7746 20588 7752
rect 19996 7305 20024 7746
rect 19982 7296 20038 7305
rect 19982 7231 20038 7240
rect 20548 6897 20576 7746
rect 20534 6888 20590 6897
rect 20534 6823 20590 6832
rect 19064 6716 19116 6722
rect 19064 6658 19116 6664
rect 20536 6716 20588 6722
rect 20536 6658 20588 6664
rect 19064 6580 19116 6586
rect 19064 6522 19116 6528
rect 19076 2273 19104 6522
rect 20548 5945 20576 6658
rect 20534 5936 20590 5945
rect 20534 5871 20590 5880
rect 20536 5628 20588 5634
rect 20536 5570 20588 5576
rect 20548 4993 20576 5570
rect 20534 4984 20590 4993
rect 20534 4919 20590 4928
rect 21100 4682 21128 17946
rect 21928 17942 21956 21856
rect 22480 18010 22508 21856
rect 22468 18004 22520 18010
rect 22468 17946 22520 17952
rect 21916 17936 21968 17942
rect 21916 17878 21968 17884
rect 21088 4676 21140 4682
rect 21088 4618 21140 4624
rect 20536 4540 20588 4546
rect 20536 4482 20588 4488
rect 20548 4177 20576 4482
rect 20534 4168 20590 4177
rect 20534 4103 20590 4112
rect 19248 3928 19300 3934
rect 19248 3870 19300 3876
rect 19260 2817 19288 3870
rect 19246 2808 19302 2817
rect 19246 2743 19302 2752
rect 19248 2296 19300 2302
rect 19062 2264 19118 2273
rect 19248 2238 19300 2244
rect 19062 2199 19118 2208
rect 19260 1865 19288 2238
rect 19246 1856 19302 1865
rect 19246 1791 19302 1800
rect 18878 1448 18934 1457
rect 18878 1383 18934 1392
rect 18786 496 18842 505
rect 18786 431 18842 440
rect 17958 88 18014 97
rect 17958 23 18014 32
<< via2 >>
rect 17958 22336 18014 22392
rect 4388 19466 4444 19468
rect 4468 19466 4524 19468
rect 4548 19466 4604 19468
rect 4628 19466 4684 19468
rect 4388 19414 4414 19466
rect 4414 19414 4444 19466
rect 4468 19414 4478 19466
rect 4478 19414 4524 19466
rect 4548 19414 4594 19466
rect 4594 19414 4604 19466
rect 4628 19414 4658 19466
rect 4658 19414 4684 19466
rect 4388 19412 4444 19414
rect 4468 19412 4524 19414
rect 4548 19412 4604 19414
rect 4628 19412 4684 19414
rect 4388 18378 4444 18380
rect 4468 18378 4524 18380
rect 4548 18378 4604 18380
rect 4628 18378 4684 18380
rect 4388 18326 4414 18378
rect 4414 18326 4444 18378
rect 4468 18326 4478 18378
rect 4478 18326 4524 18378
rect 4548 18326 4594 18378
rect 4594 18326 4604 18378
rect 4628 18326 4658 18378
rect 4658 18326 4684 18378
rect 4388 18324 4444 18326
rect 4468 18324 4524 18326
rect 4548 18324 4604 18326
rect 4628 18324 4684 18326
rect 4388 17290 4444 17292
rect 4468 17290 4524 17292
rect 4548 17290 4604 17292
rect 4628 17290 4684 17292
rect 4388 17238 4414 17290
rect 4414 17238 4444 17290
rect 4468 17238 4478 17290
rect 4478 17238 4524 17290
rect 4548 17238 4594 17290
rect 4594 17238 4604 17290
rect 4628 17238 4658 17290
rect 4658 17238 4684 17290
rect 4388 17236 4444 17238
rect 4468 17236 4524 17238
rect 4548 17236 4604 17238
rect 4628 17236 4684 17238
rect 4066 17032 4122 17088
rect 5814 18664 5870 18720
rect 4388 16202 4444 16204
rect 4468 16202 4524 16204
rect 4548 16202 4604 16204
rect 4628 16202 4684 16204
rect 4388 16150 4414 16202
rect 4414 16150 4444 16202
rect 4468 16150 4478 16202
rect 4478 16150 4524 16202
rect 4548 16150 4594 16202
rect 4594 16150 4604 16202
rect 4628 16150 4658 16202
rect 4658 16150 4684 16202
rect 4388 16148 4444 16150
rect 4468 16148 4524 16150
rect 4548 16148 4604 16150
rect 4628 16148 4684 16150
rect 4388 15114 4444 15116
rect 4468 15114 4524 15116
rect 4548 15114 4604 15116
rect 4628 15114 4684 15116
rect 4388 15062 4414 15114
rect 4414 15062 4444 15114
rect 4468 15062 4478 15114
rect 4478 15062 4524 15114
rect 4548 15062 4594 15114
rect 4594 15062 4604 15114
rect 4628 15062 4658 15114
rect 4658 15062 4684 15114
rect 4388 15060 4444 15062
rect 4468 15060 4524 15062
rect 4548 15060 4604 15062
rect 4628 15060 4684 15062
rect 7820 20010 7876 20012
rect 7900 20010 7956 20012
rect 7980 20010 8036 20012
rect 8060 20010 8116 20012
rect 7820 19958 7846 20010
rect 7846 19958 7876 20010
rect 7900 19958 7910 20010
rect 7910 19958 7956 20010
rect 7980 19958 8026 20010
rect 8026 19958 8036 20010
rect 8060 19958 8090 20010
rect 8090 19958 8116 20010
rect 7820 19956 7876 19958
rect 7900 19956 7956 19958
rect 7980 19956 8036 19958
rect 8060 19956 8116 19958
rect 7820 18922 7876 18924
rect 7900 18922 7956 18924
rect 7980 18922 8036 18924
rect 8060 18922 8116 18924
rect 7820 18870 7846 18922
rect 7846 18870 7876 18922
rect 7900 18870 7910 18922
rect 7910 18870 7956 18922
rect 7980 18870 8026 18922
rect 8026 18870 8036 18922
rect 8060 18870 8090 18922
rect 8090 18870 8116 18922
rect 7820 18868 7876 18870
rect 7900 18868 7956 18870
rect 7980 18868 8036 18870
rect 8060 18868 8116 18870
rect 8114 18664 8170 18720
rect 7820 17834 7876 17836
rect 7900 17834 7956 17836
rect 7980 17834 8036 17836
rect 8060 17834 8116 17836
rect 7820 17782 7846 17834
rect 7846 17782 7876 17834
rect 7900 17782 7910 17834
rect 7910 17782 7956 17834
rect 7980 17782 8026 17834
rect 8026 17782 8036 17834
rect 8060 17782 8090 17834
rect 8090 17782 8116 17834
rect 7820 17780 7876 17782
rect 7900 17780 7956 17782
rect 7980 17780 8036 17782
rect 8060 17780 8116 17782
rect 7820 16746 7876 16748
rect 7900 16746 7956 16748
rect 7980 16746 8036 16748
rect 8060 16746 8116 16748
rect 7820 16694 7846 16746
rect 7846 16694 7876 16746
rect 7900 16694 7910 16746
rect 7910 16694 7956 16746
rect 7980 16694 8026 16746
rect 8026 16694 8036 16746
rect 8060 16694 8090 16746
rect 8090 16694 8116 16746
rect 7820 16692 7876 16694
rect 7900 16692 7956 16694
rect 7980 16692 8036 16694
rect 8060 16692 8116 16694
rect 11252 19466 11308 19468
rect 11332 19466 11388 19468
rect 11412 19466 11468 19468
rect 11492 19466 11548 19468
rect 11252 19414 11278 19466
rect 11278 19414 11308 19466
rect 11332 19414 11342 19466
rect 11342 19414 11388 19466
rect 11412 19414 11458 19466
rect 11458 19414 11468 19466
rect 11492 19414 11522 19466
rect 11522 19414 11548 19466
rect 11252 19412 11308 19414
rect 11332 19412 11388 19414
rect 11412 19412 11468 19414
rect 11492 19412 11548 19414
rect 7820 15658 7876 15660
rect 7900 15658 7956 15660
rect 7980 15658 8036 15660
rect 8060 15658 8116 15660
rect 7820 15606 7846 15658
rect 7846 15606 7876 15658
rect 7900 15606 7910 15658
rect 7910 15606 7956 15658
rect 7980 15606 8026 15658
rect 8026 15606 8036 15658
rect 8060 15606 8090 15658
rect 8090 15606 8116 15658
rect 7820 15604 7876 15606
rect 7900 15604 7956 15606
rect 7980 15604 8036 15606
rect 8060 15604 8116 15606
rect 4388 14026 4444 14028
rect 4468 14026 4524 14028
rect 4548 14026 4604 14028
rect 4628 14026 4684 14028
rect 4388 13974 4414 14026
rect 4414 13974 4444 14026
rect 4468 13974 4478 14026
rect 4478 13974 4524 14026
rect 4548 13974 4594 14026
rect 4594 13974 4604 14026
rect 4628 13974 4658 14026
rect 4658 13974 4684 14026
rect 4388 13972 4444 13974
rect 4468 13972 4524 13974
rect 4548 13972 4604 13974
rect 4628 13972 4684 13974
rect 4388 12938 4444 12940
rect 4468 12938 4524 12940
rect 4548 12938 4604 12940
rect 4628 12938 4684 12940
rect 4388 12886 4414 12938
rect 4414 12886 4444 12938
rect 4468 12886 4478 12938
rect 4478 12886 4524 12938
rect 4548 12886 4594 12938
rect 4594 12886 4604 12938
rect 4628 12886 4658 12938
rect 4658 12886 4684 12938
rect 4388 12884 4444 12886
rect 4468 12884 4524 12886
rect 4548 12884 4604 12886
rect 4628 12884 4684 12886
rect 4388 11850 4444 11852
rect 4468 11850 4524 11852
rect 4548 11850 4604 11852
rect 4628 11850 4684 11852
rect 4388 11798 4414 11850
rect 4414 11798 4444 11850
rect 4468 11798 4478 11850
rect 4478 11798 4524 11850
rect 4548 11798 4594 11850
rect 4594 11798 4604 11850
rect 4628 11798 4658 11850
rect 4658 11798 4684 11850
rect 4388 11796 4444 11798
rect 4468 11796 4524 11798
rect 4548 11796 4604 11798
rect 4628 11796 4684 11798
rect 7820 14570 7876 14572
rect 7900 14570 7956 14572
rect 7980 14570 8036 14572
rect 8060 14570 8116 14572
rect 7820 14518 7846 14570
rect 7846 14518 7876 14570
rect 7900 14518 7910 14570
rect 7910 14518 7956 14570
rect 7980 14518 8026 14570
rect 8026 14518 8036 14570
rect 8060 14518 8090 14570
rect 8090 14518 8116 14570
rect 7820 14516 7876 14518
rect 7900 14516 7956 14518
rect 7980 14516 8036 14518
rect 8060 14516 8116 14518
rect 7820 13482 7876 13484
rect 7900 13482 7956 13484
rect 7980 13482 8036 13484
rect 8060 13482 8116 13484
rect 7820 13430 7846 13482
rect 7846 13430 7876 13482
rect 7900 13430 7910 13482
rect 7910 13430 7956 13482
rect 7980 13430 8026 13482
rect 8026 13430 8036 13482
rect 8060 13430 8090 13482
rect 8090 13430 8116 13482
rect 7820 13428 7876 13430
rect 7900 13428 7956 13430
rect 7980 13428 8036 13430
rect 8060 13428 8116 13430
rect 7820 12394 7876 12396
rect 7900 12394 7956 12396
rect 7980 12394 8036 12396
rect 8060 12394 8116 12396
rect 7820 12342 7846 12394
rect 7846 12342 7876 12394
rect 7900 12342 7910 12394
rect 7910 12342 7956 12394
rect 7980 12342 8026 12394
rect 8026 12342 8036 12394
rect 8060 12342 8090 12394
rect 8090 12342 8116 12394
rect 7820 12340 7876 12342
rect 7900 12340 7956 12342
rect 7980 12340 8036 12342
rect 8060 12340 8116 12342
rect 11252 18378 11308 18380
rect 11332 18378 11388 18380
rect 11412 18378 11468 18380
rect 11492 18378 11548 18380
rect 11252 18326 11278 18378
rect 11278 18326 11308 18378
rect 11332 18326 11342 18378
rect 11342 18326 11388 18378
rect 11412 18326 11458 18378
rect 11458 18326 11468 18378
rect 11492 18326 11522 18378
rect 11522 18326 11548 18378
rect 11252 18324 11308 18326
rect 11332 18324 11388 18326
rect 11412 18324 11468 18326
rect 11492 18324 11548 18326
rect 11252 17290 11308 17292
rect 11332 17290 11388 17292
rect 11412 17290 11468 17292
rect 11492 17290 11548 17292
rect 11252 17238 11278 17290
rect 11278 17238 11308 17290
rect 11332 17238 11342 17290
rect 11342 17238 11388 17290
rect 11412 17238 11458 17290
rect 11458 17238 11468 17290
rect 11492 17238 11522 17290
rect 11522 17238 11548 17290
rect 11252 17236 11308 17238
rect 11332 17236 11388 17238
rect 11412 17236 11468 17238
rect 11492 17236 11548 17238
rect 11252 16202 11308 16204
rect 11332 16202 11388 16204
rect 11412 16202 11468 16204
rect 11492 16202 11548 16204
rect 11252 16150 11278 16202
rect 11278 16150 11308 16202
rect 11332 16150 11342 16202
rect 11342 16150 11388 16202
rect 11412 16150 11458 16202
rect 11458 16150 11468 16202
rect 11492 16150 11522 16202
rect 11522 16150 11548 16202
rect 11252 16148 11308 16150
rect 11332 16148 11388 16150
rect 11412 16148 11468 16150
rect 11492 16148 11548 16150
rect 11252 15114 11308 15116
rect 11332 15114 11388 15116
rect 11412 15114 11468 15116
rect 11492 15114 11548 15116
rect 11252 15062 11278 15114
rect 11278 15062 11308 15114
rect 11332 15062 11342 15114
rect 11342 15062 11388 15114
rect 11412 15062 11458 15114
rect 11458 15062 11468 15114
rect 11492 15062 11522 15114
rect 11522 15062 11548 15114
rect 11252 15060 11308 15062
rect 11332 15060 11388 15062
rect 11412 15060 11468 15062
rect 11492 15060 11548 15062
rect 11252 14026 11308 14028
rect 11332 14026 11388 14028
rect 11412 14026 11468 14028
rect 11492 14026 11548 14028
rect 11252 13974 11278 14026
rect 11278 13974 11308 14026
rect 11332 13974 11342 14026
rect 11342 13974 11388 14026
rect 11412 13974 11458 14026
rect 11458 13974 11468 14026
rect 11492 13974 11522 14026
rect 11522 13974 11548 14026
rect 11252 13972 11308 13974
rect 11332 13972 11388 13974
rect 11412 13972 11468 13974
rect 11492 13972 11548 13974
rect 11252 12938 11308 12940
rect 11332 12938 11388 12940
rect 11412 12938 11468 12940
rect 11492 12938 11548 12940
rect 11252 12886 11278 12938
rect 11278 12886 11308 12938
rect 11332 12886 11342 12938
rect 11342 12886 11388 12938
rect 11412 12886 11458 12938
rect 11458 12886 11468 12938
rect 11492 12886 11522 12938
rect 11522 12886 11548 12938
rect 11252 12884 11308 12886
rect 11332 12884 11388 12886
rect 11412 12884 11468 12886
rect 11492 12884 11548 12886
rect 4388 10762 4444 10764
rect 4468 10762 4524 10764
rect 4548 10762 4604 10764
rect 4628 10762 4684 10764
rect 4388 10710 4414 10762
rect 4414 10710 4444 10762
rect 4468 10710 4478 10762
rect 4478 10710 4524 10762
rect 4548 10710 4594 10762
rect 4594 10710 4604 10762
rect 4628 10710 4658 10762
rect 4658 10710 4684 10762
rect 4388 10708 4444 10710
rect 4468 10708 4524 10710
rect 4548 10708 4604 10710
rect 4628 10708 4684 10710
rect 7820 11306 7876 11308
rect 7900 11306 7956 11308
rect 7980 11306 8036 11308
rect 8060 11306 8116 11308
rect 7820 11254 7846 11306
rect 7846 11254 7876 11306
rect 7900 11254 7910 11306
rect 7910 11254 7956 11306
rect 7980 11254 8026 11306
rect 8026 11254 8036 11306
rect 8060 11254 8090 11306
rect 8090 11254 8116 11306
rect 7820 11252 7876 11254
rect 7900 11252 7956 11254
rect 7980 11252 8036 11254
rect 8060 11252 8116 11254
rect 11252 11850 11308 11852
rect 11332 11850 11388 11852
rect 11412 11850 11468 11852
rect 11492 11850 11548 11852
rect 11252 11798 11278 11850
rect 11278 11798 11308 11850
rect 11332 11798 11342 11850
rect 11342 11798 11388 11850
rect 11412 11798 11458 11850
rect 11458 11798 11468 11850
rect 11492 11798 11522 11850
rect 11522 11798 11548 11850
rect 11252 11796 11308 11798
rect 11332 11796 11388 11798
rect 11412 11796 11468 11798
rect 11492 11796 11548 11798
rect 10598 11456 10654 11512
rect 11252 10762 11308 10764
rect 11332 10762 11388 10764
rect 11412 10762 11468 10764
rect 11492 10762 11548 10764
rect 11252 10710 11278 10762
rect 11278 10710 11308 10762
rect 11332 10710 11342 10762
rect 11342 10710 11388 10762
rect 11412 10710 11458 10762
rect 11458 10710 11468 10762
rect 11492 10710 11522 10762
rect 11522 10710 11548 10762
rect 11252 10708 11308 10710
rect 11332 10708 11388 10710
rect 11412 10708 11468 10710
rect 11492 10708 11548 10710
rect 7820 10218 7876 10220
rect 7900 10218 7956 10220
rect 7980 10218 8036 10220
rect 8060 10218 8116 10220
rect 7820 10166 7846 10218
rect 7846 10166 7876 10218
rect 7900 10166 7910 10218
rect 7910 10166 7956 10218
rect 7980 10166 8026 10218
rect 8026 10166 8036 10218
rect 8060 10166 8090 10218
rect 8090 10166 8116 10218
rect 7820 10164 7876 10166
rect 7900 10164 7956 10166
rect 7980 10164 8036 10166
rect 8060 10164 8116 10166
rect 4388 9674 4444 9676
rect 4468 9674 4524 9676
rect 4548 9674 4604 9676
rect 4628 9674 4684 9676
rect 4388 9622 4414 9674
rect 4414 9622 4444 9674
rect 4468 9622 4478 9674
rect 4478 9622 4524 9674
rect 4548 9622 4594 9674
rect 4594 9622 4604 9674
rect 4628 9622 4658 9674
rect 4658 9622 4684 9674
rect 4388 9620 4444 9622
rect 4468 9620 4524 9622
rect 4548 9620 4604 9622
rect 4628 9620 4684 9622
rect 4388 8586 4444 8588
rect 4468 8586 4524 8588
rect 4548 8586 4604 8588
rect 4628 8586 4684 8588
rect 4388 8534 4414 8586
rect 4414 8534 4444 8586
rect 4468 8534 4478 8586
rect 4478 8534 4524 8586
rect 4548 8534 4594 8586
rect 4594 8534 4604 8586
rect 4628 8534 4658 8586
rect 4658 8534 4684 8586
rect 4388 8532 4444 8534
rect 4468 8532 4524 8534
rect 4548 8532 4604 8534
rect 4628 8532 4684 8534
rect 4388 7498 4444 7500
rect 4468 7498 4524 7500
rect 4548 7498 4604 7500
rect 4628 7498 4684 7500
rect 4388 7446 4414 7498
rect 4414 7446 4444 7498
rect 4468 7446 4478 7498
rect 4478 7446 4524 7498
rect 4548 7446 4594 7498
rect 4594 7446 4604 7498
rect 4628 7446 4658 7498
rect 4658 7446 4684 7498
rect 4388 7444 4444 7446
rect 4468 7444 4524 7446
rect 4548 7444 4604 7446
rect 4628 7444 4684 7446
rect 7820 9130 7876 9132
rect 7900 9130 7956 9132
rect 7980 9130 8036 9132
rect 8060 9130 8116 9132
rect 7820 9078 7846 9130
rect 7846 9078 7876 9130
rect 7900 9078 7910 9130
rect 7910 9078 7956 9130
rect 7980 9078 8026 9130
rect 8026 9078 8036 9130
rect 8060 9078 8090 9130
rect 8090 9078 8116 9130
rect 7820 9076 7876 9078
rect 7900 9076 7956 9078
rect 7980 9076 8036 9078
rect 8060 9076 8116 9078
rect 11252 9674 11308 9676
rect 11332 9674 11388 9676
rect 11412 9674 11468 9676
rect 11492 9674 11548 9676
rect 11252 9622 11278 9674
rect 11278 9622 11308 9674
rect 11332 9622 11342 9674
rect 11342 9622 11388 9674
rect 11412 9622 11458 9674
rect 11458 9622 11468 9674
rect 11492 9622 11522 9674
rect 11522 9622 11548 9674
rect 11252 9620 11308 9622
rect 11332 9620 11388 9622
rect 11412 9620 11468 9622
rect 11492 9620 11548 9622
rect 11252 8586 11308 8588
rect 11332 8586 11388 8588
rect 11412 8586 11468 8588
rect 11492 8586 11548 8588
rect 11252 8534 11278 8586
rect 11278 8534 11308 8586
rect 11332 8534 11342 8586
rect 11342 8534 11388 8586
rect 11412 8534 11458 8586
rect 11458 8534 11468 8586
rect 11492 8534 11522 8586
rect 11522 8534 11548 8586
rect 11252 8532 11308 8534
rect 11332 8532 11388 8534
rect 11412 8532 11468 8534
rect 11492 8532 11548 8534
rect 7820 8042 7876 8044
rect 7900 8042 7956 8044
rect 7980 8042 8036 8044
rect 8060 8042 8116 8044
rect 7820 7990 7846 8042
rect 7846 7990 7876 8042
rect 7900 7990 7910 8042
rect 7910 7990 7956 8042
rect 7980 7990 8026 8042
rect 8026 7990 8036 8042
rect 8060 7990 8090 8042
rect 8090 7990 8116 8042
rect 7820 7988 7876 7990
rect 7900 7988 7956 7990
rect 7980 7988 8036 7990
rect 8060 7988 8116 7990
rect 11252 7498 11308 7500
rect 11332 7498 11388 7500
rect 11412 7498 11468 7500
rect 11492 7498 11548 7500
rect 11252 7446 11278 7498
rect 11278 7446 11308 7498
rect 11332 7446 11342 7498
rect 11342 7446 11388 7498
rect 11412 7446 11458 7498
rect 11458 7446 11468 7498
rect 11492 7446 11522 7498
rect 11522 7446 11548 7498
rect 11252 7444 11308 7446
rect 11332 7444 11388 7446
rect 11412 7444 11468 7446
rect 11492 7444 11548 7446
rect 7820 6954 7876 6956
rect 7900 6954 7956 6956
rect 7980 6954 8036 6956
rect 8060 6954 8116 6956
rect 7820 6902 7846 6954
rect 7846 6902 7876 6954
rect 7900 6902 7910 6954
rect 7910 6902 7956 6954
rect 7980 6902 8026 6954
rect 8026 6902 8036 6954
rect 8060 6902 8090 6954
rect 8090 6902 8116 6954
rect 7820 6900 7876 6902
rect 7900 6900 7956 6902
rect 7980 6900 8036 6902
rect 8060 6900 8116 6902
rect 4388 6410 4444 6412
rect 4468 6410 4524 6412
rect 4548 6410 4604 6412
rect 4628 6410 4684 6412
rect 4388 6358 4414 6410
rect 4414 6358 4444 6410
rect 4468 6358 4478 6410
rect 4478 6358 4524 6410
rect 4548 6358 4594 6410
rect 4594 6358 4604 6410
rect 4628 6358 4658 6410
rect 4658 6358 4684 6410
rect 4388 6356 4444 6358
rect 4468 6356 4524 6358
rect 4548 6356 4604 6358
rect 4628 6356 4684 6358
rect 11252 6410 11308 6412
rect 11332 6410 11388 6412
rect 11412 6410 11468 6412
rect 11492 6410 11548 6412
rect 11252 6358 11278 6410
rect 11278 6358 11308 6410
rect 11332 6358 11342 6410
rect 11342 6358 11388 6410
rect 11412 6358 11458 6410
rect 11458 6358 11468 6410
rect 11492 6358 11522 6410
rect 11522 6358 11548 6410
rect 11252 6356 11308 6358
rect 11332 6356 11388 6358
rect 11412 6356 11468 6358
rect 11492 6356 11548 6358
rect 7820 5866 7876 5868
rect 7900 5866 7956 5868
rect 7980 5866 8036 5868
rect 8060 5866 8116 5868
rect 7820 5814 7846 5866
rect 7846 5814 7876 5866
rect 7900 5814 7910 5866
rect 7910 5814 7956 5866
rect 7980 5814 8026 5866
rect 8026 5814 8036 5866
rect 8060 5814 8090 5866
rect 8090 5814 8116 5866
rect 7820 5812 7876 5814
rect 7900 5812 7956 5814
rect 7980 5812 8036 5814
rect 8060 5812 8116 5814
rect 2962 5608 3018 5664
rect 4388 5322 4444 5324
rect 4468 5322 4524 5324
rect 4548 5322 4604 5324
rect 4628 5322 4684 5324
rect 4388 5270 4414 5322
rect 4414 5270 4444 5322
rect 4468 5270 4478 5322
rect 4478 5270 4524 5322
rect 4548 5270 4594 5322
rect 4594 5270 4604 5322
rect 4628 5270 4658 5322
rect 4658 5270 4684 5322
rect 4388 5268 4444 5270
rect 4468 5268 4524 5270
rect 4548 5268 4604 5270
rect 4628 5268 4684 5270
rect 11252 5322 11308 5324
rect 11332 5322 11388 5324
rect 11412 5322 11468 5324
rect 11492 5322 11548 5324
rect 11252 5270 11278 5322
rect 11278 5270 11308 5322
rect 11332 5270 11342 5322
rect 11342 5270 11388 5322
rect 11412 5270 11458 5322
rect 11458 5270 11468 5322
rect 11492 5270 11522 5322
rect 11522 5270 11548 5322
rect 11252 5268 11308 5270
rect 11332 5268 11388 5270
rect 11412 5268 11468 5270
rect 11492 5268 11548 5270
rect 7820 4778 7876 4780
rect 7900 4778 7956 4780
rect 7980 4778 8036 4780
rect 8060 4778 8116 4780
rect 7820 4726 7846 4778
rect 7846 4726 7876 4778
rect 7900 4726 7910 4778
rect 7910 4726 7956 4778
rect 7980 4726 8026 4778
rect 8026 4726 8036 4778
rect 8060 4726 8090 4778
rect 8090 4726 8116 4778
rect 7820 4724 7876 4726
rect 7900 4724 7956 4726
rect 7980 4724 8036 4726
rect 8060 4724 8116 4726
rect 4388 4234 4444 4236
rect 4468 4234 4524 4236
rect 4548 4234 4604 4236
rect 4628 4234 4684 4236
rect 4388 4182 4414 4234
rect 4414 4182 4444 4234
rect 4468 4182 4478 4234
rect 4478 4182 4524 4234
rect 4548 4182 4594 4234
rect 4594 4182 4604 4234
rect 4628 4182 4658 4234
rect 4658 4182 4684 4234
rect 4388 4180 4444 4182
rect 4468 4180 4524 4182
rect 4548 4180 4604 4182
rect 4628 4180 4684 4182
rect 11252 4234 11308 4236
rect 11332 4234 11388 4236
rect 11412 4234 11468 4236
rect 11492 4234 11548 4236
rect 11252 4182 11278 4234
rect 11278 4182 11308 4234
rect 11332 4182 11342 4234
rect 11342 4182 11388 4234
rect 11412 4182 11458 4234
rect 11458 4182 11468 4234
rect 11492 4182 11522 4234
rect 11522 4182 11548 4234
rect 11252 4180 11308 4182
rect 11332 4180 11388 4182
rect 11412 4180 11468 4182
rect 11492 4180 11548 4182
rect 14684 20010 14740 20012
rect 14764 20010 14820 20012
rect 14844 20010 14900 20012
rect 14924 20010 14980 20012
rect 14684 19958 14710 20010
rect 14710 19958 14740 20010
rect 14764 19958 14774 20010
rect 14774 19958 14820 20010
rect 14844 19958 14890 20010
rect 14890 19958 14900 20010
rect 14924 19958 14954 20010
rect 14954 19958 14980 20010
rect 14684 19956 14740 19958
rect 14764 19956 14820 19958
rect 14844 19956 14900 19958
rect 14924 19956 14980 19958
rect 14684 18922 14740 18924
rect 14764 18922 14820 18924
rect 14844 18922 14900 18924
rect 14924 18922 14980 18924
rect 14684 18870 14710 18922
rect 14710 18870 14740 18922
rect 14764 18870 14774 18922
rect 14774 18870 14820 18922
rect 14844 18870 14890 18922
rect 14890 18870 14900 18922
rect 14924 18870 14954 18922
rect 14954 18870 14980 18922
rect 14684 18868 14740 18870
rect 14764 18868 14820 18870
rect 14844 18868 14900 18870
rect 14924 18868 14980 18870
rect 14684 17834 14740 17836
rect 14764 17834 14820 17836
rect 14844 17834 14900 17836
rect 14924 17834 14980 17836
rect 14684 17782 14710 17834
rect 14710 17782 14740 17834
rect 14764 17782 14774 17834
rect 14774 17782 14820 17834
rect 14844 17782 14890 17834
rect 14890 17782 14900 17834
rect 14924 17782 14954 17834
rect 14954 17782 14980 17834
rect 14684 17780 14740 17782
rect 14764 17780 14820 17782
rect 14844 17780 14900 17782
rect 14924 17780 14980 17782
rect 14684 16746 14740 16748
rect 14764 16746 14820 16748
rect 14844 16746 14900 16748
rect 14924 16746 14980 16748
rect 14684 16694 14710 16746
rect 14710 16694 14740 16746
rect 14764 16694 14774 16746
rect 14774 16694 14820 16746
rect 14844 16694 14890 16746
rect 14890 16694 14900 16746
rect 14924 16694 14954 16746
rect 14954 16694 14980 16746
rect 14684 16692 14740 16694
rect 14764 16692 14820 16694
rect 14844 16692 14900 16694
rect 14924 16692 14980 16694
rect 14684 15658 14740 15660
rect 14764 15658 14820 15660
rect 14844 15658 14900 15660
rect 14924 15658 14980 15660
rect 14684 15606 14710 15658
rect 14710 15606 14740 15658
rect 14764 15606 14774 15658
rect 14774 15606 14820 15658
rect 14844 15606 14890 15658
rect 14890 15606 14900 15658
rect 14924 15606 14954 15658
rect 14954 15606 14980 15658
rect 14684 15604 14740 15606
rect 14764 15604 14820 15606
rect 14844 15604 14900 15606
rect 14924 15604 14980 15606
rect 14684 14570 14740 14572
rect 14764 14570 14820 14572
rect 14844 14570 14900 14572
rect 14924 14570 14980 14572
rect 14684 14518 14710 14570
rect 14710 14518 14740 14570
rect 14764 14518 14774 14570
rect 14774 14518 14820 14570
rect 14844 14518 14890 14570
rect 14890 14518 14900 14570
rect 14924 14518 14954 14570
rect 14954 14518 14980 14570
rect 14684 14516 14740 14518
rect 14764 14516 14820 14518
rect 14844 14516 14900 14518
rect 14924 14516 14980 14518
rect 14684 13482 14740 13484
rect 14764 13482 14820 13484
rect 14844 13482 14900 13484
rect 14924 13482 14980 13484
rect 14684 13430 14710 13482
rect 14710 13430 14740 13482
rect 14764 13430 14774 13482
rect 14774 13430 14820 13482
rect 14844 13430 14890 13482
rect 14890 13430 14900 13482
rect 14924 13430 14954 13482
rect 14954 13430 14980 13482
rect 14684 13428 14740 13430
rect 14764 13428 14820 13430
rect 14844 13428 14900 13430
rect 14924 13428 14980 13430
rect 14684 12394 14740 12396
rect 14764 12394 14820 12396
rect 14844 12394 14900 12396
rect 14924 12394 14980 12396
rect 14684 12342 14710 12394
rect 14710 12342 14740 12394
rect 14764 12342 14774 12394
rect 14774 12342 14820 12394
rect 14844 12342 14890 12394
rect 14890 12342 14900 12394
rect 14924 12342 14954 12394
rect 14954 12342 14980 12394
rect 14684 12340 14740 12342
rect 14764 12340 14820 12342
rect 14844 12340 14900 12342
rect 14924 12340 14980 12342
rect 14554 11456 14610 11512
rect 14684 11306 14740 11308
rect 14764 11306 14820 11308
rect 14844 11306 14900 11308
rect 14924 11306 14980 11308
rect 14684 11254 14710 11306
rect 14710 11254 14740 11306
rect 14764 11254 14774 11306
rect 14774 11254 14820 11306
rect 14844 11254 14890 11306
rect 14890 11254 14900 11306
rect 14924 11254 14954 11306
rect 14954 11254 14980 11306
rect 14684 11252 14740 11254
rect 14764 11252 14820 11254
rect 14844 11252 14900 11254
rect 14924 11252 14980 11254
rect 14684 10218 14740 10220
rect 14764 10218 14820 10220
rect 14844 10218 14900 10220
rect 14924 10218 14980 10220
rect 14684 10166 14710 10218
rect 14710 10166 14740 10218
rect 14764 10166 14774 10218
rect 14774 10166 14820 10218
rect 14844 10166 14890 10218
rect 14890 10166 14900 10218
rect 14924 10166 14954 10218
rect 14954 10166 14980 10218
rect 14684 10164 14740 10166
rect 14764 10164 14820 10166
rect 14844 10164 14900 10166
rect 14924 10164 14980 10166
rect 14684 9130 14740 9132
rect 14764 9130 14820 9132
rect 14844 9130 14900 9132
rect 14924 9130 14980 9132
rect 14684 9078 14710 9130
rect 14710 9078 14740 9130
rect 14764 9078 14774 9130
rect 14774 9078 14820 9130
rect 14844 9078 14890 9130
rect 14890 9078 14900 9130
rect 14924 9078 14954 9130
rect 14954 9078 14980 9130
rect 14684 9076 14740 9078
rect 14764 9076 14820 9078
rect 14844 9076 14900 9078
rect 14924 9076 14980 9078
rect 14684 8042 14740 8044
rect 14764 8042 14820 8044
rect 14844 8042 14900 8044
rect 14924 8042 14980 8044
rect 14684 7990 14710 8042
rect 14710 7990 14740 8042
rect 14764 7990 14774 8042
rect 14774 7990 14820 8042
rect 14844 7990 14890 8042
rect 14890 7990 14900 8042
rect 14924 7990 14954 8042
rect 14954 7990 14980 8042
rect 14684 7988 14740 7990
rect 14764 7988 14820 7990
rect 14844 7988 14900 7990
rect 14924 7988 14980 7990
rect 14684 6954 14740 6956
rect 14764 6954 14820 6956
rect 14844 6954 14900 6956
rect 14924 6954 14980 6956
rect 14684 6902 14710 6954
rect 14710 6902 14740 6954
rect 14764 6902 14774 6954
rect 14774 6902 14820 6954
rect 14844 6902 14890 6954
rect 14890 6902 14900 6954
rect 14924 6902 14954 6954
rect 14954 6902 14980 6954
rect 14684 6900 14740 6902
rect 14764 6900 14820 6902
rect 14844 6900 14900 6902
rect 14924 6900 14980 6902
rect 14684 5866 14740 5868
rect 14764 5866 14820 5868
rect 14844 5866 14900 5868
rect 14924 5866 14980 5868
rect 14684 5814 14710 5866
rect 14710 5814 14740 5866
rect 14764 5814 14774 5866
rect 14774 5814 14820 5866
rect 14844 5814 14890 5866
rect 14890 5814 14900 5866
rect 14924 5814 14954 5866
rect 14954 5814 14980 5866
rect 14684 5812 14740 5814
rect 14764 5812 14820 5814
rect 14844 5812 14900 5814
rect 14924 5812 14980 5814
rect 14684 4778 14740 4780
rect 14764 4778 14820 4780
rect 14844 4778 14900 4780
rect 14924 4778 14980 4780
rect 14684 4726 14710 4778
rect 14710 4726 14740 4778
rect 14764 4726 14774 4778
rect 14774 4726 14820 4778
rect 14844 4726 14890 4778
rect 14890 4726 14900 4778
rect 14924 4726 14954 4778
rect 14954 4726 14980 4778
rect 14684 4724 14740 4726
rect 14764 4724 14820 4726
rect 14844 4724 14900 4726
rect 14924 4724 14980 4726
rect 17866 21384 17922 21440
rect 18694 21928 18750 21984
rect 18116 19466 18172 19468
rect 18196 19466 18252 19468
rect 18276 19466 18332 19468
rect 18356 19466 18412 19468
rect 18116 19414 18142 19466
rect 18142 19414 18172 19466
rect 18196 19414 18206 19466
rect 18206 19414 18252 19466
rect 18276 19414 18322 19466
rect 18322 19414 18332 19466
rect 18356 19414 18386 19466
rect 18386 19414 18412 19466
rect 18116 19412 18172 19414
rect 18196 19412 18252 19414
rect 18276 19412 18332 19414
rect 18356 19412 18412 19414
rect 18116 18378 18172 18380
rect 18196 18378 18252 18380
rect 18276 18378 18332 18380
rect 18356 18378 18412 18380
rect 18116 18326 18142 18378
rect 18142 18326 18172 18378
rect 18196 18326 18206 18378
rect 18206 18326 18252 18378
rect 18276 18326 18322 18378
rect 18322 18326 18332 18378
rect 18356 18326 18386 18378
rect 18386 18326 18412 18378
rect 18116 18324 18172 18326
rect 18196 18324 18252 18326
rect 18276 18324 18332 18326
rect 18356 18324 18412 18326
rect 18116 17290 18172 17292
rect 18196 17290 18252 17292
rect 18276 17290 18332 17292
rect 18356 17290 18412 17292
rect 18116 17238 18142 17290
rect 18142 17238 18172 17290
rect 18196 17238 18206 17290
rect 18206 17238 18252 17290
rect 18276 17238 18322 17290
rect 18322 17238 18332 17290
rect 18356 17238 18386 17290
rect 18386 17238 18412 17290
rect 18116 17236 18172 17238
rect 18196 17236 18252 17238
rect 18276 17236 18332 17238
rect 18356 17236 18412 17238
rect 18116 16202 18172 16204
rect 18196 16202 18252 16204
rect 18276 16202 18332 16204
rect 18356 16202 18412 16204
rect 18116 16150 18142 16202
rect 18142 16150 18172 16202
rect 18196 16150 18206 16202
rect 18206 16150 18252 16202
rect 18276 16150 18322 16202
rect 18322 16150 18332 16202
rect 18356 16150 18386 16202
rect 18386 16150 18412 16202
rect 18116 16148 18172 16150
rect 18196 16148 18252 16150
rect 18276 16148 18332 16150
rect 18356 16148 18412 16150
rect 18116 15114 18172 15116
rect 18196 15114 18252 15116
rect 18276 15114 18332 15116
rect 18356 15114 18412 15116
rect 18116 15062 18142 15114
rect 18142 15062 18172 15114
rect 18196 15062 18206 15114
rect 18206 15062 18252 15114
rect 18276 15062 18322 15114
rect 18322 15062 18332 15114
rect 18356 15062 18386 15114
rect 18386 15062 18412 15114
rect 18116 15060 18172 15062
rect 18196 15060 18252 15062
rect 18276 15060 18332 15062
rect 18356 15060 18412 15062
rect 18116 14026 18172 14028
rect 18196 14026 18252 14028
rect 18276 14026 18332 14028
rect 18356 14026 18412 14028
rect 18116 13974 18142 14026
rect 18142 13974 18172 14026
rect 18196 13974 18206 14026
rect 18206 13974 18252 14026
rect 18276 13974 18322 14026
rect 18322 13974 18332 14026
rect 18356 13974 18386 14026
rect 18386 13974 18412 14026
rect 18116 13972 18172 13974
rect 18196 13972 18252 13974
rect 18276 13972 18332 13974
rect 18356 13972 18412 13974
rect 19614 19616 19670 19672
rect 19154 19208 19210 19264
rect 18694 17848 18750 17904
rect 19246 18664 19302 18720
rect 19338 18528 19394 18584
rect 7820 3690 7876 3692
rect 7900 3690 7956 3692
rect 7980 3690 8036 3692
rect 8060 3690 8116 3692
rect 7820 3638 7846 3690
rect 7846 3638 7876 3690
rect 7900 3638 7910 3690
rect 7910 3638 7956 3690
rect 7980 3638 8026 3690
rect 8026 3638 8036 3690
rect 8060 3638 8090 3690
rect 8090 3638 8116 3690
rect 7820 3636 7876 3638
rect 7900 3636 7956 3638
rect 7980 3636 8036 3638
rect 8060 3636 8116 3638
rect 14684 3690 14740 3692
rect 14764 3690 14820 3692
rect 14844 3690 14900 3692
rect 14924 3690 14980 3692
rect 14684 3638 14710 3690
rect 14710 3638 14740 3690
rect 14764 3638 14774 3690
rect 14774 3638 14820 3690
rect 14844 3638 14890 3690
rect 14890 3638 14900 3690
rect 14924 3638 14954 3690
rect 14954 3638 14980 3690
rect 14684 3636 14740 3638
rect 14764 3636 14820 3638
rect 14844 3636 14900 3638
rect 14924 3636 14980 3638
rect 4388 3146 4444 3148
rect 4468 3146 4524 3148
rect 4548 3146 4604 3148
rect 4628 3146 4684 3148
rect 4388 3094 4414 3146
rect 4414 3094 4444 3146
rect 4468 3094 4478 3146
rect 4478 3094 4524 3146
rect 4548 3094 4594 3146
rect 4594 3094 4604 3146
rect 4628 3094 4658 3146
rect 4658 3094 4684 3146
rect 4388 3092 4444 3094
rect 4468 3092 4524 3094
rect 4548 3092 4604 3094
rect 4628 3092 4684 3094
rect 11252 3146 11308 3148
rect 11332 3146 11388 3148
rect 11412 3146 11468 3148
rect 11492 3146 11548 3148
rect 11252 3094 11278 3146
rect 11278 3094 11308 3146
rect 11332 3094 11342 3146
rect 11342 3094 11388 3146
rect 11412 3094 11458 3146
rect 11458 3094 11468 3146
rect 11492 3094 11522 3146
rect 11522 3094 11548 3146
rect 11252 3092 11308 3094
rect 11332 3092 11388 3094
rect 11412 3092 11468 3094
rect 11492 3092 11548 3094
rect 7820 2602 7876 2604
rect 7900 2602 7956 2604
rect 7980 2602 8036 2604
rect 8060 2602 8116 2604
rect 7820 2550 7846 2602
rect 7846 2550 7876 2602
rect 7900 2550 7910 2602
rect 7910 2550 7956 2602
rect 7980 2550 8026 2602
rect 8026 2550 8036 2602
rect 8060 2550 8090 2602
rect 8090 2550 8116 2602
rect 7820 2548 7876 2550
rect 7900 2548 7956 2550
rect 7980 2548 8036 2550
rect 8060 2548 8116 2550
rect 14684 2602 14740 2604
rect 14764 2602 14820 2604
rect 14844 2602 14900 2604
rect 14924 2602 14980 2604
rect 14684 2550 14710 2602
rect 14710 2550 14740 2602
rect 14764 2550 14774 2602
rect 14774 2550 14820 2602
rect 14844 2550 14890 2602
rect 14890 2550 14900 2602
rect 14924 2550 14954 2602
rect 14954 2550 14980 2602
rect 14684 2548 14740 2550
rect 14764 2548 14820 2550
rect 14844 2548 14900 2550
rect 14924 2548 14980 2550
rect 4388 2058 4444 2060
rect 4468 2058 4524 2060
rect 4548 2058 4604 2060
rect 4628 2058 4684 2060
rect 4388 2006 4414 2058
rect 4414 2006 4444 2058
rect 4468 2006 4478 2058
rect 4478 2006 4524 2058
rect 4548 2006 4594 2058
rect 4594 2006 4604 2058
rect 4628 2006 4658 2058
rect 4658 2006 4684 2058
rect 4388 2004 4444 2006
rect 4468 2004 4524 2006
rect 4548 2004 4604 2006
rect 4628 2004 4684 2006
rect 11252 2058 11308 2060
rect 11332 2058 11388 2060
rect 11412 2058 11468 2060
rect 11492 2058 11548 2060
rect 11252 2006 11278 2058
rect 11278 2006 11308 2058
rect 11332 2006 11342 2058
rect 11342 2006 11388 2058
rect 11412 2006 11458 2058
rect 11458 2006 11468 2058
rect 11492 2006 11522 2058
rect 11522 2006 11548 2058
rect 11252 2004 11308 2006
rect 11332 2004 11388 2006
rect 11412 2004 11468 2006
rect 11492 2004 11548 2006
rect 18116 12938 18172 12940
rect 18196 12938 18252 12940
rect 18276 12938 18332 12940
rect 18356 12938 18412 12940
rect 18116 12886 18142 12938
rect 18142 12886 18172 12938
rect 18196 12886 18206 12938
rect 18206 12886 18252 12938
rect 18276 12886 18322 12938
rect 18322 12886 18332 12938
rect 18356 12886 18386 12938
rect 18386 12886 18412 12938
rect 18116 12884 18172 12886
rect 18196 12884 18252 12886
rect 18276 12884 18332 12886
rect 18356 12884 18412 12886
rect 19246 12272 19302 12328
rect 18116 11850 18172 11852
rect 18196 11850 18252 11852
rect 18276 11850 18332 11852
rect 18356 11850 18412 11852
rect 18116 11798 18142 11850
rect 18142 11798 18172 11850
rect 18196 11798 18206 11850
rect 18206 11798 18252 11850
rect 18276 11798 18322 11850
rect 18322 11798 18332 11850
rect 18356 11798 18386 11850
rect 18386 11798 18412 11850
rect 18116 11796 18172 11798
rect 18196 11796 18252 11798
rect 18276 11796 18332 11798
rect 18356 11796 18412 11798
rect 18116 10762 18172 10764
rect 18196 10762 18252 10764
rect 18276 10762 18332 10764
rect 18356 10762 18412 10764
rect 18116 10710 18142 10762
rect 18142 10710 18172 10762
rect 18196 10710 18206 10762
rect 18206 10710 18252 10762
rect 18276 10710 18322 10762
rect 18322 10710 18332 10762
rect 18356 10710 18386 10762
rect 18386 10710 18412 10762
rect 18116 10708 18172 10710
rect 18196 10708 18252 10710
rect 18276 10708 18332 10710
rect 18356 10708 18412 10710
rect 18116 9674 18172 9676
rect 18196 9674 18252 9676
rect 18276 9674 18332 9676
rect 18356 9674 18412 9676
rect 18116 9622 18142 9674
rect 18142 9622 18172 9674
rect 18196 9622 18206 9674
rect 18206 9622 18252 9674
rect 18276 9622 18322 9674
rect 18322 9622 18332 9674
rect 18356 9622 18386 9674
rect 18386 9622 18412 9674
rect 18116 9620 18172 9622
rect 18196 9620 18252 9622
rect 18276 9620 18332 9622
rect 18356 9620 18412 9622
rect 18116 8586 18172 8588
rect 18196 8586 18252 8588
rect 18276 8586 18332 8588
rect 18356 8586 18412 8588
rect 18116 8534 18142 8586
rect 18142 8534 18172 8586
rect 18196 8534 18206 8586
rect 18206 8534 18252 8586
rect 18276 8534 18322 8586
rect 18322 8534 18332 8586
rect 18356 8534 18386 8586
rect 18386 8534 18412 8586
rect 18116 8532 18172 8534
rect 18196 8532 18252 8534
rect 18276 8532 18332 8534
rect 18356 8532 18412 8534
rect 18116 7498 18172 7500
rect 18196 7498 18252 7500
rect 18276 7498 18332 7500
rect 18356 7498 18412 7500
rect 18116 7446 18142 7498
rect 18142 7446 18172 7498
rect 18196 7446 18206 7498
rect 18206 7446 18252 7498
rect 18276 7446 18322 7498
rect 18322 7446 18332 7498
rect 18356 7446 18386 7498
rect 18386 7446 18412 7498
rect 18116 7444 18172 7446
rect 18196 7444 18252 7446
rect 18276 7444 18332 7446
rect 18356 7444 18412 7446
rect 18510 6424 18566 6480
rect 18116 6410 18172 6412
rect 18196 6410 18252 6412
rect 18276 6410 18332 6412
rect 18356 6410 18412 6412
rect 18116 6358 18142 6410
rect 18142 6358 18172 6410
rect 18196 6358 18206 6410
rect 18206 6358 18252 6410
rect 18276 6358 18322 6410
rect 18322 6358 18332 6410
rect 18356 6358 18386 6410
rect 18386 6358 18412 6410
rect 18116 6356 18172 6358
rect 18196 6356 18252 6358
rect 18276 6356 18332 6358
rect 18356 6356 18412 6358
rect 17958 5472 18014 5528
rect 18116 5322 18172 5324
rect 18196 5322 18252 5324
rect 18276 5322 18332 5324
rect 18356 5322 18412 5324
rect 18116 5270 18142 5322
rect 18142 5270 18172 5322
rect 18196 5270 18206 5322
rect 18206 5270 18252 5322
rect 18276 5270 18322 5322
rect 18322 5270 18332 5322
rect 18356 5270 18386 5322
rect 18386 5270 18412 5322
rect 18116 5268 18172 5270
rect 18196 5268 18252 5270
rect 18276 5268 18332 5270
rect 18356 5268 18412 5270
rect 17958 4520 18014 4576
rect 18116 4234 18172 4236
rect 18196 4234 18252 4236
rect 18276 4234 18332 4236
rect 18356 4234 18412 4236
rect 18116 4182 18142 4234
rect 18142 4182 18172 4234
rect 18196 4182 18206 4234
rect 18206 4182 18252 4234
rect 18276 4182 18322 4234
rect 18322 4182 18332 4234
rect 18356 4182 18386 4234
rect 18386 4182 18412 4234
rect 18116 4180 18172 4182
rect 18196 4180 18252 4182
rect 18276 4180 18332 4182
rect 18356 4180 18412 4182
rect 17866 3568 17922 3624
rect 18510 3160 18566 3216
rect 18116 3146 18172 3148
rect 18196 3146 18252 3148
rect 18276 3146 18332 3148
rect 18356 3146 18412 3148
rect 18116 3094 18142 3146
rect 18142 3094 18172 3146
rect 18196 3094 18206 3146
rect 18206 3094 18252 3146
rect 18276 3094 18322 3146
rect 18322 3094 18332 3146
rect 18356 3094 18386 3146
rect 18386 3094 18412 3146
rect 18116 3092 18172 3094
rect 18196 3092 18252 3094
rect 18276 3092 18332 3094
rect 18356 3092 18412 3094
rect 18116 2058 18172 2060
rect 18196 2058 18252 2060
rect 18276 2058 18332 2060
rect 18356 2058 18412 2060
rect 18116 2006 18142 2058
rect 18142 2006 18172 2058
rect 18196 2006 18206 2058
rect 18206 2006 18252 2058
rect 18276 2006 18322 2058
rect 18322 2006 18332 2058
rect 18356 2006 18386 2058
rect 18386 2006 18412 2058
rect 18116 2004 18172 2006
rect 18196 2004 18252 2006
rect 18276 2004 18332 2006
rect 18356 2004 18412 2006
rect 18694 848 18750 904
rect 20166 20976 20222 21032
rect 20626 20568 20682 20624
rect 20534 20024 20590 20080
rect 20166 18276 20222 18312
rect 20166 18256 20168 18276
rect 20168 18256 20220 18276
rect 20220 18256 20222 18276
rect 20166 15944 20222 16000
rect 20442 17304 20498 17360
rect 20350 14584 20406 14640
rect 20718 16896 20774 16952
rect 20626 16352 20682 16408
rect 20718 15556 20774 15592
rect 20718 15536 20720 15556
rect 20720 15536 20772 15556
rect 20772 15536 20774 15556
rect 20718 14992 20774 15048
rect 20810 14176 20866 14232
rect 20442 13632 20498 13688
rect 20350 13224 20406 13280
rect 20258 12816 20314 12872
rect 19982 11864 20038 11920
rect 19982 10504 20038 10560
rect 18970 9960 19026 10016
rect 20258 10912 20314 10968
rect 20258 9552 20314 9608
rect 19982 8600 20038 8656
rect 20534 11456 20590 11512
rect 20718 13632 20774 13688
rect 20534 9144 20590 9200
rect 20534 8192 20590 8248
rect 20258 7784 20314 7840
rect 19982 7240 20038 7296
rect 20534 6832 20590 6888
rect 20534 5880 20590 5936
rect 20534 4928 20590 4984
rect 20534 4112 20590 4168
rect 19246 2752 19302 2808
rect 19062 2208 19118 2264
rect 19246 1800 19302 1856
rect 18878 1392 18934 1448
rect 18786 440 18842 496
rect 17958 32 18014 88
<< metal3 >>
rect 17953 22394 18019 22397
rect 22000 22394 22800 22424
rect 17953 22392 22800 22394
rect 17953 22336 17958 22392
rect 18014 22336 22800 22392
rect 17953 22334 22800 22336
rect 17953 22331 18019 22334
rect 22000 22304 22800 22334
rect 18689 21986 18755 21989
rect 22000 21986 22800 22016
rect 18689 21984 22800 21986
rect 18689 21928 18694 21984
rect 18750 21928 22800 21984
rect 18689 21926 22800 21928
rect 18689 21923 18755 21926
rect 22000 21896 22800 21926
rect 17861 21442 17927 21445
rect 22000 21442 22800 21472
rect 17861 21440 22800 21442
rect 17861 21384 17866 21440
rect 17922 21384 22800 21440
rect 17861 21382 22800 21384
rect 17861 21379 17927 21382
rect 22000 21352 22800 21382
rect 20161 21034 20227 21037
rect 22000 21034 22800 21064
rect 20161 21032 22800 21034
rect 20161 20976 20166 21032
rect 20222 20976 22800 21032
rect 20161 20974 22800 20976
rect 20161 20971 20227 20974
rect 22000 20944 22800 20974
rect 20621 20626 20687 20629
rect 22000 20626 22800 20656
rect 20621 20624 22800 20626
rect 20621 20568 20626 20624
rect 20682 20568 22800 20624
rect 20621 20566 22800 20568
rect 20621 20563 20687 20566
rect 22000 20536 22800 20566
rect 20529 20082 20595 20085
rect 22000 20082 22800 20112
rect 20529 20080 22800 20082
rect 20529 20024 20534 20080
rect 20590 20024 22800 20080
rect 20529 20022 22800 20024
rect 20529 20019 20595 20022
rect 7808 20016 8128 20017
rect 7808 19952 7816 20016
rect 7880 19952 7896 20016
rect 7960 19952 7976 20016
rect 8040 19952 8056 20016
rect 8120 19952 8128 20016
rect 7808 19951 8128 19952
rect 14672 20016 14992 20017
rect 14672 19952 14680 20016
rect 14744 19952 14760 20016
rect 14824 19952 14840 20016
rect 14904 19952 14920 20016
rect 14984 19952 14992 20016
rect 22000 19992 22800 20022
rect 14672 19951 14992 19952
rect 19609 19674 19675 19677
rect 22000 19674 22800 19704
rect 19609 19672 22800 19674
rect 19609 19616 19614 19672
rect 19670 19616 22800 19672
rect 19609 19614 22800 19616
rect 19609 19611 19675 19614
rect 22000 19584 22800 19614
rect 4376 19472 4696 19473
rect 4376 19408 4384 19472
rect 4448 19408 4464 19472
rect 4528 19408 4544 19472
rect 4608 19408 4624 19472
rect 4688 19408 4696 19472
rect 4376 19407 4696 19408
rect 11240 19472 11560 19473
rect 11240 19408 11248 19472
rect 11312 19408 11328 19472
rect 11392 19408 11408 19472
rect 11472 19408 11488 19472
rect 11552 19408 11560 19472
rect 11240 19407 11560 19408
rect 18104 19472 18424 19473
rect 18104 19408 18112 19472
rect 18176 19408 18192 19472
rect 18256 19408 18272 19472
rect 18336 19408 18352 19472
rect 18416 19408 18424 19472
rect 18104 19407 18424 19408
rect 19149 19266 19215 19269
rect 22000 19266 22800 19296
rect 19149 19264 22800 19266
rect 19149 19208 19154 19264
rect 19210 19208 22800 19264
rect 19149 19206 22800 19208
rect 19149 19203 19215 19206
rect 22000 19176 22800 19206
rect 7808 18928 8128 18929
rect 7808 18864 7816 18928
rect 7880 18864 7896 18928
rect 7960 18864 7976 18928
rect 8040 18864 8056 18928
rect 8120 18864 8128 18928
rect 7808 18863 8128 18864
rect 14672 18928 14992 18929
rect 14672 18864 14680 18928
rect 14744 18864 14760 18928
rect 14824 18864 14840 18928
rect 14904 18864 14920 18928
rect 14984 18864 14992 18928
rect 14672 18863 14992 18864
rect 5809 18722 5875 18725
rect 8109 18722 8175 18725
rect 5809 18720 8175 18722
rect 5809 18664 5814 18720
rect 5870 18664 8114 18720
rect 8170 18664 8175 18720
rect 5809 18662 8175 18664
rect 5809 18659 5875 18662
rect 8109 18659 8175 18662
rect 19241 18722 19307 18725
rect 22000 18722 22800 18752
rect 19241 18720 22800 18722
rect 19241 18664 19246 18720
rect 19302 18664 22800 18720
rect 19241 18662 22800 18664
rect 19241 18659 19307 18662
rect 22000 18632 22800 18662
rect 19333 18588 19399 18589
rect 19333 18584 19380 18588
rect 19444 18586 19450 18588
rect 19333 18528 19338 18584
rect 19333 18524 19380 18528
rect 19444 18526 19490 18586
rect 19444 18524 19450 18526
rect 19333 18523 19399 18524
rect 4376 18384 4696 18385
rect 4376 18320 4384 18384
rect 4448 18320 4464 18384
rect 4528 18320 4544 18384
rect 4608 18320 4624 18384
rect 4688 18320 4696 18384
rect 4376 18319 4696 18320
rect 11240 18384 11560 18385
rect 11240 18320 11248 18384
rect 11312 18320 11328 18384
rect 11392 18320 11408 18384
rect 11472 18320 11488 18384
rect 11552 18320 11560 18384
rect 11240 18319 11560 18320
rect 18104 18384 18424 18385
rect 18104 18320 18112 18384
rect 18176 18320 18192 18384
rect 18256 18320 18272 18384
rect 18336 18320 18352 18384
rect 18416 18320 18424 18384
rect 18104 18319 18424 18320
rect 20161 18314 20227 18317
rect 22000 18314 22800 18344
rect 20161 18312 22800 18314
rect 20161 18256 20166 18312
rect 20222 18256 22800 18312
rect 20161 18254 22800 18256
rect 20161 18251 20227 18254
rect 22000 18224 22800 18254
rect 18689 17906 18755 17909
rect 22000 17906 22800 17936
rect 18689 17904 22800 17906
rect 18689 17848 18694 17904
rect 18750 17848 22800 17904
rect 18689 17846 22800 17848
rect 18689 17843 18755 17846
rect 7808 17840 8128 17841
rect 7808 17776 7816 17840
rect 7880 17776 7896 17840
rect 7960 17776 7976 17840
rect 8040 17776 8056 17840
rect 8120 17776 8128 17840
rect 7808 17775 8128 17776
rect 14672 17840 14992 17841
rect 14672 17776 14680 17840
rect 14744 17776 14760 17840
rect 14824 17776 14840 17840
rect 14904 17776 14920 17840
rect 14984 17776 14992 17840
rect 22000 17816 22800 17846
rect 14672 17775 14992 17776
rect 20437 17362 20503 17365
rect 22000 17362 22800 17392
rect 20437 17360 22800 17362
rect 20437 17304 20442 17360
rect 20498 17304 22800 17360
rect 20437 17302 22800 17304
rect 20437 17299 20503 17302
rect 4376 17296 4696 17297
rect 4376 17232 4384 17296
rect 4448 17232 4464 17296
rect 4528 17232 4544 17296
rect 4608 17232 4624 17296
rect 4688 17232 4696 17296
rect 4376 17231 4696 17232
rect 11240 17296 11560 17297
rect 11240 17232 11248 17296
rect 11312 17232 11328 17296
rect 11392 17232 11408 17296
rect 11472 17232 11488 17296
rect 11552 17232 11560 17296
rect 11240 17231 11560 17232
rect 18104 17296 18424 17297
rect 18104 17232 18112 17296
rect 18176 17232 18192 17296
rect 18256 17232 18272 17296
rect 18336 17232 18352 17296
rect 18416 17232 18424 17296
rect 22000 17272 22800 17302
rect 18104 17231 18424 17232
rect 0 17090 800 17120
rect 4061 17090 4127 17093
rect 0 17088 4127 17090
rect 0 17032 4066 17088
rect 4122 17032 4127 17088
rect 0 17030 4127 17032
rect 0 17000 800 17030
rect 4061 17027 4127 17030
rect 20713 16954 20779 16957
rect 22000 16954 22800 16984
rect 20713 16952 22800 16954
rect 20713 16896 20718 16952
rect 20774 16896 22800 16952
rect 20713 16894 22800 16896
rect 20713 16891 20779 16894
rect 22000 16864 22800 16894
rect 7808 16752 8128 16753
rect 7808 16688 7816 16752
rect 7880 16688 7896 16752
rect 7960 16688 7976 16752
rect 8040 16688 8056 16752
rect 8120 16688 8128 16752
rect 7808 16687 8128 16688
rect 14672 16752 14992 16753
rect 14672 16688 14680 16752
rect 14744 16688 14760 16752
rect 14824 16688 14840 16752
rect 14904 16688 14920 16752
rect 14984 16688 14992 16752
rect 14672 16687 14992 16688
rect 20621 16410 20687 16413
rect 22000 16410 22800 16440
rect 20621 16408 22800 16410
rect 20621 16352 20626 16408
rect 20682 16352 22800 16408
rect 20621 16350 22800 16352
rect 20621 16347 20687 16350
rect 22000 16320 22800 16350
rect 4376 16208 4696 16209
rect 4376 16144 4384 16208
rect 4448 16144 4464 16208
rect 4528 16144 4544 16208
rect 4608 16144 4624 16208
rect 4688 16144 4696 16208
rect 4376 16143 4696 16144
rect 11240 16208 11560 16209
rect 11240 16144 11248 16208
rect 11312 16144 11328 16208
rect 11392 16144 11408 16208
rect 11472 16144 11488 16208
rect 11552 16144 11560 16208
rect 11240 16143 11560 16144
rect 18104 16208 18424 16209
rect 18104 16144 18112 16208
rect 18176 16144 18192 16208
rect 18256 16144 18272 16208
rect 18336 16144 18352 16208
rect 18416 16144 18424 16208
rect 18104 16143 18424 16144
rect 20161 16002 20227 16005
rect 22000 16002 22800 16032
rect 20161 16000 22800 16002
rect 20161 15944 20166 16000
rect 20222 15944 22800 16000
rect 20161 15942 22800 15944
rect 20161 15939 20227 15942
rect 22000 15912 22800 15942
rect 7808 15664 8128 15665
rect 7808 15600 7816 15664
rect 7880 15600 7896 15664
rect 7960 15600 7976 15664
rect 8040 15600 8056 15664
rect 8120 15600 8128 15664
rect 7808 15599 8128 15600
rect 14672 15664 14992 15665
rect 14672 15600 14680 15664
rect 14744 15600 14760 15664
rect 14824 15600 14840 15664
rect 14904 15600 14920 15664
rect 14984 15600 14992 15664
rect 14672 15599 14992 15600
rect 20713 15594 20779 15597
rect 22000 15594 22800 15624
rect 20713 15592 22800 15594
rect 20713 15536 20718 15592
rect 20774 15536 22800 15592
rect 20713 15534 22800 15536
rect 20713 15531 20779 15534
rect 22000 15504 22800 15534
rect 4376 15120 4696 15121
rect 4376 15056 4384 15120
rect 4448 15056 4464 15120
rect 4528 15056 4544 15120
rect 4608 15056 4624 15120
rect 4688 15056 4696 15120
rect 4376 15055 4696 15056
rect 11240 15120 11560 15121
rect 11240 15056 11248 15120
rect 11312 15056 11328 15120
rect 11392 15056 11408 15120
rect 11472 15056 11488 15120
rect 11552 15056 11560 15120
rect 11240 15055 11560 15056
rect 18104 15120 18424 15121
rect 18104 15056 18112 15120
rect 18176 15056 18192 15120
rect 18256 15056 18272 15120
rect 18336 15056 18352 15120
rect 18416 15056 18424 15120
rect 18104 15055 18424 15056
rect 20713 15050 20779 15053
rect 22000 15050 22800 15080
rect 20713 15048 22800 15050
rect 20713 14992 20718 15048
rect 20774 14992 22800 15048
rect 20713 14990 22800 14992
rect 20713 14987 20779 14990
rect 22000 14960 22800 14990
rect 20345 14642 20411 14645
rect 22000 14642 22800 14672
rect 20345 14640 22800 14642
rect 20345 14584 20350 14640
rect 20406 14584 22800 14640
rect 20345 14582 22800 14584
rect 20345 14579 20411 14582
rect 7808 14576 8128 14577
rect 7808 14512 7816 14576
rect 7880 14512 7896 14576
rect 7960 14512 7976 14576
rect 8040 14512 8056 14576
rect 8120 14512 8128 14576
rect 7808 14511 8128 14512
rect 14672 14576 14992 14577
rect 14672 14512 14680 14576
rect 14744 14512 14760 14576
rect 14824 14512 14840 14576
rect 14904 14512 14920 14576
rect 14984 14512 14992 14576
rect 22000 14552 22800 14582
rect 14672 14511 14992 14512
rect 20805 14234 20871 14237
rect 22000 14234 22800 14264
rect 20805 14232 22800 14234
rect 20805 14176 20810 14232
rect 20866 14176 22800 14232
rect 20805 14174 22800 14176
rect 20805 14171 20871 14174
rect 22000 14144 22800 14174
rect 4376 14032 4696 14033
rect 4376 13968 4384 14032
rect 4448 13968 4464 14032
rect 4528 13968 4544 14032
rect 4608 13968 4624 14032
rect 4688 13968 4696 14032
rect 4376 13967 4696 13968
rect 11240 14032 11560 14033
rect 11240 13968 11248 14032
rect 11312 13968 11328 14032
rect 11392 13968 11408 14032
rect 11472 13968 11488 14032
rect 11552 13968 11560 14032
rect 11240 13967 11560 13968
rect 18104 14032 18424 14033
rect 18104 13968 18112 14032
rect 18176 13968 18192 14032
rect 18256 13968 18272 14032
rect 18336 13968 18352 14032
rect 18416 13968 18424 14032
rect 18104 13967 18424 13968
rect 19374 13628 19380 13692
rect 19444 13690 19450 13692
rect 20437 13690 20503 13693
rect 19444 13688 20503 13690
rect 19444 13632 20442 13688
rect 20498 13632 20503 13688
rect 19444 13630 20503 13632
rect 19444 13628 19450 13630
rect 20437 13627 20503 13630
rect 20713 13690 20779 13693
rect 22000 13690 22800 13720
rect 20713 13688 22800 13690
rect 20713 13632 20718 13688
rect 20774 13632 22800 13688
rect 20713 13630 22800 13632
rect 20713 13627 20779 13630
rect 22000 13600 22800 13630
rect 7808 13488 8128 13489
rect 7808 13424 7816 13488
rect 7880 13424 7896 13488
rect 7960 13424 7976 13488
rect 8040 13424 8056 13488
rect 8120 13424 8128 13488
rect 7808 13423 8128 13424
rect 14672 13488 14992 13489
rect 14672 13424 14680 13488
rect 14744 13424 14760 13488
rect 14824 13424 14840 13488
rect 14904 13424 14920 13488
rect 14984 13424 14992 13488
rect 14672 13423 14992 13424
rect 20345 13282 20411 13285
rect 22000 13282 22800 13312
rect 20345 13280 22800 13282
rect 20345 13224 20350 13280
rect 20406 13224 22800 13280
rect 20345 13222 22800 13224
rect 20345 13219 20411 13222
rect 22000 13192 22800 13222
rect 4376 12944 4696 12945
rect 4376 12880 4384 12944
rect 4448 12880 4464 12944
rect 4528 12880 4544 12944
rect 4608 12880 4624 12944
rect 4688 12880 4696 12944
rect 4376 12879 4696 12880
rect 11240 12944 11560 12945
rect 11240 12880 11248 12944
rect 11312 12880 11328 12944
rect 11392 12880 11408 12944
rect 11472 12880 11488 12944
rect 11552 12880 11560 12944
rect 11240 12879 11560 12880
rect 18104 12944 18424 12945
rect 18104 12880 18112 12944
rect 18176 12880 18192 12944
rect 18256 12880 18272 12944
rect 18336 12880 18352 12944
rect 18416 12880 18424 12944
rect 18104 12879 18424 12880
rect 20253 12874 20319 12877
rect 22000 12874 22800 12904
rect 20253 12872 22800 12874
rect 20253 12816 20258 12872
rect 20314 12816 22800 12872
rect 20253 12814 22800 12816
rect 20253 12811 20319 12814
rect 22000 12784 22800 12814
rect 7808 12400 8128 12401
rect 7808 12336 7816 12400
rect 7880 12336 7896 12400
rect 7960 12336 7976 12400
rect 8040 12336 8056 12400
rect 8120 12336 8128 12400
rect 7808 12335 8128 12336
rect 14672 12400 14992 12401
rect 14672 12336 14680 12400
rect 14744 12336 14760 12400
rect 14824 12336 14840 12400
rect 14904 12336 14920 12400
rect 14984 12336 14992 12400
rect 14672 12335 14992 12336
rect 19241 12330 19307 12333
rect 22000 12330 22800 12360
rect 19241 12328 22800 12330
rect 19241 12272 19246 12328
rect 19302 12272 22800 12328
rect 19241 12270 22800 12272
rect 19241 12267 19307 12270
rect 22000 12240 22800 12270
rect 19977 11922 20043 11925
rect 22000 11922 22800 11952
rect 19977 11920 22800 11922
rect 19977 11864 19982 11920
rect 20038 11864 22800 11920
rect 19977 11862 22800 11864
rect 19977 11859 20043 11862
rect 4376 11856 4696 11857
rect 4376 11792 4384 11856
rect 4448 11792 4464 11856
rect 4528 11792 4544 11856
rect 4608 11792 4624 11856
rect 4688 11792 4696 11856
rect 4376 11791 4696 11792
rect 11240 11856 11560 11857
rect 11240 11792 11248 11856
rect 11312 11792 11328 11856
rect 11392 11792 11408 11856
rect 11472 11792 11488 11856
rect 11552 11792 11560 11856
rect 11240 11791 11560 11792
rect 18104 11856 18424 11857
rect 18104 11792 18112 11856
rect 18176 11792 18192 11856
rect 18256 11792 18272 11856
rect 18336 11792 18352 11856
rect 18416 11792 18424 11856
rect 22000 11832 22800 11862
rect 18104 11791 18424 11792
rect 10593 11514 10659 11517
rect 14549 11514 14615 11517
rect 10593 11512 14615 11514
rect 10593 11456 10598 11512
rect 10654 11456 14554 11512
rect 14610 11456 14615 11512
rect 10593 11454 14615 11456
rect 10593 11451 10659 11454
rect 14549 11451 14615 11454
rect 20529 11514 20595 11517
rect 22000 11514 22800 11544
rect 20529 11512 22800 11514
rect 20529 11456 20534 11512
rect 20590 11456 22800 11512
rect 20529 11454 22800 11456
rect 20529 11451 20595 11454
rect 22000 11424 22800 11454
rect 7808 11312 8128 11313
rect 7808 11248 7816 11312
rect 7880 11248 7896 11312
rect 7960 11248 7976 11312
rect 8040 11248 8056 11312
rect 8120 11248 8128 11312
rect 7808 11247 8128 11248
rect 14672 11312 14992 11313
rect 14672 11248 14680 11312
rect 14744 11248 14760 11312
rect 14824 11248 14840 11312
rect 14904 11248 14920 11312
rect 14984 11248 14992 11312
rect 14672 11247 14992 11248
rect 20253 10970 20319 10973
rect 22000 10970 22800 11000
rect 20253 10968 22800 10970
rect 20253 10912 20258 10968
rect 20314 10912 22800 10968
rect 20253 10910 22800 10912
rect 20253 10907 20319 10910
rect 22000 10880 22800 10910
rect 4376 10768 4696 10769
rect 4376 10704 4384 10768
rect 4448 10704 4464 10768
rect 4528 10704 4544 10768
rect 4608 10704 4624 10768
rect 4688 10704 4696 10768
rect 4376 10703 4696 10704
rect 11240 10768 11560 10769
rect 11240 10704 11248 10768
rect 11312 10704 11328 10768
rect 11392 10704 11408 10768
rect 11472 10704 11488 10768
rect 11552 10704 11560 10768
rect 11240 10703 11560 10704
rect 18104 10768 18424 10769
rect 18104 10704 18112 10768
rect 18176 10704 18192 10768
rect 18256 10704 18272 10768
rect 18336 10704 18352 10768
rect 18416 10704 18424 10768
rect 18104 10703 18424 10704
rect 19977 10562 20043 10565
rect 22000 10562 22800 10592
rect 19977 10560 22800 10562
rect 19977 10504 19982 10560
rect 20038 10504 22800 10560
rect 19977 10502 22800 10504
rect 19977 10499 20043 10502
rect 22000 10472 22800 10502
rect 7808 10224 8128 10225
rect 7808 10160 7816 10224
rect 7880 10160 7896 10224
rect 7960 10160 7976 10224
rect 8040 10160 8056 10224
rect 8120 10160 8128 10224
rect 7808 10159 8128 10160
rect 14672 10224 14992 10225
rect 14672 10160 14680 10224
rect 14744 10160 14760 10224
rect 14824 10160 14840 10224
rect 14904 10160 14920 10224
rect 14984 10160 14992 10224
rect 14672 10159 14992 10160
rect 18965 10018 19031 10021
rect 22000 10018 22800 10048
rect 18965 10016 22800 10018
rect 18965 9960 18970 10016
rect 19026 9960 22800 10016
rect 18965 9958 22800 9960
rect 18965 9955 19031 9958
rect 22000 9928 22800 9958
rect 4376 9680 4696 9681
rect 4376 9616 4384 9680
rect 4448 9616 4464 9680
rect 4528 9616 4544 9680
rect 4608 9616 4624 9680
rect 4688 9616 4696 9680
rect 4376 9615 4696 9616
rect 11240 9680 11560 9681
rect 11240 9616 11248 9680
rect 11312 9616 11328 9680
rect 11392 9616 11408 9680
rect 11472 9616 11488 9680
rect 11552 9616 11560 9680
rect 11240 9615 11560 9616
rect 18104 9680 18424 9681
rect 18104 9616 18112 9680
rect 18176 9616 18192 9680
rect 18256 9616 18272 9680
rect 18336 9616 18352 9680
rect 18416 9616 18424 9680
rect 18104 9615 18424 9616
rect 20253 9610 20319 9613
rect 22000 9610 22800 9640
rect 20253 9608 22800 9610
rect 20253 9552 20258 9608
rect 20314 9552 22800 9608
rect 20253 9550 22800 9552
rect 20253 9547 20319 9550
rect 22000 9520 22800 9550
rect 20529 9202 20595 9205
rect 22000 9202 22800 9232
rect 20529 9200 22800 9202
rect 20529 9144 20534 9200
rect 20590 9144 22800 9200
rect 20529 9142 22800 9144
rect 20529 9139 20595 9142
rect 7808 9136 8128 9137
rect 7808 9072 7816 9136
rect 7880 9072 7896 9136
rect 7960 9072 7976 9136
rect 8040 9072 8056 9136
rect 8120 9072 8128 9136
rect 7808 9071 8128 9072
rect 14672 9136 14992 9137
rect 14672 9072 14680 9136
rect 14744 9072 14760 9136
rect 14824 9072 14840 9136
rect 14904 9072 14920 9136
rect 14984 9072 14992 9136
rect 22000 9112 22800 9142
rect 14672 9071 14992 9072
rect 19977 8658 20043 8661
rect 22000 8658 22800 8688
rect 19977 8656 22800 8658
rect 19977 8600 19982 8656
rect 20038 8600 22800 8656
rect 19977 8598 22800 8600
rect 19977 8595 20043 8598
rect 4376 8592 4696 8593
rect 4376 8528 4384 8592
rect 4448 8528 4464 8592
rect 4528 8528 4544 8592
rect 4608 8528 4624 8592
rect 4688 8528 4696 8592
rect 4376 8527 4696 8528
rect 11240 8592 11560 8593
rect 11240 8528 11248 8592
rect 11312 8528 11328 8592
rect 11392 8528 11408 8592
rect 11472 8528 11488 8592
rect 11552 8528 11560 8592
rect 11240 8527 11560 8528
rect 18104 8592 18424 8593
rect 18104 8528 18112 8592
rect 18176 8528 18192 8592
rect 18256 8528 18272 8592
rect 18336 8528 18352 8592
rect 18416 8528 18424 8592
rect 22000 8568 22800 8598
rect 18104 8527 18424 8528
rect 20529 8250 20595 8253
rect 22000 8250 22800 8280
rect 20529 8248 22800 8250
rect 20529 8192 20534 8248
rect 20590 8192 22800 8248
rect 20529 8190 22800 8192
rect 20529 8187 20595 8190
rect 22000 8160 22800 8190
rect 7808 8048 8128 8049
rect 7808 7984 7816 8048
rect 7880 7984 7896 8048
rect 7960 7984 7976 8048
rect 8040 7984 8056 8048
rect 8120 7984 8128 8048
rect 7808 7983 8128 7984
rect 14672 8048 14992 8049
rect 14672 7984 14680 8048
rect 14744 7984 14760 8048
rect 14824 7984 14840 8048
rect 14904 7984 14920 8048
rect 14984 7984 14992 8048
rect 14672 7983 14992 7984
rect 20253 7842 20319 7845
rect 22000 7842 22800 7872
rect 20253 7840 22800 7842
rect 20253 7784 20258 7840
rect 20314 7784 22800 7840
rect 20253 7782 22800 7784
rect 20253 7779 20319 7782
rect 22000 7752 22800 7782
rect 4376 7504 4696 7505
rect 4376 7440 4384 7504
rect 4448 7440 4464 7504
rect 4528 7440 4544 7504
rect 4608 7440 4624 7504
rect 4688 7440 4696 7504
rect 4376 7439 4696 7440
rect 11240 7504 11560 7505
rect 11240 7440 11248 7504
rect 11312 7440 11328 7504
rect 11392 7440 11408 7504
rect 11472 7440 11488 7504
rect 11552 7440 11560 7504
rect 11240 7439 11560 7440
rect 18104 7504 18424 7505
rect 18104 7440 18112 7504
rect 18176 7440 18192 7504
rect 18256 7440 18272 7504
rect 18336 7440 18352 7504
rect 18416 7440 18424 7504
rect 18104 7439 18424 7440
rect 19977 7298 20043 7301
rect 22000 7298 22800 7328
rect 19977 7296 22800 7298
rect 19977 7240 19982 7296
rect 20038 7240 22800 7296
rect 19977 7238 22800 7240
rect 19977 7235 20043 7238
rect 22000 7208 22800 7238
rect 7808 6960 8128 6961
rect 7808 6896 7816 6960
rect 7880 6896 7896 6960
rect 7960 6896 7976 6960
rect 8040 6896 8056 6960
rect 8120 6896 8128 6960
rect 7808 6895 8128 6896
rect 14672 6960 14992 6961
rect 14672 6896 14680 6960
rect 14744 6896 14760 6960
rect 14824 6896 14840 6960
rect 14904 6896 14920 6960
rect 14984 6896 14992 6960
rect 14672 6895 14992 6896
rect 20529 6890 20595 6893
rect 22000 6890 22800 6920
rect 20529 6888 22800 6890
rect 20529 6832 20534 6888
rect 20590 6832 22800 6888
rect 20529 6830 22800 6832
rect 20529 6827 20595 6830
rect 22000 6800 22800 6830
rect 18505 6482 18571 6485
rect 22000 6482 22800 6512
rect 18505 6480 22800 6482
rect 18505 6424 18510 6480
rect 18566 6424 22800 6480
rect 18505 6422 22800 6424
rect 18505 6419 18571 6422
rect 4376 6416 4696 6417
rect 4376 6352 4384 6416
rect 4448 6352 4464 6416
rect 4528 6352 4544 6416
rect 4608 6352 4624 6416
rect 4688 6352 4696 6416
rect 4376 6351 4696 6352
rect 11240 6416 11560 6417
rect 11240 6352 11248 6416
rect 11312 6352 11328 6416
rect 11392 6352 11408 6416
rect 11472 6352 11488 6416
rect 11552 6352 11560 6416
rect 11240 6351 11560 6352
rect 18104 6416 18424 6417
rect 18104 6352 18112 6416
rect 18176 6352 18192 6416
rect 18256 6352 18272 6416
rect 18336 6352 18352 6416
rect 18416 6352 18424 6416
rect 22000 6392 22800 6422
rect 18104 6351 18424 6352
rect 20529 5938 20595 5941
rect 22000 5938 22800 5968
rect 20529 5936 22800 5938
rect 20529 5880 20534 5936
rect 20590 5880 22800 5936
rect 20529 5878 22800 5880
rect 20529 5875 20595 5878
rect 7808 5872 8128 5873
rect 7808 5808 7816 5872
rect 7880 5808 7896 5872
rect 7960 5808 7976 5872
rect 8040 5808 8056 5872
rect 8120 5808 8128 5872
rect 7808 5807 8128 5808
rect 14672 5872 14992 5873
rect 14672 5808 14680 5872
rect 14744 5808 14760 5872
rect 14824 5808 14840 5872
rect 14904 5808 14920 5872
rect 14984 5808 14992 5872
rect 22000 5848 22800 5878
rect 14672 5807 14992 5808
rect 0 5666 800 5696
rect 2957 5666 3023 5669
rect 0 5664 3023 5666
rect 0 5608 2962 5664
rect 3018 5608 3023 5664
rect 0 5606 3023 5608
rect 0 5576 800 5606
rect 2957 5603 3023 5606
rect 17953 5530 18019 5533
rect 22000 5530 22800 5560
rect 17953 5528 22800 5530
rect 17953 5472 17958 5528
rect 18014 5472 22800 5528
rect 17953 5470 22800 5472
rect 17953 5467 18019 5470
rect 22000 5440 22800 5470
rect 4376 5328 4696 5329
rect 4376 5264 4384 5328
rect 4448 5264 4464 5328
rect 4528 5264 4544 5328
rect 4608 5264 4624 5328
rect 4688 5264 4696 5328
rect 4376 5263 4696 5264
rect 11240 5328 11560 5329
rect 11240 5264 11248 5328
rect 11312 5264 11328 5328
rect 11392 5264 11408 5328
rect 11472 5264 11488 5328
rect 11552 5264 11560 5328
rect 11240 5263 11560 5264
rect 18104 5328 18424 5329
rect 18104 5264 18112 5328
rect 18176 5264 18192 5328
rect 18256 5264 18272 5328
rect 18336 5264 18352 5328
rect 18416 5264 18424 5328
rect 18104 5263 18424 5264
rect 20529 4986 20595 4989
rect 22000 4986 22800 5016
rect 20529 4984 22800 4986
rect 20529 4928 20534 4984
rect 20590 4928 22800 4984
rect 20529 4926 22800 4928
rect 20529 4923 20595 4926
rect 22000 4896 22800 4926
rect 7808 4784 8128 4785
rect 7808 4720 7816 4784
rect 7880 4720 7896 4784
rect 7960 4720 7976 4784
rect 8040 4720 8056 4784
rect 8120 4720 8128 4784
rect 7808 4719 8128 4720
rect 14672 4784 14992 4785
rect 14672 4720 14680 4784
rect 14744 4720 14760 4784
rect 14824 4720 14840 4784
rect 14904 4720 14920 4784
rect 14984 4720 14992 4784
rect 14672 4719 14992 4720
rect 17953 4578 18019 4581
rect 22000 4578 22800 4608
rect 17953 4576 22800 4578
rect 17953 4520 17958 4576
rect 18014 4520 22800 4576
rect 17953 4518 22800 4520
rect 17953 4515 18019 4518
rect 22000 4488 22800 4518
rect 4376 4240 4696 4241
rect 4376 4176 4384 4240
rect 4448 4176 4464 4240
rect 4528 4176 4544 4240
rect 4608 4176 4624 4240
rect 4688 4176 4696 4240
rect 4376 4175 4696 4176
rect 11240 4240 11560 4241
rect 11240 4176 11248 4240
rect 11312 4176 11328 4240
rect 11392 4176 11408 4240
rect 11472 4176 11488 4240
rect 11552 4176 11560 4240
rect 11240 4175 11560 4176
rect 18104 4240 18424 4241
rect 18104 4176 18112 4240
rect 18176 4176 18192 4240
rect 18256 4176 18272 4240
rect 18336 4176 18352 4240
rect 18416 4176 18424 4240
rect 18104 4175 18424 4176
rect 20529 4170 20595 4173
rect 22000 4170 22800 4200
rect 20529 4168 22800 4170
rect 20529 4112 20534 4168
rect 20590 4112 22800 4168
rect 20529 4110 22800 4112
rect 20529 4107 20595 4110
rect 22000 4080 22800 4110
rect 7808 3696 8128 3697
rect 7808 3632 7816 3696
rect 7880 3632 7896 3696
rect 7960 3632 7976 3696
rect 8040 3632 8056 3696
rect 8120 3632 8128 3696
rect 7808 3631 8128 3632
rect 14672 3696 14992 3697
rect 14672 3632 14680 3696
rect 14744 3632 14760 3696
rect 14824 3632 14840 3696
rect 14904 3632 14920 3696
rect 14984 3632 14992 3696
rect 14672 3631 14992 3632
rect 17861 3626 17927 3629
rect 22000 3626 22800 3656
rect 17861 3624 22800 3626
rect 17861 3568 17866 3624
rect 17922 3568 22800 3624
rect 17861 3566 22800 3568
rect 17861 3563 17927 3566
rect 22000 3536 22800 3566
rect 18505 3218 18571 3221
rect 22000 3218 22800 3248
rect 18505 3216 22800 3218
rect 18505 3160 18510 3216
rect 18566 3160 22800 3216
rect 18505 3158 22800 3160
rect 18505 3155 18571 3158
rect 4376 3152 4696 3153
rect 4376 3088 4384 3152
rect 4448 3088 4464 3152
rect 4528 3088 4544 3152
rect 4608 3088 4624 3152
rect 4688 3088 4696 3152
rect 4376 3087 4696 3088
rect 11240 3152 11560 3153
rect 11240 3088 11248 3152
rect 11312 3088 11328 3152
rect 11392 3088 11408 3152
rect 11472 3088 11488 3152
rect 11552 3088 11560 3152
rect 11240 3087 11560 3088
rect 18104 3152 18424 3153
rect 18104 3088 18112 3152
rect 18176 3088 18192 3152
rect 18256 3088 18272 3152
rect 18336 3088 18352 3152
rect 18416 3088 18424 3152
rect 22000 3128 22800 3158
rect 18104 3087 18424 3088
rect 19241 2810 19307 2813
rect 22000 2810 22800 2840
rect 19241 2808 22800 2810
rect 19241 2752 19246 2808
rect 19302 2752 22800 2808
rect 19241 2750 22800 2752
rect 19241 2747 19307 2750
rect 22000 2720 22800 2750
rect 7808 2608 8128 2609
rect 7808 2544 7816 2608
rect 7880 2544 7896 2608
rect 7960 2544 7976 2608
rect 8040 2544 8056 2608
rect 8120 2544 8128 2608
rect 7808 2543 8128 2544
rect 14672 2608 14992 2609
rect 14672 2544 14680 2608
rect 14744 2544 14760 2608
rect 14824 2544 14840 2608
rect 14904 2544 14920 2608
rect 14984 2544 14992 2608
rect 14672 2543 14992 2544
rect 19057 2266 19123 2269
rect 22000 2266 22800 2296
rect 19057 2264 22800 2266
rect 19057 2208 19062 2264
rect 19118 2208 22800 2264
rect 19057 2206 22800 2208
rect 19057 2203 19123 2206
rect 22000 2176 22800 2206
rect 4376 2064 4696 2065
rect 4376 2000 4384 2064
rect 4448 2000 4464 2064
rect 4528 2000 4544 2064
rect 4608 2000 4624 2064
rect 4688 2000 4696 2064
rect 4376 1999 4696 2000
rect 11240 2064 11560 2065
rect 11240 2000 11248 2064
rect 11312 2000 11328 2064
rect 11392 2000 11408 2064
rect 11472 2000 11488 2064
rect 11552 2000 11560 2064
rect 11240 1999 11560 2000
rect 18104 2064 18424 2065
rect 18104 2000 18112 2064
rect 18176 2000 18192 2064
rect 18256 2000 18272 2064
rect 18336 2000 18352 2064
rect 18416 2000 18424 2064
rect 18104 1999 18424 2000
rect 19241 1858 19307 1861
rect 22000 1858 22800 1888
rect 19241 1856 22800 1858
rect 19241 1800 19246 1856
rect 19302 1800 22800 1856
rect 19241 1798 22800 1800
rect 19241 1795 19307 1798
rect 22000 1768 22800 1798
rect 18873 1450 18939 1453
rect 22000 1450 22800 1480
rect 18873 1448 22800 1450
rect 18873 1392 18878 1448
rect 18934 1392 22800 1448
rect 18873 1390 22800 1392
rect 18873 1387 18939 1390
rect 22000 1360 22800 1390
rect 18689 906 18755 909
rect 22000 906 22800 936
rect 18689 904 22800 906
rect 18689 848 18694 904
rect 18750 848 22800 904
rect 18689 846 22800 848
rect 18689 843 18755 846
rect 22000 816 22800 846
rect 18781 498 18847 501
rect 22000 498 22800 528
rect 18781 496 22800 498
rect 18781 440 18786 496
rect 18842 440 22800 496
rect 18781 438 22800 440
rect 18781 435 18847 438
rect 22000 408 22800 438
rect 17953 90 18019 93
rect 22000 90 22800 120
rect 17953 88 22800 90
rect 17953 32 17958 88
rect 18014 32 22800 88
rect 17953 30 22800 32
rect 17953 27 18019 30
rect 22000 0 22800 30
<< via3 >>
rect 7816 20012 7880 20016
rect 7816 19956 7820 20012
rect 7820 19956 7876 20012
rect 7876 19956 7880 20012
rect 7816 19952 7880 19956
rect 7896 20012 7960 20016
rect 7896 19956 7900 20012
rect 7900 19956 7956 20012
rect 7956 19956 7960 20012
rect 7896 19952 7960 19956
rect 7976 20012 8040 20016
rect 7976 19956 7980 20012
rect 7980 19956 8036 20012
rect 8036 19956 8040 20012
rect 7976 19952 8040 19956
rect 8056 20012 8120 20016
rect 8056 19956 8060 20012
rect 8060 19956 8116 20012
rect 8116 19956 8120 20012
rect 8056 19952 8120 19956
rect 14680 20012 14744 20016
rect 14680 19956 14684 20012
rect 14684 19956 14740 20012
rect 14740 19956 14744 20012
rect 14680 19952 14744 19956
rect 14760 20012 14824 20016
rect 14760 19956 14764 20012
rect 14764 19956 14820 20012
rect 14820 19956 14824 20012
rect 14760 19952 14824 19956
rect 14840 20012 14904 20016
rect 14840 19956 14844 20012
rect 14844 19956 14900 20012
rect 14900 19956 14904 20012
rect 14840 19952 14904 19956
rect 14920 20012 14984 20016
rect 14920 19956 14924 20012
rect 14924 19956 14980 20012
rect 14980 19956 14984 20012
rect 14920 19952 14984 19956
rect 4384 19468 4448 19472
rect 4384 19412 4388 19468
rect 4388 19412 4444 19468
rect 4444 19412 4448 19468
rect 4384 19408 4448 19412
rect 4464 19468 4528 19472
rect 4464 19412 4468 19468
rect 4468 19412 4524 19468
rect 4524 19412 4528 19468
rect 4464 19408 4528 19412
rect 4544 19468 4608 19472
rect 4544 19412 4548 19468
rect 4548 19412 4604 19468
rect 4604 19412 4608 19468
rect 4544 19408 4608 19412
rect 4624 19468 4688 19472
rect 4624 19412 4628 19468
rect 4628 19412 4684 19468
rect 4684 19412 4688 19468
rect 4624 19408 4688 19412
rect 11248 19468 11312 19472
rect 11248 19412 11252 19468
rect 11252 19412 11308 19468
rect 11308 19412 11312 19468
rect 11248 19408 11312 19412
rect 11328 19468 11392 19472
rect 11328 19412 11332 19468
rect 11332 19412 11388 19468
rect 11388 19412 11392 19468
rect 11328 19408 11392 19412
rect 11408 19468 11472 19472
rect 11408 19412 11412 19468
rect 11412 19412 11468 19468
rect 11468 19412 11472 19468
rect 11408 19408 11472 19412
rect 11488 19468 11552 19472
rect 11488 19412 11492 19468
rect 11492 19412 11548 19468
rect 11548 19412 11552 19468
rect 11488 19408 11552 19412
rect 18112 19468 18176 19472
rect 18112 19412 18116 19468
rect 18116 19412 18172 19468
rect 18172 19412 18176 19468
rect 18112 19408 18176 19412
rect 18192 19468 18256 19472
rect 18192 19412 18196 19468
rect 18196 19412 18252 19468
rect 18252 19412 18256 19468
rect 18192 19408 18256 19412
rect 18272 19468 18336 19472
rect 18272 19412 18276 19468
rect 18276 19412 18332 19468
rect 18332 19412 18336 19468
rect 18272 19408 18336 19412
rect 18352 19468 18416 19472
rect 18352 19412 18356 19468
rect 18356 19412 18412 19468
rect 18412 19412 18416 19468
rect 18352 19408 18416 19412
rect 7816 18924 7880 18928
rect 7816 18868 7820 18924
rect 7820 18868 7876 18924
rect 7876 18868 7880 18924
rect 7816 18864 7880 18868
rect 7896 18924 7960 18928
rect 7896 18868 7900 18924
rect 7900 18868 7956 18924
rect 7956 18868 7960 18924
rect 7896 18864 7960 18868
rect 7976 18924 8040 18928
rect 7976 18868 7980 18924
rect 7980 18868 8036 18924
rect 8036 18868 8040 18924
rect 7976 18864 8040 18868
rect 8056 18924 8120 18928
rect 8056 18868 8060 18924
rect 8060 18868 8116 18924
rect 8116 18868 8120 18924
rect 8056 18864 8120 18868
rect 14680 18924 14744 18928
rect 14680 18868 14684 18924
rect 14684 18868 14740 18924
rect 14740 18868 14744 18924
rect 14680 18864 14744 18868
rect 14760 18924 14824 18928
rect 14760 18868 14764 18924
rect 14764 18868 14820 18924
rect 14820 18868 14824 18924
rect 14760 18864 14824 18868
rect 14840 18924 14904 18928
rect 14840 18868 14844 18924
rect 14844 18868 14900 18924
rect 14900 18868 14904 18924
rect 14840 18864 14904 18868
rect 14920 18924 14984 18928
rect 14920 18868 14924 18924
rect 14924 18868 14980 18924
rect 14980 18868 14984 18924
rect 14920 18864 14984 18868
rect 19380 18584 19444 18588
rect 19380 18528 19394 18584
rect 19394 18528 19444 18584
rect 19380 18524 19444 18528
rect 4384 18380 4448 18384
rect 4384 18324 4388 18380
rect 4388 18324 4444 18380
rect 4444 18324 4448 18380
rect 4384 18320 4448 18324
rect 4464 18380 4528 18384
rect 4464 18324 4468 18380
rect 4468 18324 4524 18380
rect 4524 18324 4528 18380
rect 4464 18320 4528 18324
rect 4544 18380 4608 18384
rect 4544 18324 4548 18380
rect 4548 18324 4604 18380
rect 4604 18324 4608 18380
rect 4544 18320 4608 18324
rect 4624 18380 4688 18384
rect 4624 18324 4628 18380
rect 4628 18324 4684 18380
rect 4684 18324 4688 18380
rect 4624 18320 4688 18324
rect 11248 18380 11312 18384
rect 11248 18324 11252 18380
rect 11252 18324 11308 18380
rect 11308 18324 11312 18380
rect 11248 18320 11312 18324
rect 11328 18380 11392 18384
rect 11328 18324 11332 18380
rect 11332 18324 11388 18380
rect 11388 18324 11392 18380
rect 11328 18320 11392 18324
rect 11408 18380 11472 18384
rect 11408 18324 11412 18380
rect 11412 18324 11468 18380
rect 11468 18324 11472 18380
rect 11408 18320 11472 18324
rect 11488 18380 11552 18384
rect 11488 18324 11492 18380
rect 11492 18324 11548 18380
rect 11548 18324 11552 18380
rect 11488 18320 11552 18324
rect 18112 18380 18176 18384
rect 18112 18324 18116 18380
rect 18116 18324 18172 18380
rect 18172 18324 18176 18380
rect 18112 18320 18176 18324
rect 18192 18380 18256 18384
rect 18192 18324 18196 18380
rect 18196 18324 18252 18380
rect 18252 18324 18256 18380
rect 18192 18320 18256 18324
rect 18272 18380 18336 18384
rect 18272 18324 18276 18380
rect 18276 18324 18332 18380
rect 18332 18324 18336 18380
rect 18272 18320 18336 18324
rect 18352 18380 18416 18384
rect 18352 18324 18356 18380
rect 18356 18324 18412 18380
rect 18412 18324 18416 18380
rect 18352 18320 18416 18324
rect 7816 17836 7880 17840
rect 7816 17780 7820 17836
rect 7820 17780 7876 17836
rect 7876 17780 7880 17836
rect 7816 17776 7880 17780
rect 7896 17836 7960 17840
rect 7896 17780 7900 17836
rect 7900 17780 7956 17836
rect 7956 17780 7960 17836
rect 7896 17776 7960 17780
rect 7976 17836 8040 17840
rect 7976 17780 7980 17836
rect 7980 17780 8036 17836
rect 8036 17780 8040 17836
rect 7976 17776 8040 17780
rect 8056 17836 8120 17840
rect 8056 17780 8060 17836
rect 8060 17780 8116 17836
rect 8116 17780 8120 17836
rect 8056 17776 8120 17780
rect 14680 17836 14744 17840
rect 14680 17780 14684 17836
rect 14684 17780 14740 17836
rect 14740 17780 14744 17836
rect 14680 17776 14744 17780
rect 14760 17836 14824 17840
rect 14760 17780 14764 17836
rect 14764 17780 14820 17836
rect 14820 17780 14824 17836
rect 14760 17776 14824 17780
rect 14840 17836 14904 17840
rect 14840 17780 14844 17836
rect 14844 17780 14900 17836
rect 14900 17780 14904 17836
rect 14840 17776 14904 17780
rect 14920 17836 14984 17840
rect 14920 17780 14924 17836
rect 14924 17780 14980 17836
rect 14980 17780 14984 17836
rect 14920 17776 14984 17780
rect 4384 17292 4448 17296
rect 4384 17236 4388 17292
rect 4388 17236 4444 17292
rect 4444 17236 4448 17292
rect 4384 17232 4448 17236
rect 4464 17292 4528 17296
rect 4464 17236 4468 17292
rect 4468 17236 4524 17292
rect 4524 17236 4528 17292
rect 4464 17232 4528 17236
rect 4544 17292 4608 17296
rect 4544 17236 4548 17292
rect 4548 17236 4604 17292
rect 4604 17236 4608 17292
rect 4544 17232 4608 17236
rect 4624 17292 4688 17296
rect 4624 17236 4628 17292
rect 4628 17236 4684 17292
rect 4684 17236 4688 17292
rect 4624 17232 4688 17236
rect 11248 17292 11312 17296
rect 11248 17236 11252 17292
rect 11252 17236 11308 17292
rect 11308 17236 11312 17292
rect 11248 17232 11312 17236
rect 11328 17292 11392 17296
rect 11328 17236 11332 17292
rect 11332 17236 11388 17292
rect 11388 17236 11392 17292
rect 11328 17232 11392 17236
rect 11408 17292 11472 17296
rect 11408 17236 11412 17292
rect 11412 17236 11468 17292
rect 11468 17236 11472 17292
rect 11408 17232 11472 17236
rect 11488 17292 11552 17296
rect 11488 17236 11492 17292
rect 11492 17236 11548 17292
rect 11548 17236 11552 17292
rect 11488 17232 11552 17236
rect 18112 17292 18176 17296
rect 18112 17236 18116 17292
rect 18116 17236 18172 17292
rect 18172 17236 18176 17292
rect 18112 17232 18176 17236
rect 18192 17292 18256 17296
rect 18192 17236 18196 17292
rect 18196 17236 18252 17292
rect 18252 17236 18256 17292
rect 18192 17232 18256 17236
rect 18272 17292 18336 17296
rect 18272 17236 18276 17292
rect 18276 17236 18332 17292
rect 18332 17236 18336 17292
rect 18272 17232 18336 17236
rect 18352 17292 18416 17296
rect 18352 17236 18356 17292
rect 18356 17236 18412 17292
rect 18412 17236 18416 17292
rect 18352 17232 18416 17236
rect 7816 16748 7880 16752
rect 7816 16692 7820 16748
rect 7820 16692 7876 16748
rect 7876 16692 7880 16748
rect 7816 16688 7880 16692
rect 7896 16748 7960 16752
rect 7896 16692 7900 16748
rect 7900 16692 7956 16748
rect 7956 16692 7960 16748
rect 7896 16688 7960 16692
rect 7976 16748 8040 16752
rect 7976 16692 7980 16748
rect 7980 16692 8036 16748
rect 8036 16692 8040 16748
rect 7976 16688 8040 16692
rect 8056 16748 8120 16752
rect 8056 16692 8060 16748
rect 8060 16692 8116 16748
rect 8116 16692 8120 16748
rect 8056 16688 8120 16692
rect 14680 16748 14744 16752
rect 14680 16692 14684 16748
rect 14684 16692 14740 16748
rect 14740 16692 14744 16748
rect 14680 16688 14744 16692
rect 14760 16748 14824 16752
rect 14760 16692 14764 16748
rect 14764 16692 14820 16748
rect 14820 16692 14824 16748
rect 14760 16688 14824 16692
rect 14840 16748 14904 16752
rect 14840 16692 14844 16748
rect 14844 16692 14900 16748
rect 14900 16692 14904 16748
rect 14840 16688 14904 16692
rect 14920 16748 14984 16752
rect 14920 16692 14924 16748
rect 14924 16692 14980 16748
rect 14980 16692 14984 16748
rect 14920 16688 14984 16692
rect 4384 16204 4448 16208
rect 4384 16148 4388 16204
rect 4388 16148 4444 16204
rect 4444 16148 4448 16204
rect 4384 16144 4448 16148
rect 4464 16204 4528 16208
rect 4464 16148 4468 16204
rect 4468 16148 4524 16204
rect 4524 16148 4528 16204
rect 4464 16144 4528 16148
rect 4544 16204 4608 16208
rect 4544 16148 4548 16204
rect 4548 16148 4604 16204
rect 4604 16148 4608 16204
rect 4544 16144 4608 16148
rect 4624 16204 4688 16208
rect 4624 16148 4628 16204
rect 4628 16148 4684 16204
rect 4684 16148 4688 16204
rect 4624 16144 4688 16148
rect 11248 16204 11312 16208
rect 11248 16148 11252 16204
rect 11252 16148 11308 16204
rect 11308 16148 11312 16204
rect 11248 16144 11312 16148
rect 11328 16204 11392 16208
rect 11328 16148 11332 16204
rect 11332 16148 11388 16204
rect 11388 16148 11392 16204
rect 11328 16144 11392 16148
rect 11408 16204 11472 16208
rect 11408 16148 11412 16204
rect 11412 16148 11468 16204
rect 11468 16148 11472 16204
rect 11408 16144 11472 16148
rect 11488 16204 11552 16208
rect 11488 16148 11492 16204
rect 11492 16148 11548 16204
rect 11548 16148 11552 16204
rect 11488 16144 11552 16148
rect 18112 16204 18176 16208
rect 18112 16148 18116 16204
rect 18116 16148 18172 16204
rect 18172 16148 18176 16204
rect 18112 16144 18176 16148
rect 18192 16204 18256 16208
rect 18192 16148 18196 16204
rect 18196 16148 18252 16204
rect 18252 16148 18256 16204
rect 18192 16144 18256 16148
rect 18272 16204 18336 16208
rect 18272 16148 18276 16204
rect 18276 16148 18332 16204
rect 18332 16148 18336 16204
rect 18272 16144 18336 16148
rect 18352 16204 18416 16208
rect 18352 16148 18356 16204
rect 18356 16148 18412 16204
rect 18412 16148 18416 16204
rect 18352 16144 18416 16148
rect 7816 15660 7880 15664
rect 7816 15604 7820 15660
rect 7820 15604 7876 15660
rect 7876 15604 7880 15660
rect 7816 15600 7880 15604
rect 7896 15660 7960 15664
rect 7896 15604 7900 15660
rect 7900 15604 7956 15660
rect 7956 15604 7960 15660
rect 7896 15600 7960 15604
rect 7976 15660 8040 15664
rect 7976 15604 7980 15660
rect 7980 15604 8036 15660
rect 8036 15604 8040 15660
rect 7976 15600 8040 15604
rect 8056 15660 8120 15664
rect 8056 15604 8060 15660
rect 8060 15604 8116 15660
rect 8116 15604 8120 15660
rect 8056 15600 8120 15604
rect 14680 15660 14744 15664
rect 14680 15604 14684 15660
rect 14684 15604 14740 15660
rect 14740 15604 14744 15660
rect 14680 15600 14744 15604
rect 14760 15660 14824 15664
rect 14760 15604 14764 15660
rect 14764 15604 14820 15660
rect 14820 15604 14824 15660
rect 14760 15600 14824 15604
rect 14840 15660 14904 15664
rect 14840 15604 14844 15660
rect 14844 15604 14900 15660
rect 14900 15604 14904 15660
rect 14840 15600 14904 15604
rect 14920 15660 14984 15664
rect 14920 15604 14924 15660
rect 14924 15604 14980 15660
rect 14980 15604 14984 15660
rect 14920 15600 14984 15604
rect 4384 15116 4448 15120
rect 4384 15060 4388 15116
rect 4388 15060 4444 15116
rect 4444 15060 4448 15116
rect 4384 15056 4448 15060
rect 4464 15116 4528 15120
rect 4464 15060 4468 15116
rect 4468 15060 4524 15116
rect 4524 15060 4528 15116
rect 4464 15056 4528 15060
rect 4544 15116 4608 15120
rect 4544 15060 4548 15116
rect 4548 15060 4604 15116
rect 4604 15060 4608 15116
rect 4544 15056 4608 15060
rect 4624 15116 4688 15120
rect 4624 15060 4628 15116
rect 4628 15060 4684 15116
rect 4684 15060 4688 15116
rect 4624 15056 4688 15060
rect 11248 15116 11312 15120
rect 11248 15060 11252 15116
rect 11252 15060 11308 15116
rect 11308 15060 11312 15116
rect 11248 15056 11312 15060
rect 11328 15116 11392 15120
rect 11328 15060 11332 15116
rect 11332 15060 11388 15116
rect 11388 15060 11392 15116
rect 11328 15056 11392 15060
rect 11408 15116 11472 15120
rect 11408 15060 11412 15116
rect 11412 15060 11468 15116
rect 11468 15060 11472 15116
rect 11408 15056 11472 15060
rect 11488 15116 11552 15120
rect 11488 15060 11492 15116
rect 11492 15060 11548 15116
rect 11548 15060 11552 15116
rect 11488 15056 11552 15060
rect 18112 15116 18176 15120
rect 18112 15060 18116 15116
rect 18116 15060 18172 15116
rect 18172 15060 18176 15116
rect 18112 15056 18176 15060
rect 18192 15116 18256 15120
rect 18192 15060 18196 15116
rect 18196 15060 18252 15116
rect 18252 15060 18256 15116
rect 18192 15056 18256 15060
rect 18272 15116 18336 15120
rect 18272 15060 18276 15116
rect 18276 15060 18332 15116
rect 18332 15060 18336 15116
rect 18272 15056 18336 15060
rect 18352 15116 18416 15120
rect 18352 15060 18356 15116
rect 18356 15060 18412 15116
rect 18412 15060 18416 15116
rect 18352 15056 18416 15060
rect 7816 14572 7880 14576
rect 7816 14516 7820 14572
rect 7820 14516 7876 14572
rect 7876 14516 7880 14572
rect 7816 14512 7880 14516
rect 7896 14572 7960 14576
rect 7896 14516 7900 14572
rect 7900 14516 7956 14572
rect 7956 14516 7960 14572
rect 7896 14512 7960 14516
rect 7976 14572 8040 14576
rect 7976 14516 7980 14572
rect 7980 14516 8036 14572
rect 8036 14516 8040 14572
rect 7976 14512 8040 14516
rect 8056 14572 8120 14576
rect 8056 14516 8060 14572
rect 8060 14516 8116 14572
rect 8116 14516 8120 14572
rect 8056 14512 8120 14516
rect 14680 14572 14744 14576
rect 14680 14516 14684 14572
rect 14684 14516 14740 14572
rect 14740 14516 14744 14572
rect 14680 14512 14744 14516
rect 14760 14572 14824 14576
rect 14760 14516 14764 14572
rect 14764 14516 14820 14572
rect 14820 14516 14824 14572
rect 14760 14512 14824 14516
rect 14840 14572 14904 14576
rect 14840 14516 14844 14572
rect 14844 14516 14900 14572
rect 14900 14516 14904 14572
rect 14840 14512 14904 14516
rect 14920 14572 14984 14576
rect 14920 14516 14924 14572
rect 14924 14516 14980 14572
rect 14980 14516 14984 14572
rect 14920 14512 14984 14516
rect 4384 14028 4448 14032
rect 4384 13972 4388 14028
rect 4388 13972 4444 14028
rect 4444 13972 4448 14028
rect 4384 13968 4448 13972
rect 4464 14028 4528 14032
rect 4464 13972 4468 14028
rect 4468 13972 4524 14028
rect 4524 13972 4528 14028
rect 4464 13968 4528 13972
rect 4544 14028 4608 14032
rect 4544 13972 4548 14028
rect 4548 13972 4604 14028
rect 4604 13972 4608 14028
rect 4544 13968 4608 13972
rect 4624 14028 4688 14032
rect 4624 13972 4628 14028
rect 4628 13972 4684 14028
rect 4684 13972 4688 14028
rect 4624 13968 4688 13972
rect 11248 14028 11312 14032
rect 11248 13972 11252 14028
rect 11252 13972 11308 14028
rect 11308 13972 11312 14028
rect 11248 13968 11312 13972
rect 11328 14028 11392 14032
rect 11328 13972 11332 14028
rect 11332 13972 11388 14028
rect 11388 13972 11392 14028
rect 11328 13968 11392 13972
rect 11408 14028 11472 14032
rect 11408 13972 11412 14028
rect 11412 13972 11468 14028
rect 11468 13972 11472 14028
rect 11408 13968 11472 13972
rect 11488 14028 11552 14032
rect 11488 13972 11492 14028
rect 11492 13972 11548 14028
rect 11548 13972 11552 14028
rect 11488 13968 11552 13972
rect 18112 14028 18176 14032
rect 18112 13972 18116 14028
rect 18116 13972 18172 14028
rect 18172 13972 18176 14028
rect 18112 13968 18176 13972
rect 18192 14028 18256 14032
rect 18192 13972 18196 14028
rect 18196 13972 18252 14028
rect 18252 13972 18256 14028
rect 18192 13968 18256 13972
rect 18272 14028 18336 14032
rect 18272 13972 18276 14028
rect 18276 13972 18332 14028
rect 18332 13972 18336 14028
rect 18272 13968 18336 13972
rect 18352 14028 18416 14032
rect 18352 13972 18356 14028
rect 18356 13972 18412 14028
rect 18412 13972 18416 14028
rect 18352 13968 18416 13972
rect 19380 13628 19444 13692
rect 7816 13484 7880 13488
rect 7816 13428 7820 13484
rect 7820 13428 7876 13484
rect 7876 13428 7880 13484
rect 7816 13424 7880 13428
rect 7896 13484 7960 13488
rect 7896 13428 7900 13484
rect 7900 13428 7956 13484
rect 7956 13428 7960 13484
rect 7896 13424 7960 13428
rect 7976 13484 8040 13488
rect 7976 13428 7980 13484
rect 7980 13428 8036 13484
rect 8036 13428 8040 13484
rect 7976 13424 8040 13428
rect 8056 13484 8120 13488
rect 8056 13428 8060 13484
rect 8060 13428 8116 13484
rect 8116 13428 8120 13484
rect 8056 13424 8120 13428
rect 14680 13484 14744 13488
rect 14680 13428 14684 13484
rect 14684 13428 14740 13484
rect 14740 13428 14744 13484
rect 14680 13424 14744 13428
rect 14760 13484 14824 13488
rect 14760 13428 14764 13484
rect 14764 13428 14820 13484
rect 14820 13428 14824 13484
rect 14760 13424 14824 13428
rect 14840 13484 14904 13488
rect 14840 13428 14844 13484
rect 14844 13428 14900 13484
rect 14900 13428 14904 13484
rect 14840 13424 14904 13428
rect 14920 13484 14984 13488
rect 14920 13428 14924 13484
rect 14924 13428 14980 13484
rect 14980 13428 14984 13484
rect 14920 13424 14984 13428
rect 4384 12940 4448 12944
rect 4384 12884 4388 12940
rect 4388 12884 4444 12940
rect 4444 12884 4448 12940
rect 4384 12880 4448 12884
rect 4464 12940 4528 12944
rect 4464 12884 4468 12940
rect 4468 12884 4524 12940
rect 4524 12884 4528 12940
rect 4464 12880 4528 12884
rect 4544 12940 4608 12944
rect 4544 12884 4548 12940
rect 4548 12884 4604 12940
rect 4604 12884 4608 12940
rect 4544 12880 4608 12884
rect 4624 12940 4688 12944
rect 4624 12884 4628 12940
rect 4628 12884 4684 12940
rect 4684 12884 4688 12940
rect 4624 12880 4688 12884
rect 11248 12940 11312 12944
rect 11248 12884 11252 12940
rect 11252 12884 11308 12940
rect 11308 12884 11312 12940
rect 11248 12880 11312 12884
rect 11328 12940 11392 12944
rect 11328 12884 11332 12940
rect 11332 12884 11388 12940
rect 11388 12884 11392 12940
rect 11328 12880 11392 12884
rect 11408 12940 11472 12944
rect 11408 12884 11412 12940
rect 11412 12884 11468 12940
rect 11468 12884 11472 12940
rect 11408 12880 11472 12884
rect 11488 12940 11552 12944
rect 11488 12884 11492 12940
rect 11492 12884 11548 12940
rect 11548 12884 11552 12940
rect 11488 12880 11552 12884
rect 18112 12940 18176 12944
rect 18112 12884 18116 12940
rect 18116 12884 18172 12940
rect 18172 12884 18176 12940
rect 18112 12880 18176 12884
rect 18192 12940 18256 12944
rect 18192 12884 18196 12940
rect 18196 12884 18252 12940
rect 18252 12884 18256 12940
rect 18192 12880 18256 12884
rect 18272 12940 18336 12944
rect 18272 12884 18276 12940
rect 18276 12884 18332 12940
rect 18332 12884 18336 12940
rect 18272 12880 18336 12884
rect 18352 12940 18416 12944
rect 18352 12884 18356 12940
rect 18356 12884 18412 12940
rect 18412 12884 18416 12940
rect 18352 12880 18416 12884
rect 7816 12396 7880 12400
rect 7816 12340 7820 12396
rect 7820 12340 7876 12396
rect 7876 12340 7880 12396
rect 7816 12336 7880 12340
rect 7896 12396 7960 12400
rect 7896 12340 7900 12396
rect 7900 12340 7956 12396
rect 7956 12340 7960 12396
rect 7896 12336 7960 12340
rect 7976 12396 8040 12400
rect 7976 12340 7980 12396
rect 7980 12340 8036 12396
rect 8036 12340 8040 12396
rect 7976 12336 8040 12340
rect 8056 12396 8120 12400
rect 8056 12340 8060 12396
rect 8060 12340 8116 12396
rect 8116 12340 8120 12396
rect 8056 12336 8120 12340
rect 14680 12396 14744 12400
rect 14680 12340 14684 12396
rect 14684 12340 14740 12396
rect 14740 12340 14744 12396
rect 14680 12336 14744 12340
rect 14760 12396 14824 12400
rect 14760 12340 14764 12396
rect 14764 12340 14820 12396
rect 14820 12340 14824 12396
rect 14760 12336 14824 12340
rect 14840 12396 14904 12400
rect 14840 12340 14844 12396
rect 14844 12340 14900 12396
rect 14900 12340 14904 12396
rect 14840 12336 14904 12340
rect 14920 12396 14984 12400
rect 14920 12340 14924 12396
rect 14924 12340 14980 12396
rect 14980 12340 14984 12396
rect 14920 12336 14984 12340
rect 4384 11852 4448 11856
rect 4384 11796 4388 11852
rect 4388 11796 4444 11852
rect 4444 11796 4448 11852
rect 4384 11792 4448 11796
rect 4464 11852 4528 11856
rect 4464 11796 4468 11852
rect 4468 11796 4524 11852
rect 4524 11796 4528 11852
rect 4464 11792 4528 11796
rect 4544 11852 4608 11856
rect 4544 11796 4548 11852
rect 4548 11796 4604 11852
rect 4604 11796 4608 11852
rect 4544 11792 4608 11796
rect 4624 11852 4688 11856
rect 4624 11796 4628 11852
rect 4628 11796 4684 11852
rect 4684 11796 4688 11852
rect 4624 11792 4688 11796
rect 11248 11852 11312 11856
rect 11248 11796 11252 11852
rect 11252 11796 11308 11852
rect 11308 11796 11312 11852
rect 11248 11792 11312 11796
rect 11328 11852 11392 11856
rect 11328 11796 11332 11852
rect 11332 11796 11388 11852
rect 11388 11796 11392 11852
rect 11328 11792 11392 11796
rect 11408 11852 11472 11856
rect 11408 11796 11412 11852
rect 11412 11796 11468 11852
rect 11468 11796 11472 11852
rect 11408 11792 11472 11796
rect 11488 11852 11552 11856
rect 11488 11796 11492 11852
rect 11492 11796 11548 11852
rect 11548 11796 11552 11852
rect 11488 11792 11552 11796
rect 18112 11852 18176 11856
rect 18112 11796 18116 11852
rect 18116 11796 18172 11852
rect 18172 11796 18176 11852
rect 18112 11792 18176 11796
rect 18192 11852 18256 11856
rect 18192 11796 18196 11852
rect 18196 11796 18252 11852
rect 18252 11796 18256 11852
rect 18192 11792 18256 11796
rect 18272 11852 18336 11856
rect 18272 11796 18276 11852
rect 18276 11796 18332 11852
rect 18332 11796 18336 11852
rect 18272 11792 18336 11796
rect 18352 11852 18416 11856
rect 18352 11796 18356 11852
rect 18356 11796 18412 11852
rect 18412 11796 18416 11852
rect 18352 11792 18416 11796
rect 7816 11308 7880 11312
rect 7816 11252 7820 11308
rect 7820 11252 7876 11308
rect 7876 11252 7880 11308
rect 7816 11248 7880 11252
rect 7896 11308 7960 11312
rect 7896 11252 7900 11308
rect 7900 11252 7956 11308
rect 7956 11252 7960 11308
rect 7896 11248 7960 11252
rect 7976 11308 8040 11312
rect 7976 11252 7980 11308
rect 7980 11252 8036 11308
rect 8036 11252 8040 11308
rect 7976 11248 8040 11252
rect 8056 11308 8120 11312
rect 8056 11252 8060 11308
rect 8060 11252 8116 11308
rect 8116 11252 8120 11308
rect 8056 11248 8120 11252
rect 14680 11308 14744 11312
rect 14680 11252 14684 11308
rect 14684 11252 14740 11308
rect 14740 11252 14744 11308
rect 14680 11248 14744 11252
rect 14760 11308 14824 11312
rect 14760 11252 14764 11308
rect 14764 11252 14820 11308
rect 14820 11252 14824 11308
rect 14760 11248 14824 11252
rect 14840 11308 14904 11312
rect 14840 11252 14844 11308
rect 14844 11252 14900 11308
rect 14900 11252 14904 11308
rect 14840 11248 14904 11252
rect 14920 11308 14984 11312
rect 14920 11252 14924 11308
rect 14924 11252 14980 11308
rect 14980 11252 14984 11308
rect 14920 11248 14984 11252
rect 4384 10764 4448 10768
rect 4384 10708 4388 10764
rect 4388 10708 4444 10764
rect 4444 10708 4448 10764
rect 4384 10704 4448 10708
rect 4464 10764 4528 10768
rect 4464 10708 4468 10764
rect 4468 10708 4524 10764
rect 4524 10708 4528 10764
rect 4464 10704 4528 10708
rect 4544 10764 4608 10768
rect 4544 10708 4548 10764
rect 4548 10708 4604 10764
rect 4604 10708 4608 10764
rect 4544 10704 4608 10708
rect 4624 10764 4688 10768
rect 4624 10708 4628 10764
rect 4628 10708 4684 10764
rect 4684 10708 4688 10764
rect 4624 10704 4688 10708
rect 11248 10764 11312 10768
rect 11248 10708 11252 10764
rect 11252 10708 11308 10764
rect 11308 10708 11312 10764
rect 11248 10704 11312 10708
rect 11328 10764 11392 10768
rect 11328 10708 11332 10764
rect 11332 10708 11388 10764
rect 11388 10708 11392 10764
rect 11328 10704 11392 10708
rect 11408 10764 11472 10768
rect 11408 10708 11412 10764
rect 11412 10708 11468 10764
rect 11468 10708 11472 10764
rect 11408 10704 11472 10708
rect 11488 10764 11552 10768
rect 11488 10708 11492 10764
rect 11492 10708 11548 10764
rect 11548 10708 11552 10764
rect 11488 10704 11552 10708
rect 18112 10764 18176 10768
rect 18112 10708 18116 10764
rect 18116 10708 18172 10764
rect 18172 10708 18176 10764
rect 18112 10704 18176 10708
rect 18192 10764 18256 10768
rect 18192 10708 18196 10764
rect 18196 10708 18252 10764
rect 18252 10708 18256 10764
rect 18192 10704 18256 10708
rect 18272 10764 18336 10768
rect 18272 10708 18276 10764
rect 18276 10708 18332 10764
rect 18332 10708 18336 10764
rect 18272 10704 18336 10708
rect 18352 10764 18416 10768
rect 18352 10708 18356 10764
rect 18356 10708 18412 10764
rect 18412 10708 18416 10764
rect 18352 10704 18416 10708
rect 7816 10220 7880 10224
rect 7816 10164 7820 10220
rect 7820 10164 7876 10220
rect 7876 10164 7880 10220
rect 7816 10160 7880 10164
rect 7896 10220 7960 10224
rect 7896 10164 7900 10220
rect 7900 10164 7956 10220
rect 7956 10164 7960 10220
rect 7896 10160 7960 10164
rect 7976 10220 8040 10224
rect 7976 10164 7980 10220
rect 7980 10164 8036 10220
rect 8036 10164 8040 10220
rect 7976 10160 8040 10164
rect 8056 10220 8120 10224
rect 8056 10164 8060 10220
rect 8060 10164 8116 10220
rect 8116 10164 8120 10220
rect 8056 10160 8120 10164
rect 14680 10220 14744 10224
rect 14680 10164 14684 10220
rect 14684 10164 14740 10220
rect 14740 10164 14744 10220
rect 14680 10160 14744 10164
rect 14760 10220 14824 10224
rect 14760 10164 14764 10220
rect 14764 10164 14820 10220
rect 14820 10164 14824 10220
rect 14760 10160 14824 10164
rect 14840 10220 14904 10224
rect 14840 10164 14844 10220
rect 14844 10164 14900 10220
rect 14900 10164 14904 10220
rect 14840 10160 14904 10164
rect 14920 10220 14984 10224
rect 14920 10164 14924 10220
rect 14924 10164 14980 10220
rect 14980 10164 14984 10220
rect 14920 10160 14984 10164
rect 4384 9676 4448 9680
rect 4384 9620 4388 9676
rect 4388 9620 4444 9676
rect 4444 9620 4448 9676
rect 4384 9616 4448 9620
rect 4464 9676 4528 9680
rect 4464 9620 4468 9676
rect 4468 9620 4524 9676
rect 4524 9620 4528 9676
rect 4464 9616 4528 9620
rect 4544 9676 4608 9680
rect 4544 9620 4548 9676
rect 4548 9620 4604 9676
rect 4604 9620 4608 9676
rect 4544 9616 4608 9620
rect 4624 9676 4688 9680
rect 4624 9620 4628 9676
rect 4628 9620 4684 9676
rect 4684 9620 4688 9676
rect 4624 9616 4688 9620
rect 11248 9676 11312 9680
rect 11248 9620 11252 9676
rect 11252 9620 11308 9676
rect 11308 9620 11312 9676
rect 11248 9616 11312 9620
rect 11328 9676 11392 9680
rect 11328 9620 11332 9676
rect 11332 9620 11388 9676
rect 11388 9620 11392 9676
rect 11328 9616 11392 9620
rect 11408 9676 11472 9680
rect 11408 9620 11412 9676
rect 11412 9620 11468 9676
rect 11468 9620 11472 9676
rect 11408 9616 11472 9620
rect 11488 9676 11552 9680
rect 11488 9620 11492 9676
rect 11492 9620 11548 9676
rect 11548 9620 11552 9676
rect 11488 9616 11552 9620
rect 18112 9676 18176 9680
rect 18112 9620 18116 9676
rect 18116 9620 18172 9676
rect 18172 9620 18176 9676
rect 18112 9616 18176 9620
rect 18192 9676 18256 9680
rect 18192 9620 18196 9676
rect 18196 9620 18252 9676
rect 18252 9620 18256 9676
rect 18192 9616 18256 9620
rect 18272 9676 18336 9680
rect 18272 9620 18276 9676
rect 18276 9620 18332 9676
rect 18332 9620 18336 9676
rect 18272 9616 18336 9620
rect 18352 9676 18416 9680
rect 18352 9620 18356 9676
rect 18356 9620 18412 9676
rect 18412 9620 18416 9676
rect 18352 9616 18416 9620
rect 7816 9132 7880 9136
rect 7816 9076 7820 9132
rect 7820 9076 7876 9132
rect 7876 9076 7880 9132
rect 7816 9072 7880 9076
rect 7896 9132 7960 9136
rect 7896 9076 7900 9132
rect 7900 9076 7956 9132
rect 7956 9076 7960 9132
rect 7896 9072 7960 9076
rect 7976 9132 8040 9136
rect 7976 9076 7980 9132
rect 7980 9076 8036 9132
rect 8036 9076 8040 9132
rect 7976 9072 8040 9076
rect 8056 9132 8120 9136
rect 8056 9076 8060 9132
rect 8060 9076 8116 9132
rect 8116 9076 8120 9132
rect 8056 9072 8120 9076
rect 14680 9132 14744 9136
rect 14680 9076 14684 9132
rect 14684 9076 14740 9132
rect 14740 9076 14744 9132
rect 14680 9072 14744 9076
rect 14760 9132 14824 9136
rect 14760 9076 14764 9132
rect 14764 9076 14820 9132
rect 14820 9076 14824 9132
rect 14760 9072 14824 9076
rect 14840 9132 14904 9136
rect 14840 9076 14844 9132
rect 14844 9076 14900 9132
rect 14900 9076 14904 9132
rect 14840 9072 14904 9076
rect 14920 9132 14984 9136
rect 14920 9076 14924 9132
rect 14924 9076 14980 9132
rect 14980 9076 14984 9132
rect 14920 9072 14984 9076
rect 4384 8588 4448 8592
rect 4384 8532 4388 8588
rect 4388 8532 4444 8588
rect 4444 8532 4448 8588
rect 4384 8528 4448 8532
rect 4464 8588 4528 8592
rect 4464 8532 4468 8588
rect 4468 8532 4524 8588
rect 4524 8532 4528 8588
rect 4464 8528 4528 8532
rect 4544 8588 4608 8592
rect 4544 8532 4548 8588
rect 4548 8532 4604 8588
rect 4604 8532 4608 8588
rect 4544 8528 4608 8532
rect 4624 8588 4688 8592
rect 4624 8532 4628 8588
rect 4628 8532 4684 8588
rect 4684 8532 4688 8588
rect 4624 8528 4688 8532
rect 11248 8588 11312 8592
rect 11248 8532 11252 8588
rect 11252 8532 11308 8588
rect 11308 8532 11312 8588
rect 11248 8528 11312 8532
rect 11328 8588 11392 8592
rect 11328 8532 11332 8588
rect 11332 8532 11388 8588
rect 11388 8532 11392 8588
rect 11328 8528 11392 8532
rect 11408 8588 11472 8592
rect 11408 8532 11412 8588
rect 11412 8532 11468 8588
rect 11468 8532 11472 8588
rect 11408 8528 11472 8532
rect 11488 8588 11552 8592
rect 11488 8532 11492 8588
rect 11492 8532 11548 8588
rect 11548 8532 11552 8588
rect 11488 8528 11552 8532
rect 18112 8588 18176 8592
rect 18112 8532 18116 8588
rect 18116 8532 18172 8588
rect 18172 8532 18176 8588
rect 18112 8528 18176 8532
rect 18192 8588 18256 8592
rect 18192 8532 18196 8588
rect 18196 8532 18252 8588
rect 18252 8532 18256 8588
rect 18192 8528 18256 8532
rect 18272 8588 18336 8592
rect 18272 8532 18276 8588
rect 18276 8532 18332 8588
rect 18332 8532 18336 8588
rect 18272 8528 18336 8532
rect 18352 8588 18416 8592
rect 18352 8532 18356 8588
rect 18356 8532 18412 8588
rect 18412 8532 18416 8588
rect 18352 8528 18416 8532
rect 7816 8044 7880 8048
rect 7816 7988 7820 8044
rect 7820 7988 7876 8044
rect 7876 7988 7880 8044
rect 7816 7984 7880 7988
rect 7896 8044 7960 8048
rect 7896 7988 7900 8044
rect 7900 7988 7956 8044
rect 7956 7988 7960 8044
rect 7896 7984 7960 7988
rect 7976 8044 8040 8048
rect 7976 7988 7980 8044
rect 7980 7988 8036 8044
rect 8036 7988 8040 8044
rect 7976 7984 8040 7988
rect 8056 8044 8120 8048
rect 8056 7988 8060 8044
rect 8060 7988 8116 8044
rect 8116 7988 8120 8044
rect 8056 7984 8120 7988
rect 14680 8044 14744 8048
rect 14680 7988 14684 8044
rect 14684 7988 14740 8044
rect 14740 7988 14744 8044
rect 14680 7984 14744 7988
rect 14760 8044 14824 8048
rect 14760 7988 14764 8044
rect 14764 7988 14820 8044
rect 14820 7988 14824 8044
rect 14760 7984 14824 7988
rect 14840 8044 14904 8048
rect 14840 7988 14844 8044
rect 14844 7988 14900 8044
rect 14900 7988 14904 8044
rect 14840 7984 14904 7988
rect 14920 8044 14984 8048
rect 14920 7988 14924 8044
rect 14924 7988 14980 8044
rect 14980 7988 14984 8044
rect 14920 7984 14984 7988
rect 4384 7500 4448 7504
rect 4384 7444 4388 7500
rect 4388 7444 4444 7500
rect 4444 7444 4448 7500
rect 4384 7440 4448 7444
rect 4464 7500 4528 7504
rect 4464 7444 4468 7500
rect 4468 7444 4524 7500
rect 4524 7444 4528 7500
rect 4464 7440 4528 7444
rect 4544 7500 4608 7504
rect 4544 7444 4548 7500
rect 4548 7444 4604 7500
rect 4604 7444 4608 7500
rect 4544 7440 4608 7444
rect 4624 7500 4688 7504
rect 4624 7444 4628 7500
rect 4628 7444 4684 7500
rect 4684 7444 4688 7500
rect 4624 7440 4688 7444
rect 11248 7500 11312 7504
rect 11248 7444 11252 7500
rect 11252 7444 11308 7500
rect 11308 7444 11312 7500
rect 11248 7440 11312 7444
rect 11328 7500 11392 7504
rect 11328 7444 11332 7500
rect 11332 7444 11388 7500
rect 11388 7444 11392 7500
rect 11328 7440 11392 7444
rect 11408 7500 11472 7504
rect 11408 7444 11412 7500
rect 11412 7444 11468 7500
rect 11468 7444 11472 7500
rect 11408 7440 11472 7444
rect 11488 7500 11552 7504
rect 11488 7444 11492 7500
rect 11492 7444 11548 7500
rect 11548 7444 11552 7500
rect 11488 7440 11552 7444
rect 18112 7500 18176 7504
rect 18112 7444 18116 7500
rect 18116 7444 18172 7500
rect 18172 7444 18176 7500
rect 18112 7440 18176 7444
rect 18192 7500 18256 7504
rect 18192 7444 18196 7500
rect 18196 7444 18252 7500
rect 18252 7444 18256 7500
rect 18192 7440 18256 7444
rect 18272 7500 18336 7504
rect 18272 7444 18276 7500
rect 18276 7444 18332 7500
rect 18332 7444 18336 7500
rect 18272 7440 18336 7444
rect 18352 7500 18416 7504
rect 18352 7444 18356 7500
rect 18356 7444 18412 7500
rect 18412 7444 18416 7500
rect 18352 7440 18416 7444
rect 7816 6956 7880 6960
rect 7816 6900 7820 6956
rect 7820 6900 7876 6956
rect 7876 6900 7880 6956
rect 7816 6896 7880 6900
rect 7896 6956 7960 6960
rect 7896 6900 7900 6956
rect 7900 6900 7956 6956
rect 7956 6900 7960 6956
rect 7896 6896 7960 6900
rect 7976 6956 8040 6960
rect 7976 6900 7980 6956
rect 7980 6900 8036 6956
rect 8036 6900 8040 6956
rect 7976 6896 8040 6900
rect 8056 6956 8120 6960
rect 8056 6900 8060 6956
rect 8060 6900 8116 6956
rect 8116 6900 8120 6956
rect 8056 6896 8120 6900
rect 14680 6956 14744 6960
rect 14680 6900 14684 6956
rect 14684 6900 14740 6956
rect 14740 6900 14744 6956
rect 14680 6896 14744 6900
rect 14760 6956 14824 6960
rect 14760 6900 14764 6956
rect 14764 6900 14820 6956
rect 14820 6900 14824 6956
rect 14760 6896 14824 6900
rect 14840 6956 14904 6960
rect 14840 6900 14844 6956
rect 14844 6900 14900 6956
rect 14900 6900 14904 6956
rect 14840 6896 14904 6900
rect 14920 6956 14984 6960
rect 14920 6900 14924 6956
rect 14924 6900 14980 6956
rect 14980 6900 14984 6956
rect 14920 6896 14984 6900
rect 4384 6412 4448 6416
rect 4384 6356 4388 6412
rect 4388 6356 4444 6412
rect 4444 6356 4448 6412
rect 4384 6352 4448 6356
rect 4464 6412 4528 6416
rect 4464 6356 4468 6412
rect 4468 6356 4524 6412
rect 4524 6356 4528 6412
rect 4464 6352 4528 6356
rect 4544 6412 4608 6416
rect 4544 6356 4548 6412
rect 4548 6356 4604 6412
rect 4604 6356 4608 6412
rect 4544 6352 4608 6356
rect 4624 6412 4688 6416
rect 4624 6356 4628 6412
rect 4628 6356 4684 6412
rect 4684 6356 4688 6412
rect 4624 6352 4688 6356
rect 11248 6412 11312 6416
rect 11248 6356 11252 6412
rect 11252 6356 11308 6412
rect 11308 6356 11312 6412
rect 11248 6352 11312 6356
rect 11328 6412 11392 6416
rect 11328 6356 11332 6412
rect 11332 6356 11388 6412
rect 11388 6356 11392 6412
rect 11328 6352 11392 6356
rect 11408 6412 11472 6416
rect 11408 6356 11412 6412
rect 11412 6356 11468 6412
rect 11468 6356 11472 6412
rect 11408 6352 11472 6356
rect 11488 6412 11552 6416
rect 11488 6356 11492 6412
rect 11492 6356 11548 6412
rect 11548 6356 11552 6412
rect 11488 6352 11552 6356
rect 18112 6412 18176 6416
rect 18112 6356 18116 6412
rect 18116 6356 18172 6412
rect 18172 6356 18176 6412
rect 18112 6352 18176 6356
rect 18192 6412 18256 6416
rect 18192 6356 18196 6412
rect 18196 6356 18252 6412
rect 18252 6356 18256 6412
rect 18192 6352 18256 6356
rect 18272 6412 18336 6416
rect 18272 6356 18276 6412
rect 18276 6356 18332 6412
rect 18332 6356 18336 6412
rect 18272 6352 18336 6356
rect 18352 6412 18416 6416
rect 18352 6356 18356 6412
rect 18356 6356 18412 6412
rect 18412 6356 18416 6412
rect 18352 6352 18416 6356
rect 7816 5868 7880 5872
rect 7816 5812 7820 5868
rect 7820 5812 7876 5868
rect 7876 5812 7880 5868
rect 7816 5808 7880 5812
rect 7896 5868 7960 5872
rect 7896 5812 7900 5868
rect 7900 5812 7956 5868
rect 7956 5812 7960 5868
rect 7896 5808 7960 5812
rect 7976 5868 8040 5872
rect 7976 5812 7980 5868
rect 7980 5812 8036 5868
rect 8036 5812 8040 5868
rect 7976 5808 8040 5812
rect 8056 5868 8120 5872
rect 8056 5812 8060 5868
rect 8060 5812 8116 5868
rect 8116 5812 8120 5868
rect 8056 5808 8120 5812
rect 14680 5868 14744 5872
rect 14680 5812 14684 5868
rect 14684 5812 14740 5868
rect 14740 5812 14744 5868
rect 14680 5808 14744 5812
rect 14760 5868 14824 5872
rect 14760 5812 14764 5868
rect 14764 5812 14820 5868
rect 14820 5812 14824 5868
rect 14760 5808 14824 5812
rect 14840 5868 14904 5872
rect 14840 5812 14844 5868
rect 14844 5812 14900 5868
rect 14900 5812 14904 5868
rect 14840 5808 14904 5812
rect 14920 5868 14984 5872
rect 14920 5812 14924 5868
rect 14924 5812 14980 5868
rect 14980 5812 14984 5868
rect 14920 5808 14984 5812
rect 4384 5324 4448 5328
rect 4384 5268 4388 5324
rect 4388 5268 4444 5324
rect 4444 5268 4448 5324
rect 4384 5264 4448 5268
rect 4464 5324 4528 5328
rect 4464 5268 4468 5324
rect 4468 5268 4524 5324
rect 4524 5268 4528 5324
rect 4464 5264 4528 5268
rect 4544 5324 4608 5328
rect 4544 5268 4548 5324
rect 4548 5268 4604 5324
rect 4604 5268 4608 5324
rect 4544 5264 4608 5268
rect 4624 5324 4688 5328
rect 4624 5268 4628 5324
rect 4628 5268 4684 5324
rect 4684 5268 4688 5324
rect 4624 5264 4688 5268
rect 11248 5324 11312 5328
rect 11248 5268 11252 5324
rect 11252 5268 11308 5324
rect 11308 5268 11312 5324
rect 11248 5264 11312 5268
rect 11328 5324 11392 5328
rect 11328 5268 11332 5324
rect 11332 5268 11388 5324
rect 11388 5268 11392 5324
rect 11328 5264 11392 5268
rect 11408 5324 11472 5328
rect 11408 5268 11412 5324
rect 11412 5268 11468 5324
rect 11468 5268 11472 5324
rect 11408 5264 11472 5268
rect 11488 5324 11552 5328
rect 11488 5268 11492 5324
rect 11492 5268 11548 5324
rect 11548 5268 11552 5324
rect 11488 5264 11552 5268
rect 18112 5324 18176 5328
rect 18112 5268 18116 5324
rect 18116 5268 18172 5324
rect 18172 5268 18176 5324
rect 18112 5264 18176 5268
rect 18192 5324 18256 5328
rect 18192 5268 18196 5324
rect 18196 5268 18252 5324
rect 18252 5268 18256 5324
rect 18192 5264 18256 5268
rect 18272 5324 18336 5328
rect 18272 5268 18276 5324
rect 18276 5268 18332 5324
rect 18332 5268 18336 5324
rect 18272 5264 18336 5268
rect 18352 5324 18416 5328
rect 18352 5268 18356 5324
rect 18356 5268 18412 5324
rect 18412 5268 18416 5324
rect 18352 5264 18416 5268
rect 7816 4780 7880 4784
rect 7816 4724 7820 4780
rect 7820 4724 7876 4780
rect 7876 4724 7880 4780
rect 7816 4720 7880 4724
rect 7896 4780 7960 4784
rect 7896 4724 7900 4780
rect 7900 4724 7956 4780
rect 7956 4724 7960 4780
rect 7896 4720 7960 4724
rect 7976 4780 8040 4784
rect 7976 4724 7980 4780
rect 7980 4724 8036 4780
rect 8036 4724 8040 4780
rect 7976 4720 8040 4724
rect 8056 4780 8120 4784
rect 8056 4724 8060 4780
rect 8060 4724 8116 4780
rect 8116 4724 8120 4780
rect 8056 4720 8120 4724
rect 14680 4780 14744 4784
rect 14680 4724 14684 4780
rect 14684 4724 14740 4780
rect 14740 4724 14744 4780
rect 14680 4720 14744 4724
rect 14760 4780 14824 4784
rect 14760 4724 14764 4780
rect 14764 4724 14820 4780
rect 14820 4724 14824 4780
rect 14760 4720 14824 4724
rect 14840 4780 14904 4784
rect 14840 4724 14844 4780
rect 14844 4724 14900 4780
rect 14900 4724 14904 4780
rect 14840 4720 14904 4724
rect 14920 4780 14984 4784
rect 14920 4724 14924 4780
rect 14924 4724 14980 4780
rect 14980 4724 14984 4780
rect 14920 4720 14984 4724
rect 4384 4236 4448 4240
rect 4384 4180 4388 4236
rect 4388 4180 4444 4236
rect 4444 4180 4448 4236
rect 4384 4176 4448 4180
rect 4464 4236 4528 4240
rect 4464 4180 4468 4236
rect 4468 4180 4524 4236
rect 4524 4180 4528 4236
rect 4464 4176 4528 4180
rect 4544 4236 4608 4240
rect 4544 4180 4548 4236
rect 4548 4180 4604 4236
rect 4604 4180 4608 4236
rect 4544 4176 4608 4180
rect 4624 4236 4688 4240
rect 4624 4180 4628 4236
rect 4628 4180 4684 4236
rect 4684 4180 4688 4236
rect 4624 4176 4688 4180
rect 11248 4236 11312 4240
rect 11248 4180 11252 4236
rect 11252 4180 11308 4236
rect 11308 4180 11312 4236
rect 11248 4176 11312 4180
rect 11328 4236 11392 4240
rect 11328 4180 11332 4236
rect 11332 4180 11388 4236
rect 11388 4180 11392 4236
rect 11328 4176 11392 4180
rect 11408 4236 11472 4240
rect 11408 4180 11412 4236
rect 11412 4180 11468 4236
rect 11468 4180 11472 4236
rect 11408 4176 11472 4180
rect 11488 4236 11552 4240
rect 11488 4180 11492 4236
rect 11492 4180 11548 4236
rect 11548 4180 11552 4236
rect 11488 4176 11552 4180
rect 18112 4236 18176 4240
rect 18112 4180 18116 4236
rect 18116 4180 18172 4236
rect 18172 4180 18176 4236
rect 18112 4176 18176 4180
rect 18192 4236 18256 4240
rect 18192 4180 18196 4236
rect 18196 4180 18252 4236
rect 18252 4180 18256 4236
rect 18192 4176 18256 4180
rect 18272 4236 18336 4240
rect 18272 4180 18276 4236
rect 18276 4180 18332 4236
rect 18332 4180 18336 4236
rect 18272 4176 18336 4180
rect 18352 4236 18416 4240
rect 18352 4180 18356 4236
rect 18356 4180 18412 4236
rect 18412 4180 18416 4236
rect 18352 4176 18416 4180
rect 7816 3692 7880 3696
rect 7816 3636 7820 3692
rect 7820 3636 7876 3692
rect 7876 3636 7880 3692
rect 7816 3632 7880 3636
rect 7896 3692 7960 3696
rect 7896 3636 7900 3692
rect 7900 3636 7956 3692
rect 7956 3636 7960 3692
rect 7896 3632 7960 3636
rect 7976 3692 8040 3696
rect 7976 3636 7980 3692
rect 7980 3636 8036 3692
rect 8036 3636 8040 3692
rect 7976 3632 8040 3636
rect 8056 3692 8120 3696
rect 8056 3636 8060 3692
rect 8060 3636 8116 3692
rect 8116 3636 8120 3692
rect 8056 3632 8120 3636
rect 14680 3692 14744 3696
rect 14680 3636 14684 3692
rect 14684 3636 14740 3692
rect 14740 3636 14744 3692
rect 14680 3632 14744 3636
rect 14760 3692 14824 3696
rect 14760 3636 14764 3692
rect 14764 3636 14820 3692
rect 14820 3636 14824 3692
rect 14760 3632 14824 3636
rect 14840 3692 14904 3696
rect 14840 3636 14844 3692
rect 14844 3636 14900 3692
rect 14900 3636 14904 3692
rect 14840 3632 14904 3636
rect 14920 3692 14984 3696
rect 14920 3636 14924 3692
rect 14924 3636 14980 3692
rect 14980 3636 14984 3692
rect 14920 3632 14984 3636
rect 4384 3148 4448 3152
rect 4384 3092 4388 3148
rect 4388 3092 4444 3148
rect 4444 3092 4448 3148
rect 4384 3088 4448 3092
rect 4464 3148 4528 3152
rect 4464 3092 4468 3148
rect 4468 3092 4524 3148
rect 4524 3092 4528 3148
rect 4464 3088 4528 3092
rect 4544 3148 4608 3152
rect 4544 3092 4548 3148
rect 4548 3092 4604 3148
rect 4604 3092 4608 3148
rect 4544 3088 4608 3092
rect 4624 3148 4688 3152
rect 4624 3092 4628 3148
rect 4628 3092 4684 3148
rect 4684 3092 4688 3148
rect 4624 3088 4688 3092
rect 11248 3148 11312 3152
rect 11248 3092 11252 3148
rect 11252 3092 11308 3148
rect 11308 3092 11312 3148
rect 11248 3088 11312 3092
rect 11328 3148 11392 3152
rect 11328 3092 11332 3148
rect 11332 3092 11388 3148
rect 11388 3092 11392 3148
rect 11328 3088 11392 3092
rect 11408 3148 11472 3152
rect 11408 3092 11412 3148
rect 11412 3092 11468 3148
rect 11468 3092 11472 3148
rect 11408 3088 11472 3092
rect 11488 3148 11552 3152
rect 11488 3092 11492 3148
rect 11492 3092 11548 3148
rect 11548 3092 11552 3148
rect 11488 3088 11552 3092
rect 18112 3148 18176 3152
rect 18112 3092 18116 3148
rect 18116 3092 18172 3148
rect 18172 3092 18176 3148
rect 18112 3088 18176 3092
rect 18192 3148 18256 3152
rect 18192 3092 18196 3148
rect 18196 3092 18252 3148
rect 18252 3092 18256 3148
rect 18192 3088 18256 3092
rect 18272 3148 18336 3152
rect 18272 3092 18276 3148
rect 18276 3092 18332 3148
rect 18332 3092 18336 3148
rect 18272 3088 18336 3092
rect 18352 3148 18416 3152
rect 18352 3092 18356 3148
rect 18356 3092 18412 3148
rect 18412 3092 18416 3148
rect 18352 3088 18416 3092
rect 7816 2604 7880 2608
rect 7816 2548 7820 2604
rect 7820 2548 7876 2604
rect 7876 2548 7880 2604
rect 7816 2544 7880 2548
rect 7896 2604 7960 2608
rect 7896 2548 7900 2604
rect 7900 2548 7956 2604
rect 7956 2548 7960 2604
rect 7896 2544 7960 2548
rect 7976 2604 8040 2608
rect 7976 2548 7980 2604
rect 7980 2548 8036 2604
rect 8036 2548 8040 2604
rect 7976 2544 8040 2548
rect 8056 2604 8120 2608
rect 8056 2548 8060 2604
rect 8060 2548 8116 2604
rect 8116 2548 8120 2604
rect 8056 2544 8120 2548
rect 14680 2604 14744 2608
rect 14680 2548 14684 2604
rect 14684 2548 14740 2604
rect 14740 2548 14744 2604
rect 14680 2544 14744 2548
rect 14760 2604 14824 2608
rect 14760 2548 14764 2604
rect 14764 2548 14820 2604
rect 14820 2548 14824 2604
rect 14760 2544 14824 2548
rect 14840 2604 14904 2608
rect 14840 2548 14844 2604
rect 14844 2548 14900 2604
rect 14900 2548 14904 2604
rect 14840 2544 14904 2548
rect 14920 2604 14984 2608
rect 14920 2548 14924 2604
rect 14924 2548 14980 2604
rect 14980 2548 14984 2604
rect 14920 2544 14984 2548
rect 4384 2060 4448 2064
rect 4384 2004 4388 2060
rect 4388 2004 4444 2060
rect 4444 2004 4448 2060
rect 4384 2000 4448 2004
rect 4464 2060 4528 2064
rect 4464 2004 4468 2060
rect 4468 2004 4524 2060
rect 4524 2004 4528 2060
rect 4464 2000 4528 2004
rect 4544 2060 4608 2064
rect 4544 2004 4548 2060
rect 4548 2004 4604 2060
rect 4604 2004 4608 2060
rect 4544 2000 4608 2004
rect 4624 2060 4688 2064
rect 4624 2004 4628 2060
rect 4628 2004 4684 2060
rect 4684 2004 4688 2060
rect 4624 2000 4688 2004
rect 11248 2060 11312 2064
rect 11248 2004 11252 2060
rect 11252 2004 11308 2060
rect 11308 2004 11312 2060
rect 11248 2000 11312 2004
rect 11328 2060 11392 2064
rect 11328 2004 11332 2060
rect 11332 2004 11388 2060
rect 11388 2004 11392 2060
rect 11328 2000 11392 2004
rect 11408 2060 11472 2064
rect 11408 2004 11412 2060
rect 11412 2004 11468 2060
rect 11468 2004 11472 2060
rect 11408 2000 11472 2004
rect 11488 2060 11552 2064
rect 11488 2004 11492 2060
rect 11492 2004 11548 2060
rect 11548 2004 11552 2060
rect 11488 2000 11552 2004
rect 18112 2060 18176 2064
rect 18112 2004 18116 2060
rect 18116 2004 18172 2060
rect 18172 2004 18176 2060
rect 18112 2000 18176 2004
rect 18192 2060 18256 2064
rect 18192 2004 18196 2060
rect 18196 2004 18252 2060
rect 18252 2004 18256 2060
rect 18192 2000 18256 2004
rect 18272 2060 18336 2064
rect 18272 2004 18276 2060
rect 18276 2004 18332 2060
rect 18332 2004 18336 2060
rect 18272 2000 18336 2004
rect 18352 2060 18416 2064
rect 18352 2004 18356 2060
rect 18356 2004 18412 2060
rect 18412 2004 18416 2060
rect 18352 2000 18416 2004
<< metal4 >>
rect 4376 19472 4696 20032
rect 4376 19408 4384 19472
rect 4448 19408 4464 19472
rect 4528 19408 4544 19472
rect 4608 19408 4624 19472
rect 4688 19408 4696 19472
rect 4376 18384 4696 19408
rect 4376 18320 4384 18384
rect 4448 18320 4464 18384
rect 4528 18320 4544 18384
rect 4608 18320 4624 18384
rect 4688 18320 4696 18384
rect 4376 17296 4696 18320
rect 4376 17232 4384 17296
rect 4448 17232 4464 17296
rect 4528 17232 4544 17296
rect 4608 17232 4624 17296
rect 4688 17232 4696 17296
rect 4376 16208 4696 17232
rect 4376 16144 4384 16208
rect 4448 16144 4464 16208
rect 4528 16144 4544 16208
rect 4608 16144 4624 16208
rect 4688 16144 4696 16208
rect 4376 15120 4696 16144
rect 4376 15056 4384 15120
rect 4448 15056 4464 15120
rect 4528 15056 4544 15120
rect 4608 15056 4624 15120
rect 4688 15056 4696 15120
rect 4376 14032 4696 15056
rect 4376 13968 4384 14032
rect 4448 13968 4464 14032
rect 4528 13968 4544 14032
rect 4608 13968 4624 14032
rect 4688 13968 4696 14032
rect 4376 12944 4696 13968
rect 4376 12880 4384 12944
rect 4448 12880 4464 12944
rect 4528 12880 4544 12944
rect 4608 12880 4624 12944
rect 4688 12880 4696 12944
rect 4376 11856 4696 12880
rect 4376 11792 4384 11856
rect 4448 11792 4464 11856
rect 4528 11792 4544 11856
rect 4608 11792 4624 11856
rect 4688 11792 4696 11856
rect 4376 10768 4696 11792
rect 4376 10704 4384 10768
rect 4448 10704 4464 10768
rect 4528 10704 4544 10768
rect 4608 10704 4624 10768
rect 4688 10704 4696 10768
rect 4376 9680 4696 10704
rect 4376 9616 4384 9680
rect 4448 9616 4464 9680
rect 4528 9616 4544 9680
rect 4608 9616 4624 9680
rect 4688 9616 4696 9680
rect 4376 8592 4696 9616
rect 4376 8528 4384 8592
rect 4448 8528 4464 8592
rect 4528 8528 4544 8592
rect 4608 8528 4624 8592
rect 4688 8528 4696 8592
rect 4376 7504 4696 8528
rect 4376 7440 4384 7504
rect 4448 7440 4464 7504
rect 4528 7440 4544 7504
rect 4608 7440 4624 7504
rect 4688 7440 4696 7504
rect 4376 6416 4696 7440
rect 4376 6352 4384 6416
rect 4448 6352 4464 6416
rect 4528 6352 4544 6416
rect 4608 6352 4624 6416
rect 4688 6352 4696 6416
rect 4376 5328 4696 6352
rect 4376 5264 4384 5328
rect 4448 5264 4464 5328
rect 4528 5264 4544 5328
rect 4608 5264 4624 5328
rect 4688 5264 4696 5328
rect 4376 4240 4696 5264
rect 4376 4176 4384 4240
rect 4448 4176 4464 4240
rect 4528 4176 4544 4240
rect 4608 4176 4624 4240
rect 4688 4176 4696 4240
rect 4376 3152 4696 4176
rect 4376 3088 4384 3152
rect 4448 3088 4464 3152
rect 4528 3088 4544 3152
rect 4608 3088 4624 3152
rect 4688 3088 4696 3152
rect 4376 2064 4696 3088
rect 4376 2000 4384 2064
rect 4448 2000 4464 2064
rect 4528 2000 4544 2064
rect 4608 2000 4624 2064
rect 4688 2000 4696 2064
rect 4376 1984 4696 2000
rect 7808 20016 8128 20032
rect 7808 19952 7816 20016
rect 7880 19952 7896 20016
rect 7960 19952 7976 20016
rect 8040 19952 8056 20016
rect 8120 19952 8128 20016
rect 7808 18928 8128 19952
rect 7808 18864 7816 18928
rect 7880 18864 7896 18928
rect 7960 18864 7976 18928
rect 8040 18864 8056 18928
rect 8120 18864 8128 18928
rect 7808 17840 8128 18864
rect 7808 17776 7816 17840
rect 7880 17776 7896 17840
rect 7960 17776 7976 17840
rect 8040 17776 8056 17840
rect 8120 17776 8128 17840
rect 7808 16752 8128 17776
rect 7808 16688 7816 16752
rect 7880 16688 7896 16752
rect 7960 16688 7976 16752
rect 8040 16688 8056 16752
rect 8120 16688 8128 16752
rect 7808 15664 8128 16688
rect 7808 15600 7816 15664
rect 7880 15600 7896 15664
rect 7960 15600 7976 15664
rect 8040 15600 8056 15664
rect 8120 15600 8128 15664
rect 7808 14576 8128 15600
rect 7808 14512 7816 14576
rect 7880 14512 7896 14576
rect 7960 14512 7976 14576
rect 8040 14512 8056 14576
rect 8120 14512 8128 14576
rect 7808 13488 8128 14512
rect 7808 13424 7816 13488
rect 7880 13424 7896 13488
rect 7960 13424 7976 13488
rect 8040 13424 8056 13488
rect 8120 13424 8128 13488
rect 7808 12400 8128 13424
rect 7808 12336 7816 12400
rect 7880 12336 7896 12400
rect 7960 12336 7976 12400
rect 8040 12336 8056 12400
rect 8120 12336 8128 12400
rect 7808 11312 8128 12336
rect 7808 11248 7816 11312
rect 7880 11248 7896 11312
rect 7960 11248 7976 11312
rect 8040 11248 8056 11312
rect 8120 11248 8128 11312
rect 7808 10224 8128 11248
rect 7808 10160 7816 10224
rect 7880 10160 7896 10224
rect 7960 10160 7976 10224
rect 8040 10160 8056 10224
rect 8120 10160 8128 10224
rect 7808 9136 8128 10160
rect 7808 9072 7816 9136
rect 7880 9072 7896 9136
rect 7960 9072 7976 9136
rect 8040 9072 8056 9136
rect 8120 9072 8128 9136
rect 7808 8048 8128 9072
rect 7808 7984 7816 8048
rect 7880 7984 7896 8048
rect 7960 7984 7976 8048
rect 8040 7984 8056 8048
rect 8120 7984 8128 8048
rect 7808 6960 8128 7984
rect 7808 6896 7816 6960
rect 7880 6896 7896 6960
rect 7960 6896 7976 6960
rect 8040 6896 8056 6960
rect 8120 6896 8128 6960
rect 7808 5872 8128 6896
rect 7808 5808 7816 5872
rect 7880 5808 7896 5872
rect 7960 5808 7976 5872
rect 8040 5808 8056 5872
rect 8120 5808 8128 5872
rect 7808 4784 8128 5808
rect 7808 4720 7816 4784
rect 7880 4720 7896 4784
rect 7960 4720 7976 4784
rect 8040 4720 8056 4784
rect 8120 4720 8128 4784
rect 7808 3696 8128 4720
rect 7808 3632 7816 3696
rect 7880 3632 7896 3696
rect 7960 3632 7976 3696
rect 8040 3632 8056 3696
rect 8120 3632 8128 3696
rect 7808 2608 8128 3632
rect 7808 2544 7816 2608
rect 7880 2544 7896 2608
rect 7960 2544 7976 2608
rect 8040 2544 8056 2608
rect 8120 2544 8128 2608
rect 7808 1984 8128 2544
rect 11240 19472 11560 20032
rect 11240 19408 11248 19472
rect 11312 19408 11328 19472
rect 11392 19408 11408 19472
rect 11472 19408 11488 19472
rect 11552 19408 11560 19472
rect 11240 18384 11560 19408
rect 11240 18320 11248 18384
rect 11312 18320 11328 18384
rect 11392 18320 11408 18384
rect 11472 18320 11488 18384
rect 11552 18320 11560 18384
rect 11240 17296 11560 18320
rect 11240 17232 11248 17296
rect 11312 17232 11328 17296
rect 11392 17232 11408 17296
rect 11472 17232 11488 17296
rect 11552 17232 11560 17296
rect 11240 16208 11560 17232
rect 11240 16144 11248 16208
rect 11312 16144 11328 16208
rect 11392 16144 11408 16208
rect 11472 16144 11488 16208
rect 11552 16144 11560 16208
rect 11240 15120 11560 16144
rect 11240 15056 11248 15120
rect 11312 15056 11328 15120
rect 11392 15056 11408 15120
rect 11472 15056 11488 15120
rect 11552 15056 11560 15120
rect 11240 14032 11560 15056
rect 11240 13968 11248 14032
rect 11312 13968 11328 14032
rect 11392 13968 11408 14032
rect 11472 13968 11488 14032
rect 11552 13968 11560 14032
rect 11240 12944 11560 13968
rect 11240 12880 11248 12944
rect 11312 12880 11328 12944
rect 11392 12880 11408 12944
rect 11472 12880 11488 12944
rect 11552 12880 11560 12944
rect 11240 11856 11560 12880
rect 11240 11792 11248 11856
rect 11312 11792 11328 11856
rect 11392 11792 11408 11856
rect 11472 11792 11488 11856
rect 11552 11792 11560 11856
rect 11240 10768 11560 11792
rect 11240 10704 11248 10768
rect 11312 10704 11328 10768
rect 11392 10704 11408 10768
rect 11472 10704 11488 10768
rect 11552 10704 11560 10768
rect 11240 9680 11560 10704
rect 11240 9616 11248 9680
rect 11312 9616 11328 9680
rect 11392 9616 11408 9680
rect 11472 9616 11488 9680
rect 11552 9616 11560 9680
rect 11240 8592 11560 9616
rect 11240 8528 11248 8592
rect 11312 8528 11328 8592
rect 11392 8528 11408 8592
rect 11472 8528 11488 8592
rect 11552 8528 11560 8592
rect 11240 7504 11560 8528
rect 11240 7440 11248 7504
rect 11312 7440 11328 7504
rect 11392 7440 11408 7504
rect 11472 7440 11488 7504
rect 11552 7440 11560 7504
rect 11240 6416 11560 7440
rect 11240 6352 11248 6416
rect 11312 6352 11328 6416
rect 11392 6352 11408 6416
rect 11472 6352 11488 6416
rect 11552 6352 11560 6416
rect 11240 5328 11560 6352
rect 11240 5264 11248 5328
rect 11312 5264 11328 5328
rect 11392 5264 11408 5328
rect 11472 5264 11488 5328
rect 11552 5264 11560 5328
rect 11240 4240 11560 5264
rect 11240 4176 11248 4240
rect 11312 4176 11328 4240
rect 11392 4176 11408 4240
rect 11472 4176 11488 4240
rect 11552 4176 11560 4240
rect 11240 3152 11560 4176
rect 11240 3088 11248 3152
rect 11312 3088 11328 3152
rect 11392 3088 11408 3152
rect 11472 3088 11488 3152
rect 11552 3088 11560 3152
rect 11240 2064 11560 3088
rect 11240 2000 11248 2064
rect 11312 2000 11328 2064
rect 11392 2000 11408 2064
rect 11472 2000 11488 2064
rect 11552 2000 11560 2064
rect 11240 1984 11560 2000
rect 14672 20016 14992 20032
rect 14672 19952 14680 20016
rect 14744 19952 14760 20016
rect 14824 19952 14840 20016
rect 14904 19952 14920 20016
rect 14984 19952 14992 20016
rect 14672 18928 14992 19952
rect 14672 18864 14680 18928
rect 14744 18864 14760 18928
rect 14824 18864 14840 18928
rect 14904 18864 14920 18928
rect 14984 18864 14992 18928
rect 14672 17840 14992 18864
rect 14672 17776 14680 17840
rect 14744 17776 14760 17840
rect 14824 17776 14840 17840
rect 14904 17776 14920 17840
rect 14984 17776 14992 17840
rect 14672 16752 14992 17776
rect 14672 16688 14680 16752
rect 14744 16688 14760 16752
rect 14824 16688 14840 16752
rect 14904 16688 14920 16752
rect 14984 16688 14992 16752
rect 14672 15664 14992 16688
rect 14672 15600 14680 15664
rect 14744 15600 14760 15664
rect 14824 15600 14840 15664
rect 14904 15600 14920 15664
rect 14984 15600 14992 15664
rect 14672 14576 14992 15600
rect 14672 14512 14680 14576
rect 14744 14512 14760 14576
rect 14824 14512 14840 14576
rect 14904 14512 14920 14576
rect 14984 14512 14992 14576
rect 14672 13488 14992 14512
rect 14672 13424 14680 13488
rect 14744 13424 14760 13488
rect 14824 13424 14840 13488
rect 14904 13424 14920 13488
rect 14984 13424 14992 13488
rect 14672 12400 14992 13424
rect 14672 12336 14680 12400
rect 14744 12336 14760 12400
rect 14824 12336 14840 12400
rect 14904 12336 14920 12400
rect 14984 12336 14992 12400
rect 14672 11312 14992 12336
rect 14672 11248 14680 11312
rect 14744 11248 14760 11312
rect 14824 11248 14840 11312
rect 14904 11248 14920 11312
rect 14984 11248 14992 11312
rect 14672 10224 14992 11248
rect 14672 10160 14680 10224
rect 14744 10160 14760 10224
rect 14824 10160 14840 10224
rect 14904 10160 14920 10224
rect 14984 10160 14992 10224
rect 14672 9136 14992 10160
rect 14672 9072 14680 9136
rect 14744 9072 14760 9136
rect 14824 9072 14840 9136
rect 14904 9072 14920 9136
rect 14984 9072 14992 9136
rect 14672 8048 14992 9072
rect 14672 7984 14680 8048
rect 14744 7984 14760 8048
rect 14824 7984 14840 8048
rect 14904 7984 14920 8048
rect 14984 7984 14992 8048
rect 14672 6960 14992 7984
rect 14672 6896 14680 6960
rect 14744 6896 14760 6960
rect 14824 6896 14840 6960
rect 14904 6896 14920 6960
rect 14984 6896 14992 6960
rect 14672 5872 14992 6896
rect 14672 5808 14680 5872
rect 14744 5808 14760 5872
rect 14824 5808 14840 5872
rect 14904 5808 14920 5872
rect 14984 5808 14992 5872
rect 14672 4784 14992 5808
rect 14672 4720 14680 4784
rect 14744 4720 14760 4784
rect 14824 4720 14840 4784
rect 14904 4720 14920 4784
rect 14984 4720 14992 4784
rect 14672 3696 14992 4720
rect 14672 3632 14680 3696
rect 14744 3632 14760 3696
rect 14824 3632 14840 3696
rect 14904 3632 14920 3696
rect 14984 3632 14992 3696
rect 14672 2608 14992 3632
rect 14672 2544 14680 2608
rect 14744 2544 14760 2608
rect 14824 2544 14840 2608
rect 14904 2544 14920 2608
rect 14984 2544 14992 2608
rect 14672 1984 14992 2544
rect 18104 19472 18424 20032
rect 18104 19408 18112 19472
rect 18176 19408 18192 19472
rect 18256 19408 18272 19472
rect 18336 19408 18352 19472
rect 18416 19408 18424 19472
rect 18104 18384 18424 19408
rect 19379 18588 19445 18589
rect 19379 18524 19380 18588
rect 19444 18524 19445 18588
rect 19379 18523 19445 18524
rect 18104 18320 18112 18384
rect 18176 18320 18192 18384
rect 18256 18320 18272 18384
rect 18336 18320 18352 18384
rect 18416 18320 18424 18384
rect 18104 17296 18424 18320
rect 18104 17232 18112 17296
rect 18176 17232 18192 17296
rect 18256 17232 18272 17296
rect 18336 17232 18352 17296
rect 18416 17232 18424 17296
rect 18104 16208 18424 17232
rect 18104 16144 18112 16208
rect 18176 16144 18192 16208
rect 18256 16144 18272 16208
rect 18336 16144 18352 16208
rect 18416 16144 18424 16208
rect 18104 15120 18424 16144
rect 18104 15056 18112 15120
rect 18176 15056 18192 15120
rect 18256 15056 18272 15120
rect 18336 15056 18352 15120
rect 18416 15056 18424 15120
rect 18104 14032 18424 15056
rect 18104 13968 18112 14032
rect 18176 13968 18192 14032
rect 18256 13968 18272 14032
rect 18336 13968 18352 14032
rect 18416 13968 18424 14032
rect 18104 12944 18424 13968
rect 19382 13693 19442 18523
rect 19379 13692 19445 13693
rect 19379 13628 19380 13692
rect 19444 13628 19445 13692
rect 19379 13627 19445 13628
rect 18104 12880 18112 12944
rect 18176 12880 18192 12944
rect 18256 12880 18272 12944
rect 18336 12880 18352 12944
rect 18416 12880 18424 12944
rect 18104 11856 18424 12880
rect 18104 11792 18112 11856
rect 18176 11792 18192 11856
rect 18256 11792 18272 11856
rect 18336 11792 18352 11856
rect 18416 11792 18424 11856
rect 18104 10768 18424 11792
rect 18104 10704 18112 10768
rect 18176 10704 18192 10768
rect 18256 10704 18272 10768
rect 18336 10704 18352 10768
rect 18416 10704 18424 10768
rect 18104 9680 18424 10704
rect 18104 9616 18112 9680
rect 18176 9616 18192 9680
rect 18256 9616 18272 9680
rect 18336 9616 18352 9680
rect 18416 9616 18424 9680
rect 18104 8592 18424 9616
rect 18104 8528 18112 8592
rect 18176 8528 18192 8592
rect 18256 8528 18272 8592
rect 18336 8528 18352 8592
rect 18416 8528 18424 8592
rect 18104 7504 18424 8528
rect 18104 7440 18112 7504
rect 18176 7440 18192 7504
rect 18256 7440 18272 7504
rect 18336 7440 18352 7504
rect 18416 7440 18424 7504
rect 18104 6416 18424 7440
rect 18104 6352 18112 6416
rect 18176 6352 18192 6416
rect 18256 6352 18272 6416
rect 18336 6352 18352 6416
rect 18416 6352 18424 6416
rect 18104 5328 18424 6352
rect 18104 5264 18112 5328
rect 18176 5264 18192 5328
rect 18256 5264 18272 5328
rect 18336 5264 18352 5328
rect 18416 5264 18424 5328
rect 18104 4240 18424 5264
rect 18104 4176 18112 4240
rect 18176 4176 18192 4240
rect 18256 4176 18272 4240
rect 18336 4176 18352 4240
rect 18416 4176 18424 4240
rect 18104 3152 18424 4176
rect 18104 3088 18112 3152
rect 18176 3088 18192 3152
rect 18256 3088 18272 3152
rect 18336 3088 18352 3152
rect 18416 3088 18424 3152
rect 18104 2064 18424 3088
rect 18104 2000 18112 2064
rect 18176 2000 18192 2064
rect 18256 2000 18272 2064
rect 18336 2000 18352 2064
rect 18416 2000 18424 2064
rect 18104 1984 18424 2000
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1608761684
transform 1 0 20516 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1608761684
transform -1 0 21620 0 -1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1608761684
transform 1 0 21068 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_209
timestamp 1608761684
transform 1 0 20332 0 -1 19984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1608761684
transform 1 0 20884 0 -1 19984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1608761684
transform 1 0 21160 0 -1 19984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1608761684
transform 1 0 19964 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_199
timestamp 1608761684
transform 1 0 19412 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1608761684
transform 1 0 18216 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_168
timestamp 1608761684
transform 1 0 16560 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_180
timestamp 1608761684
transform 1 0 17664 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_187
timestamp 1608761684
transform 1 0 18308 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1608761684
transform 1 0 15364 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_149
timestamp 1608761684
transform 1 0 14812 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_156
timestamp 1608761684
transform 1 0 15456 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_137
timestamp 1608761684
transform 1 0 13708 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1608761684
transform 1 0 12512 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_106
timestamp 1608761684
transform 1 0 10856 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_118
timestamp 1608761684
transform 1 0 11960 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_125
timestamp 1608761684
transform 1 0 12604 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1608761684
transform 1 0 9660 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_87
timestamp 1608761684
transform 1 0 9108 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_94
timestamp 1608761684
transform 1 0 9752 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1608761684
transform 1 0 6900 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_75
timestamp 1608761684
transform 1 0 8004 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1608761684
transform 1 0 6808 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1608761684
transform 1 0 5152 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_56
timestamp 1608761684
transform 1 0 6256 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1608761684
transform 1 0 3956 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1608761684
transform 1 0 3588 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1608761684
transform 1 0 4048 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1608761684
transform 1 0 1104 0 -1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1608761684
transform 1 0 1380 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1608761684
transform 1 0 2484 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1608761684
transform -1 0 21620 0 1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1608761684
transform 1 0 20792 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_212
timestamp 1608761684
transform 1 0 20608 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1608761684
transform 1 0 20884 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_219
timestamp 1608761684
transform 1 0 21252 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1608761684
transform 1 0 20240 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761684
transform 1 0 19412 0 1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_195
timestamp 1608761684
transform 1 0 19044 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_205
timestamp 1608761684
transform 1 0 19964 0 1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1608761684
transform 1 0 17388 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00
timestamp 1608761684
transform 1 0 17940 0 1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_174
timestamp 1608761684
transform 1 0 17112 0 1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1608761684
transform 1 0 17756 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1608761684
transform 1 0 15272 0 1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1608761684
transform 1 0 16284 0 1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1608761684
transform 1 0 15180 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_163
timestamp 1608761684
transform 1 0 16100 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1608761684
transform 1 0 13616 0 1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_31_126
timestamp 1608761684
transform 1 0 12696 0 1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_134
timestamp 1608761684
transform 1 0 13432 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_145
timestamp 1608761684
transform 1 0 14444 0 1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761684
transform 1 0 11224 0 1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1608761684
transform 1 0 9660 0 1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1608761684
transform 1 0 9568 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_86
timestamp 1608761684
transform 1 0 9016 0 1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_102
timestamp 1608761684
transform 1 0 10488 0 1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1608761684
transform 1 0 8740 0 1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1608761684
transform 1 0 7728 0 1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_81
timestamp 1608761684
transform 1 0 8556 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_48
timestamp 1608761684
transform 1 0 5520 0 1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_60
timestamp 1608761684
transform 1 0 6624 0 1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1608761684
transform 1 0 4692 0 1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1608761684
transform 1 0 3956 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_27
timestamp 1608761684
transform 1 0 3588 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_32
timestamp 1608761684
transform 1 0 4048 0 1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_38
timestamp 1608761684
transform 1 0 4600 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1608761684
transform 1 0 1104 0 1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1608761684
transform 1 0 1380 0 1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1608761684
transform 1 0 2484 0 1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1608761684
transform -1 0 21620 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_213
timestamp 1608761684
transform 1 0 20700 0 -1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1608761684
transform 1 0 21252 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761684
transform 1 0 19412 0 -1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761684
transform 1 0 20148 0 -1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_205
timestamp 1608761684
transform 1 0 19964 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1608761684
transform 1 0 18032 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1608761684
transform 1 0 17940 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_177
timestamp 1608761684
transform 1 0 17388 0 -1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_187
timestamp 1608761684
transform 1 0 18308 0 -1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761684
transform 1 0 15916 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_159
timestamp 1608761684
transform 1 0 15732 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761684
transform 1 0 14260 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1608761684
transform 1 0 14076 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1608761684
transform 1 0 11776 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761684
transform 1 0 12604 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1608761684
transform 1 0 12328 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_114
timestamp 1608761684
transform 1 0 11592 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_119
timestamp 1608761684
transform 1 0 12052 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_123
timestamp 1608761684
transform 1 0 12420 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761684
transform 1 0 10120 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_96
timestamp 1608761684
transform 1 0 9936 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761684
transform 1 0 8464 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_78
timestamp 1608761684
transform 1 0 8280 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761684
transform 1 0 6808 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1608761684
transform 1 0 5428 0 -1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1608761684
transform 1 0 6716 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_45
timestamp 1608761684
transform 1 0 5244 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_56
timestamp 1608761684
transform 1 0 6256 0 -1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_60
timestamp 1608761684
transform 1 0 6624 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761684
transform 1 0 3772 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_27
timestamp 1608761684
transform 1 0 3588 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761684
transform 1 0 2116 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1608761684
transform 1 0 1104 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1608761684
transform 1 0 1380 0 -1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1608761684
transform -1 0 21620 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1608761684
transform 1 0 20792 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_209
timestamp 1608761684
transform 1 0 20332 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_213
timestamp 1608761684
transform 1 0 20700 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_215
timestamp 1608761684
transform 1 0 20884 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_219
timestamp 1608761684
transform 1 0 21252 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1608761684
transform 1 0 19964 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1608761684
transform 1 0 19412 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1608761684
transform 1 0 18492 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_188
timestamp 1608761684
transform 1 0 18400 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_193
timestamp 1608761684
transform 1 0 18860 0 1 17808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_203
timestamp 1608761684
transform 1 0 19780 0 1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761684
transform 1 0 17112 0 1 17808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_180
timestamp 1608761684
transform 1 0 17664 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1608761684
transform 1 0 15180 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_150
timestamp 1608761684
transform 1 0 14904 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_154
timestamp 1608761684
transform 1 0 15272 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_166
timestamp 1608761684
transform 1 0 16376 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1608761684
transform 1 0 13892 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_131
timestamp 1608761684
transform 1 0 13156 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_142
timestamp 1608761684
transform 1 0 14168 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1608761684
transform 1 0 10856 0 1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1608761684
transform 1 0 12328 0 1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_29_105
timestamp 1608761684
transform 1 0 10764 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_115
timestamp 1608761684
transform 1 0 11684 0 1 17808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_121
timestamp 1608761684
transform 1 0 12236 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1608761684
transform 1 0 9568 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_89
timestamp 1608761684
transform 1 0 9292 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1608761684
transform 1 0 9660 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1608761684
transform 1 0 7728 0 1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_29_68
timestamp 1608761684
transform 1 0 7360 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_81
timestamp 1608761684
transform 1 0 8556 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1608761684
transform 1 0 5060 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761684
transform 1 0 5888 0 1 17808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_29_46
timestamp 1608761684
transform 1 0 5336 0 1 17808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1608761684
transform 1 0 3956 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_27
timestamp 1608761684
transform 1 0 3588 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_32
timestamp 1608761684
transform 1 0 4048 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_40
timestamp 1608761684
transform 1 0 4784 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1608761684
transform 1 0 2760 0 1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1608761684
transform 1 0 1104 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1608761684
transform 1 0 1380 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_15
timestamp 1608761684
transform 1 0 2484 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1608761684
transform 1 0 20516 0 -1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1608761684
transform -1 0 21620 0 -1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1608761684
transform 1 0 20884 0 -1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1608761684
transform 1 0 21252 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761684
transform 1 0 19412 0 -1 17808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_190
timestamp 1608761684
transform 1 0 18584 0 -1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_198
timestamp 1608761684
transform 1 0 19320 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_205
timestamp 1608761684
transform 1 0 19964 0 -1 17808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761684
transform 1 0 18032 0 -1 17808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1608761684
transform 1 0 17940 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_171
timestamp 1608761684
transform 1 0 16836 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_147
timestamp 1608761684
transform 1 0 14628 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_159
timestamp 1608761684
transform 1 0 15732 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_135
timestamp 1608761684
transform 1 0 13524 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1608761684
transform 1 0 12328 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_110
timestamp 1608761684
transform 1 0 11224 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_123
timestamp 1608761684
transform 1 0 12420 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_86
timestamp 1608761684
transform 1 0 9016 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_98
timestamp 1608761684
transform 1 0 10120 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_74
timestamp 1608761684
transform 1 0 7912 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1608761684
transform 1 0 6716 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_46
timestamp 1608761684
transform 1 0 5336 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_58
timestamp 1608761684
transform 1 0 6440 0 -1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_62
timestamp 1608761684
transform 1 0 6808 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1608761684
transform 1 0 3404 0 -1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_28_34
timestamp 1608761684
transform 1 0 4232 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761684
transform 1 0 1380 0 -1 17808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1608761684
transform 1 0 1104 0 -1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_19
timestamp 1608761684
transform 1 0 2852 0 -1 17808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1608761684
transform 1 0 20700 0 -1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608761684
transform -1 0 21620 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608761684
transform -1 0 21620 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1608761684
transform 1 0 20792 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_211
timestamp 1608761684
transform 1 0 20516 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_217
timestamp 1608761684
transform 1 0 21068 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_212
timestamp 1608761684
transform 1 0 20608 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_215
timestamp 1608761684
transform 1 0 20884 0 1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_219
timestamp 1608761684
transform 1 0 21252 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1608761684
transform 1 0 20240 0 1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761684
transform 1 0 19964 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_203
timestamp 1608761684
transform 1 0 19780 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_207
timestamp 1608761684
transform 1 0 20148 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761684
transform 1 0 19228 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761684
transform 1 0 19044 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_195
timestamp 1608761684
transform 1 0 19044 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_201
timestamp 1608761684
transform 1 0 19596 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1608761684
transform 1 0 18492 0 1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_188
timestamp 1608761684
transform 1 0 18400 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_193
timestamp 1608761684
transform 1 0 18860 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1608761684
transform 1 0 18032 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1608761684
transform 1 0 17940 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_172
timestamp 1608761684
transform 1 0 16928 0 -1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_180
timestamp 1608761684
transform 1 0 17664 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_187
timestamp 1608761684
transform 1 0 18308 0 -1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_182
timestamp 1608761684
transform 1 0 17848 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761684
transform 1 0 15456 0 -1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761684
transform 1 0 16376 0 1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1608761684
transform 1 0 15180 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_148
timestamp 1608761684
transform 1 0 14720 0 -1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_146
timestamp 1608761684
transform 1 0 14536 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_152
timestamp 1608761684
transform 1 0 15088 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_154
timestamp 1608761684
transform 1 0 15272 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1608761684
transform 1 0 13432 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1608761684
transform 1 0 13892 0 -1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_132
timestamp 1608761684
transform 1 0 13248 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_137
timestamp 1608761684
transform 1 0 13708 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_134
timestamp 1608761684
transform 1 0 13432 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1608761684
transform 1 0 11316 0 -1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1608761684
transform 1 0 12420 0 -1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1608761684
transform 1 0 12328 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_107
timestamp 1608761684
transform 1 0 10948 0 -1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_120
timestamp 1608761684
transform 1 0 12144 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_110
timestamp 1608761684
transform 1 0 11224 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_122
timestamp 1608761684
transform 1 0 12328 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1608761684
transform 1 0 9844 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1608761684
transform 1 0 10120 0 -1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1608761684
transform 1 0 9568 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_96
timestamp 1608761684
transform 1 0 9936 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_87
timestamp 1608761684
transform 1 0 9108 0 1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_91
timestamp 1608761684
transform 1 0 9476 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_93
timestamp 1608761684
transform 1 0 9660 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1608761684
transform 1 0 10120 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1608761684
transform 1 0 7820 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761684
transform 1 0 8464 0 -1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1608761684
transform 1 0 8280 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761684
transform 1 0 7268 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_71
timestamp 1608761684
transform 1 0 7636 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_76
timestamp 1608761684
transform 1 0 8096 0 -1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_64
timestamp 1608761684
transform 1 0 6992 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_73
timestamp 1608761684
transform 1 0 7820 0 1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_77
timestamp 1608761684
transform 1 0 8188 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1608761684
transform 1 0 6808 0 -1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1608761684
transform 1 0 6716 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_51
timestamp 1608761684
transform 1 0 5796 0 -1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_59
timestamp 1608761684
transform 1 0 6532 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_56
timestamp 1608761684
transform 1 0 6256 0 1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1608761684
transform 1 0 3128 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761684
transform 1 0 4784 0 1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761684
transform 1 0 4048 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1608761684
transform 1 0 3956 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_27
timestamp 1608761684
transform 1 0 3588 0 -1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_39
timestamp 1608761684
transform 1 0 4692 0 -1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_21
timestamp 1608761684
transform 1 0 3036 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_25
timestamp 1608761684
transform 1 0 3404 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_38
timestamp 1608761684
transform 1 0 4600 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608761684
transform 1 0 1104 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608761684
transform 1 0 1104 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1608761684
transform 1 0 1380 0 -1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1608761684
transform 1 0 2484 0 -1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1608761684
transform 1 0 1380 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_15
timestamp 1608761684
transform 1 0 2484 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608761684
transform -1 0 21620 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1608761684
transform 1 0 20792 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_212
timestamp 1608761684
transform 1 0 20608 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_215
timestamp 1608761684
transform 1 0 20884 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_219
timestamp 1608761684
transform 1 0 21252 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1608761684
transform 1 0 20240 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1608761684
transform 1 0 19688 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_198
timestamp 1608761684
transform 1 0 19320 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_206
timestamp 1608761684
transform 1 0 20056 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l2_in_0_
timestamp 1608761684
transform 1 0 17388 0 1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_175
timestamp 1608761684
transform 1 0 17204 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_186
timestamp 1608761684
transform 1 0 18216 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1608761684
transform 1 0 15272 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l1_in_0_
timestamp 1608761684
transform 1 0 16376 0 1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1608761684
transform 1 0 15180 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_148
timestamp 1608761684
transform 1 0 14720 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_152
timestamp 1608761684
transform 1 0 15088 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_157
timestamp 1608761684
transform 1 0 15548 0 1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_165
timestamp 1608761684
transform 1 0 16284 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761684
transform 1 0 13248 0 1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_130
timestamp 1608761684
transform 1 0 13064 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761684
transform 1 0 11592 0 1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_112
timestamp 1608761684
transform 1 0 11408 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761684
transform 1 0 9936 0 1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1608761684
transform 1 0 9568 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_85
timestamp 1608761684
transform 1 0 8924 0 1 15632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_91
timestamp 1608761684
transform 1 0 9476 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_93
timestamp 1608761684
transform 1 0 9660 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1608761684
transform 1 0 6992 0 1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_25_73
timestamp 1608761684
transform 1 0 7820 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761684
transform 1 0 4968 0 1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_25_58
timestamp 1608761684
transform 1 0 6440 0 1 15632
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1608761684
transform 1 0 3956 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_25
timestamp 1608761684
transform 1 0 3404 0 1 15632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_32
timestamp 1608761684
transform 1 0 4048 0 1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_40
timestamp 1608761684
transform 1 0 4784 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761684
transform 1 0 1932 0 1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608761684
transform 1 0 1104 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp 1608761684
transform 1 0 1380 0 1 15632
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1608761684
transform 1 0 20516 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608761684
transform -1 0 21620 0 -1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_209
timestamp 1608761684
transform 1 0 20332 0 -1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1608761684
transform 1 0 20884 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1608761684
transform 1 0 21252 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1608761684
transform 1 0 19964 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761684
transform 1 0 18952 0 -1 15632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_192
timestamp 1608761684
transform 1 0 18768 0 -1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_200
timestamp 1608761684
transform 1 0 19504 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_204
timestamp 1608761684
transform 1 0 19872 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1608761684
transform 1 0 17940 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_177
timestamp 1608761684
transform 1 0 17388 0 -1 15632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_184
timestamp 1608761684
transform 1 0 18032 0 -1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1608761684
transform 1 0 15180 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_165
timestamp 1608761684
transform 1 0 16284 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1608761684
transform 1 0 14352 0 -1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_24_135
timestamp 1608761684
transform 1 0 13524 0 -1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_143
timestamp 1608761684
transform 1 0 14260 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1608761684
transform 1 0 12328 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_110
timestamp 1608761684
transform 1 0 11224 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_123
timestamp 1608761684
transform 1 0 12420 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_86
timestamp 1608761684
transform 1 0 9016 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_98
timestamp 1608761684
transform 1 0 10120 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_74
timestamp 1608761684
transform 1 0 7912 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1608761684
transform 1 0 6716 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_45
timestamp 1608761684
transform 1 0 5244 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_57
timestamp 1608761684
transform 1 0 6348 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_62
timestamp 1608761684
transform 1 0 6808 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1608761684
transform 1 0 3312 0 -1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_22
timestamp 1608761684
transform 1 0 3128 0 -1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_33
timestamp 1608761684
transform 1 0 4140 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1608761684
transform 1 0 2300 0 -1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608761684
transform 1 0 1104 0 -1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1608761684
transform 1 0 1380 0 -1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_11
timestamp 1608761684
transform 1 0 2116 0 -1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608761684
transform -1 0 21620 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1608761684
transform 1 0 20792 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_213
timestamp 1608761684
transform 1 0 20700 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_215
timestamp 1608761684
transform 1 0 20884 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_219
timestamp 1608761684
transform 1 0 21252 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761684
transform 1 0 18860 0 1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761684
transform 1 0 19596 0 1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_191
timestamp 1608761684
transform 1 0 18676 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_199
timestamp 1608761684
transform 1 0 19412 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_207
timestamp 1608761684
transform 1 0 20148 0 1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1608761684
transform 1 0 17112 0 1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_172
timestamp 1608761684
transform 1 0 16928 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_183
timestamp 1608761684
transform 1 0 17940 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761684
transform 1 0 15456 0 1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1608761684
transform 1 0 15180 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_146
timestamp 1608761684
transform 1 0 14536 0 1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_152
timestamp 1608761684
transform 1 0 15088 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_154
timestamp 1608761684
transform 1 0 15272 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_right_track_0.prog_clk
timestamp 1608761684
transform 1 0 13156 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_128
timestamp 1608761684
transform 1 0 12880 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_134
timestamp 1608761684
transform 1 0 13432 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_108
timestamp 1608761684
transform 1 0 11040 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_120
timestamp 1608761684
transform 1 0 12144 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1608761684
transform 1 0 9660 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1608761684
transform 1 0 9568 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_90
timestamp 1608761684
transform 1 0 9384 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_96
timestamp 1608761684
transform 1 0 9936 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1608761684
transform 1 0 7820 0 1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_23_65
timestamp 1608761684
transform 1 0 7084 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_82
timestamp 1608761684
transform 1 0 8648 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761684
transform 1 0 4968 0 1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_right_track_0.prog_clk
timestamp 1608761684
transform 1 0 6808 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_58
timestamp 1608761684
transform 1 0 6440 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1608761684
transform 1 0 3312 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1608761684
transform 1 0 3956 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_27
timestamp 1608761684
transform 1 0 3588 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_32
timestamp 1608761684
transform 1 0 4048 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_40
timestamp 1608761684
transform 1 0 4784 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761684
transform 1 0 1472 0 1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608761684
transform 1 0 1104 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_3
timestamp 1608761684
transform 1 0 1380 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_20
timestamp 1608761684
transform 1 0 2944 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1608761684
transform 1 0 20516 0 -1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608761684
transform -1 0 21620 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_209
timestamp 1608761684
transform 1 0 20332 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1608761684
transform 1 0 20884 0 -1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1608761684
transform 1 0 21252 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761684
transform 1 0 19044 0 -1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761684
transform 1 0 19780 0 -1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_22_192
timestamp 1608761684
transform 1 0 18768 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_201
timestamp 1608761684
transform 1 0 19596 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1608761684
transform 1 0 16744 0 -1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1608761684
transform 1 0 17940 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_168
timestamp 1608761684
transform 1 0 16560 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_179
timestamp 1608761684
transform 1 0 17572 0 -1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_184
timestamp 1608761684
transform 1 0 18032 0 -1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761684
transform 1 0 15088 0 -1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_150
timestamp 1608761684
transform 1 0 14904 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761684
transform 1 0 13432 0 -1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_132
timestamp 1608761684
transform 1 0 13248 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1608761684
transform 1 0 12420 0 -1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1608761684
transform 1 0 12328 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_115
timestamp 1608761684
transform 1 0 11684 0 -1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_121
timestamp 1608761684
transform 1 0 12236 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1608761684
transform 1 0 9752 0 -1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_92
timestamp 1608761684
transform 1 0 9568 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_103
timestamp 1608761684
transform 1 0 10580 0 -1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761684
transform 1 0 8096 0 -1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_74
timestamp 1608761684
transform 1 0 7912 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1608761684
transform 1 0 5152 0 -1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1608761684
transform 1 0 6716 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_42
timestamp 1608761684
transform 1 0 4968 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_53
timestamp 1608761684
transform 1 0 5980 0 -1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_62
timestamp 1608761684
transform 1 0 6808 0 -1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761684
transform 1 0 3496 0 -1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_22_23
timestamp 1608761684
transform 1 0 3220 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608761684
transform 1 0 1104 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1608761684
transform 1 0 1380 0 -1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_15
timestamp 1608761684
transform 1 0 2484 0 -1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608761684
transform -1 0 21620 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1608761684
transform 1 0 20792 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_212
timestamp 1608761684
transform 1 0 20608 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_215
timestamp 1608761684
transform 1 0 20884 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_219
timestamp 1608761684
transform 1 0 21252 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1608761684
transform 1 0 20240 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_191
timestamp 1608761684
transform 1 0 18676 0 1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_203
timestamp 1608761684
transform 1 0 19780 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_207
timestamp 1608761684
transform 1 0 20148 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1608761684
transform 1 0 17664 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1608761684
transform 1 0 18308 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1608761684
transform 1 0 16652 0 1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_178
timestamp 1608761684
transform 1 0 17480 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_183
timestamp 1608761684
transform 1 0 17940 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1608761684
transform 1 0 15180 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_148
timestamp 1608761684
transform 1 0 14720 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_152
timestamp 1608761684
transform 1 0 15088 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_154
timestamp 1608761684
transform 1 0 15272 0 1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_166
timestamp 1608761684
transform 1 0 16376 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1608761684
transform 1 0 13340 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_131
timestamp 1608761684
transform 1 0 13156 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_136
timestamp 1608761684
transform 1 0 13616 0 1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1608761684
transform 1 0 12328 0 1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_120
timestamp 1608761684
transform 1 0 12144 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761684
transform 1 0 10672 0 1 13456
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1608761684
transform 1 0 9568 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_right_track_0.prog_clk
timestamp 1608761684
transform 1 0 8924 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_88
timestamp 1608761684
transform 1 0 9200 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_93
timestamp 1608761684
transform 1 0 9660 0 1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_101
timestamp 1608761684
transform 1 0 10396 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761684
transform 1 0 7268 0 1 13456
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_65
timestamp 1608761684
transform 1 0 7084 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_83
timestamp 1608761684
transform 1 0 8740 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761684
transform 1 0 5612 0 1 13456
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_47
timestamp 1608761684
transform 1 0 5428 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1608761684
transform 1 0 4600 0 1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1608761684
transform 1 0 3956 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_26
timestamp 1608761684
transform 1 0 3496 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_30
timestamp 1608761684
transform 1 0 3864 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_32
timestamp 1608761684
transform 1 0 4048 0 1 13456
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761684
transform 1 0 2024 0 1 13456
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608761684
transform 1 0 1104 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_3
timestamp 1608761684
transform 1 0 1380 0 1 13456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_9
timestamp 1608761684
transform 1 0 1932 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608761684
transform -1 0 21620 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608761684
transform -1 0 21620 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_219
timestamp 1608761684
transform 1 0 21252 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1608761684
transform 1 0 21252 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1608761684
transform 1 0 20792 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_215
timestamp 1608761684
transform 1 0 20884 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1608761684
transform 1 0 20884 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1608761684
transform 1 0 20516 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_211
timestamp 1608761684
transform 1 0 20516 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_209
timestamp 1608761684
transform 1 0 20332 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1608761684
transform 1 0 20148 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1608761684
transform 1 0 19964 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1608761684
transform 1 0 19596 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761684
transform 1 0 18584 0 -1 13456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_197
timestamp 1608761684
transform 1 0 19228 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_205
timestamp 1608761684
transform 1 0 19964 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_196
timestamp 1608761684
transform 1 0 19136 0 -1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_204
timestamp 1608761684
transform 1 0 19872 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761684
transform 1 0 16652 0 1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1608761684
transform 1 0 17940 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_168
timestamp 1608761684
transform 1 0 16560 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_185
timestamp 1608761684
transform 1 0 18124 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_168
timestamp 1608761684
transform 1 0 16560 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_180
timestamp 1608761684
transform 1 0 17664 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_184
timestamp 1608761684
transform 1 0 18032 0 -1 13456
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761684
transform 1 0 15272 0 1 12368
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1608761684
transform 1 0 15180 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_150
timestamp 1608761684
transform 1 0 14904 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_160
timestamp 1608761684
transform 1 0 15824 0 1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_156
timestamp 1608761684
transform 1 0 15456 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1608761684
transform 1 0 13340 0 1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_19_126
timestamp 1608761684
transform 1 0 12696 0 1 12368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_132
timestamp 1608761684
transform 1 0 13248 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_142
timestamp 1608761684
transform 1 0 14168 0 1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_132
timestamp 1608761684
transform 1 0 13248 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_144
timestamp 1608761684
transform 1 0 14352 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761684
transform 1 0 11132 0 1 12368
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1608761684
transform 1 0 12420 0 -1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1608761684
transform 1 0 12328 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_right_track_0.prog_clk
timestamp 1608761684
transform 1 0 12420 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_115
timestamp 1608761684
transform 1 0 11684 0 1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_116
timestamp 1608761684
transform 1 0 11776 0 -1 13456
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761684
transform 1 0 9660 0 1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1608761684
transform 1 0 9568 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_right_track_0.prog_clk
timestamp 1608761684
transform 1 0 9936 0 -1 13456
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_20_86
timestamp 1608761684
transform 1 0 9016 0 -1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_94
timestamp 1608761684
transform 1 0 9752 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_68
timestamp 1608761684
transform 1 0 7360 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_80
timestamp 1608761684
transform 1 0 8464 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_74
timestamp 1608761684
transform 1 0 7912 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1608761684
transform 1 0 4968 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1608761684
transform 1 0 6716 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_44
timestamp 1608761684
transform 1 0 5152 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_56
timestamp 1608761684
transform 1 0 6256 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_45
timestamp 1608761684
transform 1 0 5244 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_57
timestamp 1608761684
transform 1 0 6348 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_62
timestamp 1608761684
transform 1 0 6808 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1608761684
transform 1 0 3956 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_27
timestamp 1608761684
transform 1 0 3588 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_32
timestamp 1608761684
transform 1 0 4048 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_27
timestamp 1608761684
transform 1 0 3588 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_39
timestamp 1608761684
transform 1 0 4692 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608761684
transform 1 0 1104 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608761684
transform 1 0 1104 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1608761684
transform 1 0 1380 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1608761684
transform 1 0 2484 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1608761684
transform 1 0 1380 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1608761684
transform 1 0 2484 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1608761684
transform 1 0 20516 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608761684
transform -1 0 21620 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_209
timestamp 1608761684
transform 1 0 20332 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1608761684
transform 1 0 20884 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1608761684
transform 1 0 21252 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1608761684
transform 1 0 19964 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761684
transform 1 0 19228 0 -1 12368
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_193
timestamp 1608761684
transform 1 0 18860 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_203
timestamp 1608761684
transform 1 0 19780 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1608761684
transform 1 0 18032 0 -1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1608761684
transform 1 0 17940 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_168
timestamp 1608761684
transform 1 0 16560 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_180
timestamp 1608761684
transform 1 0 17664 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761684
transform 1 0 15088 0 -1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_18_149
timestamp 1608761684
transform 1 0 14812 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1608761684
transform 1 0 12696 0 -1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1608761684
transform 1 0 13984 0 -1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_right_track_0.prog_clk
timestamp 1608761684
transform 1 0 13708 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_135
timestamp 1608761684
transform 1 0 13524 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1608761684
transform 1 0 12328 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1608761684
transform 1 0 10764 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_117
timestamp 1608761684
transform 1 0 11868 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_121
timestamp 1608761684
transform 1 0 12236 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_123
timestamp 1608761684
transform 1 0 12420 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1608761684
transform 1 0 9936 0 -1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_94
timestamp 1608761684
transform 1 0 9752 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761684
transform 1 0 8280 0 -1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_right_track_0.prog_clk
timestamp 1608761684
transform 1 0 7820 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_71
timestamp 1608761684
transform 1 0 7636 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_76
timestamp 1608761684
transform 1 0 8096 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1608761684
transform 1 0 6808 0 -1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1608761684
transform 1 0 6716 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_51
timestamp 1608761684
transform 1 0 5796 0 -1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_59
timestamp 1608761684
transform 1 0 6532 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_27
timestamp 1608761684
transform 1 0 3588 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_39
timestamp 1608761684
transform 1 0 4692 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608761684
transform 1 0 1104 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1608761684
transform 1 0 1380 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1608761684
transform 1 0 2484 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608761684
transform -1 0 21620 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1608761684
transform 1 0 20792 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_212
timestamp 1608761684
transform 1 0 20608 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_215
timestamp 1608761684
transform 1 0 20884 0 1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_219
timestamp 1608761684
transform 1 0 21252 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1608761684
transform 1 0 19044 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1608761684
transform 1 0 20240 0 1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_193
timestamp 1608761684
transform 1 0 18860 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_198
timestamp 1608761684
transform 1 0 19320 0 1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_206
timestamp 1608761684
transform 1 0 20056 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1608761684
transform 1 0 18032 0 1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_17_178
timestamp 1608761684
transform 1 0 17480 0 1 11280
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1608761684
transform 1 0 15180 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_154
timestamp 1608761684
transform 1 0 15272 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_166
timestamp 1608761684
transform 1 0 16376 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1608761684
transform 1 0 13616 0 1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_134
timestamp 1608761684
transform 1 0 13432 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_145
timestamp 1608761684
transform 1 0 14444 0 1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1608761684
transform 1 0 11316 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761684
transform 1 0 11960 0 1 11280
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_109
timestamp 1608761684
transform 1 0 11132 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_114
timestamp 1608761684
transform 1 0 11592 0 1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1608761684
transform 1 0 10304 0 1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608761684
transform 1 0 9568 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_85
timestamp 1608761684
transform 1 0 8924 0 1 11280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_91
timestamp 1608761684
transform 1 0 9476 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_93
timestamp 1608761684
transform 1 0 9660 0 1 11280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_99
timestamp 1608761684
transform 1 0 10212 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1608761684
transform 1 0 8096 0 1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_74
timestamp 1608761684
transform 1 0 7912 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761684
transform 1 0 6440 0 1 11280
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_17_44
timestamp 1608761684
transform 1 0 5152 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_56
timestamp 1608761684
transform 1 0 6256 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608761684
transform 1 0 3956 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_27
timestamp 1608761684
transform 1 0 3588 0 1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_32
timestamp 1608761684
transform 1 0 4048 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608761684
transform 1 0 1104 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1608761684
transform 1 0 1380 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1608761684
transform 1 0 2484 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1608761684
transform 1 0 20516 0 -1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608761684
transform -1 0 21620 0 -1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_209
timestamp 1608761684
transform 1 0 20332 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1608761684
transform 1 0 20884 0 -1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1608761684
transform 1 0 21252 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1608761684
transform 1 0 19964 0 -1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1608761684
transform 1 0 18860 0 -1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_192
timestamp 1608761684
transform 1 0 18768 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_202
timestamp 1608761684
transform 1 0 19688 0 -1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1608761684
transform 1 0 16928 0 -1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608761684
transform 1 0 17940 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_170
timestamp 1608761684
transform 1 0 16744 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_181
timestamp 1608761684
transform 1 0 17756 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_184
timestamp 1608761684
transform 1 0 18032 0 -1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1608761684
transform 1 0 14628 0 -1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1608761684
transform 1 0 15916 0 -1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_150
timestamp 1608761684
transform 1 0 14904 0 -1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_158
timestamp 1608761684
transform 1 0 15640 0 -1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1608761684
transform 1 0 13616 0 -1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_135
timestamp 1608761684
transform 1 0 13524 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_145
timestamp 1608761684
transform 1 0 14444 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608761684
transform 1 0 12328 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1608761684
transform 1 0 10764 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_117
timestamp 1608761684
transform 1 0 11868 0 -1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_121
timestamp 1608761684
transform 1 0 12236 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_123
timestamp 1608761684
transform 1 0 12420 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1608761684
transform 1 0 9660 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1608761684
transform 1 0 7728 0 -1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_70
timestamp 1608761684
transform 1 0 7544 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_81
timestamp 1608761684
transform 1 0 8556 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608761684
transform 1 0 6716 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_51
timestamp 1608761684
transform 1 0 5796 0 -1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_59
timestamp 1608761684
transform 1 0 6532 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_62
timestamp 1608761684
transform 1 0 6808 0 -1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_27
timestamp 1608761684
transform 1 0 3588 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_39
timestamp 1608761684
transform 1 0 4692 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608761684
transform 1 0 1104 0 -1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1608761684
transform 1 0 1380 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1608761684
transform 1 0 2484 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608761684
transform -1 0 21620 0 1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608761684
transform 1 0 20792 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_212
timestamp 1608761684
transform 1 0 20608 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_215
timestamp 1608761684
transform 1 0 20884 0 1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_219
timestamp 1608761684
transform 1 0 21252 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1608761684
transform 1 0 20240 0 1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_188
timestamp 1608761684
transform 1 0 18400 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_200
timestamp 1608761684
transform 1 0 19504 0 1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1608761684
transform 1 0 16468 0 1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_15_176
timestamp 1608761684
transform 1 0 17296 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608761684
transform 1 0 15180 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_150
timestamp 1608761684
transform 1 0 14904 0 1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_154
timestamp 1608761684
transform 1 0 15272 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_166
timestamp 1608761684
transform 1 0 16376 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_126
timestamp 1608761684
transform 1 0 12696 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_138
timestamp 1608761684
transform 1 0 13800 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761684
transform 1 0 11040 0 1 10192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_106
timestamp 1608761684
transform 1 0 10856 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_114
timestamp 1608761684
transform 1 0 11592 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1608761684
transform 1 0 10028 0 1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608761684
transform 1 0 9568 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_90
timestamp 1608761684
transform 1 0 9384 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_93
timestamp 1608761684
transform 1 0 9660 0 1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761684
transform 1 0 7176 0 1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_64
timestamp 1608761684
transform 1 0 6992 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_82
timestamp 1608761684
transform 1 0 8648 0 1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_44
timestamp 1608761684
transform 1 0 5152 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_56
timestamp 1608761684
transform 1 0 6256 0 1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608761684
transform 1 0 3956 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1608761684
transform 1 0 3588 0 1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_32
timestamp 1608761684
transform 1 0 4048 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608761684
transform 1 0 1104 0 1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1608761684
transform 1 0 1380 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1608761684
transform 1 0 2484 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1608761684
transform 1 0 20516 0 -1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608761684
transform -1 0 21620 0 1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608761684
transform -1 0 21620 0 -1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608761684
transform 1 0 20792 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_212
timestamp 1608761684
transform 1 0 20608 0 1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_215
timestamp 1608761684
transform 1 0 20884 0 1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_219
timestamp 1608761684
transform 1 0 21252 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1608761684
transform 1 0 20884 0 -1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1608761684
transform 1 0 21252 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1608761684
transform 1 0 19596 0 1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761684
transform 1 0 18492 0 -1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1608761684
transform 1 0 18584 0 1 9104
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_188
timestamp 1608761684
transform 1 0 18400 0 1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_199
timestamp 1608761684
transform 1 0 19412 0 1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_204
timestamp 1608761684
transform 1 0 19872 0 1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_188
timestamp 1608761684
transform 1 0 18400 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_205
timestamp 1608761684
transform 1 0 19964 0 -1 10192
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1608761684
transform 1 0 17572 0 1 9104
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608761684
transform 1 0 17940 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_178
timestamp 1608761684
transform 1 0 17480 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_177
timestamp 1608761684
transform 1 0 17388 0 -1 10192
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_184
timestamp 1608761684
transform 1 0 18032 0 -1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761684
transform 1 0 15916 0 -1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608761684
transform 1 0 15180 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_151
timestamp 1608761684
transform 1 0 14996 0 1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_154
timestamp 1608761684
transform 1 0 15272 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_166
timestamp 1608761684
transform 1 0 16376 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_155
timestamp 1608761684
transform 1 0 15364 0 -1 10192
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761684
transform 1 0 12788 0 -1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761684
transform 1 0 13524 0 1 9104
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_13_128
timestamp 1608761684
transform 1 0 12880 0 1 9104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_134
timestamp 1608761684
transform 1 0 13432 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_143
timestamp 1608761684
transform 1 0 14260 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1608761684
transform 1 0 10948 0 1 9104
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1608761684
transform 1 0 10856 0 -1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1608761684
transform 1 0 12052 0 1 9104
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608761684
transform 1 0 12328 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_105
timestamp 1608761684
transform 1 0 10764 0 1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_116
timestamp 1608761684
transform 1 0 11776 0 1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_115
timestamp 1608761684
transform 1 0 11684 0 -1 10192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_121
timestamp 1608761684
transform 1 0 12236 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_123
timestamp 1608761684
transform 1 0 12420 0 -1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1608761684
transform 1 0 9936 0 1 9104
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608761684
transform 1 0 9568 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_86
timestamp 1608761684
transform 1 0 9016 0 1 9104
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_13_93
timestamp 1608761684
transform 1 0 9660 0 1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_96
timestamp 1608761684
transform 1 0 9936 0 -1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_104
timestamp 1608761684
transform 1 0 10672 0 -1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761684
transform 1 0 7544 0 1 9104
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761684
transform 1 0 8464 0 -1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_13_68
timestamp 1608761684
transform 1 0 7360 0 1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_74
timestamp 1608761684
transform 1 0 7912 0 -1 10192
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608761684
transform 1 0 6716 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_44
timestamp 1608761684
transform 1 0 5152 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_56
timestamp 1608761684
transform 1 0 6256 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_51
timestamp 1608761684
transform 1 0 5796 0 -1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_59
timestamp 1608761684
transform 1 0 6532 0 -1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_62
timestamp 1608761684
transform 1 0 6808 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608761684
transform 1 0 3956 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_27
timestamp 1608761684
transform 1 0 3588 0 1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_32
timestamp 1608761684
transform 1 0 4048 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_27
timestamp 1608761684
transform 1 0 3588 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_39
timestamp 1608761684
transform 1 0 4692 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608761684
transform 1 0 1104 0 1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608761684
transform 1 0 1104 0 -1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1608761684
transform 1 0 1380 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1608761684
transform 1 0 2484 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1608761684
transform 1 0 1380 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1608761684
transform 1 0 2484 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1608761684
transform 1 0 20516 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608761684
transform -1 0 21620 0 -1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_209
timestamp 1608761684
transform 1 0 20332 0 -1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1608761684
transform 1 0 20884 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1608761684
transform 1 0 21252 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1608761684
transform 1 0 19964 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_201
timestamp 1608761684
transform 1 0 19596 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761684
transform 1 0 18124 0 -1 9104
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608761684
transform 1 0 17940 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_168
timestamp 1608761684
transform 1 0 16560 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_180
timestamp 1608761684
transform 1 0 17664 0 -1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_184
timestamp 1608761684
transform 1 0 18032 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1608761684
transform 1 0 15088 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_147
timestamp 1608761684
transform 1 0 14628 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_151
timestamp 1608761684
transform 1 0 14996 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_156
timestamp 1608761684
transform 1 0 15456 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1608761684
transform 1 0 13156 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_135
timestamp 1608761684
transform 1 0 13524 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1608761684
transform 1 0 11592 0 -1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608761684
transform 1 0 12328 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_112
timestamp 1608761684
transform 1 0 11408 0 -1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_117
timestamp 1608761684
transform 1 0 11868 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_121
timestamp 1608761684
transform 1 0 12236 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_123
timestamp 1608761684
transform 1 0 12420 0 -1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1608761684
transform 1 0 10580 0 -1 9104
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_86
timestamp 1608761684
transform 1 0 9016 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_98
timestamp 1608761684
transform 1 0 10120 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_102
timestamp 1608761684
transform 1 0 10488 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_74
timestamp 1608761684
transform 1 0 7912 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608761684
transform 1 0 6716 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_51
timestamp 1608761684
transform 1 0 5796 0 -1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_59
timestamp 1608761684
transform 1 0 6532 0 -1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_62
timestamp 1608761684
transform 1 0 6808 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_27
timestamp 1608761684
transform 1 0 3588 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_39
timestamp 1608761684
transform 1 0 4692 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608761684
transform 1 0 1104 0 -1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1608761684
transform 1 0 1380 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1608761684
transform 1 0 2484 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608761684
transform -1 0 21620 0 1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608761684
transform 1 0 20792 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_212
timestamp 1608761684
transform 1 0 20608 0 1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_215
timestamp 1608761684
transform 1 0 20884 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_219
timestamp 1608761684
transform 1 0 21252 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1608761684
transform 1 0 20240 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_190
timestamp 1608761684
transform 1 0 18584 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_202
timestamp 1608761684
transform 1 0 19688 0 1 8016
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1608761684
transform 1 0 17204 0 1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_173
timestamp 1608761684
transform 1 0 17020 0 1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_178
timestamp 1608761684
transform 1 0 17480 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1608761684
transform 1 0 16192 0 1 8016
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761684
transform 1 0 15456 0 1 8016
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608761684
transform 1 0 15180 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_150
timestamp 1608761684
transform 1 0 14904 0 1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_154
timestamp 1608761684
transform 1 0 15272 0 1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_162
timestamp 1608761684
transform 1 0 16008 0 1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761684
transform 1 0 13248 0 1 8016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_127
timestamp 1608761684
transform 1 0 12788 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_131
timestamp 1608761684
transform 1 0 13156 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_138
timestamp 1608761684
transform 1 0 13800 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1608761684
transform 1 0 11316 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1608761684
transform 1 0 10764 0 1 8016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_115
timestamp 1608761684
transform 1 0 11684 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608761684
transform 1 0 9568 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1608761684
transform 1 0 9660 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_68
timestamp 1608761684
transform 1 0 7360 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_80
timestamp 1608761684
transform 1 0 8464 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_44
timestamp 1608761684
transform 1 0 5152 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_56
timestamp 1608761684
transform 1 0 6256 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608761684
transform 1 0 3956 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1608761684
transform 1 0 3588 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_32
timestamp 1608761684
transform 1 0 4048 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608761684
transform 1 0 1104 0 1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1608761684
transform 1 0 1380 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1608761684
transform 1 0 2484 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1608761684
transform 1 0 20516 0 -1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608761684
transform -1 0 21620 0 -1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_209
timestamp 1608761684
transform 1 0 20332 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1608761684
transform 1 0 20884 0 -1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1608761684
transform 1 0 21252 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1608761684
transform 1 0 19964 0 -1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_200
timestamp 1608761684
transform 1 0 19504 0 -1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_204
timestamp 1608761684
transform 1 0 19872 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761684
transform 1 0 18032 0 -1 8016
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608761684
transform 1 0 17940 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_178
timestamp 1608761684
transform 1 0 17480 0 -1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_182
timestamp 1608761684
transform 1 0 17848 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761684
transform 1 0 16008 0 -1 8016
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_157
timestamp 1608761684
transform 1 0 15548 0 -1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_161
timestamp 1608761684
transform 1 0 15916 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1608761684
transform 1 0 13616 0 -1 8016
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_135
timestamp 1608761684
transform 1 0 13524 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_145
timestamp 1608761684
transform 1 0 14444 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608761684
transform 1 0 12328 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1608761684
transform 1 0 11132 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_121
timestamp 1608761684
transform 1 0 12236 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_123
timestamp 1608761684
transform 1 0 12420 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761684
transform 1 0 10580 0 -1 8016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_86
timestamp 1608761684
transform 1 0 9016 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_98
timestamp 1608761684
transform 1 0 10120 0 -1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_102
timestamp 1608761684
transform 1 0 10488 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_74
timestamp 1608761684
transform 1 0 7912 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608761684
transform 1 0 6716 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_51
timestamp 1608761684
transform 1 0 5796 0 -1 8016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_59
timestamp 1608761684
transform 1 0 6532 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_62
timestamp 1608761684
transform 1 0 6808 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_27
timestamp 1608761684
transform 1 0 3588 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_39
timestamp 1608761684
transform 1 0 4692 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608761684
transform 1 0 1104 0 -1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1608761684
transform 1 0 1380 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1608761684
transform 1 0 2484 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608761684
transform -1 0 21620 0 1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608761684
transform 1 0 20792 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_215
timestamp 1608761684
transform 1 0 20884 0 1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_219
timestamp 1608761684
transform 1 0 21252 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_194
timestamp 1608761684
transform 1 0 18952 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_206
timestamp 1608761684
transform 1 0 20056 0 1 6928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_170
timestamp 1608761684
transform 1 0 16744 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_182
timestamp 1608761684
transform 1 0 17848 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1608761684
transform 1 0 14628 0 1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761684
transform 1 0 15272 0 1 6928
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608761684
transform 1 0 15180 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_150
timestamp 1608761684
transform 1 0 14904 0 1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761684
transform 1 0 12972 0 1 6928
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_127
timestamp 1608761684
transform 1 0 12788 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_145
timestamp 1608761684
transform 1 0 14444 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761684
transform 1 0 11316 0 1 6928
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_109
timestamp 1608761684
transform 1 0 11132 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1608761684
transform 1 0 9844 0 1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1608761684
transform 1 0 10304 0 1 6928
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608761684
transform 1 0 9568 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_93
timestamp 1608761684
transform 1 0 9660 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_98
timestamp 1608761684
transform 1 0 10120 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_68
timestamp 1608761684
transform 1 0 7360 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_80
timestamp 1608761684
transform 1 0 8464 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_44
timestamp 1608761684
transform 1 0 5152 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_56
timestamp 1608761684
transform 1 0 6256 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608761684
transform 1 0 3956 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_27
timestamp 1608761684
transform 1 0 3588 0 1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_32
timestamp 1608761684
transform 1 0 4048 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608761684
transform 1 0 1104 0 1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1608761684
transform 1 0 1380 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1608761684
transform 1 0 2484 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1608761684
transform 1 0 20516 0 -1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608761684
transform -1 0 21620 0 -1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1608761684
transform 1 0 20884 0 -1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1608761684
transform 1 0 21252 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_196
timestamp 1608761684
transform 1 0 19136 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_208
timestamp 1608761684
transform 1 0 20240 0 -1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1608761684
transform 1 0 16652 0 -1 6928
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608761684
transform 1 0 17940 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_178
timestamp 1608761684
transform 1 0 17480 0 -1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_182
timestamp 1608761684
transform 1 0 17848 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_184
timestamp 1608761684
transform 1 0 18032 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_149
timestamp 1608761684
transform 1 0 14812 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_161
timestamp 1608761684
transform 1 0 15916 0 -1 6928
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1608761684
transform 1 0 13984 0 -1 6928
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_135
timestamp 1608761684
transform 1 0 13524 0 -1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1608761684
transform 1 0 13892 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1608761684
transform 1 0 10856 0 -1 6928
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608761684
transform 1 0 12328 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_115
timestamp 1608761684
transform 1 0 11684 0 -1 6928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_121
timestamp 1608761684
transform 1 0 12236 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_123
timestamp 1608761684
transform 1 0 12420 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761684
transform 1 0 9200 0 -1 6928
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_87
timestamp 1608761684
transform 1 0 9108 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_104
timestamp 1608761684
transform 1 0 10672 0 -1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761684
transform 1 0 7268 0 -1 6928
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_66
timestamp 1608761684
transform 1 0 7176 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_83
timestamp 1608761684
transform 1 0 8740 0 -1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608761684
transform 1 0 6716 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_51
timestamp 1608761684
transform 1 0 5796 0 -1 6928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_59
timestamp 1608761684
transform 1 0 6532 0 -1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_62
timestamp 1608761684
transform 1 0 6808 0 -1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_27
timestamp 1608761684
transform 1 0 3588 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_39
timestamp 1608761684
transform 1 0 4692 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608761684
transform 1 0 1104 0 -1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1608761684
transform 1 0 1380 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1608761684
transform 1 0 2484 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1608761684
transform 1 0 20516 0 -1 5840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608761684
transform -1 0 21620 0 -1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608761684
transform -1 0 21620 0 1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608761684
transform 1 0 20792 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1608761684
transform 1 0 20884 0 -1 5840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1608761684
transform 1 0 21252 0 -1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_215
timestamp 1608761684
transform 1 0 20884 0 1 5840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_219
timestamp 1608761684
transform 1 0 21252 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_196
timestamp 1608761684
transform 1 0 19136 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_208
timestamp 1608761684
transform 1 0 20240 0 -1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_190
timestamp 1608761684
transform 1 0 18584 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_202
timestamp 1608761684
transform 1 0 19688 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608761684
transform 1 0 17940 0 -1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_171
timestamp 1608761684
transform 1 0 16836 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_184
timestamp 1608761684
transform 1 0 18032 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_178
timestamp 1608761684
transform 1 0 17480 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608761684
transform 1 0 15180 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_147
timestamp 1608761684
transform 1 0 14628 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_159
timestamp 1608761684
transform 1 0 15732 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_154
timestamp 1608761684
transform 1 0 15272 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_166
timestamp 1608761684
transform 1 0 16376 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_135
timestamp 1608761684
transform 1 0 13524 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_129
timestamp 1608761684
transform 1 0 12972 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_141
timestamp 1608761684
transform 1 0 14076 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608761684
transform 1 0 12328 0 -1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_110
timestamp 1608761684
transform 1 0 11224 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_123
timestamp 1608761684
transform 1 0 12420 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_105
timestamp 1608761684
transform 1 0 10764 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_117
timestamp 1608761684
transform 1 0 11868 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608761684
transform 1 0 9568 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_86
timestamp 1608761684
transform 1 0 9016 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_98
timestamp 1608761684
transform 1 0 10120 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1608761684
transform 1 0 9660 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_74
timestamp 1608761684
transform 1 0 7912 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_68
timestamp 1608761684
transform 1 0 7360 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_80
timestamp 1608761684
transform 1 0 8464 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608761684
transform 1 0 6716 0 -1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_51
timestamp 1608761684
transform 1 0 5796 0 -1 5840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_59
timestamp 1608761684
transform 1 0 6532 0 -1 5840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_62
timestamp 1608761684
transform 1 0 6808 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_44
timestamp 1608761684
transform 1 0 5152 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_56
timestamp 1608761684
transform 1 0 6256 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608761684
transform 1 0 3956 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_27
timestamp 1608761684
transform 1 0 3588 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_39
timestamp 1608761684
transform 1 0 4692 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1608761684
transform 1 0 3588 0 1 5840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_32
timestamp 1608761684
transform 1 0 4048 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608761684
transform 1 0 1104 0 -1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608761684
transform 1 0 1104 0 1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1608761684
transform 1 0 1380 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1608761684
transform 1 0 2484 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1608761684
transform 1 0 1380 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1608761684
transform 1 0 2484 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608761684
transform -1 0 21620 0 1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608761684
transform 1 0 20792 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_215
timestamp 1608761684
transform 1 0 20884 0 1 4752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_219
timestamp 1608761684
transform 1 0 21252 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_190
timestamp 1608761684
transform 1 0 18584 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_202
timestamp 1608761684
transform 1 0 19688 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_178
timestamp 1608761684
transform 1 0 17480 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608761684
transform 1 0 15180 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_154
timestamp 1608761684
transform 1 0 15272 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_166
timestamp 1608761684
transform 1 0 16376 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_129
timestamp 1608761684
transform 1 0 12972 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_141
timestamp 1608761684
transform 1 0 14076 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_105
timestamp 1608761684
transform 1 0 10764 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_117
timestamp 1608761684
transform 1 0 11868 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608761684
transform 1 0 9568 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1608761684
transform 1 0 9660 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_68
timestamp 1608761684
transform 1 0 7360 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_80
timestamp 1608761684
transform 1 0 8464 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_44
timestamp 1608761684
transform 1 0 5152 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_56
timestamp 1608761684
transform 1 0 6256 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608761684
transform 1 0 3956 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1608761684
transform 1 0 3588 0 1 4752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_32
timestamp 1608761684
transform 1 0 4048 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608761684
transform 1 0 1104 0 1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1608761684
transform 1 0 1380 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1608761684
transform 1 0 2484 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _87_
timestamp 1608761684
transform 1 0 20516 0 -1 4752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608761684
transform -1 0 21620 0 -1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1608761684
transform 1 0 20884 0 -1 4752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1608761684
transform 1 0 21252 0 -1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_196
timestamp 1608761684
transform 1 0 19136 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_208
timestamp 1608761684
transform 1 0 20240 0 -1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608761684
transform 1 0 17940 0 -1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_171
timestamp 1608761684
transform 1 0 16836 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_184
timestamp 1608761684
transform 1 0 18032 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_147
timestamp 1608761684
transform 1 0 14628 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_159
timestamp 1608761684
transform 1 0 15732 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_135
timestamp 1608761684
transform 1 0 13524 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608761684
transform 1 0 12328 0 -1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_110
timestamp 1608761684
transform 1 0 11224 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_123
timestamp 1608761684
transform 1 0 12420 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_86
timestamp 1608761684
transform 1 0 9016 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_98
timestamp 1608761684
transform 1 0 10120 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_74
timestamp 1608761684
transform 1 0 7912 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608761684
transform 1 0 6716 0 -1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_51
timestamp 1608761684
transform 1 0 5796 0 -1 4752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_59
timestamp 1608761684
transform 1 0 6532 0 -1 4752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_62
timestamp 1608761684
transform 1 0 6808 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_27
timestamp 1608761684
transform 1 0 3588 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_39
timestamp 1608761684
transform 1 0 4692 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608761684
transform 1 0 1104 0 -1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1608761684
transform 1 0 1380 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1608761684
transform 1 0 2484 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608761684
transform -1 0 21620 0 1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608761684
transform 1 0 20792 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_215
timestamp 1608761684
transform 1 0 20884 0 1 3664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_219
timestamp 1608761684
transform 1 0 21252 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_190
timestamp 1608761684
transform 1 0 18584 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_202
timestamp 1608761684
transform 1 0 19688 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_178
timestamp 1608761684
transform 1 0 17480 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608761684
transform 1 0 15180 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_154
timestamp 1608761684
transform 1 0 15272 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_166
timestamp 1608761684
transform 1 0 16376 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_129
timestamp 1608761684
transform 1 0 12972 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_141
timestamp 1608761684
transform 1 0 14076 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_105
timestamp 1608761684
transform 1 0 10764 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_117
timestamp 1608761684
transform 1 0 11868 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608761684
transform 1 0 9568 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1608761684
transform 1 0 9660 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_68
timestamp 1608761684
transform 1 0 7360 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_80
timestamp 1608761684
transform 1 0 8464 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_44
timestamp 1608761684
transform 1 0 5152 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_56
timestamp 1608761684
transform 1 0 6256 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608761684
transform 1 0 3956 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1608761684
transform 1 0 3588 0 1 3664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_32
timestamp 1608761684
transform 1 0 4048 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608761684
transform 1 0 1104 0 1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1608761684
transform 1 0 1380 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1608761684
transform 1 0 2484 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608761684
transform -1 0 21620 0 -1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_196
timestamp 1608761684
transform 1 0 19136 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_208
timestamp 1608761684
transform 1 0 20240 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608761684
transform 1 0 17940 0 -1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_171
timestamp 1608761684
transform 1 0 16836 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_184
timestamp 1608761684
transform 1 0 18032 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_147
timestamp 1608761684
transform 1 0 14628 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_159
timestamp 1608761684
transform 1 0 15732 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_135
timestamp 1608761684
transform 1 0 13524 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608761684
transform 1 0 12328 0 -1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_110
timestamp 1608761684
transform 1 0 11224 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_123
timestamp 1608761684
transform 1 0 12420 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_86
timestamp 1608761684
transform 1 0 9016 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_98
timestamp 1608761684
transform 1 0 10120 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_74
timestamp 1608761684
transform 1 0 7912 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608761684
transform 1 0 6716 0 -1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_51
timestamp 1608761684
transform 1 0 5796 0 -1 3664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_59
timestamp 1608761684
transform 1 0 6532 0 -1 3664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_62
timestamp 1608761684
transform 1 0 6808 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_27
timestamp 1608761684
transform 1 0 3588 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_39
timestamp 1608761684
transform 1 0 4692 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608761684
transform 1 0 1104 0 -1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1608761684
transform 1 0 1380 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1608761684
transform 1 0 2484 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608761684
transform -1 0 21620 0 -1 2576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608761684
transform -1 0 21620 0 1 2576
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608761684
transform 1 0 21068 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608761684
transform 1 0 20792 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1608761684
transform 1 0 20516 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1608761684
transform 1 0 21160 0 -1 2576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1608761684
transform 1 0 20884 0 1 2576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_219
timestamp 1608761684
transform 1 0 21252 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1608761684
transform 1 0 19412 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_190
timestamp 1608761684
transform 1 0 18584 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_202
timestamp 1608761684
transform 1 0 19688 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608761684
transform 1 0 18216 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1608761684
transform 1 0 16560 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1608761684
transform 1 0 17664 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1608761684
transform 1 0 18308 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_178
timestamp 1608761684
transform 1 0 17480 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608761684
transform 1 0 15364 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608761684
transform 1 0 15180 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1608761684
transform 1 0 14812 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1608761684
transform 1 0 15456 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_154
timestamp 1608761684
transform 1 0 15272 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_166
timestamp 1608761684
transform 1 0 16376 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1608761684
transform 1 0 13708 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_129
timestamp 1608761684
transform 1 0 12972 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_141
timestamp 1608761684
transform 1 0 14076 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608761684
transform 1 0 12512 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1608761684
transform 1 0 10856 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1608761684
transform 1 0 11960 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1608761684
transform 1 0 12604 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_105
timestamp 1608761684
transform 1 0 10764 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_117
timestamp 1608761684
transform 1 0 11868 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1608761684
transform 1 0 9660 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608761684
transform 1 0 9568 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1608761684
transform 1 0 9108 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1608761684
transform 1 0 9752 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_93
timestamp 1608761684
transform 1 0 9660 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1608761684
transform 1 0 6900 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1608761684
transform 1 0 8004 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_68
timestamp 1608761684
transform 1 0 7360 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_80
timestamp 1608761684
transform 1 0 8464 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1608761684
transform 1 0 6808 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1608761684
transform 1 0 5152 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56
timestamp 1608761684
transform 1 0 6256 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_44
timestamp 1608761684
transform 1 0 5152 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_56
timestamp 1608761684
transform 1 0 6256 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1608761684
transform 1 0 3956 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608761684
transform 1 0 3956 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1608761684
transform 1 0 3588 0 -1 2576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1608761684
transform 1 0 4048 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1608761684
transform 1 0 3588 0 1 2576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_32
timestamp 1608761684
transform 1 0 4048 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608761684
transform 1 0 1104 0 -1 2576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1608761684
transform 1 0 1104 0 1 2576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1608761684
transform 1 0 1380 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1608761684
transform 1 0 2484 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1608761684
transform 1 0 1380 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1608761684
transform 1 0 2484 0 1 2576
box -38 -48 1142 592
<< labels >>
rlabel metal3 s 0 5576 800 5696 4 ccff_head
port 1 nsew
rlabel metal3 s 0 17000 800 17120 4 ccff_tail
port 2 nsew
rlabel metal3 s 22000 4080 22800 4200 4 chanx_right_in[0]
port 3 nsew
rlabel metal3 s 22000 8568 22800 8688 4 chanx_right_in[10]
port 4 nsew
rlabel metal3 s 22000 9112 22800 9232 4 chanx_right_in[11]
port 5 nsew
rlabel metal3 s 22000 9520 22800 9640 4 chanx_right_in[12]
port 6 nsew
rlabel metal3 s 22000 9928 22800 10048 4 chanx_right_in[13]
port 7 nsew
rlabel metal3 s 22000 10472 22800 10592 4 chanx_right_in[14]
port 8 nsew
rlabel metal3 s 22000 10880 22800 11000 4 chanx_right_in[15]
port 9 nsew
rlabel metal3 s 22000 11424 22800 11544 4 chanx_right_in[16]
port 10 nsew
rlabel metal3 s 22000 11832 22800 11952 4 chanx_right_in[17]
port 11 nsew
rlabel metal3 s 22000 12240 22800 12360 4 chanx_right_in[18]
port 12 nsew
rlabel metal3 s 22000 12784 22800 12904 4 chanx_right_in[19]
port 13 nsew
rlabel metal3 s 22000 4488 22800 4608 4 chanx_right_in[1]
port 14 nsew
rlabel metal3 s 22000 4896 22800 5016 4 chanx_right_in[2]
port 15 nsew
rlabel metal3 s 22000 5440 22800 5560 4 chanx_right_in[3]
port 16 nsew
rlabel metal3 s 22000 5848 22800 5968 4 chanx_right_in[4]
port 17 nsew
rlabel metal3 s 22000 6392 22800 6512 4 chanx_right_in[5]
port 18 nsew
rlabel metal3 s 22000 6800 22800 6920 4 chanx_right_in[6]
port 19 nsew
rlabel metal3 s 22000 7208 22800 7328 4 chanx_right_in[7]
port 20 nsew
rlabel metal3 s 22000 7752 22800 7872 4 chanx_right_in[8]
port 21 nsew
rlabel metal3 s 22000 8160 22800 8280 4 chanx_right_in[9]
port 22 nsew
rlabel metal3 s 22000 13192 22800 13312 4 chanx_right_out[0]
port 23 nsew
rlabel metal3 s 22000 17816 22800 17936 4 chanx_right_out[10]
port 24 nsew
rlabel metal3 s 22000 18224 22800 18344 4 chanx_right_out[11]
port 25 nsew
rlabel metal3 s 22000 18632 22800 18752 4 chanx_right_out[12]
port 26 nsew
rlabel metal3 s 22000 19176 22800 19296 4 chanx_right_out[13]
port 27 nsew
rlabel metal3 s 22000 19584 22800 19704 4 chanx_right_out[14]
port 28 nsew
rlabel metal3 s 22000 19992 22800 20112 4 chanx_right_out[15]
port 29 nsew
rlabel metal3 s 22000 20536 22800 20656 4 chanx_right_out[16]
port 30 nsew
rlabel metal3 s 22000 20944 22800 21064 4 chanx_right_out[17]
port 31 nsew
rlabel metal3 s 22000 21352 22800 21472 4 chanx_right_out[18]
port 32 nsew
rlabel metal3 s 22000 21896 22800 22016 4 chanx_right_out[19]
port 33 nsew
rlabel metal3 s 22000 13600 22800 13720 4 chanx_right_out[1]
port 34 nsew
rlabel metal3 s 22000 14144 22800 14264 4 chanx_right_out[2]
port 35 nsew
rlabel metal3 s 22000 14552 22800 14672 4 chanx_right_out[3]
port 36 nsew
rlabel metal3 s 22000 14960 22800 15080 4 chanx_right_out[4]
port 37 nsew
rlabel metal3 s 22000 15504 22800 15624 4 chanx_right_out[5]
port 38 nsew
rlabel metal3 s 22000 15912 22800 16032 4 chanx_right_out[6]
port 39 nsew
rlabel metal3 s 22000 16320 22800 16440 4 chanx_right_out[7]
port 40 nsew
rlabel metal3 s 22000 16864 22800 16984 4 chanx_right_out[8]
port 41 nsew
rlabel metal3 s 22000 17272 22800 17392 4 chanx_right_out[9]
port 42 nsew
rlabel metal2 s 846 21856 902 22656 4 chany_top_in[0]
port 43 nsew
rlabel metal2 s 6366 21856 6422 22656 4 chany_top_in[10]
port 44 nsew
rlabel metal2 s 6918 21856 6974 22656 4 chany_top_in[11]
port 45 nsew
rlabel metal2 s 7470 21856 7526 22656 4 chany_top_in[12]
port 46 nsew
rlabel metal2 s 8022 21856 8078 22656 4 chany_top_in[13]
port 47 nsew
rlabel metal2 s 8574 21856 8630 22656 4 chany_top_in[14]
port 48 nsew
rlabel metal2 s 9126 21856 9182 22656 4 chany_top_in[15]
port 49 nsew
rlabel metal2 s 9678 21856 9734 22656 4 chany_top_in[16]
port 50 nsew
rlabel metal2 s 10230 21856 10286 22656 4 chany_top_in[17]
port 51 nsew
rlabel metal2 s 10782 21856 10838 22656 4 chany_top_in[18]
port 52 nsew
rlabel metal2 s 11334 21856 11390 22656 4 chany_top_in[19]
port 53 nsew
rlabel metal2 s 1398 21856 1454 22656 4 chany_top_in[1]
port 54 nsew
rlabel metal2 s 1950 21856 2006 22656 4 chany_top_in[2]
port 55 nsew
rlabel metal2 s 2502 21856 2558 22656 4 chany_top_in[3]
port 56 nsew
rlabel metal2 s 3054 21856 3110 22656 4 chany_top_in[4]
port 57 nsew
rlabel metal2 s 3606 21856 3662 22656 4 chany_top_in[5]
port 58 nsew
rlabel metal2 s 4158 21856 4214 22656 4 chany_top_in[6]
port 59 nsew
rlabel metal2 s 4710 21856 4766 22656 4 chany_top_in[7]
port 60 nsew
rlabel metal2 s 5262 21856 5318 22656 4 chany_top_in[8]
port 61 nsew
rlabel metal2 s 5814 21856 5870 22656 4 chany_top_in[9]
port 62 nsew
rlabel metal2 s 11978 21856 12034 22656 4 chany_top_out[0]
port 63 nsew
rlabel metal2 s 17498 21856 17554 22656 4 chany_top_out[10]
port 64 nsew
rlabel metal2 s 18050 21856 18106 22656 4 chany_top_out[11]
port 65 nsew
rlabel metal2 s 18602 21856 18658 22656 4 chany_top_out[12]
port 66 nsew
rlabel metal2 s 19154 21856 19210 22656 4 chany_top_out[13]
port 67 nsew
rlabel metal2 s 19706 21856 19762 22656 4 chany_top_out[14]
port 68 nsew
rlabel metal2 s 20258 21856 20314 22656 4 chany_top_out[15]
port 69 nsew
rlabel metal2 s 20810 21856 20866 22656 4 chany_top_out[16]
port 70 nsew
rlabel metal2 s 21362 21856 21418 22656 4 chany_top_out[17]
port 71 nsew
rlabel metal2 s 21914 21856 21970 22656 4 chany_top_out[18]
port 72 nsew
rlabel metal2 s 22466 21856 22522 22656 4 chany_top_out[19]
port 73 nsew
rlabel metal2 s 12530 21856 12586 22656 4 chany_top_out[1]
port 74 nsew
rlabel metal2 s 13082 21856 13138 22656 4 chany_top_out[2]
port 75 nsew
rlabel metal2 s 13634 21856 13690 22656 4 chany_top_out[3]
port 76 nsew
rlabel metal2 s 14186 21856 14242 22656 4 chany_top_out[4]
port 77 nsew
rlabel metal2 s 14738 21856 14794 22656 4 chany_top_out[5]
port 78 nsew
rlabel metal2 s 15290 21856 15346 22656 4 chany_top_out[6]
port 79 nsew
rlabel metal2 s 15842 21856 15898 22656 4 chany_top_out[7]
port 80 nsew
rlabel metal2 s 16394 21856 16450 22656 4 chany_top_out[8]
port 81 nsew
rlabel metal2 s 16946 21856 17002 22656 4 chany_top_out[9]
port 82 nsew
rlabel metal3 s 22000 22304 22800 22424 4 prog_clk_0_E_in
port 83 nsew
rlabel metal3 s 22000 2176 22800 2296 4 right_bottom_grid_pin_11_
port 84 nsew
rlabel metal3 s 22000 2720 22800 2840 4 right_bottom_grid_pin_13_
port 85 nsew
rlabel metal3 s 22000 3128 22800 3248 4 right_bottom_grid_pin_15_
port 86 nsew
rlabel metal3 s 22000 3536 22800 3656 4 right_bottom_grid_pin_17_
port 87 nsew
rlabel metal3 s 22000 0 22800 120 4 right_bottom_grid_pin_1_
port 88 nsew
rlabel metal3 s 22000 408 22800 528 4 right_bottom_grid_pin_3_
port 89 nsew
rlabel metal3 s 22000 816 22800 936 4 right_bottom_grid_pin_5_
port 90 nsew
rlabel metal3 s 22000 1360 22800 1480 4 right_bottom_grid_pin_7_
port 91 nsew
rlabel metal3 s 22000 1768 22800 1888 4 right_bottom_grid_pin_9_
port 92 nsew
rlabel metal2 s 294 21856 350 22656 4 top_left_grid_pin_1_
port 93 nsew
rlabel metal4 s 4376 1984 4696 20032 4 VPWR
port 94 nsew
rlabel metal4 s 7808 1984 8128 20032 4 VGND
port 95 nsew
<< properties >>
string FIXED_BBOX 0 0 22800 22656
string GDS_FILE /ef/openfpga/openlane/runs/sb_0__0_/results/magic/sb_0__0_.gds
string GDS_END 646960
string GDS_START 78430
<< end >>
