magic
tech sky130A
magscale 1 2
timestamp 1608134833
<< obsli1 >>
rect 1104 2159 15824 17425
<< obsm1 >>
rect 750 1096 16822 18080
<< metal2 >>
rect 110 19200 166 20000
rect 386 19200 442 20000
rect 754 19200 810 20000
rect 1122 19200 1178 20000
rect 1398 19200 1454 20000
rect 1766 19200 1822 20000
rect 2134 19200 2190 20000
rect 2410 19200 2466 20000
rect 2778 19200 2834 20000
rect 3146 19200 3202 20000
rect 3514 19200 3570 20000
rect 3790 19200 3846 20000
rect 4158 19200 4214 20000
rect 4526 19200 4582 20000
rect 4802 19200 4858 20000
rect 5170 19200 5226 20000
rect 5538 19200 5594 20000
rect 5814 19200 5870 20000
rect 6182 19200 6238 20000
rect 6550 19200 6606 20000
rect 6918 19200 6974 20000
rect 7194 19200 7250 20000
rect 7562 19200 7618 20000
rect 7930 19200 7986 20000
rect 8206 19200 8262 20000
rect 8574 19200 8630 20000
rect 8942 19200 8998 20000
rect 9218 19200 9274 20000
rect 9586 19200 9642 20000
rect 9954 19200 10010 20000
rect 10322 19200 10378 20000
rect 10598 19200 10654 20000
rect 10966 19200 11022 20000
rect 11334 19200 11390 20000
rect 11610 19200 11666 20000
rect 11978 19200 12034 20000
rect 12346 19200 12402 20000
rect 12622 19200 12678 20000
rect 12990 19200 13046 20000
rect 13358 19200 13414 20000
rect 13726 19200 13782 20000
rect 14002 19200 14058 20000
rect 14370 19200 14426 20000
rect 14738 19200 14794 20000
rect 15014 19200 15070 20000
rect 15382 19200 15438 20000
rect 15750 19200 15806 20000
rect 16026 19200 16082 20000
rect 16394 19200 16450 20000
rect 16762 19200 16818 20000
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1122 0 1178 800
rect 1398 0 1454 800
rect 1766 0 1822 800
rect 2134 0 2190 800
rect 2410 0 2466 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3514 0 3570 800
rect 3790 0 3846 800
rect 4158 0 4214 800
rect 4526 0 4582 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5814 0 5870 800
rect 6182 0 6238 800
rect 6550 0 6606 800
rect 6918 0 6974 800
rect 7194 0 7250 800
rect 7562 0 7618 800
rect 7930 0 7986 800
rect 8206 0 8262 800
rect 8574 0 8630 800
rect 8942 0 8998 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10598 0 10654 800
rect 10966 0 11022 800
rect 11334 0 11390 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12622 0 12678 800
rect 12990 0 13046 800
rect 13358 0 13414 800
rect 13726 0 13782 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15014 0 15070 800
rect 15382 0 15438 800
rect 15750 0 15806 800
rect 16026 0 16082 800
rect 16394 0 16450 800
rect 16762 0 16818 800
<< obsm2 >>
rect 222 19144 330 19417
rect 498 19144 698 19417
rect 866 19144 1066 19417
rect 1234 19144 1342 19417
rect 1510 19144 1710 19417
rect 1878 19144 2078 19417
rect 2246 19144 2354 19417
rect 2522 19144 2722 19417
rect 2890 19144 3090 19417
rect 3258 19144 3458 19417
rect 3626 19144 3734 19417
rect 3902 19144 4102 19417
rect 4270 19144 4470 19417
rect 4638 19144 4746 19417
rect 4914 19144 5114 19417
rect 5282 19144 5482 19417
rect 5650 19144 5758 19417
rect 5926 19144 6126 19417
rect 6294 19144 6494 19417
rect 6662 19144 6862 19417
rect 7030 19144 7138 19417
rect 7306 19144 7506 19417
rect 7674 19144 7874 19417
rect 8042 19144 8150 19417
rect 8318 19144 8518 19417
rect 8686 19144 8886 19417
rect 9054 19144 9162 19417
rect 9330 19144 9530 19417
rect 9698 19144 9898 19417
rect 10066 19144 10266 19417
rect 10434 19144 10542 19417
rect 10710 19144 10910 19417
rect 11078 19144 11278 19417
rect 11446 19144 11554 19417
rect 11722 19144 11922 19417
rect 12090 19144 12290 19417
rect 12458 19144 12566 19417
rect 12734 19144 12934 19417
rect 13102 19144 13302 19417
rect 13470 19144 13670 19417
rect 13838 19144 13946 19417
rect 14114 19144 14314 19417
rect 14482 19144 14682 19417
rect 14850 19144 14958 19417
rect 15126 19144 15326 19417
rect 15494 19144 15694 19417
rect 15862 19144 15970 19417
rect 16138 19144 16338 19417
rect 16506 19144 16706 19417
rect 110 856 16816 19144
rect 222 439 330 856
rect 498 439 698 856
rect 866 439 1066 856
rect 1234 439 1342 856
rect 1510 439 1710 856
rect 1878 439 2078 856
rect 2246 439 2354 856
rect 2522 439 2722 856
rect 2890 439 3090 856
rect 3258 439 3458 856
rect 3626 439 3734 856
rect 3902 439 4102 856
rect 4270 439 4470 856
rect 4638 439 4746 856
rect 4914 439 5114 856
rect 5282 439 5482 856
rect 5650 439 5758 856
rect 5926 439 6126 856
rect 6294 439 6494 856
rect 6662 439 6862 856
rect 7030 439 7138 856
rect 7306 439 7506 856
rect 7674 439 7874 856
rect 8042 439 8150 856
rect 8318 439 8518 856
rect 8686 439 8886 856
rect 9054 439 9162 856
rect 9330 439 9530 856
rect 9698 439 9898 856
rect 10066 439 10266 856
rect 10434 439 10542 856
rect 10710 439 10910 856
rect 11078 439 11278 856
rect 11446 439 11554 856
rect 11722 439 11922 856
rect 12090 439 12290 856
rect 12458 439 12566 856
rect 12734 439 12934 856
rect 13102 439 13302 856
rect 13470 439 13670 856
rect 13838 439 13946 856
rect 14114 439 14314 856
rect 14482 439 14682 856
rect 14850 439 14958 856
rect 15126 439 15326 856
rect 15494 439 15694 856
rect 15862 439 15970 856
rect 16138 439 16338 856
rect 16506 439 16706 856
<< metal3 >>
rect 0 19320 800 19440
rect 0 18368 800 18488
rect 0 17280 800 17400
rect 16200 16600 17000 16720
rect 0 16328 800 16448
rect 0 15376 800 15496
rect 0 14288 800 14408
rect 0 13336 800 13456
rect 0 12384 800 12504
rect 0 11296 800 11416
rect 0 10344 800 10464
rect 16200 9936 17000 10056
rect 0 9392 800 9512
rect 0 8304 800 8424
rect 0 7352 800 7472
rect 0 6400 800 6520
rect 0 5312 800 5432
rect 0 4360 800 4480
rect 0 3408 800 3528
rect 16200 3272 17000 3392
rect 0 2320 800 2440
rect 0 1368 800 1488
rect 0 416 800 536
<< obsm3 >>
rect 880 19240 16200 19413
rect 105 18568 16200 19240
rect 880 18288 16200 18568
rect 105 17480 16200 18288
rect 880 17200 16200 17480
rect 105 16800 16200 17200
rect 105 16528 16120 16800
rect 880 16520 16120 16528
rect 880 16248 16200 16520
rect 105 15576 16200 16248
rect 880 15296 16200 15576
rect 105 14488 16200 15296
rect 880 14208 16200 14488
rect 105 13536 16200 14208
rect 880 13256 16200 13536
rect 105 12584 16200 13256
rect 880 12304 16200 12584
rect 105 11496 16200 12304
rect 880 11216 16200 11496
rect 105 10544 16200 11216
rect 880 10264 16200 10544
rect 105 10136 16200 10264
rect 105 9856 16120 10136
rect 105 9592 16200 9856
rect 880 9312 16200 9592
rect 105 8504 16200 9312
rect 880 8224 16200 8504
rect 105 7552 16200 8224
rect 880 7272 16200 7552
rect 105 6600 16200 7272
rect 880 6320 16200 6600
rect 105 5512 16200 6320
rect 880 5232 16200 5512
rect 105 4560 16200 5232
rect 880 4280 16200 4560
rect 105 3608 16200 4280
rect 880 3472 16200 3608
rect 880 3328 16120 3472
rect 105 3192 16120 3328
rect 105 2520 16200 3192
rect 880 2240 16200 2520
rect 105 1568 16200 2240
rect 880 1288 16200 1568
rect 105 616 16200 1288
rect 880 443 16200 616
<< metal4 >>
rect 3409 2128 3729 17456
rect 5875 2128 6195 17456
<< obsm4 >>
rect 4659 2048 5795 17456
rect 6275 2048 14845 17456
rect 4659 1531 14845 2048
<< labels >>
rlabel metal3 s 16200 16600 17000 16720 6 Test_en_E_in
port 1 nsew default input
rlabel metal3 s 16200 9936 17000 10056 6 Test_en_E_out
port 2 nsew default output
rlabel metal2 s 3146 19200 3202 20000 6 Test_en_N_out
port 3 nsew default output
rlabel metal2 s 13726 0 13782 800 6 Test_en_S_in
port 4 nsew default input
rlabel metal3 s 0 17280 800 17400 6 Test_en_W_in
port 5 nsew default input
rlabel metal3 s 0 18368 800 18488 6 Test_en_W_out
port 6 nsew default output
rlabel metal3 s 0 416 800 536 6 ccff_head
port 7 nsew default input
rlabel metal3 s 16200 3272 17000 3392 6 ccff_tail
port 8 nsew default output
rlabel metal2 s 6918 0 6974 800 6 chany_bottom_in[0]
port 9 nsew default input
rlabel metal2 s 10322 0 10378 800 6 chany_bottom_in[10]
port 10 nsew default input
rlabel metal2 s 10598 0 10654 800 6 chany_bottom_in[11]
port 11 nsew default input
rlabel metal2 s 10966 0 11022 800 6 chany_bottom_in[12]
port 12 nsew default input
rlabel metal2 s 11334 0 11390 800 6 chany_bottom_in[13]
port 13 nsew default input
rlabel metal2 s 11610 0 11666 800 6 chany_bottom_in[14]
port 14 nsew default input
rlabel metal2 s 11978 0 12034 800 6 chany_bottom_in[15]
port 15 nsew default input
rlabel metal2 s 12346 0 12402 800 6 chany_bottom_in[16]
port 16 nsew default input
rlabel metal2 s 12622 0 12678 800 6 chany_bottom_in[17]
port 17 nsew default input
rlabel metal2 s 12990 0 13046 800 6 chany_bottom_in[18]
port 18 nsew default input
rlabel metal2 s 13358 0 13414 800 6 chany_bottom_in[19]
port 19 nsew default input
rlabel metal2 s 7194 0 7250 800 6 chany_bottom_in[1]
port 20 nsew default input
rlabel metal2 s 7562 0 7618 800 6 chany_bottom_in[2]
port 21 nsew default input
rlabel metal2 s 7930 0 7986 800 6 chany_bottom_in[3]
port 22 nsew default input
rlabel metal2 s 8206 0 8262 800 6 chany_bottom_in[4]
port 23 nsew default input
rlabel metal2 s 8574 0 8630 800 6 chany_bottom_in[5]
port 24 nsew default input
rlabel metal2 s 8942 0 8998 800 6 chany_bottom_in[6]
port 25 nsew default input
rlabel metal2 s 9218 0 9274 800 6 chany_bottom_in[7]
port 26 nsew default input
rlabel metal2 s 9586 0 9642 800 6 chany_bottom_in[8]
port 27 nsew default input
rlabel metal2 s 9954 0 10010 800 6 chany_bottom_in[9]
port 28 nsew default input
rlabel metal2 s 110 0 166 800 6 chany_bottom_out[0]
port 29 nsew default output
rlabel metal2 s 3514 0 3570 800 6 chany_bottom_out[10]
port 30 nsew default output
rlabel metal2 s 3790 0 3846 800 6 chany_bottom_out[11]
port 31 nsew default output
rlabel metal2 s 4158 0 4214 800 6 chany_bottom_out[12]
port 32 nsew default output
rlabel metal2 s 4526 0 4582 800 6 chany_bottom_out[13]
port 33 nsew default output
rlabel metal2 s 4802 0 4858 800 6 chany_bottom_out[14]
port 34 nsew default output
rlabel metal2 s 5170 0 5226 800 6 chany_bottom_out[15]
port 35 nsew default output
rlabel metal2 s 5538 0 5594 800 6 chany_bottom_out[16]
port 36 nsew default output
rlabel metal2 s 5814 0 5870 800 6 chany_bottom_out[17]
port 37 nsew default output
rlabel metal2 s 6182 0 6238 800 6 chany_bottom_out[18]
port 38 nsew default output
rlabel metal2 s 6550 0 6606 800 6 chany_bottom_out[19]
port 39 nsew default output
rlabel metal2 s 386 0 442 800 6 chany_bottom_out[1]
port 40 nsew default output
rlabel metal2 s 754 0 810 800 6 chany_bottom_out[2]
port 41 nsew default output
rlabel metal2 s 1122 0 1178 800 6 chany_bottom_out[3]
port 42 nsew default output
rlabel metal2 s 1398 0 1454 800 6 chany_bottom_out[4]
port 43 nsew default output
rlabel metal2 s 1766 0 1822 800 6 chany_bottom_out[5]
port 44 nsew default output
rlabel metal2 s 2134 0 2190 800 6 chany_bottom_out[6]
port 45 nsew default output
rlabel metal2 s 2410 0 2466 800 6 chany_bottom_out[7]
port 46 nsew default output
rlabel metal2 s 2778 0 2834 800 6 chany_bottom_out[8]
port 47 nsew default output
rlabel metal2 s 3146 0 3202 800 6 chany_bottom_out[9]
port 48 nsew default output
rlabel metal2 s 10322 19200 10378 20000 6 chany_top_in[0]
port 49 nsew default input
rlabel metal2 s 13726 19200 13782 20000 6 chany_top_in[10]
port 50 nsew default input
rlabel metal2 s 14002 19200 14058 20000 6 chany_top_in[11]
port 51 nsew default input
rlabel metal2 s 14370 19200 14426 20000 6 chany_top_in[12]
port 52 nsew default input
rlabel metal2 s 14738 19200 14794 20000 6 chany_top_in[13]
port 53 nsew default input
rlabel metal2 s 15014 19200 15070 20000 6 chany_top_in[14]
port 54 nsew default input
rlabel metal2 s 15382 19200 15438 20000 6 chany_top_in[15]
port 55 nsew default input
rlabel metal2 s 15750 19200 15806 20000 6 chany_top_in[16]
port 56 nsew default input
rlabel metal2 s 16026 19200 16082 20000 6 chany_top_in[17]
port 57 nsew default input
rlabel metal2 s 16394 19200 16450 20000 6 chany_top_in[18]
port 58 nsew default input
rlabel metal2 s 16762 19200 16818 20000 6 chany_top_in[19]
port 59 nsew default input
rlabel metal2 s 10598 19200 10654 20000 6 chany_top_in[1]
port 60 nsew default input
rlabel metal2 s 10966 19200 11022 20000 6 chany_top_in[2]
port 61 nsew default input
rlabel metal2 s 11334 19200 11390 20000 6 chany_top_in[3]
port 62 nsew default input
rlabel metal2 s 11610 19200 11666 20000 6 chany_top_in[4]
port 63 nsew default input
rlabel metal2 s 11978 19200 12034 20000 6 chany_top_in[5]
port 64 nsew default input
rlabel metal2 s 12346 19200 12402 20000 6 chany_top_in[6]
port 65 nsew default input
rlabel metal2 s 12622 19200 12678 20000 6 chany_top_in[7]
port 66 nsew default input
rlabel metal2 s 12990 19200 13046 20000 6 chany_top_in[8]
port 67 nsew default input
rlabel metal2 s 13358 19200 13414 20000 6 chany_top_in[9]
port 68 nsew default input
rlabel metal2 s 3514 19200 3570 20000 6 chany_top_out[0]
port 69 nsew default output
rlabel metal2 s 6918 19200 6974 20000 6 chany_top_out[10]
port 70 nsew default output
rlabel metal2 s 7194 19200 7250 20000 6 chany_top_out[11]
port 71 nsew default output
rlabel metal2 s 7562 19200 7618 20000 6 chany_top_out[12]
port 72 nsew default output
rlabel metal2 s 7930 19200 7986 20000 6 chany_top_out[13]
port 73 nsew default output
rlabel metal2 s 8206 19200 8262 20000 6 chany_top_out[14]
port 74 nsew default output
rlabel metal2 s 8574 19200 8630 20000 6 chany_top_out[15]
port 75 nsew default output
rlabel metal2 s 8942 19200 8998 20000 6 chany_top_out[16]
port 76 nsew default output
rlabel metal2 s 9218 19200 9274 20000 6 chany_top_out[17]
port 77 nsew default output
rlabel metal2 s 9586 19200 9642 20000 6 chany_top_out[18]
port 78 nsew default output
rlabel metal2 s 9954 19200 10010 20000 6 chany_top_out[19]
port 79 nsew default output
rlabel metal2 s 3790 19200 3846 20000 6 chany_top_out[1]
port 80 nsew default output
rlabel metal2 s 4158 19200 4214 20000 6 chany_top_out[2]
port 81 nsew default output
rlabel metal2 s 4526 19200 4582 20000 6 chany_top_out[3]
port 82 nsew default output
rlabel metal2 s 4802 19200 4858 20000 6 chany_top_out[4]
port 83 nsew default output
rlabel metal2 s 5170 19200 5226 20000 6 chany_top_out[5]
port 84 nsew default output
rlabel metal2 s 5538 19200 5594 20000 6 chany_top_out[6]
port 85 nsew default output
rlabel metal2 s 5814 19200 5870 20000 6 chany_top_out[7]
port 86 nsew default output
rlabel metal2 s 6182 19200 6238 20000 6 chany_top_out[8]
port 87 nsew default output
rlabel metal2 s 6550 19200 6606 20000 6 chany_top_out[9]
port 88 nsew default output
rlabel metal2 s 110 19200 166 20000 6 clk_2_N_in
port 89 nsew default input
rlabel metal2 s 1398 19200 1454 20000 6 clk_2_N_out
port 90 nsew default output
rlabel metal2 s 14002 0 14058 800 6 clk_2_S_in
port 91 nsew default input
rlabel metal2 s 15382 0 15438 800 6 clk_2_S_out
port 92 nsew default output
rlabel metal2 s 386 19200 442 20000 6 clk_3_N_in
port 93 nsew default input
rlabel metal2 s 1766 19200 1822 20000 6 clk_3_N_out
port 94 nsew default output
rlabel metal2 s 14370 0 14426 800 6 clk_3_S_in
port 95 nsew default input
rlabel metal2 s 15750 0 15806 800 6 clk_3_S_out
port 96 nsew default output
rlabel metal3 s 0 1368 800 1488 6 left_grid_pin_16_
port 97 nsew default output
rlabel metal3 s 0 2320 800 2440 6 left_grid_pin_17_
port 98 nsew default output
rlabel metal3 s 0 3408 800 3528 6 left_grid_pin_18_
port 99 nsew default output
rlabel metal3 s 0 4360 800 4480 6 left_grid_pin_19_
port 100 nsew default output
rlabel metal3 s 0 5312 800 5432 6 left_grid_pin_20_
port 101 nsew default output
rlabel metal3 s 0 6400 800 6520 6 left_grid_pin_21_
port 102 nsew default output
rlabel metal3 s 0 7352 800 7472 6 left_grid_pin_22_
port 103 nsew default output
rlabel metal3 s 0 8304 800 8424 6 left_grid_pin_23_
port 104 nsew default output
rlabel metal3 s 0 9392 800 9512 6 left_grid_pin_24_
port 105 nsew default output
rlabel metal3 s 0 10344 800 10464 6 left_grid_pin_25_
port 106 nsew default output
rlabel metal3 s 0 11296 800 11416 6 left_grid_pin_26_
port 107 nsew default output
rlabel metal3 s 0 12384 800 12504 6 left_grid_pin_27_
port 108 nsew default output
rlabel metal3 s 0 13336 800 13456 6 left_grid_pin_28_
port 109 nsew default output
rlabel metal3 s 0 14288 800 14408 6 left_grid_pin_29_
port 110 nsew default output
rlabel metal3 s 0 15376 800 15496 6 left_grid_pin_30_
port 111 nsew default output
rlabel metal3 s 0 16328 800 16448 6 left_grid_pin_31_
port 112 nsew default output
rlabel metal2 s 2134 19200 2190 20000 6 prog_clk_0_N_out
port 113 nsew default output
rlabel metal2 s 16026 0 16082 800 6 prog_clk_0_S_out
port 114 nsew default output
rlabel metal3 s 0 19320 800 19440 6 prog_clk_0_W_in
port 115 nsew default input
rlabel metal2 s 754 19200 810 20000 6 prog_clk_2_N_in
port 116 nsew default input
rlabel metal2 s 2410 19200 2466 20000 6 prog_clk_2_N_out
port 117 nsew default output
rlabel metal2 s 14738 0 14794 800 6 prog_clk_2_S_in
port 118 nsew default input
rlabel metal2 s 16394 0 16450 800 6 prog_clk_2_S_out
port 119 nsew default output
rlabel metal2 s 1122 19200 1178 20000 6 prog_clk_3_N_in
port 120 nsew default input
rlabel metal2 s 2778 19200 2834 20000 6 prog_clk_3_N_out
port 121 nsew default output
rlabel metal2 s 15014 0 15070 800 6 prog_clk_3_S_in
port 122 nsew default input
rlabel metal2 s 16762 0 16818 800 6 prog_clk_3_S_out
port 123 nsew default output
rlabel metal4 s 3409 2128 3729 17456 6 VPWR
port 124 nsew power input
rlabel metal4 s 5875 2128 6195 17456 6 VGND
port 125 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 17000 20000
string LEFview TRUE
<< end >>
