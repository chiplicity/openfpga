version https://git-lfs.github.com/spec/v1
oid sha256:bc199ee8a5c7ab44636d4e6f185b21ecd54835de4f9438dc6685bc8495316f58
size 36407428
