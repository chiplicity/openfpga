magic
tech EFS8A
magscale 1 2
timestamp 1604437673
<< locali >>
rect 31769 33371 31803 33609
rect 31861 32215 31895 32521
rect 29101 18139 29135 18309
rect 28917 16983 28951 17085
rect 6469 14807 6503 14909
rect 21557 2975 21591 3145
<< viali >>
rect 35633 35785 35667 35819
rect 30205 35581 30239 35615
rect 35449 35581 35483 35615
rect 36001 35581 36035 35615
rect 30472 35513 30506 35547
rect 30021 35445 30055 35479
rect 31585 35445 31619 35479
rect 29929 35241 29963 35275
rect 30849 35241 30883 35275
rect 36185 35241 36219 35275
rect 30297 35105 30331 35139
rect 30941 35105 30975 35139
rect 34345 35105 34379 35139
rect 34805 35105 34839 35139
rect 36001 35105 36035 35139
rect 31125 35037 31159 35071
rect 34897 35037 34931 35071
rect 34989 35037 35023 35071
rect 30481 34901 30515 34935
rect 33333 34901 33367 34935
rect 34437 34901 34471 34935
rect 35541 34901 35575 34935
rect 29101 34697 29135 34731
rect 31401 34697 31435 34731
rect 32781 34697 32815 34731
rect 34345 34697 34379 34731
rect 37565 34697 37599 34731
rect 32045 34629 32079 34663
rect 36277 34629 36311 34663
rect 29561 34561 29595 34595
rect 33149 34561 33183 34595
rect 33701 34561 33735 34595
rect 33885 34561 33919 34595
rect 30021 34493 30055 34527
rect 30288 34493 30322 34527
rect 33609 34493 33643 34527
rect 34897 34493 34931 34527
rect 35153 34493 35187 34527
rect 36829 34493 36863 34527
rect 37381 34493 37415 34527
rect 37933 34493 37967 34527
rect 29837 34357 29871 34391
rect 33241 34357 33275 34391
rect 34621 34357 34655 34391
rect 28365 34153 28399 34187
rect 34161 34153 34195 34187
rect 36093 34153 36127 34187
rect 34958 34085 34992 34119
rect 28457 34017 28491 34051
rect 29828 34017 29862 34051
rect 32393 34017 32427 34051
rect 28641 33949 28675 33983
rect 29561 33949 29595 33983
rect 32137 33949 32171 33983
rect 34713 33949 34747 33983
rect 27997 33813 28031 33847
rect 30941 33813 30975 33847
rect 31953 33813 31987 33847
rect 33517 33813 33551 33847
rect 34621 33813 34655 33847
rect 27721 33609 27755 33643
rect 28089 33609 28123 33643
rect 28733 33609 28767 33643
rect 31769 33609 31803 33643
rect 32045 33609 32079 33643
rect 33885 33609 33919 33643
rect 36277 33609 36311 33643
rect 29653 33405 29687 33439
rect 29920 33405 29954 33439
rect 34253 33541 34287 33575
rect 34621 33541 34655 33575
rect 32597 33473 32631 33507
rect 32781 33473 32815 33507
rect 34897 33473 34931 33507
rect 33149 33405 33183 33439
rect 33701 33405 33735 33439
rect 31769 33337 31803 33371
rect 32505 33337 32539 33371
rect 35164 33337 35198 33371
rect 29101 33269 29135 33303
rect 29469 33269 29503 33303
rect 31033 33269 31067 33303
rect 31585 33269 31619 33303
rect 32137 33269 32171 33303
rect 33609 33269 33643 33303
rect 28089 33065 28123 33099
rect 29469 33065 29503 33099
rect 31861 33065 31895 33099
rect 33241 33065 33275 33099
rect 34253 33065 34287 33099
rect 36093 33065 36127 33099
rect 29828 32997 29862 33031
rect 32505 32929 32539 32963
rect 34621 32929 34655 32963
rect 34980 32929 35014 32963
rect 29561 32861 29595 32895
rect 32597 32861 32631 32895
rect 32781 32861 32815 32895
rect 34713 32861 34747 32895
rect 32137 32793 32171 32827
rect 30941 32725 30975 32759
rect 29101 32521 29135 32555
rect 31861 32521 31895 32555
rect 32045 32521 32079 32555
rect 32689 32521 32723 32555
rect 34253 32521 34287 32555
rect 34621 32521 34655 32555
rect 36277 32521 36311 32555
rect 37565 32521 37599 32555
rect 29653 32317 29687 32351
rect 31677 32317 31711 32351
rect 28733 32249 28767 32283
rect 29898 32249 29932 32283
rect 33149 32385 33183 32419
rect 33701 32385 33735 32419
rect 33793 32385 33827 32419
rect 34897 32385 34931 32419
rect 32137 32317 32171 32351
rect 33609 32317 33643 32351
rect 37381 32317 37415 32351
rect 37933 32317 37967 32351
rect 35164 32249 35198 32283
rect 29469 32181 29503 32215
rect 31033 32181 31067 32215
rect 31861 32181 31895 32215
rect 32321 32181 32355 32215
rect 33241 32181 33275 32215
rect 29101 31977 29135 32011
rect 30021 31977 30055 32011
rect 33425 31977 33459 32011
rect 36001 31977 36035 32011
rect 31125 31909 31159 31943
rect 32413 31909 32447 31943
rect 34069 31909 34103 31943
rect 28917 31841 28951 31875
rect 30389 31841 30423 31875
rect 32873 31841 32907 31875
rect 34621 31841 34655 31875
rect 35265 31841 35299 31875
rect 35817 31841 35851 31875
rect 30481 31773 30515 31807
rect 30665 31773 30699 31807
rect 34713 31773 34747 31807
rect 34805 31773 34839 31807
rect 29561 31705 29595 31739
rect 31677 31637 31711 31671
rect 33057 31637 33091 31671
rect 34253 31637 34287 31671
rect 29009 31433 29043 31467
rect 29561 31433 29595 31467
rect 29929 31433 29963 31467
rect 32965 31433 32999 31467
rect 33609 31433 33643 31467
rect 34621 31433 34655 31467
rect 36277 31433 36311 31467
rect 36829 31433 36863 31467
rect 30021 31365 30055 31399
rect 31033 31365 31067 31399
rect 30481 31297 30515 31331
rect 30573 31297 30607 31331
rect 31493 31297 31527 31331
rect 32045 31297 32079 31331
rect 32137 31297 32171 31331
rect 34897 31297 34931 31331
rect 28273 31229 28307 31263
rect 28641 31161 28675 31195
rect 30389 31161 30423 31195
rect 33977 31161 34011 31195
rect 34345 31161 34379 31195
rect 35164 31161 35198 31195
rect 31585 31093 31619 31127
rect 31953 31093 31987 31127
rect 31585 30889 31619 30923
rect 32597 30889 32631 30923
rect 33333 30889 33367 30923
rect 35817 30889 35851 30923
rect 29828 30821 29862 30855
rect 34682 30821 34716 30855
rect 29561 30753 29595 30787
rect 34437 30753 34471 30787
rect 32689 30685 32723 30719
rect 32873 30685 32907 30719
rect 29469 30549 29503 30583
rect 30941 30549 30975 30583
rect 32229 30549 32263 30583
rect 34345 30549 34379 30583
rect 32321 30345 32355 30379
rect 32689 30345 32723 30379
rect 33057 30345 33091 30379
rect 34529 30345 34563 30379
rect 28273 30277 28307 30311
rect 31677 30277 31711 30311
rect 32045 30277 32079 30311
rect 33241 30277 33275 30311
rect 28733 30209 28767 30243
rect 29101 30209 29135 30243
rect 29377 30209 29411 30243
rect 33885 30209 33919 30243
rect 34897 30209 34931 30243
rect 28089 30141 28123 30175
rect 32137 30141 32171 30175
rect 33609 30141 33643 30175
rect 29622 30073 29656 30107
rect 35142 30073 35176 30107
rect 27997 30005 28031 30039
rect 30757 30005 30791 30039
rect 33701 30005 33735 30039
rect 36277 30005 36311 30039
rect 30113 29801 30147 29835
rect 33333 29801 33367 29835
rect 34253 29801 34287 29835
rect 35265 29801 35299 29835
rect 36001 29801 36035 29835
rect 28448 29733 28482 29767
rect 30665 29733 30699 29767
rect 34161 29733 34195 29767
rect 28181 29665 28215 29699
rect 30849 29665 30883 29699
rect 31033 29665 31067 29699
rect 32137 29665 32171 29699
rect 34621 29665 34655 29699
rect 35817 29665 35851 29699
rect 34713 29597 34747 29631
rect 34805 29597 34839 29631
rect 35633 29529 35667 29563
rect 27721 29461 27755 29495
rect 29561 29461 29595 29495
rect 32321 29461 32355 29495
rect 33701 29461 33735 29495
rect 30021 29257 30055 29291
rect 31033 29257 31067 29291
rect 32137 29257 32171 29291
rect 33609 29257 33643 29291
rect 34713 29257 34747 29291
rect 36277 29257 36311 29291
rect 28733 29189 28767 29223
rect 29101 29189 29135 29223
rect 31401 29189 31435 29223
rect 33885 29189 33919 29223
rect 28273 29121 28307 29155
rect 29561 29121 29595 29155
rect 30665 29121 30699 29155
rect 34345 29121 34379 29155
rect 34897 29121 34931 29155
rect 28089 29053 28123 29087
rect 29929 29053 29963 29087
rect 30481 29053 30515 29087
rect 33701 29053 33735 29087
rect 27537 28985 27571 29019
rect 27997 28985 28031 29019
rect 30389 28985 30423 29019
rect 35142 28985 35176 29019
rect 27629 28917 27663 28951
rect 30113 28713 30147 28747
rect 34345 28713 34379 28747
rect 34989 28713 35023 28747
rect 35633 28713 35667 28747
rect 36737 28713 36771 28747
rect 27721 28645 27755 28679
rect 28264 28645 28298 28679
rect 27997 28577 28031 28611
rect 30481 28577 30515 28611
rect 35449 28577 35483 28611
rect 36553 28577 36587 28611
rect 32413 28509 32447 28543
rect 29377 28373 29411 28407
rect 30665 28373 30699 28407
rect 36001 28373 36035 28407
rect 27997 28169 28031 28203
rect 28641 28169 28675 28203
rect 29285 28169 29319 28203
rect 30665 28169 30699 28203
rect 32229 28169 32263 28203
rect 32321 28169 32355 28203
rect 35633 28169 35667 28203
rect 30297 28101 30331 28135
rect 28181 28033 28215 28067
rect 29745 28033 29779 28067
rect 29837 28033 29871 28067
rect 31861 28033 31895 28067
rect 32873 28033 32907 28067
rect 29101 27965 29135 27999
rect 29653 27965 29687 27999
rect 32689 27965 32723 27999
rect 35449 27965 35483 27999
rect 36645 27965 36679 27999
rect 31493 27897 31527 27931
rect 32781 27897 32815 27931
rect 35357 27829 35391 27863
rect 36001 27829 36035 27863
rect 29929 27625 29963 27659
rect 32137 27625 32171 27659
rect 34152 27557 34186 27591
rect 23121 27489 23155 27523
rect 24409 27489 24443 27523
rect 24961 27489 24995 27523
rect 28917 27489 28951 27523
rect 32505 27489 32539 27523
rect 28457 27421 28491 27455
rect 29009 27421 29043 27455
rect 29101 27421 29135 27455
rect 30113 27421 30147 27455
rect 32597 27421 32631 27455
rect 32689 27421 32723 27455
rect 33885 27421 33919 27455
rect 36369 27421 36403 27455
rect 28089 27353 28123 27387
rect 29561 27353 29595 27387
rect 31953 27353 31987 27387
rect 21925 27285 21959 27319
rect 23305 27285 23339 27319
rect 24593 27285 24627 27319
rect 28549 27285 28583 27319
rect 35265 27285 35299 27319
rect 35817 27285 35851 27319
rect 31309 27081 31343 27115
rect 33149 27081 33183 27115
rect 36369 27081 36403 27115
rect 21373 26945 21407 26979
rect 22385 26945 22419 26979
rect 29285 26945 29319 26979
rect 22201 26877 22235 26911
rect 24593 26877 24627 26911
rect 24685 26877 24719 26911
rect 27997 26877 28031 26911
rect 29552 26877 29586 26911
rect 31769 26877 31803 26911
rect 32036 26877 32070 26911
rect 34989 26877 35023 26911
rect 35256 26877 35290 26911
rect 21741 26809 21775 26843
rect 24225 26809 24259 26843
rect 24930 26809 24964 26843
rect 27905 26809 27939 26843
rect 28181 26809 28215 26843
rect 31677 26809 31711 26843
rect 33977 26809 34011 26843
rect 21833 26741 21867 26775
rect 22293 26741 22327 26775
rect 23121 26741 23155 26775
rect 26065 26741 26099 26775
rect 28365 26741 28399 26775
rect 28733 26741 28767 26775
rect 29101 26741 29135 26775
rect 30665 26741 30699 26775
rect 34253 26741 34287 26775
rect 34621 26741 34655 26775
rect 22845 26537 22879 26571
rect 23765 26537 23799 26571
rect 27905 26537 27939 26571
rect 30389 26537 30423 26571
rect 34437 26537 34471 26571
rect 36277 26537 36311 26571
rect 21732 26469 21766 26503
rect 24194 26469 24228 26503
rect 29254 26469 29288 26503
rect 31585 26469 31619 26503
rect 32680 26469 32714 26503
rect 35164 26469 35198 26503
rect 23949 26401 23983 26435
rect 26525 26401 26559 26435
rect 26792 26401 26826 26435
rect 29009 26401 29043 26435
rect 21465 26333 21499 26367
rect 32413 26333 32447 26367
rect 34897 26333 34931 26367
rect 25329 26265 25363 26299
rect 28549 26265 28583 26299
rect 31861 26265 31895 26299
rect 33793 26265 33827 26299
rect 21189 26197 21223 26231
rect 34713 26197 34747 26231
rect 20453 25993 20487 26027
rect 20821 25993 20855 26027
rect 22293 25993 22327 26027
rect 22845 25993 22879 26027
rect 25329 25993 25363 26027
rect 28641 25993 28675 26027
rect 29469 25993 29503 26027
rect 31769 25993 31803 26027
rect 34897 25925 34931 25959
rect 20913 25857 20947 25891
rect 33885 25857 33919 25891
rect 35449 25857 35483 25891
rect 35909 25857 35943 25891
rect 36277 25857 36311 25891
rect 23489 25789 23523 25823
rect 23949 25789 23983 25823
rect 25973 25789 26007 25823
rect 26341 25789 26375 25823
rect 26433 25789 26467 25823
rect 29285 25789 29319 25823
rect 30389 25789 30423 25823
rect 30656 25789 30690 25823
rect 34621 25789 34655 25823
rect 35357 25789 35391 25823
rect 21180 25721 21214 25755
rect 24216 25721 24250 25755
rect 26678 25721 26712 25755
rect 29929 25721 29963 25755
rect 33149 25721 33183 25755
rect 33609 25721 33643 25755
rect 34345 25721 34379 25755
rect 35265 25721 35299 25755
rect 36461 25721 36495 25755
rect 27813 25653 27847 25687
rect 29101 25653 29135 25687
rect 30205 25653 30239 25687
rect 32413 25653 32447 25687
rect 33241 25653 33275 25687
rect 33701 25653 33735 25687
rect 24041 25449 24075 25483
rect 24501 25449 24535 25483
rect 26249 25449 26283 25483
rect 26985 25449 27019 25483
rect 27905 25449 27939 25483
rect 29285 25449 29319 25483
rect 29561 25449 29595 25483
rect 29929 25449 29963 25483
rect 32689 25449 32723 25483
rect 33701 25449 33735 25483
rect 23673 25381 23707 25415
rect 24593 25381 24627 25415
rect 25237 25381 25271 25415
rect 30021 25381 30055 25415
rect 32505 25381 32539 25415
rect 20913 25313 20947 25347
rect 21180 25313 21214 25347
rect 26801 25313 26835 25347
rect 28273 25313 28307 25347
rect 33057 25313 33091 25347
rect 34345 25313 34379 25347
rect 24685 25245 24719 25279
rect 25513 25245 25547 25279
rect 28365 25245 28399 25279
rect 28549 25245 28583 25279
rect 30205 25245 30239 25279
rect 33149 25245 33183 25279
rect 33333 25245 33367 25279
rect 34437 25245 34471 25279
rect 34760 25245 34794 25279
rect 34897 25245 34931 25279
rect 35173 25245 35207 25279
rect 36277 25245 36311 25279
rect 31953 25177 31987 25211
rect 20637 25109 20671 25143
rect 22293 25109 22327 25143
rect 24133 25109 24167 25143
rect 27353 25109 27387 25143
rect 20453 24905 20487 24939
rect 24685 24905 24719 24939
rect 27629 24905 27663 24939
rect 27997 24905 28031 24939
rect 29653 24905 29687 24939
rect 31769 24905 31803 24939
rect 34529 24905 34563 24939
rect 34897 24905 34931 24939
rect 24317 24837 24351 24871
rect 30021 24837 30055 24871
rect 20545 24769 20579 24803
rect 25605 24769 25639 24803
rect 26433 24769 26467 24803
rect 27169 24769 27203 24803
rect 32184 24769 32218 24803
rect 32321 24769 32355 24803
rect 32597 24769 32631 24803
rect 35357 24769 35391 24803
rect 35541 24769 35575 24803
rect 35909 24769 35943 24803
rect 23673 24701 23707 24735
rect 26065 24701 26099 24735
rect 27077 24701 27111 24735
rect 30205 24701 30239 24735
rect 30757 24701 30791 24735
rect 31861 24701 31895 24735
rect 36277 24701 36311 24735
rect 20790 24633 20824 24667
rect 28365 24633 28399 24667
rect 31309 24633 31343 24667
rect 35265 24633 35299 24667
rect 20085 24565 20119 24599
rect 21925 24565 21959 24599
rect 23489 24565 23523 24599
rect 23857 24565 23891 24599
rect 25053 24565 25087 24599
rect 25421 24565 25455 24599
rect 25513 24565 25547 24599
rect 26617 24565 26651 24599
rect 26985 24565 27019 24599
rect 28733 24565 28767 24599
rect 30389 24565 30423 24599
rect 33701 24565 33735 24599
rect 20545 24361 20579 24395
rect 22753 24361 22787 24395
rect 24317 24361 24351 24395
rect 24685 24361 24719 24395
rect 25421 24361 25455 24395
rect 26801 24361 26835 24395
rect 27537 24361 27571 24395
rect 31953 24361 31987 24395
rect 33057 24361 33091 24395
rect 33425 24361 33459 24395
rect 34989 24361 35023 24395
rect 35357 24361 35391 24395
rect 21649 24293 21683 24327
rect 23121 24293 23155 24327
rect 24777 24293 24811 24327
rect 27997 24293 28031 24327
rect 30481 24293 30515 24327
rect 21557 24225 21591 24259
rect 27353 24225 27387 24259
rect 28457 24225 28491 24259
rect 28724 24225 28758 24259
rect 35725 24225 35759 24259
rect 21833 24157 21867 24191
rect 23213 24157 23247 24191
rect 23397 24157 23431 24191
rect 24961 24157 24995 24191
rect 35817 24157 35851 24191
rect 36001 24157 36035 24191
rect 21189 24021 21223 24055
rect 24133 24021 24167 24055
rect 29837 24021 29871 24055
rect 32689 24021 32723 24055
rect 34069 24021 34103 24055
rect 34529 24021 34563 24055
rect 20269 23817 20303 23851
rect 20729 23817 20763 23851
rect 22201 23817 22235 23851
rect 22845 23817 22879 23851
rect 23121 23817 23155 23851
rect 23949 23817 23983 23851
rect 25881 23817 25915 23851
rect 26157 23817 26191 23851
rect 26617 23817 26651 23851
rect 27445 23817 27479 23851
rect 28641 23817 28675 23851
rect 29285 23817 29319 23851
rect 34897 23817 34931 23851
rect 36645 23817 36679 23851
rect 24409 23749 24443 23783
rect 27629 23749 27663 23783
rect 30665 23749 30699 23783
rect 21833 23681 21867 23715
rect 25053 23681 25087 23715
rect 28273 23681 28307 23715
rect 29745 23681 29779 23715
rect 29837 23681 29871 23715
rect 30297 23681 30331 23715
rect 34345 23681 34379 23715
rect 35449 23681 35483 23715
rect 21557 23613 21591 23647
rect 24777 23613 24811 23647
rect 25973 23613 26007 23647
rect 27077 23613 27111 23647
rect 27997 23613 28031 23647
rect 35909 23613 35943 23647
rect 21649 23545 21683 23579
rect 24317 23545 24351 23579
rect 24869 23545 24903 23579
rect 29101 23545 29135 23579
rect 29653 23545 29687 23579
rect 30849 23545 30883 23579
rect 35265 23545 35299 23579
rect 19993 23477 20027 23511
rect 21005 23477 21039 23511
rect 21189 23477 21223 23511
rect 25421 23477 25455 23511
rect 28089 23477 28123 23511
rect 34713 23477 34747 23511
rect 35357 23477 35391 23511
rect 36277 23477 36311 23511
rect 20729 23273 20763 23307
rect 22293 23273 22327 23307
rect 23397 23273 23431 23307
rect 23765 23273 23799 23307
rect 24409 23273 24443 23307
rect 25145 23273 25179 23307
rect 26985 23273 27019 23307
rect 28457 23273 28491 23307
rect 34161 23273 34195 23307
rect 36553 23273 36587 23307
rect 21169 23137 21203 23171
rect 22937 23137 22971 23171
rect 23305 23137 23339 23171
rect 24961 23137 24995 23171
rect 27905 23137 27939 23171
rect 29265 23137 29299 23171
rect 35440 23137 35474 23171
rect 20913 23069 20947 23103
rect 23857 23069 23891 23103
rect 24041 23069 24075 23103
rect 24869 23069 24903 23103
rect 29009 23069 29043 23103
rect 35173 23069 35207 23103
rect 27721 23001 27755 23035
rect 28089 22933 28123 22967
rect 28917 22933 28951 22967
rect 30389 22933 30423 22967
rect 34897 22933 34931 22967
rect 20913 22729 20947 22763
rect 21557 22729 21591 22763
rect 24685 22729 24719 22763
rect 25421 22729 25455 22763
rect 27905 22729 27939 22763
rect 28365 22729 28399 22763
rect 28641 22729 28675 22763
rect 29009 22729 29043 22763
rect 36737 22729 36771 22763
rect 23673 22661 23707 22695
rect 20269 22593 20303 22627
rect 22109 22593 22143 22627
rect 24317 22593 24351 22627
rect 25881 22593 25915 22627
rect 26433 22593 26467 22627
rect 27445 22593 27479 22627
rect 29285 22593 29319 22627
rect 22017 22525 22051 22559
rect 23489 22525 23523 22559
rect 24133 22525 24167 22559
rect 25237 22525 25271 22559
rect 27353 22525 27387 22559
rect 29541 22525 29575 22559
rect 32229 22525 32263 22559
rect 35357 22525 35391 22559
rect 35624 22525 35658 22559
rect 22569 22457 22603 22491
rect 24041 22457 24075 22491
rect 26801 22457 26835 22491
rect 27261 22457 27295 22491
rect 31769 22457 31803 22491
rect 32474 22457 32508 22491
rect 34345 22457 34379 22491
rect 20637 22389 20671 22423
rect 21373 22389 21407 22423
rect 21925 22389 21959 22423
rect 23121 22389 23155 22423
rect 25053 22389 25087 22423
rect 26893 22389 26927 22423
rect 30665 22389 30699 22423
rect 32137 22389 32171 22423
rect 33609 22389 33643 22423
rect 34621 22389 34655 22423
rect 35173 22389 35207 22423
rect 22293 22185 22327 22219
rect 23397 22185 23431 22219
rect 24961 22185 24995 22219
rect 27263 22185 27297 22219
rect 34807 22185 34841 22219
rect 36737 22185 36771 22219
rect 23305 22117 23339 22151
rect 23765 22117 23799 22151
rect 21169 22049 21203 22083
rect 25329 22049 25363 22083
rect 30113 22049 30147 22083
rect 32505 22049 32539 22083
rect 33885 22049 33919 22083
rect 35081 22049 35115 22083
rect 20913 21981 20947 22015
rect 23857 21981 23891 22015
rect 23949 21981 23983 22015
rect 24409 21981 24443 22015
rect 26801 21981 26835 22015
rect 27261 21981 27295 22015
rect 27537 21981 27571 22015
rect 28641 21981 28675 22015
rect 29193 21981 29227 22015
rect 30205 21981 30239 22015
rect 30389 21981 30423 22015
rect 31953 21981 31987 22015
rect 32597 21981 32631 22015
rect 32689 21981 32723 22015
rect 34345 21981 34379 22015
rect 34805 21981 34839 22015
rect 36185 21981 36219 22015
rect 25513 21913 25547 21947
rect 30757 21913 30791 21947
rect 26341 21845 26375 21879
rect 29561 21845 29595 21879
rect 29745 21845 29779 21879
rect 32137 21845 32171 21879
rect 33425 21845 33459 21879
rect 34161 21845 34195 21879
rect 20913 21641 20947 21675
rect 22385 21641 22419 21675
rect 23673 21641 23707 21675
rect 25053 21641 25087 21675
rect 25697 21641 25731 21675
rect 27629 21641 27663 21675
rect 28641 21641 28675 21675
rect 31769 21641 31803 21675
rect 34345 21641 34379 21675
rect 36277 21641 36311 21675
rect 20545 21505 20579 21539
rect 21005 21505 21039 21539
rect 24225 21505 24259 21539
rect 29285 21505 29319 21539
rect 29745 21505 29779 21539
rect 30021 21505 30055 21539
rect 32229 21505 32263 21539
rect 26249 21437 26283 21471
rect 32496 21437 32530 21471
rect 34897 21437 34931 21471
rect 20177 21369 20211 21403
rect 21272 21369 21306 21403
rect 23121 21369 23155 21403
rect 24041 21369 24075 21403
rect 26516 21369 26550 21403
rect 28181 21369 28215 21403
rect 32137 21369 32171 21403
rect 35164 21369 35198 21403
rect 36829 21369 36863 21403
rect 23489 21301 23523 21335
rect 24133 21301 24167 21335
rect 24685 21301 24719 21335
rect 25237 21301 25271 21335
rect 26065 21301 26099 21335
rect 29101 21301 29135 21335
rect 29747 21301 29781 21335
rect 31125 21301 31159 21335
rect 33609 21301 33643 21335
rect 37381 21301 37415 21335
rect 20729 21097 20763 21131
rect 22293 21097 22327 21131
rect 23213 21097 23247 21131
rect 24777 21097 24811 21131
rect 25973 21097 26007 21131
rect 26985 21097 27019 21131
rect 27629 21097 27663 21131
rect 29745 21097 29779 21131
rect 30665 21097 30699 21131
rect 31953 21097 31987 21131
rect 32967 21097 33001 21131
rect 34345 21097 34379 21131
rect 34897 21097 34931 21131
rect 35357 21097 35391 21131
rect 35817 21097 35851 21131
rect 21180 21029 21214 21063
rect 23664 21029 23698 21063
rect 26341 21029 26375 21063
rect 20913 20961 20947 20995
rect 26893 20961 26927 20995
rect 28365 20961 28399 20995
rect 28632 20961 28666 20995
rect 23397 20893 23431 20927
rect 27169 20893 27203 20927
rect 30849 20893 30883 20927
rect 32321 20893 32355 20927
rect 32505 20893 32539 20927
rect 32965 20893 32999 20927
rect 33241 20893 33275 20927
rect 35909 20893 35943 20927
rect 36093 20893 36127 20927
rect 26525 20825 26559 20859
rect 35449 20825 35483 20859
rect 30297 20757 30331 20791
rect 20913 20553 20947 20587
rect 21373 20553 21407 20587
rect 22753 20553 22787 20587
rect 25697 20553 25731 20587
rect 27537 20553 27571 20587
rect 32597 20553 32631 20587
rect 33609 20553 33643 20587
rect 34621 20553 34655 20587
rect 35909 20553 35943 20587
rect 36277 20553 36311 20587
rect 29377 20485 29411 20519
rect 30389 20485 30423 20519
rect 32505 20485 32539 20519
rect 34897 20485 34931 20519
rect 36645 20485 36679 20519
rect 26065 20417 26099 20451
rect 26157 20417 26191 20451
rect 29837 20417 29871 20451
rect 30021 20417 30055 20451
rect 31585 20417 31619 20451
rect 33241 20417 33275 20451
rect 35449 20417 35483 20451
rect 23673 20349 23707 20383
rect 23940 20349 23974 20383
rect 26413 20349 26447 20383
rect 23121 20281 23155 20315
rect 23489 20281 23523 20315
rect 29101 20281 29135 20315
rect 29745 20281 29779 20315
rect 32137 20281 32171 20315
rect 35357 20281 35391 20315
rect 25053 20213 25087 20247
rect 28457 20213 28491 20247
rect 32965 20213 32999 20247
rect 33057 20213 33091 20247
rect 34345 20213 34379 20247
rect 35265 20213 35299 20247
rect 23857 20009 23891 20043
rect 24409 20009 24443 20043
rect 26249 20009 26283 20043
rect 26709 20009 26743 20043
rect 27077 20009 27111 20043
rect 28457 20009 28491 20043
rect 29469 20009 29503 20043
rect 33057 20009 33091 20043
rect 33333 20009 33367 20043
rect 36093 20009 36127 20043
rect 22744 19873 22778 19907
rect 34980 19873 35014 19907
rect 22477 19805 22511 19839
rect 33701 19805 33735 19839
rect 34713 19805 34747 19839
rect 29837 19669 29871 19703
rect 32689 19669 32723 19703
rect 34621 19669 34655 19703
rect 22845 19465 22879 19499
rect 33885 19465 33919 19499
rect 34897 19465 34931 19499
rect 22569 19397 22603 19431
rect 34345 19397 34379 19431
rect 35357 19329 35391 19363
rect 35541 19329 35575 19363
rect 29745 19261 29779 19295
rect 33701 19261 33735 19295
rect 36461 19261 36495 19295
rect 37197 19261 37231 19295
rect 30012 19193 30046 19227
rect 35265 19193 35299 19227
rect 36645 19193 36679 19227
rect 29561 19125 29595 19159
rect 31125 19125 31159 19159
rect 32505 19125 32539 19159
rect 33517 19125 33551 19159
rect 34621 19125 34655 19159
rect 36001 19125 36035 19159
rect 36277 19125 36311 19159
rect 36829 19125 36863 19159
rect 25881 18921 25915 18955
rect 34897 18921 34931 18955
rect 35173 18921 35207 18955
rect 28733 18853 28767 18887
rect 29081 18785 29115 18819
rect 32689 18785 32723 18819
rect 32956 18785 32990 18819
rect 35541 18785 35575 18819
rect 28825 18717 28859 18751
rect 35633 18717 35667 18751
rect 35725 18717 35759 18751
rect 36185 18717 36219 18751
rect 30205 18581 30239 18615
rect 31033 18581 31067 18615
rect 34069 18581 34103 18615
rect 25697 18377 25731 18411
rect 36277 18377 36311 18411
rect 36829 18377 36863 18411
rect 29101 18309 29135 18343
rect 30757 18309 30791 18343
rect 33885 18309 33919 18343
rect 25789 18241 25823 18275
rect 18889 18173 18923 18207
rect 26045 18173 26079 18207
rect 28549 18173 28583 18207
rect 29929 18241 29963 18275
rect 30941 18241 30975 18275
rect 29745 18173 29779 18207
rect 32873 18173 32907 18207
rect 33701 18173 33735 18207
rect 34897 18173 34931 18207
rect 18705 18105 18739 18139
rect 19134 18105 19168 18139
rect 28825 18105 28859 18139
rect 29101 18105 29135 18139
rect 29653 18105 29687 18139
rect 31208 18105 31242 18139
rect 33241 18105 33275 18139
rect 34621 18105 34655 18139
rect 35142 18105 35176 18139
rect 20269 18037 20303 18071
rect 27169 18037 27203 18071
rect 28181 18037 28215 18071
rect 29285 18037 29319 18071
rect 30297 18037 30331 18071
rect 32321 18037 32355 18071
rect 34253 18037 34287 18071
rect 29561 17833 29595 17867
rect 30205 17833 30239 17867
rect 31125 17833 31159 17867
rect 33241 17833 33275 17867
rect 33885 17833 33919 17867
rect 34345 17833 34379 17867
rect 35817 17833 35851 17867
rect 28448 17765 28482 17799
rect 11612 17697 11646 17731
rect 21732 17697 21766 17731
rect 24205 17697 24239 17731
rect 30941 17697 30975 17731
rect 34693 17697 34727 17731
rect 11345 17629 11379 17663
rect 21465 17629 21499 17663
rect 23949 17629 23983 17663
rect 28181 17629 28215 17663
rect 33333 17629 33367 17663
rect 33425 17629 33459 17663
rect 34437 17629 34471 17663
rect 32781 17561 32815 17595
rect 8033 17493 8067 17527
rect 10885 17493 10919 17527
rect 12725 17493 12759 17527
rect 13277 17493 13311 17527
rect 18889 17493 18923 17527
rect 22845 17493 22879 17527
rect 23673 17493 23707 17527
rect 25329 17493 25363 17527
rect 27721 17493 27755 17527
rect 31861 17493 31895 17527
rect 32873 17493 32907 17527
rect 11805 17289 11839 17323
rect 22661 17289 22695 17323
rect 23121 17289 23155 17323
rect 25053 17289 25087 17323
rect 31217 17289 31251 17323
rect 31769 17289 31803 17323
rect 32965 17289 32999 17323
rect 33609 17289 33643 17323
rect 33885 17289 33919 17323
rect 37105 17289 37139 17323
rect 27537 17221 27571 17255
rect 11437 17153 11471 17187
rect 13093 17153 13127 17187
rect 27169 17153 27203 17187
rect 28273 17153 28307 17187
rect 32413 17153 32447 17187
rect 34437 17153 34471 17187
rect 35449 17153 35483 17187
rect 7941 17085 7975 17119
rect 8197 17085 8231 17119
rect 10701 17085 10735 17119
rect 11253 17085 11287 17119
rect 12265 17085 12299 17119
rect 12909 17085 12943 17119
rect 13553 17085 13587 17119
rect 20637 17085 20671 17119
rect 20729 17085 20763 17119
rect 23489 17085 23523 17119
rect 23673 17085 23707 17119
rect 23929 17085 23963 17119
rect 27997 17085 28031 17119
rect 28089 17085 28123 17119
rect 28917 17085 28951 17119
rect 29285 17085 29319 17119
rect 29552 17085 29586 17119
rect 33701 17085 33735 17119
rect 35265 17085 35299 17119
rect 35909 17085 35943 17119
rect 36461 17085 36495 17119
rect 20269 17017 20303 17051
rect 20996 17017 21030 17051
rect 31585 17017 31619 17051
rect 32229 17017 32263 17051
rect 7757 16949 7791 16983
rect 9321 16949 9355 16983
rect 10793 16949 10827 16983
rect 11161 16949 11195 16983
rect 12449 16949 12483 16983
rect 12817 16949 12851 16983
rect 22109 16949 22143 16983
rect 27629 16949 27663 16983
rect 28641 16949 28675 16983
rect 28917 16949 28951 16983
rect 29009 16949 29043 16983
rect 30665 16949 30699 16983
rect 32137 16949 32171 16983
rect 34897 16949 34931 16983
rect 35357 16949 35391 16983
rect 36645 16949 36679 16983
rect 7297 16745 7331 16779
rect 8309 16745 8343 16779
rect 12725 16745 12759 16779
rect 23121 16745 23155 16779
rect 24225 16745 24259 16779
rect 28273 16745 28307 16779
rect 29745 16745 29779 16779
rect 30389 16745 30423 16779
rect 31125 16745 31159 16779
rect 31861 16745 31895 16779
rect 32137 16745 32171 16779
rect 33149 16745 33183 16779
rect 33793 16745 33827 16779
rect 34253 16745 34287 16779
rect 35357 16745 35391 16779
rect 35633 16745 35667 16779
rect 9413 16677 9447 16711
rect 10057 16677 10091 16711
rect 10885 16677 10919 16711
rect 22008 16677 22042 16711
rect 24593 16677 24627 16711
rect 32597 16677 32631 16711
rect 34069 16677 34103 16711
rect 7757 16609 7791 16643
rect 8217 16609 8251 16643
rect 11601 16609 11635 16643
rect 13277 16609 13311 16643
rect 24685 16609 24719 16643
rect 25237 16609 25271 16643
rect 26525 16609 26559 16643
rect 27077 16609 27111 16643
rect 28632 16609 28666 16643
rect 30941 16609 30975 16643
rect 32505 16609 32539 16643
rect 34621 16609 34655 16643
rect 35817 16609 35851 16643
rect 8493 16541 8527 16575
rect 10149 16541 10183 16575
rect 10333 16541 10367 16575
rect 11345 16541 11379 16575
rect 21741 16541 21775 16575
rect 24777 16541 24811 16575
rect 27445 16541 27479 16575
rect 28365 16541 28399 16575
rect 32689 16541 32723 16575
rect 34713 16541 34747 16575
rect 34805 16541 34839 16575
rect 24041 16473 24075 16507
rect 7849 16405 7883 16439
rect 9689 16405 9723 16439
rect 21465 16405 21499 16439
rect 26709 16405 26743 16439
rect 36001 16405 36035 16439
rect 7113 16201 7147 16235
rect 11161 16201 11195 16235
rect 23949 16201 23983 16235
rect 28733 16201 28767 16235
rect 29561 16201 29595 16235
rect 31861 16201 31895 16235
rect 32229 16201 32263 16235
rect 32781 16201 32815 16235
rect 33885 16201 33919 16235
rect 34345 16201 34379 16235
rect 34621 16201 34655 16235
rect 35633 16201 35667 16235
rect 36001 16201 36035 16235
rect 25881 16133 25915 16167
rect 30113 16133 30147 16167
rect 31125 16133 31159 16167
rect 33241 16133 33275 16167
rect 35357 16133 35391 16167
rect 7205 16065 7239 16099
rect 22477 16065 22511 16099
rect 22661 16065 22695 16099
rect 23029 16065 23063 16099
rect 23397 16065 23431 16099
rect 27537 16065 27571 16099
rect 30665 16065 30699 16099
rect 7472 15997 7506 16031
rect 9689 15997 9723 16031
rect 9781 15997 9815 16031
rect 11713 15997 11747 16031
rect 12173 15997 12207 16031
rect 12449 15997 12483 16031
rect 12705 15997 12739 16031
rect 21465 15997 21499 16031
rect 22385 15997 22419 16031
rect 24409 15997 24443 16031
rect 24501 15997 24535 16031
rect 26893 15997 26927 16031
rect 27445 15997 27479 16031
rect 30481 15997 30515 16031
rect 32597 15997 32631 16031
rect 33701 15997 33735 16031
rect 35449 15997 35483 16031
rect 9321 15929 9355 15963
rect 10048 15929 10082 15963
rect 24746 15929 24780 15963
rect 27353 15929 27387 15963
rect 30573 15929 30607 15963
rect 8585 15861 8619 15895
rect 13829 15861 13863 15895
rect 21741 15861 21775 15895
rect 22017 15861 22051 15895
rect 26433 15861 26467 15895
rect 26985 15861 27019 15895
rect 28457 15861 28491 15895
rect 29929 15861 29963 15895
rect 33609 15861 33643 15895
rect 8309 15657 8343 15691
rect 9137 15657 9171 15691
rect 9505 15657 9539 15691
rect 10057 15657 10091 15691
rect 11253 15657 11287 15691
rect 12725 15657 12759 15691
rect 13277 15657 13311 15691
rect 22385 15657 22419 15691
rect 23305 15657 23339 15691
rect 24317 15657 24351 15691
rect 24869 15657 24903 15691
rect 30573 15657 30607 15691
rect 34253 15657 34287 15691
rect 6285 15589 6319 15623
rect 6622 15589 6656 15623
rect 8677 15589 8711 15623
rect 11612 15589 11646 15623
rect 23213 15589 23247 15623
rect 32873 15589 32907 15623
rect 11345 15521 11379 15555
rect 22109 15521 22143 15555
rect 24777 15521 24811 15555
rect 26893 15521 26927 15555
rect 29193 15521 29227 15555
rect 29460 15521 29494 15555
rect 34069 15521 34103 15555
rect 35541 15521 35575 15555
rect 6377 15453 6411 15487
rect 10149 15453 10183 15487
rect 10241 15453 10275 15487
rect 23397 15453 23431 15487
rect 24961 15453 24995 15487
rect 25421 15453 25455 15487
rect 26985 15453 27019 15487
rect 27077 15453 27111 15487
rect 32965 15453 32999 15487
rect 33057 15453 33091 15487
rect 35633 15453 35667 15487
rect 35817 15453 35851 15487
rect 22845 15385 22879 15419
rect 23949 15385 23983 15419
rect 31953 15385 31987 15419
rect 34989 15385 35023 15419
rect 5273 15317 5307 15351
rect 7757 15317 7791 15351
rect 9689 15317 9723 15351
rect 19257 15317 19291 15351
rect 24409 15317 24443 15351
rect 26341 15317 26375 15351
rect 26525 15317 26559 15351
rect 27629 15317 27663 15351
rect 32413 15317 32447 15351
rect 32505 15317 32539 15351
rect 33517 15317 33551 15351
rect 33977 15317 34011 15351
rect 35173 15317 35207 15351
rect 36185 15317 36219 15351
rect 9413 15113 9447 15147
rect 11345 15113 11379 15147
rect 11713 15113 11747 15147
rect 18981 15113 19015 15147
rect 22845 15113 22879 15147
rect 23489 15113 23523 15147
rect 24041 15113 24075 15147
rect 26525 15113 26559 15147
rect 27629 15113 27663 15147
rect 29469 15113 29503 15147
rect 30297 15113 30331 15147
rect 34897 15113 34931 15147
rect 37105 15113 37139 15147
rect 22569 15045 22603 15079
rect 24317 15045 24351 15079
rect 32965 15045 32999 15079
rect 5825 14977 5859 15011
rect 10793 14977 10827 15011
rect 19165 14977 19199 15011
rect 24501 14977 24535 15011
rect 30481 14977 30515 15011
rect 33425 14977 33459 15011
rect 33609 14977 33643 15011
rect 35541 14977 35575 15011
rect 6469 14909 6503 14943
rect 6837 14909 6871 14943
rect 9781 14909 9815 14943
rect 10609 14909 10643 14943
rect 19421 14909 19455 14943
rect 24768 14909 24802 14943
rect 26985 14909 27019 14943
rect 27905 14909 27939 14943
rect 29101 14909 29135 14943
rect 33333 14909 33367 14943
rect 35265 14909 35299 14943
rect 36277 14909 36311 14943
rect 36461 14909 36495 14943
rect 5089 14841 5123 14875
rect 5641 14841 5675 14875
rect 7104 14841 7138 14875
rect 8953 14841 8987 14875
rect 10149 14841 10183 14875
rect 28273 14841 28307 14875
rect 30021 14841 30055 14875
rect 30748 14841 30782 14875
rect 5181 14773 5215 14807
rect 5549 14773 5583 14807
rect 6193 14773 6227 14807
rect 6469 14773 6503 14807
rect 6561 14773 6595 14807
rect 8217 14773 8251 14807
rect 10241 14773 10275 14807
rect 10701 14773 10735 14807
rect 20545 14773 20579 14807
rect 25881 14773 25915 14807
rect 27169 14773 27203 14807
rect 31861 14773 31895 14807
rect 32505 14773 32539 14807
rect 33977 14773 34011 14807
rect 34621 14773 34655 14807
rect 35357 14773 35391 14807
rect 35909 14773 35943 14807
rect 36645 14773 36679 14807
rect 7757 14569 7791 14603
rect 9965 14569 9999 14603
rect 19349 14569 19383 14603
rect 22937 14569 22971 14603
rect 23765 14569 23799 14603
rect 27169 14569 27203 14603
rect 28457 14569 28491 14603
rect 29837 14569 29871 14603
rect 30297 14569 30331 14603
rect 32965 14569 32999 14603
rect 34069 14569 34103 14603
rect 36461 14569 36495 14603
rect 10609 14501 10643 14535
rect 16865 14501 16899 14535
rect 30205 14501 30239 14535
rect 31953 14501 31987 14535
rect 5273 14433 5307 14467
rect 6092 14433 6126 14467
rect 8493 14433 8527 14467
rect 10057 14433 10091 14467
rect 11161 14433 11195 14467
rect 16313 14433 16347 14467
rect 16773 14433 16807 14467
rect 18225 14433 18259 14467
rect 24133 14433 24167 14467
rect 27077 14433 27111 14467
rect 33333 14433 33367 14467
rect 34785 14433 34819 14467
rect 5825 14365 5859 14399
rect 17049 14365 17083 14399
rect 17969 14365 18003 14399
rect 27353 14365 27387 14399
rect 30481 14365 30515 14399
rect 33425 14365 33459 14399
rect 33609 14365 33643 14399
rect 34529 14365 34563 14399
rect 7205 14229 7239 14263
rect 8677 14229 8711 14263
rect 10241 14229 10275 14263
rect 11345 14229 11379 14263
rect 15577 14229 15611 14263
rect 16405 14229 16439 14263
rect 17877 14229 17911 14263
rect 25421 14229 25455 14263
rect 26341 14229 26375 14263
rect 26709 14229 26743 14263
rect 27721 14229 27755 14263
rect 28089 14229 28123 14263
rect 32505 14229 32539 14263
rect 32873 14229 32907 14263
rect 35909 14229 35943 14263
rect 6653 14025 6687 14059
rect 8769 14025 8803 14059
rect 9229 14025 9263 14059
rect 9505 14025 9539 14059
rect 9965 14025 9999 14059
rect 17877 14025 17911 14059
rect 28457 14025 28491 14059
rect 29929 14025 29963 14059
rect 30665 14025 30699 14059
rect 31861 14025 31895 14059
rect 32137 14025 32171 14059
rect 33701 14025 33735 14059
rect 36737 14025 36771 14059
rect 5181 13957 5215 13991
rect 11069 13957 11103 13991
rect 25421 13957 25455 13991
rect 28089 13957 28123 13991
rect 30205 13957 30239 13991
rect 4721 13889 4755 13923
rect 5825 13889 5859 13923
rect 7389 13889 7423 13923
rect 7573 13889 7607 13923
rect 10517 13889 10551 13923
rect 10609 13889 10643 13923
rect 18797 13889 18831 13923
rect 19165 13889 19199 13923
rect 23121 13889 23155 13923
rect 25973 13889 26007 13923
rect 26709 13889 26743 13923
rect 26801 13889 26835 13923
rect 27629 13889 27663 13923
rect 32321 13889 32355 13923
rect 5089 13821 5123 13855
rect 7941 13821 7975 13855
rect 8309 13821 8343 13855
rect 11437 13821 11471 13855
rect 15485 13821 15519 13855
rect 15752 13821 15786 13855
rect 17509 13821 17543 13855
rect 18613 13821 18647 13855
rect 19717 13821 19751 13855
rect 19984 13821 20018 13855
rect 23489 13821 23523 13855
rect 23673 13821 23707 13855
rect 23929 13821 23963 13855
rect 27537 13821 27571 13855
rect 28825 13821 28859 13855
rect 34529 13821 34563 13855
rect 35173 13821 35207 13855
rect 35357 13821 35391 13855
rect 5641 13753 5675 13787
rect 7297 13753 7331 13787
rect 10425 13753 10459 13787
rect 18521 13753 18555 13787
rect 27445 13753 27479 13787
rect 32588 13753 32622 13787
rect 35624 13753 35658 13787
rect 5549 13685 5583 13719
rect 6193 13685 6227 13719
rect 6929 13685 6963 13719
rect 10057 13685 10091 13719
rect 15301 13685 15335 13719
rect 16865 13685 16899 13719
rect 18153 13685 18187 13719
rect 19625 13685 19659 13719
rect 21097 13685 21131 13719
rect 25053 13685 25087 13719
rect 25789 13685 25823 13719
rect 25881 13685 25915 13719
rect 26249 13685 26283 13719
rect 26617 13685 26651 13719
rect 27077 13685 27111 13719
rect 5273 13481 5307 13515
rect 7113 13481 7147 13515
rect 7665 13481 7699 13515
rect 18061 13481 18095 13515
rect 18613 13481 18647 13515
rect 19073 13481 19107 13515
rect 25513 13481 25547 13515
rect 26249 13481 26283 13515
rect 26617 13481 26651 13515
rect 27721 13481 27755 13515
rect 32413 13481 32447 13515
rect 34069 13481 34103 13515
rect 34621 13481 34655 13515
rect 35081 13481 35115 13515
rect 36553 13481 36587 13515
rect 6000 13413 6034 13447
rect 19717 13413 19751 13447
rect 21158 13413 21192 13447
rect 32956 13413 32990 13447
rect 8217 13345 8251 13379
rect 9873 13345 9907 13379
rect 11713 13345 11747 13379
rect 11805 13345 11839 13379
rect 16497 13345 16531 13379
rect 16948 13345 16982 13379
rect 19625 13345 19659 13379
rect 23489 13345 23523 13379
rect 23756 13345 23790 13379
rect 26065 13345 26099 13379
rect 26985 13345 27019 13379
rect 28089 13345 28123 13379
rect 29929 13345 29963 13379
rect 32689 13345 32723 13379
rect 35440 13345 35474 13379
rect 5733 13277 5767 13311
rect 11989 13277 12023 13311
rect 16681 13277 16715 13311
rect 19901 13277 19935 13311
rect 20913 13277 20947 13311
rect 27077 13277 27111 13311
rect 27169 13277 27203 13311
rect 28181 13277 28215 13311
rect 28365 13277 28399 13311
rect 28733 13277 28767 13311
rect 35173 13277 35207 13311
rect 16037 13209 16071 13243
rect 8033 13141 8067 13175
rect 8401 13141 8435 13175
rect 10057 13141 10091 13175
rect 10701 13141 10735 13175
rect 11345 13141 11379 13175
rect 14013 13141 14047 13175
rect 15577 13141 15611 13175
rect 19257 13141 19291 13175
rect 22293 13141 22327 13175
rect 24869 13141 24903 13175
rect 25789 13141 25823 13175
rect 29377 13141 29411 13175
rect 29653 13141 29687 13175
rect 30113 13141 30147 13175
rect 30573 13141 30607 13175
rect 6101 12937 6135 12971
rect 8769 12937 8803 12971
rect 10425 12937 10459 12971
rect 11713 12937 11747 12971
rect 12633 12937 12667 12971
rect 17785 12937 17819 12971
rect 18429 12937 18463 12971
rect 20085 12937 20119 12971
rect 24317 12937 24351 12971
rect 25145 12937 25179 12971
rect 25513 12937 25547 12971
rect 27445 12937 27479 12971
rect 28733 12937 28767 12971
rect 31217 12937 31251 12971
rect 31585 12937 31619 12971
rect 32137 12937 32171 12971
rect 33609 12937 33643 12971
rect 34621 12937 34655 12971
rect 35173 12937 35207 12971
rect 36829 12937 36863 12971
rect 17509 12869 17543 12903
rect 23949 12869 23983 12903
rect 28365 12869 28399 12903
rect 30297 12869 30331 12903
rect 11253 12801 11287 12835
rect 14473 12801 14507 12835
rect 19441 12801 19475 12835
rect 19533 12801 19567 12835
rect 29745 12801 29779 12835
rect 29837 12801 29871 12835
rect 32229 12801 32263 12835
rect 35449 12801 35483 12835
rect 6837 12733 6871 12767
rect 7104 12733 7138 12767
rect 9321 12733 9355 12767
rect 10977 12733 11011 12767
rect 12449 12733 12483 12767
rect 13001 12733 13035 12767
rect 15485 12733 15519 12767
rect 19349 12733 19383 12767
rect 20545 12733 20579 12767
rect 20812 12733 20846 12767
rect 25973 12733 26007 12767
rect 27997 12733 28031 12767
rect 29653 12733 29687 12767
rect 30849 12733 30883 12767
rect 34345 12733 34379 12767
rect 9137 12665 9171 12699
rect 11069 12665 11103 12699
rect 13829 12665 13863 12699
rect 14381 12665 14415 12699
rect 15752 12665 15786 12699
rect 18889 12665 18923 12699
rect 25881 12665 25915 12699
rect 31033 12665 31067 12699
rect 32474 12665 32508 12699
rect 35716 12665 35750 12699
rect 5825 12597 5859 12631
rect 6653 12597 6687 12631
rect 8217 12597 8251 12631
rect 9505 12597 9539 12631
rect 9965 12597 9999 12631
rect 10609 12597 10643 12631
rect 12081 12597 12115 12631
rect 13921 12597 13955 12631
rect 14289 12597 14323 12631
rect 15301 12597 15335 12631
rect 16865 12597 16899 12631
rect 18981 12597 19015 12631
rect 20453 12597 20487 12631
rect 21925 12597 21959 12631
rect 29285 12597 29319 12631
rect 30665 12597 30699 12631
rect 9689 12393 9723 12427
rect 10793 12393 10827 12427
rect 14013 12393 14047 12427
rect 16773 12393 16807 12427
rect 18337 12393 18371 12427
rect 19625 12393 19659 12427
rect 20637 12393 20671 12427
rect 26249 12393 26283 12427
rect 27905 12393 27939 12427
rect 28457 12393 28491 12427
rect 30389 12393 30423 12427
rect 32413 12393 32447 12427
rect 33149 12393 33183 12427
rect 35265 12393 35299 12427
rect 35633 12393 35667 12427
rect 6920 12325 6954 12359
rect 10149 12325 10183 12359
rect 26792 12325 26826 12359
rect 29254 12325 29288 12359
rect 32689 12325 32723 12359
rect 6653 12257 6687 12291
rect 10057 12257 10091 12291
rect 11437 12257 11471 12291
rect 11805 12257 11839 12291
rect 12164 12257 12198 12291
rect 15649 12257 15683 12291
rect 18245 12257 18279 12291
rect 19349 12257 19383 12291
rect 24021 12257 24055 12291
rect 29009 12257 29043 12291
rect 10333 12189 10367 12223
rect 11897 12189 11931 12223
rect 15393 12189 15427 12223
rect 18429 12189 18463 12223
rect 18889 12189 18923 12223
rect 23765 12189 23799 12223
rect 26525 12189 26559 12223
rect 35725 12189 35759 12223
rect 35909 12189 35943 12223
rect 8033 12053 8067 12087
rect 13277 12053 13311 12087
rect 17877 12053 17911 12087
rect 19993 12053 20027 12087
rect 21097 12053 21131 12087
rect 25145 12053 25179 12087
rect 25697 12053 25731 12087
rect 28825 12053 28859 12087
rect 36369 12053 36403 12087
rect 5917 11849 5951 11883
rect 8217 11849 8251 11883
rect 8769 11849 8803 11883
rect 11253 11849 11287 11883
rect 11897 11849 11931 11883
rect 12173 11849 12207 11883
rect 14841 11849 14875 11883
rect 17785 11849 17819 11883
rect 18613 11849 18647 11883
rect 25329 11849 25363 11883
rect 27077 11849 27111 11883
rect 27629 11849 27663 11883
rect 28273 11849 28307 11883
rect 28733 11849 28767 11883
rect 29009 11849 29043 11883
rect 35633 11849 35667 11883
rect 36001 11849 36035 11883
rect 12449 11713 12483 11747
rect 16497 11713 16531 11747
rect 17325 11713 17359 11747
rect 20913 11713 20947 11747
rect 29285 11713 29319 11747
rect 35357 11713 35391 11747
rect 6561 11645 6595 11679
rect 6837 11645 6871 11679
rect 9229 11645 9263 11679
rect 9321 11645 9355 11679
rect 14933 11645 14967 11679
rect 16313 11645 16347 11679
rect 18061 11645 18095 11679
rect 20269 11645 20303 11679
rect 20821 11645 20855 11679
rect 23489 11645 23523 11679
rect 23956 11645 23990 11679
rect 25697 11645 25731 11679
rect 25953 11645 25987 11679
rect 28089 11645 28123 11679
rect 6285 11577 6319 11611
rect 7082 11577 7116 11611
rect 9566 11577 9600 11611
rect 12716 11577 12750 11611
rect 16405 11577 16439 11611
rect 19901 11577 19935 11611
rect 23121 11577 23155 11611
rect 24216 11577 24250 11611
rect 29530 11577 29564 11611
rect 10701 11509 10735 11543
rect 13829 11509 13863 11543
rect 15393 11509 15427 11543
rect 15761 11509 15795 11543
rect 15945 11509 15979 11543
rect 16957 11509 16991 11543
rect 18245 11509 18279 11543
rect 20361 11509 20395 11543
rect 20729 11509 20763 11543
rect 21373 11509 21407 11543
rect 30665 11509 30699 11543
rect 8493 11305 8527 11339
rect 9413 11305 9447 11339
rect 10517 11305 10551 11339
rect 12449 11305 12483 11339
rect 13093 11305 13127 11339
rect 16865 11305 16899 11339
rect 18061 11305 18095 11339
rect 19349 11305 19383 11339
rect 22293 11305 22327 11339
rect 23673 11305 23707 11339
rect 24409 11305 24443 11339
rect 24777 11305 24811 11339
rect 28549 11305 28583 11339
rect 29285 11305 29319 11339
rect 30113 11305 30147 11339
rect 32321 11305 32355 11339
rect 7380 11237 7414 11271
rect 11314 11237 11348 11271
rect 21180 11237 21214 11271
rect 24041 11237 24075 11271
rect 27436 11237 27470 11271
rect 7113 11169 7147 11203
rect 9965 11169 9999 11203
rect 11069 11169 11103 11203
rect 13553 11169 13587 11203
rect 15752 11169 15786 11203
rect 18705 11169 18739 11203
rect 24869 11169 24903 11203
rect 25789 11169 25823 11203
rect 26801 11169 26835 11203
rect 27169 11169 27203 11203
rect 30021 11169 30055 11203
rect 32137 11169 32171 11203
rect 6837 11101 6871 11135
rect 15485 11101 15519 11135
rect 20913 11101 20947 11135
rect 25053 11101 25087 11135
rect 30205 11101 30239 11135
rect 10149 11033 10183 11067
rect 13737 11033 13771 11067
rect 18889 11033 18923 11067
rect 20361 11033 20395 11067
rect 29653 11033 29687 11067
rect 18429 10965 18463 10999
rect 19625 10965 19659 10999
rect 19993 10965 20027 10999
rect 35541 10965 35575 10999
rect 6653 10761 6687 10795
rect 7941 10761 7975 10795
rect 8309 10761 8343 10795
rect 9965 10761 9999 10795
rect 10517 10761 10551 10795
rect 10977 10761 11011 10795
rect 11713 10761 11747 10795
rect 13553 10761 13587 10795
rect 16865 10761 16899 10795
rect 18981 10761 19015 10795
rect 20269 10761 20303 10795
rect 24501 10761 24535 10795
rect 24869 10761 24903 10795
rect 25237 10761 25271 10795
rect 25881 10761 25915 10795
rect 26249 10761 26283 10795
rect 26893 10761 26927 10795
rect 27169 10761 27203 10795
rect 27905 10761 27939 10795
rect 28365 10761 28399 10795
rect 29101 10761 29135 10795
rect 29653 10761 29687 10795
rect 32137 10761 32171 10795
rect 36829 10761 36863 10795
rect 6285 10693 6319 10727
rect 27629 10693 27663 10727
rect 28733 10693 28767 10727
rect 7297 10625 7331 10659
rect 7389 10625 7423 10659
rect 8861 10625 8895 10659
rect 8953 10625 8987 10659
rect 12909 10625 12943 10659
rect 13093 10625 13127 10659
rect 15485 10625 15519 10659
rect 19717 10625 19751 10659
rect 19809 10625 19843 10659
rect 29837 10625 29871 10659
rect 8769 10557 8803 10591
rect 10793 10557 10827 10591
rect 12265 10557 12299 10591
rect 12817 10557 12851 10591
rect 18061 10557 18095 10591
rect 19625 10557 19659 10591
rect 20821 10557 20855 10591
rect 25697 10557 25731 10591
rect 26985 10557 27019 10591
rect 32321 10557 32355 10591
rect 32873 10557 32907 10591
rect 35449 10557 35483 10591
rect 35705 10557 35739 10591
rect 7205 10489 7239 10523
rect 10609 10489 10643 10523
rect 15025 10489 15059 10523
rect 15730 10489 15764 10523
rect 30104 10489 30138 10523
rect 6837 10421 6871 10455
rect 8401 10421 8435 10455
rect 11345 10421 11379 10455
rect 12449 10421 12483 10455
rect 15301 10421 15335 10455
rect 18245 10421 18279 10455
rect 18705 10421 18739 10455
rect 19257 10421 19291 10455
rect 20729 10421 20763 10455
rect 22109 10421 22143 10455
rect 31217 10421 31251 10455
rect 32505 10421 32539 10455
rect 33333 10421 33367 10455
rect 35265 10421 35299 10455
rect 6561 10217 6595 10251
rect 7665 10217 7699 10251
rect 8493 10217 8527 10251
rect 11069 10217 11103 10251
rect 12909 10217 12943 10251
rect 15485 10217 15519 10251
rect 15853 10217 15887 10251
rect 16405 10217 16439 10251
rect 17969 10217 18003 10251
rect 29469 10217 29503 10251
rect 29929 10217 29963 10251
rect 30481 10217 30515 10251
rect 33701 10217 33735 10251
rect 36553 10217 36587 10251
rect 7757 10149 7791 10183
rect 11805 10149 11839 10183
rect 13185 10149 13219 10183
rect 21250 10149 21284 10183
rect 9689 10081 9723 10115
rect 14105 10081 14139 10115
rect 19165 10081 19199 10115
rect 28917 10081 28951 10115
rect 30389 10081 30423 10115
rect 33609 10081 33643 10115
rect 35173 10081 35207 10115
rect 35440 10081 35474 10115
rect 6929 10013 6963 10047
rect 7849 10013 7883 10047
rect 10793 10013 10827 10047
rect 11897 10013 11931 10047
rect 12081 10013 12115 10047
rect 16497 10013 16531 10047
rect 16589 10013 16623 10047
rect 18061 10013 18095 10047
rect 18153 10013 18187 10047
rect 21005 10013 21039 10047
rect 30573 10013 30607 10047
rect 31033 10013 31067 10047
rect 33793 10013 33827 10047
rect 34897 10013 34931 10047
rect 8769 9945 8803 9979
rect 14289 9945 14323 9979
rect 16037 9945 16071 9979
rect 29101 9945 29135 9979
rect 33241 9945 33275 9979
rect 7297 9877 7331 9911
rect 9873 9877 9907 9911
rect 11437 9877 11471 9911
rect 12541 9877 12575 9911
rect 17601 9877 17635 9911
rect 18981 9877 19015 9911
rect 19349 9877 19383 9911
rect 19809 9877 19843 9911
rect 20177 9877 20211 9911
rect 20729 9877 20763 9911
rect 22385 9877 22419 9911
rect 25421 9877 25455 9911
rect 30021 9877 30055 9911
rect 32873 9877 32907 9911
rect 7297 9673 7331 9707
rect 7941 9673 7975 9707
rect 10793 9673 10827 9707
rect 14197 9673 14231 9707
rect 18245 9673 18279 9707
rect 20085 9673 20119 9707
rect 28917 9673 28951 9707
rect 29837 9673 29871 9707
rect 32597 9673 32631 9707
rect 33793 9673 33827 9707
rect 6653 9605 6687 9639
rect 8677 9605 8711 9639
rect 13921 9605 13955 9639
rect 14657 9605 14691 9639
rect 17601 9605 17635 9639
rect 18797 9605 18831 9639
rect 19993 9605 20027 9639
rect 11437 9537 11471 9571
rect 12909 9537 12943 9571
rect 13093 9537 13127 9571
rect 19349 9537 19383 9571
rect 19441 9537 19475 9571
rect 20637 9537 20671 9571
rect 33425 9537 33459 9571
rect 34161 9537 34195 9571
rect 7757 9469 7791 9503
rect 10701 9469 10735 9503
rect 11161 9469 11195 9503
rect 15485 9469 15519 9503
rect 19257 9469 19291 9503
rect 20913 9469 20947 9503
rect 21180 9469 21214 9503
rect 25329 9469 25363 9503
rect 25585 9469 25619 9503
rect 30297 9469 30331 9503
rect 32321 9469 32355 9503
rect 33149 9469 33183 9503
rect 34897 9469 34931 9503
rect 8401 9401 8435 9435
rect 9781 9401 9815 9435
rect 12817 9401 12851 9435
rect 13461 9401 13495 9435
rect 15752 9401 15786 9435
rect 20545 9401 20579 9435
rect 30542 9401 30576 9435
rect 35142 9401 35176 9435
rect 10333 9333 10367 9367
rect 11253 9333 11287 9367
rect 11897 9333 11931 9367
rect 12173 9333 12207 9367
rect 12449 9333 12483 9367
rect 15025 9333 15059 9367
rect 15301 9333 15335 9367
rect 16865 9333 16899 9367
rect 18889 9333 18923 9367
rect 20453 9333 20487 9367
rect 22293 9333 22327 9367
rect 25237 9333 25271 9367
rect 26709 9333 26743 9367
rect 30205 9333 30239 9367
rect 31677 9333 31711 9367
rect 32781 9333 32815 9367
rect 33241 9333 33275 9367
rect 34713 9333 34747 9367
rect 36277 9333 36311 9367
rect 36829 9333 36863 9367
rect 37381 9333 37415 9367
rect 10885 9129 10919 9163
rect 13645 9129 13679 9163
rect 14197 9129 14231 9163
rect 15945 9129 15979 9163
rect 16957 9129 16991 9163
rect 18705 9129 18739 9163
rect 19349 9129 19383 9163
rect 20269 9129 20303 9163
rect 25329 9129 25363 9163
rect 29745 9129 29779 9163
rect 30113 9129 30147 9163
rect 30481 9129 30515 9163
rect 33059 9129 33093 9163
rect 34437 9129 34471 9163
rect 36001 9129 36035 9163
rect 11621 9061 11655 9095
rect 11980 9061 12014 9095
rect 16313 9061 16347 9095
rect 19993 9061 20027 9095
rect 21180 9061 21214 9095
rect 25237 9061 25271 9095
rect 26770 9061 26804 9095
rect 30941 9061 30975 9095
rect 6929 8993 6963 9027
rect 7196 8993 7230 9027
rect 11713 8993 11747 9027
rect 18613 8993 18647 9027
rect 30849 8993 30883 9027
rect 32413 8993 32447 9027
rect 32597 8993 32631 9027
rect 35909 8993 35943 9027
rect 9965 8925 9999 8959
rect 15577 8925 15611 8959
rect 16405 8925 16439 8959
rect 16589 8925 16623 8959
rect 18797 8925 18831 8959
rect 20729 8925 20763 8959
rect 20913 8925 20947 8959
rect 25421 8925 25455 8959
rect 26525 8925 26559 8959
rect 31125 8925 31159 8959
rect 33057 8925 33091 8959
rect 33333 8925 33367 8959
rect 36185 8925 36219 8959
rect 18245 8857 18279 8891
rect 8309 8789 8343 8823
rect 11253 8789 11287 8823
rect 13093 8789 13127 8823
rect 17693 8789 17727 8823
rect 18153 8789 18187 8823
rect 22293 8789 22327 8823
rect 24317 8789 24351 8823
rect 24777 8789 24811 8823
rect 24869 8789 24903 8823
rect 26341 8789 26375 8823
rect 27905 8789 27939 8823
rect 35173 8789 35207 8823
rect 35541 8789 35575 8823
rect 6285 8585 6319 8619
rect 11253 8585 11287 8619
rect 14565 8585 14599 8619
rect 16313 8585 16347 8619
rect 18337 8585 18371 8619
rect 20453 8585 20487 8619
rect 21373 8585 21407 8619
rect 25605 8585 25639 8619
rect 28089 8585 28123 8619
rect 30021 8585 30055 8619
rect 30665 8585 30699 8619
rect 32505 8585 32539 8619
rect 33425 8585 33459 8619
rect 36461 8585 36495 8619
rect 37105 8585 37139 8619
rect 12265 8517 12299 8551
rect 15669 8517 15703 8551
rect 16957 8517 16991 8551
rect 4721 8449 4755 8483
rect 12725 8449 12759 8483
rect 13185 8449 13219 8483
rect 13461 8449 13495 8483
rect 30113 8449 30147 8483
rect 31033 8449 31067 8483
rect 31125 8449 31159 8483
rect 34345 8449 34379 8483
rect 3985 8381 4019 8415
rect 4537 8381 4571 8415
rect 6837 8381 6871 8415
rect 9781 8381 9815 8415
rect 9873 8381 9907 8415
rect 11805 8381 11839 8415
rect 13048 8381 13082 8415
rect 16773 8381 16807 8415
rect 17877 8381 17911 8415
rect 18981 8381 19015 8415
rect 19073 8381 19107 8415
rect 24225 8381 24259 8415
rect 24481 8381 24515 8415
rect 26709 8381 26743 8415
rect 35081 8381 35115 8415
rect 35348 8381 35382 8415
rect 3617 8313 3651 8347
rect 4445 8313 4479 8347
rect 7104 8313 7138 8347
rect 10140 8313 10174 8347
rect 16037 8313 16071 8347
rect 17417 8313 17451 8347
rect 19340 8313 19374 8347
rect 21097 8313 21131 8347
rect 24133 8313 24167 8347
rect 26954 8313 26988 8347
rect 31370 8313 31404 8347
rect 33149 8313 33183 8347
rect 34621 8313 34655 8347
rect 4077 8245 4111 8279
rect 6561 8245 6595 8279
rect 8217 8245 8251 8279
rect 26249 8245 26283 8279
rect 26525 8245 26559 8279
rect 33609 8245 33643 8279
rect 6377 8041 6411 8075
rect 7941 8041 7975 8075
rect 9965 8041 9999 8075
rect 12817 8041 12851 8075
rect 16681 8041 16715 8075
rect 21097 8041 21131 8075
rect 24777 8041 24811 8075
rect 25421 8041 25455 8075
rect 25789 8041 25823 8075
rect 26341 8041 26375 8075
rect 27077 8041 27111 8075
rect 30573 8041 30607 8075
rect 31125 8041 31159 8075
rect 34345 8041 34379 8075
rect 34989 8041 35023 8075
rect 35357 8041 35391 8075
rect 35909 8041 35943 8075
rect 36461 8041 36495 8075
rect 13461 7973 13495 8007
rect 15546 7973 15580 8007
rect 17417 7973 17451 8007
rect 19165 7973 19199 8007
rect 19717 7973 19751 8007
rect 23305 7973 23339 8007
rect 23642 7973 23676 8007
rect 26985 7973 27019 8007
rect 5264 7905 5298 7939
rect 7849 7905 7883 7939
rect 10425 7905 10459 7939
rect 10784 7905 10818 7939
rect 13369 7905 13403 7939
rect 18245 7905 18279 7939
rect 19533 7905 19567 7939
rect 19901 7905 19935 7939
rect 20913 7905 20947 7939
rect 23397 7905 23431 7939
rect 28540 7905 28574 7939
rect 33232 7905 33266 7939
rect 35817 7905 35851 7939
rect 4997 7837 5031 7871
rect 8033 7837 8067 7871
rect 10517 7837 10551 7871
rect 13645 7837 13679 7871
rect 15301 7837 15335 7871
rect 17785 7837 17819 7871
rect 18337 7837 18371 7871
rect 18521 7837 18555 7871
rect 27169 7837 27203 7871
rect 28273 7837 28307 7871
rect 32689 7837 32723 7871
rect 32965 7837 32999 7871
rect 36001 7837 36035 7871
rect 8493 7769 8527 7803
rect 14013 7769 14047 7803
rect 14381 7769 14415 7803
rect 3065 7701 3099 7735
rect 4353 7701 4387 7735
rect 6929 7701 6963 7735
rect 7297 7701 7331 7735
rect 7481 7701 7515 7735
rect 11897 7701 11931 7735
rect 13001 7701 13035 7735
rect 17877 7701 17911 7735
rect 26617 7701 26651 7735
rect 29653 7701 29687 7735
rect 35449 7701 35483 7735
rect 5365 7497 5399 7531
rect 8769 7497 8803 7531
rect 9689 7497 9723 7531
rect 12173 7497 12207 7531
rect 12817 7497 12851 7531
rect 17049 7497 17083 7531
rect 17509 7497 17543 7531
rect 19993 7497 20027 7531
rect 20453 7497 20487 7531
rect 20729 7497 20763 7531
rect 21465 7497 21499 7531
rect 23121 7497 23155 7531
rect 23489 7497 23523 7531
rect 26249 7497 26283 7531
rect 33517 7497 33551 7531
rect 37289 7497 37323 7531
rect 11713 7429 11747 7463
rect 16773 7429 16807 7463
rect 9781 7361 9815 7395
rect 13232 7361 13266 7395
rect 13369 7361 13403 7395
rect 17785 7361 17819 7395
rect 18061 7361 18095 7395
rect 23673 7361 23707 7395
rect 25881 7361 25915 7395
rect 32045 7361 32079 7395
rect 32137 7361 32171 7395
rect 35449 7361 35483 7395
rect 35909 7361 35943 7395
rect 2973 7293 3007 7327
rect 3229 7293 3263 7327
rect 5641 7293 5675 7327
rect 6837 7293 6871 7327
rect 10048 7293 10082 7327
rect 12909 7293 12943 7327
rect 13645 7293 13679 7327
rect 16865 7293 16899 7327
rect 20545 7293 20579 7327
rect 21097 7293 21131 7327
rect 22477 7293 22511 7327
rect 26709 7293 26743 7327
rect 26976 7293 27010 7327
rect 28641 7293 28675 7327
rect 34713 7293 34747 7327
rect 36185 7293 36219 7327
rect 4997 7225 5031 7259
rect 6285 7225 6319 7259
rect 7104 7225 7138 7259
rect 9321 7225 9355 7259
rect 15301 7225 15335 7259
rect 18328 7225 18362 7259
rect 23940 7225 23974 7259
rect 26617 7225 26651 7259
rect 29009 7225 29043 7259
rect 31677 7225 31711 7259
rect 32404 7225 32438 7259
rect 2513 7157 2547 7191
rect 2789 7157 2823 7191
rect 4353 7157 4387 7191
rect 5825 7157 5859 7191
rect 6561 7157 6595 7191
rect 8217 7157 8251 7191
rect 11161 7157 11195 7191
rect 14749 7157 14783 7191
rect 15669 7157 15703 7191
rect 19441 7157 19475 7191
rect 22385 7157 22419 7191
rect 22661 7157 22695 7191
rect 25053 7157 25087 7191
rect 28089 7157 28123 7191
rect 29285 7157 29319 7191
rect 34069 7157 34103 7191
rect 35265 7157 35299 7191
rect 35911 7157 35945 7191
rect 2789 6953 2823 6987
rect 5457 6953 5491 6987
rect 11437 6953 11471 6987
rect 12449 6953 12483 6987
rect 13001 6953 13035 6987
rect 25237 6953 25271 6987
rect 27077 6953 27111 6987
rect 33241 6953 33275 6987
rect 34805 6953 34839 6987
rect 35725 6953 35759 6987
rect 18061 6885 18095 6919
rect 2329 6817 2363 6851
rect 2881 6817 2915 6851
rect 4344 6817 4378 6851
rect 6817 6817 6851 6851
rect 10057 6817 10091 6851
rect 10324 6817 10358 6851
rect 12909 6817 12943 6851
rect 13553 6817 13587 6851
rect 13921 6817 13955 6851
rect 16681 6817 16715 6851
rect 19257 6817 19291 6851
rect 22376 6817 22410 6851
rect 25329 6817 25363 6851
rect 26525 6817 26559 6851
rect 28540 6817 28574 6851
rect 33333 6817 33367 6851
rect 35633 6817 35667 6851
rect 36645 6817 36679 6851
rect 1961 6749 1995 6783
rect 3065 6749 3099 6783
rect 4077 6749 4111 6783
rect 6561 6749 6595 6783
rect 13093 6749 13127 6783
rect 14105 6749 14139 6783
rect 15301 6749 15335 6783
rect 17233 6749 17267 6783
rect 17601 6749 17635 6783
rect 18153 6749 18187 6783
rect 18337 6749 18371 6783
rect 18705 6749 18739 6783
rect 22109 6749 22143 6783
rect 25421 6749 25455 6783
rect 25881 6749 25915 6783
rect 28273 6749 28307 6783
rect 33517 6749 33551 6783
rect 35817 6749 35851 6783
rect 6377 6681 6411 6715
rect 26249 6681 26283 6715
rect 27537 6681 27571 6715
rect 32781 6681 32815 6715
rect 2421 6613 2455 6647
rect 3525 6613 3559 6647
rect 6009 6613 6043 6647
rect 7941 6613 7975 6647
rect 8493 6613 8527 6647
rect 12081 6613 12115 6647
rect 12541 6613 12575 6647
rect 17693 6613 17727 6647
rect 19441 6613 19475 6647
rect 22017 6613 22051 6647
rect 23489 6613 23523 6647
rect 24041 6613 24075 6647
rect 24409 6613 24443 6647
rect 24869 6613 24903 6647
rect 26709 6613 26743 6647
rect 29653 6613 29687 6647
rect 32873 6613 32907 6647
rect 35173 6613 35207 6647
rect 35265 6613 35299 6647
rect 36277 6613 36311 6647
rect 2237 6409 2271 6443
rect 3709 6409 3743 6443
rect 4261 6409 4295 6443
rect 4721 6409 4755 6443
rect 7941 6409 7975 6443
rect 10057 6409 10091 6443
rect 11805 6409 11839 6443
rect 13461 6409 13495 6443
rect 13921 6409 13955 6443
rect 17509 6409 17543 6443
rect 19993 6409 20027 6443
rect 21925 6409 21959 6443
rect 23489 6409 23523 6443
rect 24685 6409 24719 6443
rect 25145 6409 25179 6443
rect 25513 6409 25547 6443
rect 29009 6409 29043 6443
rect 32965 6409 32999 6443
rect 33333 6409 33367 6443
rect 33609 6409 33643 6443
rect 35357 6409 35391 6443
rect 6561 6341 6595 6375
rect 9321 6341 9355 6375
rect 27537 6341 27571 6375
rect 35909 6341 35943 6375
rect 1869 6273 1903 6307
rect 7389 6273 7423 6307
rect 10609 6273 10643 6307
rect 10701 6273 10735 6307
rect 13001 6273 13035 6307
rect 14013 6273 14047 6307
rect 17877 6273 17911 6307
rect 18061 6273 18095 6307
rect 21189 6273 21223 6307
rect 21557 6273 21591 6307
rect 22477 6273 22511 6307
rect 22569 6273 22603 6307
rect 24133 6273 24167 6307
rect 24225 6273 24259 6307
rect 25881 6273 25915 6307
rect 26433 6273 26467 6307
rect 26525 6273 26559 6307
rect 27445 6273 27479 6307
rect 27997 6273 28031 6307
rect 28089 6273 28123 6307
rect 35449 6273 35483 6307
rect 2329 6205 2363 6239
rect 2596 6205 2630 6239
rect 5273 6205 5307 6239
rect 5825 6205 5859 6239
rect 7205 6205 7239 6239
rect 8401 6205 8435 6239
rect 9689 6205 9723 6239
rect 10517 6205 10551 6239
rect 12265 6205 12299 6239
rect 24041 6205 24075 6239
rect 27905 6205 27939 6239
rect 29285 6205 29319 6239
rect 29837 6205 29871 6239
rect 6285 6137 6319 6171
rect 12909 6137 12943 6171
rect 14280 6137 14314 6171
rect 16865 6137 16899 6171
rect 18306 6137 18340 6171
rect 22385 6137 22419 6171
rect 23029 6137 23063 6171
rect 30573 6137 30607 6171
rect 5089 6069 5123 6103
rect 5457 6069 5491 6103
rect 6837 6069 6871 6103
rect 7297 6069 7331 6103
rect 8217 6069 8251 6103
rect 8585 6069 8619 6103
rect 10149 6069 10183 6103
rect 11437 6069 11471 6103
rect 12449 6069 12483 6103
rect 12817 6069 12851 6103
rect 15393 6069 15427 6103
rect 16957 6069 16991 6103
rect 19441 6069 19475 6103
rect 22017 6069 22051 6103
rect 23673 6069 23707 6103
rect 25973 6069 26007 6103
rect 26341 6069 26375 6103
rect 26985 6069 27019 6103
rect 28549 6069 28583 6103
rect 29469 6069 29503 6103
rect 30297 6069 30331 6103
rect 4077 5865 4111 5899
rect 4537 5865 4571 5899
rect 6009 5865 6043 5899
rect 6561 5865 6595 5899
rect 7573 5865 7607 5899
rect 8309 5865 8343 5899
rect 10609 5865 10643 5899
rect 11713 5865 11747 5899
rect 12817 5865 12851 5899
rect 13185 5865 13219 5899
rect 14381 5865 14415 5899
rect 16497 5865 16531 5899
rect 17693 5865 17727 5899
rect 22293 5865 22327 5899
rect 23305 5865 23339 5899
rect 23765 5865 23799 5899
rect 23857 5865 23891 5899
rect 25513 5865 25547 5899
rect 26525 5865 26559 5899
rect 27629 5865 27663 5899
rect 27905 5865 27939 5899
rect 30389 5865 30423 5899
rect 30757 5865 30791 5899
rect 35357 5865 35391 5899
rect 1676 5797 1710 5831
rect 4445 5797 4479 5831
rect 6469 5797 6503 5831
rect 10333 5797 10367 5831
rect 12265 5797 12299 5831
rect 16865 5797 16899 5831
rect 17325 5797 17359 5831
rect 18245 5797 18279 5831
rect 28356 5797 28390 5831
rect 1409 5729 1443 5763
rect 6929 5729 6963 5763
rect 8125 5729 8159 5763
rect 9689 5729 9723 5763
rect 10793 5729 10827 5763
rect 12173 5729 12207 5763
rect 13737 5729 13771 5763
rect 15669 5729 15703 5763
rect 18153 5729 18187 5763
rect 18889 5729 18923 5763
rect 21169 5729 21203 5763
rect 25329 5729 25363 5763
rect 26893 5729 26927 5763
rect 30573 5729 30607 5763
rect 4721 5661 4755 5695
rect 7021 5661 7055 5695
rect 7113 5661 7147 5695
rect 12357 5661 12391 5695
rect 13829 5661 13863 5695
rect 14013 5661 14047 5695
rect 15761 5661 15795 5695
rect 15853 5661 15887 5695
rect 18337 5661 18371 5695
rect 19441 5661 19475 5695
rect 20913 5661 20947 5695
rect 24041 5661 24075 5695
rect 25145 5661 25179 5695
rect 26985 5661 27019 5695
rect 27169 5661 27203 5695
rect 28089 5661 28123 5695
rect 32137 5661 32171 5695
rect 3709 5593 3743 5627
rect 9873 5593 9907 5627
rect 14749 5593 14783 5627
rect 23397 5593 23431 5627
rect 2789 5525 2823 5559
rect 3341 5525 3375 5559
rect 5089 5525 5123 5559
rect 5457 5525 5491 5559
rect 7941 5525 7975 5559
rect 11805 5525 11839 5559
rect 13369 5525 13403 5559
rect 15301 5525 15335 5559
rect 17785 5525 17819 5559
rect 19901 5525 19935 5559
rect 22845 5525 22879 5559
rect 24409 5525 24443 5559
rect 24869 5525 24903 5559
rect 26065 5525 26099 5559
rect 29469 5525 29503 5559
rect 30113 5525 30147 5559
rect 31217 5525 31251 5559
rect 31769 5525 31803 5559
rect 1593 5321 1627 5355
rect 1961 5321 1995 5355
rect 3249 5321 3283 5355
rect 4629 5321 4663 5355
rect 5733 5321 5767 5355
rect 6285 5321 6319 5355
rect 10057 5321 10091 5355
rect 11805 5321 11839 5355
rect 12725 5321 12759 5355
rect 15025 5321 15059 5355
rect 15669 5321 15703 5355
rect 15945 5321 15979 5355
rect 17509 5321 17543 5355
rect 18429 5321 18463 5355
rect 19165 5321 19199 5355
rect 20729 5321 20763 5355
rect 21649 5321 21683 5355
rect 23489 5321 23523 5355
rect 25053 5321 25087 5355
rect 27353 5321 27387 5355
rect 28733 5321 28767 5355
rect 31677 5321 31711 5355
rect 6653 5253 6687 5287
rect 22017 5253 22051 5287
rect 23673 5253 23707 5287
rect 25237 5253 25271 5287
rect 26433 5253 26467 5287
rect 27261 5253 27295 5287
rect 31585 5253 31619 5287
rect 2697 5185 2731 5219
rect 5457 5185 5491 5219
rect 7297 5185 7331 5219
rect 7481 5185 7515 5219
rect 12265 5185 12299 5219
rect 13645 5185 13679 5219
rect 13921 5185 13955 5219
rect 16957 5185 16991 5219
rect 19349 5185 19383 5219
rect 22569 5185 22603 5219
rect 24133 5185 24167 5219
rect 24225 5185 24259 5219
rect 25789 5185 25823 5219
rect 27813 5185 27847 5219
rect 27905 5185 27939 5219
rect 32137 5185 32171 5219
rect 32321 5185 32355 5219
rect 3525 5117 3559 5151
rect 3709 5117 3743 5151
rect 4813 5117 4847 5151
rect 7205 5117 7239 5151
rect 8401 5117 8435 5151
rect 9505 5117 9539 5151
rect 10609 5117 10643 5151
rect 11161 5117 11195 5151
rect 13185 5117 13219 5151
rect 18245 5117 18279 5151
rect 21281 5117 21315 5151
rect 22385 5117 22419 5151
rect 25697 5117 25731 5151
rect 26893 5117 26927 5151
rect 27721 5117 27755 5151
rect 29285 5117 29319 5151
rect 29837 5117 29871 5151
rect 30389 5117 30423 5151
rect 32045 5117 32079 5151
rect 2513 5049 2547 5083
rect 4353 5049 4387 5083
rect 10517 5049 10551 5083
rect 16773 5049 16807 5083
rect 19616 5049 19650 5083
rect 24777 5049 24811 5083
rect 25605 5049 25639 5083
rect 2145 4981 2179 5015
rect 2605 4981 2639 5015
rect 3893 4981 3927 5015
rect 4997 4981 5031 5015
rect 6837 4981 6871 5015
rect 8125 4981 8159 5015
rect 8585 4981 8619 5015
rect 9045 4981 9079 5015
rect 9321 4981 9355 5015
rect 9689 4981 9723 5015
rect 10793 4981 10827 5015
rect 13093 4981 13127 5015
rect 13647 4981 13681 5015
rect 16405 4981 16439 5015
rect 16865 4981 16899 5015
rect 17785 4981 17819 5015
rect 18889 4981 18923 5015
rect 22477 4981 22511 5015
rect 23121 4981 23155 5015
rect 24041 4981 24075 5015
rect 28457 4981 28491 5015
rect 29469 4981 29503 5015
rect 30205 4981 30239 5015
rect 30573 4981 30607 5015
rect 30941 4981 30975 5015
rect 32781 4981 32815 5015
rect 33241 4981 33275 5015
rect 3341 4777 3375 4811
rect 6377 4777 6411 4811
rect 7481 4777 7515 4811
rect 8033 4777 8067 4811
rect 9505 4777 9539 4811
rect 10149 4777 10183 4811
rect 11529 4777 11563 4811
rect 14013 4777 14047 4811
rect 14749 4777 14783 4811
rect 15761 4777 15795 4811
rect 16865 4777 16899 4811
rect 17233 4777 17267 4811
rect 19809 4777 19843 4811
rect 20361 4777 20395 4811
rect 21833 4777 21867 4811
rect 25329 4777 25363 4811
rect 25697 4777 25731 4811
rect 27169 4777 27203 4811
rect 30665 4777 30699 4811
rect 32137 4777 32171 4811
rect 33609 4777 33643 4811
rect 35357 4777 35391 4811
rect 1676 4709 1710 4743
rect 4721 4709 4755 4743
rect 7941 4709 7975 4743
rect 12234 4709 12268 4743
rect 16497 4709 16531 4743
rect 19533 4709 19567 4743
rect 23664 4709 23698 4743
rect 31769 4709 31803 4743
rect 1409 4641 1443 4675
rect 4629 4641 4663 4675
rect 5825 4641 5859 4675
rect 6837 4641 6871 4675
rect 6929 4641 6963 4675
rect 8401 4641 8435 4675
rect 8493 4641 8527 4675
rect 10057 4641 10091 4675
rect 11989 4641 12023 4675
rect 15669 4641 15703 4675
rect 17581 4641 17615 4675
rect 22201 4641 22235 4675
rect 27813 4641 27847 4675
rect 27905 4641 27939 4675
rect 29541 4641 29575 4675
rect 32505 4641 32539 4675
rect 32597 4641 32631 4675
rect 33241 4641 33275 4675
rect 34244 4641 34278 4675
rect 4813 4573 4847 4607
rect 8677 4573 8711 4607
rect 10241 4573 10275 4607
rect 14381 4573 14415 4607
rect 15853 4573 15887 4607
rect 17325 4573 17359 4607
rect 22293 4573 22327 4607
rect 22385 4573 22419 4607
rect 23397 4573 23431 4607
rect 27997 4573 28031 4607
rect 29285 4573 29319 4607
rect 32781 4573 32815 4607
rect 33977 4573 34011 4607
rect 6009 4505 6043 4539
rect 15301 4505 15335 4539
rect 22937 4505 22971 4539
rect 26157 4505 26191 4539
rect 28825 4505 28859 4539
rect 2789 4437 2823 4471
rect 3801 4437 3835 4471
rect 4261 4437 4295 4471
rect 5273 4437 5307 4471
rect 5641 4437 5675 4471
rect 7113 4437 7147 4471
rect 9137 4437 9171 4471
rect 9689 4437 9723 4471
rect 11897 4437 11931 4471
rect 13369 4437 13403 4471
rect 15025 4437 15059 4471
rect 18705 4437 18739 4471
rect 21281 4437 21315 4471
rect 21649 4437 21683 4471
rect 23213 4437 23247 4471
rect 24777 4437 24811 4471
rect 26709 4437 26743 4471
rect 27445 4437 27479 4471
rect 28457 4437 28491 4471
rect 31217 4437 31251 4471
rect 2789 4233 2823 4267
rect 6193 4233 6227 4267
rect 11989 4233 12023 4267
rect 16221 4233 16255 4267
rect 17417 4233 17451 4267
rect 17785 4233 17819 4267
rect 18613 4233 18647 4267
rect 22385 4233 22419 4267
rect 23397 4233 23431 4267
rect 26157 4233 26191 4267
rect 27537 4233 27571 4267
rect 27905 4233 27939 4267
rect 25605 4165 25639 4199
rect 5549 4097 5583 4131
rect 5641 4097 5675 4131
rect 7481 4097 7515 4131
rect 17049 4097 17083 4131
rect 18337 4097 18371 4131
rect 19993 4097 20027 4131
rect 22017 4097 22051 4131
rect 26709 4097 26743 4131
rect 29101 4097 29135 4131
rect 30113 4097 30147 4131
rect 31493 4097 31527 4131
rect 33425 4097 33459 4131
rect 1409 4029 1443 4063
rect 1676 4029 1710 4063
rect 3341 4029 3375 4063
rect 3893 4029 3927 4063
rect 6653 4029 6687 4063
rect 7205 4029 7239 4063
rect 8493 4029 8527 4063
rect 8585 4029 8619 4063
rect 11069 4029 11103 4063
rect 12449 4029 12483 4063
rect 13001 4029 13035 4063
rect 13829 4029 13863 4063
rect 14096 4029 14130 4063
rect 16773 4029 16807 4063
rect 18429 4029 18463 4063
rect 19533 4029 19567 4063
rect 20269 4029 20303 4063
rect 22477 4029 22511 4063
rect 23673 4029 23707 4063
rect 23940 4029 23974 4063
rect 26525 4029 26559 4063
rect 27721 4029 27755 4063
rect 29837 4029 29871 4063
rect 31033 4029 31067 4063
rect 31769 4029 31803 4063
rect 7297 3961 7331 3995
rect 8125 3961 8159 3995
rect 8830 3961 8864 3995
rect 10885 3961 10919 3995
rect 13645 3961 13679 3995
rect 16865 3961 16899 3995
rect 26065 3961 26099 3995
rect 28733 3961 28767 3995
rect 3801 3893 3835 3927
rect 4077 3893 4111 3927
rect 4537 3893 4571 3927
rect 4813 3893 4847 3927
rect 5089 3893 5123 3927
rect 5457 3893 5491 3927
rect 6837 3893 6871 3927
rect 9965 3893 9999 3927
rect 10609 3893 10643 3927
rect 11253 3893 11287 3927
rect 11713 3893 11747 3927
rect 12633 3893 12667 3927
rect 15209 3893 15243 3927
rect 15761 3893 15795 3927
rect 16405 3893 16439 3927
rect 19073 3893 19107 3927
rect 19441 3893 19475 3927
rect 19995 3893 20029 3927
rect 21373 3893 21407 3927
rect 22661 3893 22695 3927
rect 23121 3893 23155 3927
rect 25053 3893 25087 3927
rect 26617 3893 26651 3927
rect 28365 3893 28399 3927
rect 29469 3893 29503 3927
rect 29929 3893 29963 3927
rect 30481 3893 30515 3927
rect 30941 3893 30975 3927
rect 31495 3893 31529 3927
rect 32873 3893 32907 3927
rect 33977 3893 34011 3927
rect 34437 3893 34471 3927
rect 3801 3689 3835 3723
rect 4537 3689 4571 3723
rect 9045 3689 9079 3723
rect 9505 3689 9539 3723
rect 9689 3689 9723 3723
rect 10241 3689 10275 3723
rect 12081 3689 12115 3723
rect 12633 3689 12667 3723
rect 13185 3689 13219 3723
rect 13553 3689 13587 3723
rect 14565 3689 14599 3723
rect 14933 3689 14967 3723
rect 15577 3689 15611 3723
rect 16221 3689 16255 3723
rect 16313 3689 16347 3723
rect 17233 3689 17267 3723
rect 19257 3689 19291 3723
rect 19809 3689 19843 3723
rect 20637 3689 20671 3723
rect 21281 3689 21315 3723
rect 23213 3689 23247 3723
rect 26249 3689 26283 3723
rect 27997 3689 28031 3723
rect 28365 3689 28399 3723
rect 29377 3689 29411 3723
rect 31493 3689 31527 3723
rect 31953 3689 31987 3723
rect 32321 3689 32355 3723
rect 32689 3689 32723 3723
rect 34621 3689 34655 3723
rect 1768 3621 1802 3655
rect 10517 3621 10551 3655
rect 14289 3621 14323 3655
rect 16957 3621 16991 3655
rect 23550 3621 23584 3655
rect 25237 3621 25271 3655
rect 29828 3621 29862 3655
rect 33149 3621 33183 3655
rect 1501 3553 1535 3587
rect 4445 3553 4479 3587
rect 5457 3553 5491 3587
rect 5917 3553 5951 3587
rect 6276 3553 6310 3587
rect 8493 3553 8527 3587
rect 10701 3553 10735 3587
rect 10957 3553 10991 3587
rect 17417 3553 17451 3587
rect 17740 3553 17774 3587
rect 21373 3553 21407 3587
rect 23305 3553 23339 3587
rect 26525 3553 26559 3587
rect 26709 3553 26743 3587
rect 27169 3553 27203 3587
rect 27905 3553 27939 3587
rect 29561 3553 29595 3587
rect 32137 3553 32171 3587
rect 33508 3553 33542 3587
rect 35173 3553 35207 3587
rect 4721 3485 4755 3519
rect 6009 3485 6043 3519
rect 13645 3485 13679 3519
rect 13829 3485 13863 3519
rect 16497 3485 16531 3519
rect 17877 3485 17911 3519
rect 18153 3485 18187 3519
rect 21465 3485 21499 3519
rect 22385 3485 22419 3519
rect 28457 3485 28491 3519
rect 28641 3485 28675 3519
rect 33241 3485 33275 3519
rect 4077 3417 4111 3451
rect 20269 3417 20303 3451
rect 22017 3417 22051 3451
rect 26893 3417 26927 3451
rect 2881 3349 2915 3383
rect 3433 3349 3467 3383
rect 5181 3349 5215 3383
rect 7389 3349 7423 3383
rect 8033 3349 8067 3383
rect 8309 3349 8343 3383
rect 8677 3349 8711 3383
rect 13001 3349 13035 3383
rect 15853 3349 15887 3383
rect 20913 3349 20947 3383
rect 22661 3349 22695 3383
rect 24685 3349 24719 3383
rect 25605 3349 25639 3383
rect 30941 3349 30975 3383
rect 35541 3349 35575 3383
rect 1593 3145 1627 3179
rect 5641 3145 5675 3179
rect 8309 3145 8343 3179
rect 10793 3145 10827 3179
rect 11437 3145 11471 3179
rect 12633 3145 12667 3179
rect 13461 3145 13495 3179
rect 15761 3145 15795 3179
rect 16313 3145 16347 3179
rect 16681 3145 16715 3179
rect 17049 3145 17083 3179
rect 17509 3145 17543 3179
rect 17877 3145 17911 3179
rect 18429 3145 18463 3179
rect 19165 3145 19199 3179
rect 21557 3145 21591 3179
rect 21649 3145 21683 3179
rect 25053 3145 25087 3179
rect 26525 3145 26559 3179
rect 27997 3145 28031 3179
rect 31033 3145 31067 3179
rect 33885 3145 33919 3179
rect 34253 3145 34287 3179
rect 34621 3145 34655 3179
rect 6193 3077 6227 3111
rect 6561 3077 6595 3111
rect 21373 3077 21407 3111
rect 1777 3009 1811 3043
rect 13829 3009 13863 3043
rect 14244 3009 14278 3043
rect 14381 3009 14415 3043
rect 14657 3009 14691 3043
rect 18889 3009 18923 3043
rect 19349 3009 19383 3043
rect 28641 3077 28675 3111
rect 22477 3009 22511 3043
rect 30021 3009 30055 3043
rect 30113 3009 30147 3043
rect 31448 3009 31482 3043
rect 31585 3009 31619 3043
rect 31861 3009 31895 3043
rect 32965 3009 32999 3043
rect 35357 3009 35391 3043
rect 35449 3009 35483 3043
rect 35909 3009 35943 3043
rect 4169 2941 4203 2975
rect 4261 2941 4295 2975
rect 4528 2941 4562 2975
rect 6929 2941 6963 2975
rect 7196 2941 7230 2975
rect 8953 2941 8987 2975
rect 9321 2941 9355 2975
rect 9413 2941 9447 2975
rect 9680 2941 9714 2975
rect 12449 2941 12483 2975
rect 13921 2941 13955 2975
rect 16865 2941 16899 2975
rect 18245 2941 18279 2975
rect 19616 2941 19650 2975
rect 21557 2941 21591 2975
rect 22201 2941 22235 2975
rect 22293 2941 22327 2975
rect 23121 2941 23155 2975
rect 23489 2941 23523 2975
rect 23673 2941 23707 2975
rect 26157 2941 26191 2975
rect 26624 2941 26658 2975
rect 26884 2941 26918 2975
rect 31125 2941 31159 2975
rect 35265 2941 35299 2975
rect 2044 2873 2078 2907
rect 11713 2873 11747 2907
rect 23918 2873 23952 2907
rect 25789 2873 25823 2907
rect 29101 2873 29135 2907
rect 29929 2873 29963 2907
rect 30573 2873 30607 2907
rect 3157 2805 3191 2839
rect 3709 2805 3743 2839
rect 12265 2805 12299 2839
rect 13093 2805 13127 2839
rect 20729 2805 20763 2839
rect 21833 2805 21867 2839
rect 29561 2805 29595 2839
rect 33609 2805 33643 2839
rect 34897 2805 34931 2839
rect 1777 2601 1811 2635
rect 2145 2601 2179 2635
rect 2421 2601 2455 2635
rect 2881 2601 2915 2635
rect 3433 2601 3467 2635
rect 5457 2601 5491 2635
rect 6929 2601 6963 2635
rect 7297 2601 7331 2635
rect 8309 2601 8343 2635
rect 8861 2601 8895 2635
rect 10333 2601 10367 2635
rect 10885 2601 10919 2635
rect 11253 2601 11287 2635
rect 14289 2601 14323 2635
rect 16865 2601 16899 2635
rect 17509 2601 17543 2635
rect 18153 2601 18187 2635
rect 19993 2601 20027 2635
rect 20913 2601 20947 2635
rect 22569 2601 22603 2635
rect 23121 2601 23155 2635
rect 23765 2601 23799 2635
rect 25697 2601 25731 2635
rect 26249 2601 26283 2635
rect 26617 2601 26651 2635
rect 28549 2601 28583 2635
rect 31401 2601 31435 2635
rect 34161 2601 34195 2635
rect 34805 2601 34839 2635
rect 35173 2601 35207 2635
rect 35449 2601 35483 2635
rect 37013 2601 37047 2635
rect 6009 2533 6043 2567
rect 8677 2533 8711 2567
rect 9597 2533 9631 2567
rect 10241 2533 10275 2567
rect 13154 2533 13188 2567
rect 18880 2533 18914 2567
rect 20637 2533 20671 2567
rect 21434 2533 21468 2567
rect 24584 2533 24618 2567
rect 27436 2533 27470 2567
rect 30266 2533 30300 2567
rect 33048 2533 33082 2567
rect 2789 2465 2823 2499
rect 4344 2465 4378 2499
rect 6377 2465 6411 2499
rect 7389 2465 7423 2499
rect 7941 2465 7975 2499
rect 8493 2465 8527 2499
rect 11437 2465 11471 2499
rect 12081 2465 12115 2499
rect 15301 2465 15335 2499
rect 15485 2465 15519 2499
rect 15741 2465 15775 2499
rect 18613 2465 18647 2499
rect 21189 2465 21223 2499
rect 24317 2465 24351 2499
rect 27169 2465 27203 2499
rect 29561 2465 29595 2499
rect 30021 2465 30055 2499
rect 32413 2465 32447 2499
rect 32781 2465 32815 2499
rect 35817 2465 35851 2499
rect 3065 2397 3099 2431
rect 4077 2397 4111 2431
rect 7573 2397 7607 2431
rect 9229 2397 9263 2431
rect 10517 2397 10551 2431
rect 12449 2397 12483 2431
rect 12909 2397 12943 2431
rect 14933 2397 14967 2431
rect 35909 2397 35943 2431
rect 36093 2397 36127 2431
rect 36553 2397 36587 2431
rect 36829 2397 36863 2431
rect 3801 2329 3835 2363
rect 9873 2329 9907 2363
rect 29193 2329 29227 2363
rect 11621 2261 11655 2295
rect 31953 2261 31987 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 38824 37562
rect 1104 37488 38824 37510
rect 1104 37018 38824 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 38824 37018
rect 1104 36944 38824 36966
rect 1104 36474 38824 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 38824 36474
rect 1104 36400 38824 36422
rect 1104 35930 38824 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 38824 35930
rect 1104 35856 38824 35878
rect 35618 35816 35624 35828
rect 35579 35788 35624 35816
rect 35618 35776 35624 35788
rect 35676 35776 35682 35828
rect 30193 35615 30251 35621
rect 30193 35612 30205 35615
rect 30024 35584 30205 35612
rect 30024 35488 30052 35584
rect 30193 35581 30205 35584
rect 30239 35581 30251 35615
rect 35434 35612 35440 35624
rect 35395 35584 35440 35612
rect 30193 35575 30251 35581
rect 35434 35572 35440 35584
rect 35492 35612 35498 35624
rect 35989 35615 36047 35621
rect 35989 35612 36001 35615
rect 35492 35584 36001 35612
rect 35492 35572 35498 35584
rect 35989 35581 36001 35584
rect 36035 35581 36047 35615
rect 35989 35575 36047 35581
rect 30466 35553 30472 35556
rect 30460 35544 30472 35553
rect 30427 35516 30472 35544
rect 30460 35507 30472 35516
rect 30466 35504 30472 35507
rect 30524 35504 30530 35556
rect 30006 35476 30012 35488
rect 29967 35448 30012 35476
rect 30006 35436 30012 35448
rect 30064 35436 30070 35488
rect 30834 35436 30840 35488
rect 30892 35476 30898 35488
rect 31573 35479 31631 35485
rect 31573 35476 31585 35479
rect 30892 35448 31585 35476
rect 30892 35436 30898 35448
rect 31573 35445 31585 35448
rect 31619 35445 31631 35479
rect 31573 35439 31631 35445
rect 1104 35386 38824 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 38824 35386
rect 1104 35312 38824 35334
rect 29917 35275 29975 35281
rect 29917 35241 29929 35275
rect 29963 35272 29975 35275
rect 30282 35272 30288 35284
rect 29963 35244 30288 35272
rect 29963 35241 29975 35244
rect 29917 35235 29975 35241
rect 30282 35232 30288 35244
rect 30340 35272 30346 35284
rect 30834 35272 30840 35284
rect 30340 35244 30840 35272
rect 30340 35232 30346 35244
rect 30834 35232 30840 35244
rect 30892 35232 30898 35284
rect 36170 35272 36176 35284
rect 36131 35244 36176 35272
rect 36170 35232 36176 35244
rect 36228 35232 36234 35284
rect 30285 35139 30343 35145
rect 30285 35105 30297 35139
rect 30331 35136 30343 35139
rect 30466 35136 30472 35148
rect 30331 35108 30472 35136
rect 30331 35105 30343 35108
rect 30285 35099 30343 35105
rect 30466 35096 30472 35108
rect 30524 35136 30530 35148
rect 30929 35139 30987 35145
rect 30929 35136 30941 35139
rect 30524 35108 30941 35136
rect 30524 35096 30530 35108
rect 30929 35105 30941 35108
rect 30975 35136 30987 35139
rect 32030 35136 32036 35148
rect 30975 35108 32036 35136
rect 30975 35105 30987 35108
rect 30929 35099 30987 35105
rect 32030 35096 32036 35108
rect 32088 35096 32094 35148
rect 34333 35139 34391 35145
rect 34333 35105 34345 35139
rect 34379 35136 34391 35139
rect 34698 35136 34704 35148
rect 34379 35108 34704 35136
rect 34379 35105 34391 35108
rect 34333 35099 34391 35105
rect 34698 35096 34704 35108
rect 34756 35136 34762 35148
rect 34793 35139 34851 35145
rect 34793 35136 34805 35139
rect 34756 35108 34805 35136
rect 34756 35096 34762 35108
rect 34793 35105 34805 35108
rect 34839 35105 34851 35139
rect 34793 35099 34851 35105
rect 35989 35139 36047 35145
rect 35989 35105 36001 35139
rect 36035 35136 36047 35139
rect 36170 35136 36176 35148
rect 36035 35108 36176 35136
rect 36035 35105 36047 35108
rect 35989 35099 36047 35105
rect 36170 35096 36176 35108
rect 36228 35096 36234 35148
rect 29086 35028 29092 35080
rect 29144 35068 29150 35080
rect 31113 35071 31171 35077
rect 31113 35068 31125 35071
rect 29144 35040 31125 35068
rect 29144 35028 29150 35040
rect 31113 35037 31125 35040
rect 31159 35068 31171 35071
rect 32766 35068 32772 35080
rect 31159 35040 32772 35068
rect 31159 35037 31171 35040
rect 31113 35031 31171 35037
rect 32766 35028 32772 35040
rect 32824 35028 32830 35080
rect 34885 35071 34943 35077
rect 34885 35037 34897 35071
rect 34931 35037 34943 35071
rect 34885 35031 34943 35037
rect 34977 35071 35035 35077
rect 34977 35037 34989 35071
rect 35023 35037 35035 35071
rect 34977 35031 35035 35037
rect 34790 34960 34796 35012
rect 34848 35000 34854 35012
rect 34900 35000 34928 35031
rect 34848 34972 34928 35000
rect 34848 34960 34854 34972
rect 30469 34935 30527 34941
rect 30469 34901 30481 34935
rect 30515 34932 30527 34935
rect 31662 34932 31668 34944
rect 30515 34904 31668 34932
rect 30515 34901 30527 34904
rect 30469 34895 30527 34901
rect 31662 34892 31668 34904
rect 31720 34892 31726 34944
rect 33318 34932 33324 34944
rect 33279 34904 33324 34932
rect 33318 34892 33324 34904
rect 33376 34892 33382 34944
rect 33686 34892 33692 34944
rect 33744 34932 33750 34944
rect 34425 34935 34483 34941
rect 34425 34932 34437 34935
rect 33744 34904 34437 34932
rect 33744 34892 33750 34904
rect 34425 34901 34437 34904
rect 34471 34901 34483 34935
rect 34425 34895 34483 34901
rect 34514 34892 34520 34944
rect 34572 34932 34578 34944
rect 34992 34932 35020 35031
rect 35526 34932 35532 34944
rect 34572 34904 35020 34932
rect 35487 34904 35532 34932
rect 34572 34892 34578 34904
rect 35526 34892 35532 34904
rect 35584 34892 35590 34944
rect 1104 34842 38824 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 38824 34842
rect 1104 34768 38824 34790
rect 29086 34728 29092 34740
rect 29047 34700 29092 34728
rect 29086 34688 29092 34700
rect 29144 34688 29150 34740
rect 30374 34688 30380 34740
rect 30432 34728 30438 34740
rect 31389 34731 31447 34737
rect 31389 34728 31401 34731
rect 30432 34700 31401 34728
rect 30432 34688 30438 34700
rect 31389 34697 31401 34700
rect 31435 34697 31447 34731
rect 32766 34728 32772 34740
rect 32679 34700 32772 34728
rect 31389 34691 31447 34697
rect 32766 34688 32772 34700
rect 32824 34728 32830 34740
rect 33134 34728 33140 34740
rect 32824 34700 33140 34728
rect 32824 34688 32830 34700
rect 33134 34688 33140 34700
rect 33192 34728 33198 34740
rect 34146 34728 34152 34740
rect 33192 34700 34152 34728
rect 33192 34688 33198 34700
rect 34146 34688 34152 34700
rect 34204 34688 34210 34740
rect 34333 34731 34391 34737
rect 34333 34697 34345 34731
rect 34379 34728 34391 34731
rect 34790 34728 34796 34740
rect 34379 34700 34796 34728
rect 34379 34697 34391 34700
rect 34333 34691 34391 34697
rect 34790 34688 34796 34700
rect 34848 34688 34854 34740
rect 37550 34728 37556 34740
rect 37511 34700 37556 34728
rect 37550 34688 37556 34700
rect 37608 34688 37614 34740
rect 32030 34660 32036 34672
rect 31991 34632 32036 34660
rect 32030 34620 32036 34632
rect 32088 34620 32094 34672
rect 34422 34660 34428 34672
rect 33704 34632 34428 34660
rect 33704 34601 33732 34632
rect 34422 34620 34428 34632
rect 34480 34620 34486 34672
rect 36262 34660 36268 34672
rect 36223 34632 36268 34660
rect 36262 34620 36268 34632
rect 36320 34620 36326 34672
rect 29549 34595 29607 34601
rect 29549 34561 29561 34595
rect 29595 34592 29607 34595
rect 33137 34595 33195 34601
rect 29595 34564 30144 34592
rect 29595 34561 29607 34564
rect 29549 34555 29607 34561
rect 30006 34524 30012 34536
rect 29840 34496 30012 34524
rect 29362 34348 29368 34400
rect 29420 34388 29426 34400
rect 29840 34397 29868 34496
rect 30006 34484 30012 34496
rect 30064 34484 30070 34536
rect 30116 34524 30144 34564
rect 33137 34561 33149 34595
rect 33183 34592 33195 34595
rect 33689 34595 33747 34601
rect 33689 34592 33701 34595
rect 33183 34564 33701 34592
rect 33183 34561 33195 34564
rect 33137 34555 33195 34561
rect 33689 34561 33701 34564
rect 33735 34561 33747 34595
rect 33689 34555 33747 34561
rect 33873 34595 33931 34601
rect 33873 34561 33885 34595
rect 33919 34592 33931 34595
rect 34146 34592 34152 34604
rect 33919 34564 34152 34592
rect 33919 34561 33931 34564
rect 33873 34555 33931 34561
rect 34146 34552 34152 34564
rect 34204 34592 34210 34604
rect 34514 34592 34520 34604
rect 34204 34564 34520 34592
rect 34204 34552 34210 34564
rect 34514 34552 34520 34564
rect 34572 34552 34578 34604
rect 34808 34564 35020 34592
rect 30282 34533 30288 34536
rect 30276 34524 30288 34533
rect 30116 34496 30288 34524
rect 30276 34487 30288 34496
rect 30282 34484 30288 34487
rect 30340 34484 30346 34536
rect 33318 34484 33324 34536
rect 33376 34524 33382 34536
rect 33597 34527 33655 34533
rect 33597 34524 33609 34527
rect 33376 34496 33609 34524
rect 33376 34484 33382 34496
rect 33597 34493 33609 34496
rect 33643 34524 33655 34527
rect 34808 34524 34836 34564
rect 33643 34496 34836 34524
rect 34885 34527 34943 34533
rect 33643 34493 33655 34496
rect 33597 34487 33655 34493
rect 34885 34493 34897 34527
rect 34931 34493 34943 34527
rect 34992 34524 35020 34564
rect 35141 34527 35199 34533
rect 35141 34524 35153 34527
rect 34992 34496 35153 34524
rect 34885 34487 34943 34493
rect 35141 34493 35153 34496
rect 35187 34524 35199 34527
rect 35526 34524 35532 34536
rect 35187 34496 35532 34524
rect 35187 34493 35199 34496
rect 35141 34487 35199 34493
rect 34900 34456 34928 34487
rect 35526 34484 35532 34496
rect 35584 34524 35590 34536
rect 35894 34524 35900 34536
rect 35584 34496 35900 34524
rect 35584 34484 35590 34496
rect 35894 34484 35900 34496
rect 35952 34484 35958 34536
rect 36170 34484 36176 34536
rect 36228 34524 36234 34536
rect 36817 34527 36875 34533
rect 36817 34524 36829 34527
rect 36228 34496 36829 34524
rect 36228 34484 36234 34496
rect 36817 34493 36829 34496
rect 36863 34493 36875 34527
rect 36817 34487 36875 34493
rect 37369 34527 37427 34533
rect 37369 34493 37381 34527
rect 37415 34524 37427 34527
rect 37918 34524 37924 34536
rect 37415 34496 37924 34524
rect 37415 34493 37427 34496
rect 37369 34487 37427 34493
rect 37918 34484 37924 34496
rect 37976 34484 37982 34536
rect 34624 34428 34928 34456
rect 34624 34400 34652 34428
rect 29825 34391 29883 34397
rect 29825 34388 29837 34391
rect 29420 34360 29837 34388
rect 29420 34348 29426 34360
rect 29825 34357 29837 34360
rect 29871 34357 29883 34391
rect 33226 34388 33232 34400
rect 33187 34360 33232 34388
rect 29825 34351 29883 34357
rect 33226 34348 33232 34360
rect 33284 34348 33290 34400
rect 34606 34388 34612 34400
rect 34567 34360 34612 34388
rect 34606 34348 34612 34360
rect 34664 34348 34670 34400
rect 1104 34298 38824 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 38824 34298
rect 1104 34224 38824 34246
rect 27706 34144 27712 34196
rect 27764 34184 27770 34196
rect 28353 34187 28411 34193
rect 28353 34184 28365 34187
rect 27764 34156 28365 34184
rect 27764 34144 27770 34156
rect 28353 34153 28365 34156
rect 28399 34184 28411 34187
rect 29730 34184 29736 34196
rect 28399 34156 29736 34184
rect 28399 34153 28411 34156
rect 28353 34147 28411 34153
rect 29730 34144 29736 34156
rect 29788 34144 29794 34196
rect 34146 34184 34152 34196
rect 34107 34156 34152 34184
rect 34146 34144 34152 34156
rect 34204 34144 34210 34196
rect 35894 34144 35900 34196
rect 35952 34184 35958 34196
rect 36081 34187 36139 34193
rect 36081 34184 36093 34187
rect 35952 34156 36093 34184
rect 35952 34144 35958 34156
rect 36081 34153 36093 34156
rect 36127 34153 36139 34187
rect 36081 34147 36139 34153
rect 34514 34076 34520 34128
rect 34572 34116 34578 34128
rect 34946 34119 35004 34125
rect 34946 34116 34958 34119
rect 34572 34088 34958 34116
rect 34572 34076 34578 34088
rect 34946 34085 34958 34088
rect 34992 34116 35004 34119
rect 36262 34116 36268 34128
rect 34992 34088 36268 34116
rect 34992 34085 35004 34088
rect 34946 34079 35004 34085
rect 36262 34076 36268 34088
rect 36320 34076 36326 34128
rect 28445 34051 28503 34057
rect 28445 34017 28457 34051
rect 28491 34048 28503 34051
rect 28718 34048 28724 34060
rect 28491 34020 28724 34048
rect 28491 34017 28503 34020
rect 28445 34011 28503 34017
rect 28718 34008 28724 34020
rect 28776 34048 28782 34060
rect 29816 34051 29874 34057
rect 29816 34048 29828 34051
rect 28776 34020 29828 34048
rect 28776 34008 28782 34020
rect 29816 34017 29828 34020
rect 29862 34048 29874 34051
rect 30282 34048 30288 34060
rect 29862 34020 30288 34048
rect 29862 34017 29874 34020
rect 29816 34011 29874 34017
rect 30282 34008 30288 34020
rect 30340 34008 30346 34060
rect 31570 34008 31576 34060
rect 31628 34048 31634 34060
rect 32381 34051 32439 34057
rect 32381 34048 32393 34051
rect 31628 34020 32393 34048
rect 31628 34008 31634 34020
rect 32381 34017 32393 34020
rect 32427 34017 32439 34051
rect 32381 34011 32439 34017
rect 28629 33983 28687 33989
rect 28629 33949 28641 33983
rect 28675 33980 28687 33983
rect 28902 33980 28908 33992
rect 28675 33952 28908 33980
rect 28675 33949 28687 33952
rect 28629 33943 28687 33949
rect 28902 33940 28908 33952
rect 28960 33940 28966 33992
rect 29362 33940 29368 33992
rect 29420 33980 29426 33992
rect 29549 33983 29607 33989
rect 29549 33980 29561 33983
rect 29420 33952 29561 33980
rect 29420 33940 29426 33952
rect 29549 33949 29561 33952
rect 29595 33949 29607 33983
rect 32122 33980 32128 33992
rect 32083 33952 32128 33980
rect 29549 33943 29607 33949
rect 32122 33940 32128 33952
rect 32180 33940 32186 33992
rect 34606 33940 34612 33992
rect 34664 33980 34670 33992
rect 34701 33983 34759 33989
rect 34701 33980 34713 33983
rect 34664 33952 34713 33980
rect 34664 33940 34670 33952
rect 34701 33949 34713 33952
rect 34747 33949 34759 33983
rect 34701 33943 34759 33949
rect 27982 33844 27988 33856
rect 27943 33816 27988 33844
rect 27982 33804 27988 33816
rect 28040 33804 28046 33856
rect 30926 33844 30932 33856
rect 30887 33816 30932 33844
rect 30926 33804 30932 33816
rect 30984 33804 30990 33856
rect 31941 33847 31999 33853
rect 31941 33813 31953 33847
rect 31987 33844 31999 33847
rect 32766 33844 32772 33856
rect 31987 33816 32772 33844
rect 31987 33813 31999 33816
rect 31941 33807 31999 33813
rect 32766 33804 32772 33816
rect 32824 33804 32830 33856
rect 33502 33844 33508 33856
rect 33463 33816 33508 33844
rect 33502 33804 33508 33816
rect 33560 33804 33566 33856
rect 34609 33847 34667 33853
rect 34609 33813 34621 33847
rect 34655 33844 34667 33847
rect 34698 33844 34704 33856
rect 34655 33816 34704 33844
rect 34655 33813 34667 33816
rect 34609 33807 34667 33813
rect 34698 33804 34704 33816
rect 34756 33804 34762 33856
rect 1104 33754 38824 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 34966 33754
rect 35018 33702 35030 33754
rect 35082 33702 35094 33754
rect 35146 33702 35158 33754
rect 35210 33702 38824 33754
rect 1104 33680 38824 33702
rect 27706 33640 27712 33652
rect 27667 33612 27712 33640
rect 27706 33600 27712 33612
rect 27764 33600 27770 33652
rect 28077 33643 28135 33649
rect 28077 33609 28089 33643
rect 28123 33640 28135 33643
rect 28718 33640 28724 33652
rect 28123 33612 28724 33640
rect 28123 33609 28135 33612
rect 28077 33603 28135 33609
rect 28718 33600 28724 33612
rect 28776 33600 28782 33652
rect 31757 33643 31815 33649
rect 31757 33609 31769 33643
rect 31803 33640 31815 33643
rect 32033 33643 32091 33649
rect 32033 33640 32045 33643
rect 31803 33612 32045 33640
rect 31803 33609 31815 33612
rect 31757 33603 31815 33609
rect 32033 33609 32045 33612
rect 32079 33640 32091 33643
rect 32122 33640 32128 33652
rect 32079 33612 32128 33640
rect 32079 33609 32091 33612
rect 32033 33603 32091 33609
rect 32122 33600 32128 33612
rect 32180 33600 32186 33652
rect 33870 33640 33876 33652
rect 33831 33612 33876 33640
rect 33870 33600 33876 33612
rect 33928 33600 33934 33652
rect 36262 33640 36268 33652
rect 36223 33612 36268 33640
rect 36262 33600 36268 33612
rect 36320 33600 36326 33652
rect 32140 33572 32168 33600
rect 34238 33572 34244 33584
rect 32140 33544 34244 33572
rect 34238 33532 34244 33544
rect 34296 33572 34302 33584
rect 34606 33572 34612 33584
rect 34296 33544 34612 33572
rect 34296 33532 34302 33544
rect 34606 33532 34612 33544
rect 34664 33572 34670 33584
rect 34664 33544 34928 33572
rect 34664 33532 34670 33544
rect 31754 33464 31760 33516
rect 31812 33504 31818 33516
rect 32585 33507 32643 33513
rect 32585 33504 32597 33507
rect 31812 33476 32597 33504
rect 31812 33464 31818 33476
rect 32585 33473 32597 33476
rect 32631 33473 32643 33507
rect 32766 33504 32772 33516
rect 32727 33476 32772 33504
rect 32585 33467 32643 33473
rect 29641 33439 29699 33445
rect 29641 33436 29653 33439
rect 29472 33408 29653 33436
rect 29472 33368 29500 33408
rect 29641 33405 29653 33408
rect 29687 33405 29699 33439
rect 29641 33399 29699 33405
rect 29730 33396 29736 33448
rect 29788 33436 29794 33448
rect 29908 33439 29966 33445
rect 29908 33436 29920 33439
rect 29788 33408 29920 33436
rect 29788 33396 29794 33408
rect 29908 33405 29920 33408
rect 29954 33436 29966 33439
rect 30926 33436 30932 33448
rect 29954 33408 30932 33436
rect 29954 33405 29966 33408
rect 29908 33399 29966 33405
rect 30926 33396 30932 33408
rect 30984 33396 30990 33448
rect 32600 33436 32628 33467
rect 32766 33464 32772 33476
rect 32824 33464 32830 33516
rect 34900 33513 34928 33544
rect 34885 33507 34943 33513
rect 34885 33473 34897 33507
rect 34931 33473 34943 33507
rect 34885 33467 34943 33473
rect 33137 33439 33195 33445
rect 33137 33436 33149 33439
rect 32600 33408 33149 33436
rect 33137 33405 33149 33408
rect 33183 33405 33195 33439
rect 33137 33399 33195 33405
rect 33689 33439 33747 33445
rect 33689 33405 33701 33439
rect 33735 33405 33747 33439
rect 33689 33399 33747 33405
rect 31757 33371 31815 33377
rect 31757 33368 31769 33371
rect 29472 33340 31769 33368
rect 29089 33303 29147 33309
rect 29089 33269 29101 33303
rect 29135 33300 29147 33303
rect 29362 33300 29368 33312
rect 29135 33272 29368 33300
rect 29135 33269 29147 33272
rect 29089 33263 29147 33269
rect 29362 33260 29368 33272
rect 29420 33300 29426 33312
rect 29472 33309 29500 33340
rect 31757 33337 31769 33340
rect 31803 33337 31815 33371
rect 31757 33331 31815 33337
rect 31846 33328 31852 33380
rect 31904 33368 31910 33380
rect 32493 33371 32551 33377
rect 32493 33368 32505 33371
rect 31904 33340 32505 33368
rect 31904 33328 31910 33340
rect 32493 33337 32505 33340
rect 32539 33337 32551 33371
rect 32493 33331 32551 33337
rect 29457 33303 29515 33309
rect 29457 33300 29469 33303
rect 29420 33272 29469 33300
rect 29420 33260 29426 33272
rect 29457 33269 29469 33272
rect 29503 33269 29515 33303
rect 29457 33263 29515 33269
rect 30466 33260 30472 33312
rect 30524 33300 30530 33312
rect 31021 33303 31079 33309
rect 31021 33300 31033 33303
rect 30524 33272 31033 33300
rect 30524 33260 30530 33272
rect 31021 33269 31033 33272
rect 31067 33300 31079 33303
rect 31570 33300 31576 33312
rect 31067 33272 31576 33300
rect 31067 33269 31079 33272
rect 31021 33263 31079 33269
rect 31570 33260 31576 33272
rect 31628 33260 31634 33312
rect 32122 33300 32128 33312
rect 32083 33272 32128 33300
rect 32122 33260 32128 33272
rect 32180 33260 32186 33312
rect 33597 33303 33655 33309
rect 33597 33269 33609 33303
rect 33643 33300 33655 33303
rect 33704 33300 33732 33399
rect 34698 33328 34704 33380
rect 34756 33368 34762 33380
rect 35152 33371 35210 33377
rect 35152 33368 35164 33371
rect 34756 33340 35164 33368
rect 34756 33328 34762 33340
rect 35152 33337 35164 33340
rect 35198 33368 35210 33371
rect 35802 33368 35808 33380
rect 35198 33340 35808 33368
rect 35198 33337 35210 33340
rect 35152 33331 35210 33337
rect 35802 33328 35808 33340
rect 35860 33328 35866 33380
rect 34790 33300 34796 33312
rect 33643 33272 34796 33300
rect 33643 33269 33655 33272
rect 33597 33263 33655 33269
rect 34790 33260 34796 33272
rect 34848 33260 34854 33312
rect 1104 33210 38824 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 38824 33210
rect 1104 33136 38824 33158
rect 28077 33099 28135 33105
rect 28077 33065 28089 33099
rect 28123 33096 28135 33099
rect 28902 33096 28908 33108
rect 28123 33068 28908 33096
rect 28123 33065 28135 33068
rect 28077 33059 28135 33065
rect 28902 33056 28908 33068
rect 28960 33056 28966 33108
rect 29457 33099 29515 33105
rect 29457 33065 29469 33099
rect 29503 33096 29515 33099
rect 29730 33096 29736 33108
rect 29503 33068 29736 33096
rect 29503 33065 29515 33068
rect 29457 33059 29515 33065
rect 29730 33056 29736 33068
rect 29788 33056 29794 33108
rect 31846 33096 31852 33108
rect 31807 33068 31852 33096
rect 31846 33056 31852 33068
rect 31904 33056 31910 33108
rect 33226 33096 33232 33108
rect 33187 33068 33232 33096
rect 33226 33056 33232 33068
rect 33284 33056 33290 33108
rect 34241 33099 34299 33105
rect 34241 33065 34253 33099
rect 34287 33096 34299 33099
rect 34330 33096 34336 33108
rect 34287 33068 34336 33096
rect 34287 33065 34299 33068
rect 34241 33059 34299 33065
rect 34330 33056 34336 33068
rect 34388 33056 34394 33108
rect 35802 33056 35808 33108
rect 35860 33096 35866 33108
rect 36081 33099 36139 33105
rect 36081 33096 36093 33099
rect 35860 33068 36093 33096
rect 35860 33056 35866 33068
rect 36081 33065 36093 33068
rect 36127 33065 36139 33099
rect 36081 33059 36139 33065
rect 29822 33037 29828 33040
rect 29816 33028 29828 33037
rect 29783 33000 29828 33028
rect 29816 32991 29828 33000
rect 29822 32988 29828 32991
rect 29880 32988 29886 33040
rect 34882 32988 34888 33040
rect 34940 32988 34946 33040
rect 32030 32920 32036 32972
rect 32088 32960 32094 32972
rect 32493 32963 32551 32969
rect 32493 32960 32505 32963
rect 32088 32932 32505 32960
rect 32088 32920 32094 32932
rect 32493 32929 32505 32932
rect 32539 32929 32551 32963
rect 32493 32923 32551 32929
rect 34609 32963 34667 32969
rect 34609 32929 34621 32963
rect 34655 32960 34667 32963
rect 34900 32960 34928 32988
rect 34968 32963 35026 32969
rect 34968 32960 34980 32963
rect 34655 32932 34980 32960
rect 34655 32929 34667 32932
rect 34609 32923 34667 32929
rect 34968 32929 34980 32932
rect 35014 32960 35026 32963
rect 36262 32960 36268 32972
rect 35014 32932 36268 32960
rect 35014 32929 35026 32932
rect 34968 32923 35026 32929
rect 36262 32920 36268 32932
rect 36320 32920 36326 32972
rect 29362 32852 29368 32904
rect 29420 32892 29426 32904
rect 29549 32895 29607 32901
rect 29549 32892 29561 32895
rect 29420 32864 29561 32892
rect 29420 32852 29426 32864
rect 29549 32861 29561 32864
rect 29595 32861 29607 32895
rect 32582 32892 32588 32904
rect 32543 32864 32588 32892
rect 29549 32855 29607 32861
rect 32582 32852 32588 32864
rect 32640 32852 32646 32904
rect 32769 32895 32827 32901
rect 32769 32861 32781 32895
rect 32815 32892 32827 32895
rect 33134 32892 33140 32904
rect 32815 32864 33140 32892
rect 32815 32861 32827 32864
rect 32769 32855 32827 32861
rect 33134 32852 33140 32864
rect 33192 32852 33198 32904
rect 34238 32852 34244 32904
rect 34296 32892 34302 32904
rect 34701 32895 34759 32901
rect 34701 32892 34713 32895
rect 34296 32864 34713 32892
rect 34296 32852 34302 32864
rect 34701 32861 34713 32864
rect 34747 32861 34759 32895
rect 34701 32855 34759 32861
rect 31754 32784 31760 32836
rect 31812 32824 31818 32836
rect 32125 32827 32183 32833
rect 32125 32824 32137 32827
rect 31812 32796 32137 32824
rect 31812 32784 31818 32796
rect 32125 32793 32137 32796
rect 32171 32793 32183 32827
rect 32125 32787 32183 32793
rect 30926 32756 30932 32768
rect 30887 32728 30932 32756
rect 30926 32716 30932 32728
rect 30984 32716 30990 32768
rect 1104 32666 38824 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 34966 32666
rect 35018 32614 35030 32666
rect 35082 32614 35094 32666
rect 35146 32614 35158 32666
rect 35210 32614 38824 32666
rect 1104 32592 38824 32614
rect 29089 32555 29147 32561
rect 29089 32521 29101 32555
rect 29135 32552 29147 32555
rect 29822 32552 29828 32564
rect 29135 32524 29828 32552
rect 29135 32521 29147 32524
rect 29089 32515 29147 32521
rect 29822 32512 29828 32524
rect 29880 32512 29886 32564
rect 31849 32555 31907 32561
rect 31849 32521 31861 32555
rect 31895 32552 31907 32555
rect 32030 32552 32036 32564
rect 31895 32524 32036 32552
rect 31895 32521 31907 32524
rect 31849 32515 31907 32521
rect 32030 32512 32036 32524
rect 32088 32512 32094 32564
rect 32582 32512 32588 32564
rect 32640 32552 32646 32564
rect 32677 32555 32735 32561
rect 32677 32552 32689 32555
rect 32640 32524 32689 32552
rect 32640 32512 32646 32524
rect 32677 32521 32689 32524
rect 32723 32521 32735 32555
rect 34238 32552 34244 32564
rect 34199 32524 34244 32552
rect 32677 32515 32735 32521
rect 34238 32512 34244 32524
rect 34296 32552 34302 32564
rect 34422 32552 34428 32564
rect 34296 32524 34428 32552
rect 34296 32512 34302 32524
rect 34422 32512 34428 32524
rect 34480 32552 34486 32564
rect 34609 32555 34667 32561
rect 34609 32552 34621 32555
rect 34480 32524 34621 32552
rect 34480 32512 34486 32524
rect 34609 32521 34621 32524
rect 34655 32521 34667 32555
rect 36262 32552 36268 32564
rect 36223 32524 36268 32552
rect 34609 32515 34667 32521
rect 32766 32444 32772 32496
rect 32824 32484 32830 32496
rect 33410 32484 33416 32496
rect 32824 32456 33416 32484
rect 32824 32444 32830 32456
rect 33410 32444 33416 32456
rect 33468 32484 33474 32496
rect 33468 32456 33824 32484
rect 33468 32444 33474 32456
rect 33137 32419 33195 32425
rect 33137 32385 33149 32419
rect 33183 32416 33195 32419
rect 33686 32416 33692 32428
rect 33183 32388 33692 32416
rect 33183 32385 33195 32388
rect 33137 32379 33195 32385
rect 33686 32376 33692 32388
rect 33744 32376 33750 32428
rect 33796 32425 33824 32456
rect 33781 32419 33839 32425
rect 33781 32385 33793 32419
rect 33827 32385 33839 32419
rect 34624 32416 34652 32515
rect 36262 32512 36268 32524
rect 36320 32512 36326 32564
rect 37550 32552 37556 32564
rect 37511 32524 37556 32552
rect 37550 32512 37556 32524
rect 37608 32512 37614 32564
rect 34885 32419 34943 32425
rect 34885 32416 34897 32419
rect 34624 32388 34897 32416
rect 33781 32379 33839 32385
rect 34885 32385 34897 32388
rect 34931 32385 34943 32419
rect 34885 32379 34943 32385
rect 29362 32308 29368 32360
rect 29420 32348 29426 32360
rect 29641 32351 29699 32357
rect 29641 32348 29653 32351
rect 29420 32320 29653 32348
rect 29420 32308 29426 32320
rect 29641 32317 29653 32320
rect 29687 32317 29699 32351
rect 29641 32311 29699 32317
rect 31665 32351 31723 32357
rect 31665 32317 31677 32351
rect 31711 32348 31723 32351
rect 32122 32348 32128 32360
rect 31711 32320 32128 32348
rect 31711 32317 31723 32320
rect 31665 32311 31723 32317
rect 32122 32308 32128 32320
rect 32180 32308 32186 32360
rect 33226 32308 33232 32360
rect 33284 32348 33290 32360
rect 33597 32351 33655 32357
rect 33597 32348 33609 32351
rect 33284 32320 33609 32348
rect 33284 32308 33290 32320
rect 33597 32317 33609 32320
rect 33643 32317 33655 32351
rect 37366 32348 37372 32360
rect 37279 32320 37372 32348
rect 33597 32311 33655 32317
rect 37366 32308 37372 32320
rect 37424 32348 37430 32360
rect 37921 32351 37979 32357
rect 37921 32348 37933 32351
rect 37424 32320 37933 32348
rect 37424 32308 37430 32320
rect 37921 32317 37933 32320
rect 37967 32317 37979 32351
rect 37921 32311 37979 32317
rect 28721 32283 28779 32289
rect 28721 32249 28733 32283
rect 28767 32280 28779 32283
rect 29886 32283 29944 32289
rect 29886 32280 29898 32283
rect 28767 32252 29898 32280
rect 28767 32249 28779 32252
rect 28721 32243 28779 32249
rect 29886 32249 29898 32252
rect 29932 32280 29944 32283
rect 30926 32280 30932 32292
rect 29932 32252 30932 32280
rect 29932 32249 29944 32252
rect 29886 32243 29944 32249
rect 30926 32240 30932 32252
rect 30984 32280 30990 32292
rect 32582 32280 32588 32292
rect 30984 32252 32588 32280
rect 30984 32240 30990 32252
rect 32582 32240 32588 32252
rect 32640 32240 32646 32292
rect 35158 32289 35164 32292
rect 35152 32280 35164 32289
rect 35119 32252 35164 32280
rect 35152 32243 35164 32252
rect 35158 32240 35164 32243
rect 35216 32240 35222 32292
rect 29362 32172 29368 32224
rect 29420 32212 29426 32224
rect 29457 32215 29515 32221
rect 29457 32212 29469 32215
rect 29420 32184 29469 32212
rect 29420 32172 29426 32184
rect 29457 32181 29469 32184
rect 29503 32181 29515 32215
rect 29457 32175 29515 32181
rect 30098 32172 30104 32224
rect 30156 32212 30162 32224
rect 31021 32215 31079 32221
rect 31021 32212 31033 32215
rect 30156 32184 31033 32212
rect 30156 32172 30162 32184
rect 31021 32181 31033 32184
rect 31067 32212 31079 32215
rect 31849 32215 31907 32221
rect 31849 32212 31861 32215
rect 31067 32184 31861 32212
rect 31067 32181 31079 32184
rect 31021 32175 31079 32181
rect 31849 32181 31861 32184
rect 31895 32181 31907 32215
rect 31849 32175 31907 32181
rect 32030 32172 32036 32224
rect 32088 32212 32094 32224
rect 32309 32215 32367 32221
rect 32309 32212 32321 32215
rect 32088 32184 32321 32212
rect 32088 32172 32094 32184
rect 32309 32181 32321 32184
rect 32355 32181 32367 32215
rect 33226 32212 33232 32224
rect 33187 32184 33232 32212
rect 32309 32175 32367 32181
rect 33226 32172 33232 32184
rect 33284 32172 33290 32224
rect 1104 32122 38824 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 38824 32122
rect 1104 32048 38824 32070
rect 29089 32011 29147 32017
rect 29089 31977 29101 32011
rect 29135 31977 29147 32011
rect 29089 31971 29147 31977
rect 30009 32011 30067 32017
rect 30009 31977 30021 32011
rect 30055 32008 30067 32011
rect 30374 32008 30380 32020
rect 30055 31980 30380 32008
rect 30055 31977 30067 31980
rect 30009 31971 30067 31977
rect 29104 31940 29132 31971
rect 30374 31968 30380 31980
rect 30432 31968 30438 32020
rect 33410 32008 33416 32020
rect 33371 31980 33416 32008
rect 33410 31968 33416 31980
rect 33468 32008 33474 32020
rect 33778 32008 33784 32020
rect 33468 31980 33784 32008
rect 33468 31968 33474 31980
rect 33778 31968 33784 31980
rect 33836 31968 33842 32020
rect 35986 32008 35992 32020
rect 35947 31980 35992 32008
rect 35986 31968 35992 31980
rect 36044 31968 36050 32020
rect 30282 31940 30288 31952
rect 29104 31912 30288 31940
rect 30282 31900 30288 31912
rect 30340 31900 30346 31952
rect 31113 31943 31171 31949
rect 31113 31909 31125 31943
rect 31159 31940 31171 31943
rect 32401 31943 32459 31949
rect 32401 31940 32413 31943
rect 31159 31912 32413 31940
rect 31159 31909 31171 31912
rect 31113 31903 31171 31909
rect 32401 31909 32413 31912
rect 32447 31940 32459 31943
rect 33134 31940 33140 31952
rect 32447 31912 33140 31940
rect 32447 31909 32459 31912
rect 32401 31903 32459 31909
rect 28902 31872 28908 31884
rect 28863 31844 28908 31872
rect 28902 31832 28908 31844
rect 28960 31832 28966 31884
rect 29822 31832 29828 31884
rect 29880 31872 29886 31884
rect 30377 31875 30435 31881
rect 30377 31872 30389 31875
rect 29880 31844 30389 31872
rect 29880 31832 29886 31844
rect 30377 31841 30389 31844
rect 30423 31841 30435 31875
rect 30377 31835 30435 31841
rect 30466 31804 30472 31816
rect 30300 31776 30472 31804
rect 29362 31696 29368 31748
rect 29420 31736 29426 31748
rect 29549 31739 29607 31745
rect 29549 31736 29561 31739
rect 29420 31708 29561 31736
rect 29420 31696 29426 31708
rect 29549 31705 29561 31708
rect 29595 31705 29607 31739
rect 29549 31699 29607 31705
rect 29914 31696 29920 31748
rect 29972 31736 29978 31748
rect 30300 31736 30328 31776
rect 30466 31764 30472 31776
rect 30524 31764 30530 31816
rect 30653 31807 30711 31813
rect 30653 31773 30665 31807
rect 30699 31804 30711 31807
rect 31128 31804 31156 31903
rect 33134 31900 33140 31912
rect 33192 31940 33198 31952
rect 34057 31943 34115 31949
rect 34057 31940 34069 31943
rect 33192 31912 34069 31940
rect 33192 31900 33198 31912
rect 34057 31909 34069 31912
rect 34103 31940 34115 31943
rect 34146 31940 34152 31952
rect 34103 31912 34152 31940
rect 34103 31909 34115 31912
rect 34057 31903 34115 31909
rect 34146 31900 34152 31912
rect 34204 31900 34210 31952
rect 32861 31875 32919 31881
rect 32861 31841 32873 31875
rect 32907 31872 32919 31875
rect 32950 31872 32956 31884
rect 32907 31844 32956 31872
rect 32907 31841 32919 31844
rect 32861 31835 32919 31841
rect 32950 31832 32956 31844
rect 33008 31872 33014 31884
rect 33226 31872 33232 31884
rect 33008 31844 33232 31872
rect 33008 31832 33014 31844
rect 33226 31832 33232 31844
rect 33284 31832 33290 31884
rect 34514 31832 34520 31884
rect 34572 31872 34578 31884
rect 34609 31875 34667 31881
rect 34609 31872 34621 31875
rect 34572 31844 34621 31872
rect 34572 31832 34578 31844
rect 34609 31841 34621 31844
rect 34655 31872 34667 31875
rect 35158 31872 35164 31884
rect 34655 31844 35164 31872
rect 34655 31841 34667 31844
rect 34609 31835 34667 31841
rect 35158 31832 35164 31844
rect 35216 31872 35222 31884
rect 35253 31875 35311 31881
rect 35253 31872 35265 31875
rect 35216 31844 35265 31872
rect 35216 31832 35222 31844
rect 35253 31841 35265 31844
rect 35299 31841 35311 31875
rect 35253 31835 35311 31841
rect 30699 31776 31156 31804
rect 30699 31773 30711 31776
rect 30653 31767 30711 31773
rect 34146 31764 34152 31816
rect 34204 31804 34210 31816
rect 34698 31804 34704 31816
rect 34204 31776 34468 31804
rect 34659 31776 34704 31804
rect 34204 31764 34210 31776
rect 29972 31708 30328 31736
rect 34440 31736 34468 31776
rect 34698 31764 34704 31776
rect 34756 31764 34762 31816
rect 34793 31807 34851 31813
rect 34793 31773 34805 31807
rect 34839 31804 34851 31807
rect 35268 31804 35296 31835
rect 35342 31832 35348 31884
rect 35400 31872 35406 31884
rect 35805 31875 35863 31881
rect 35805 31872 35817 31875
rect 35400 31844 35817 31872
rect 35400 31832 35406 31844
rect 35805 31841 35817 31844
rect 35851 31841 35863 31875
rect 35805 31835 35863 31841
rect 34839 31776 34873 31804
rect 35268 31776 35756 31804
rect 34839 31773 34851 31776
rect 34793 31767 34851 31773
rect 34808 31736 34836 31767
rect 34440 31708 34836 31736
rect 29972 31696 29978 31708
rect 31665 31671 31723 31677
rect 31665 31637 31677 31671
rect 31711 31668 31723 31671
rect 32122 31668 32128 31680
rect 31711 31640 32128 31668
rect 31711 31637 31723 31640
rect 31665 31631 31723 31637
rect 32122 31628 32128 31640
rect 32180 31628 32186 31680
rect 33042 31668 33048 31680
rect 33003 31640 33048 31668
rect 33042 31628 33048 31640
rect 33100 31628 33106 31680
rect 34238 31668 34244 31680
rect 34199 31640 34244 31668
rect 34238 31628 34244 31640
rect 34296 31628 34302 31680
rect 34422 31628 34428 31680
rect 34480 31668 34486 31680
rect 34606 31668 34612 31680
rect 34480 31640 34612 31668
rect 34480 31628 34486 31640
rect 34606 31628 34612 31640
rect 34664 31628 34670 31680
rect 35728 31668 35756 31776
rect 35820 31736 35848 31835
rect 36814 31736 36820 31748
rect 35820 31708 36820 31736
rect 36814 31696 36820 31708
rect 36872 31696 36878 31748
rect 36262 31668 36268 31680
rect 35728 31640 36268 31668
rect 36262 31628 36268 31640
rect 36320 31628 36326 31680
rect 1104 31578 38824 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 34966 31578
rect 35018 31526 35030 31578
rect 35082 31526 35094 31578
rect 35146 31526 35158 31578
rect 35210 31526 38824 31578
rect 1104 31504 38824 31526
rect 28994 31464 29000 31476
rect 28955 31436 29000 31464
rect 28994 31424 29000 31436
rect 29052 31424 29058 31476
rect 29549 31467 29607 31473
rect 29549 31433 29561 31467
rect 29595 31464 29607 31467
rect 29822 31464 29828 31476
rect 29595 31436 29828 31464
rect 29595 31433 29607 31436
rect 29549 31427 29607 31433
rect 29822 31424 29828 31436
rect 29880 31424 29886 31476
rect 29914 31424 29920 31476
rect 29972 31464 29978 31476
rect 32950 31464 32956 31476
rect 29972 31436 30017 31464
rect 32911 31436 32956 31464
rect 29972 31424 29978 31436
rect 32950 31424 32956 31436
rect 33008 31424 33014 31476
rect 33597 31467 33655 31473
rect 33597 31433 33609 31467
rect 33643 31464 33655 31467
rect 34422 31464 34428 31476
rect 33643 31436 34428 31464
rect 33643 31433 33655 31436
rect 33597 31427 33655 31433
rect 34422 31424 34428 31436
rect 34480 31424 34486 31476
rect 34606 31464 34612 31476
rect 34567 31436 34612 31464
rect 34606 31424 34612 31436
rect 34664 31424 34670 31476
rect 36262 31464 36268 31476
rect 36223 31436 36268 31464
rect 36262 31424 36268 31436
rect 36320 31424 36326 31476
rect 36814 31464 36820 31476
rect 36775 31436 36820 31464
rect 36814 31424 36820 31436
rect 36872 31424 36878 31476
rect 29012 31396 29040 31424
rect 30009 31399 30067 31405
rect 30009 31396 30021 31399
rect 29012 31368 30021 31396
rect 30009 31365 30021 31368
rect 30055 31365 30067 31399
rect 31021 31399 31079 31405
rect 31021 31396 31033 31399
rect 30009 31359 30067 31365
rect 30484 31368 31033 31396
rect 30374 31288 30380 31340
rect 30432 31328 30438 31340
rect 30484 31337 30512 31368
rect 31021 31365 31033 31368
rect 31067 31365 31079 31399
rect 31021 31359 31079 31365
rect 30469 31331 30527 31337
rect 30469 31328 30481 31331
rect 30432 31300 30481 31328
rect 30432 31288 30438 31300
rect 30469 31297 30481 31300
rect 30515 31297 30527 31331
rect 30469 31291 30527 31297
rect 30558 31288 30564 31340
rect 30616 31328 30622 31340
rect 31481 31331 31539 31337
rect 30616 31300 30709 31328
rect 30616 31288 30622 31300
rect 31481 31297 31493 31331
rect 31527 31328 31539 31331
rect 32030 31328 32036 31340
rect 31527 31300 32036 31328
rect 31527 31297 31539 31300
rect 31481 31291 31539 31297
rect 32030 31288 32036 31300
rect 32088 31288 32094 31340
rect 32122 31288 32128 31340
rect 32180 31328 32186 31340
rect 34624 31328 34652 31424
rect 34885 31331 34943 31337
rect 34885 31328 34897 31331
rect 32180 31300 32225 31328
rect 34624 31300 34897 31328
rect 32180 31288 32186 31300
rect 34885 31297 34897 31300
rect 34931 31297 34943 31331
rect 34885 31291 34943 31297
rect 28261 31263 28319 31269
rect 28261 31229 28273 31263
rect 28307 31260 28319 31263
rect 30576 31260 30604 31288
rect 28307 31232 30604 31260
rect 28307 31229 28319 31232
rect 28261 31223 28319 31229
rect 28629 31195 28687 31201
rect 28629 31161 28641 31195
rect 28675 31192 28687 31195
rect 30377 31195 30435 31201
rect 30377 31192 30389 31195
rect 28675 31164 30389 31192
rect 28675 31161 28687 31164
rect 28629 31155 28687 31161
rect 30377 31161 30389 31164
rect 30423 31192 30435 31195
rect 31662 31192 31668 31204
rect 30423 31164 31668 31192
rect 30423 31161 30435 31164
rect 30377 31155 30435 31161
rect 31662 31152 31668 31164
rect 31720 31152 31726 31204
rect 33965 31195 34023 31201
rect 33965 31161 33977 31195
rect 34011 31192 34023 31195
rect 34333 31195 34391 31201
rect 34333 31192 34345 31195
rect 34011 31164 34345 31192
rect 34011 31161 34023 31164
rect 33965 31155 34023 31161
rect 34333 31161 34345 31164
rect 34379 31192 34391 31195
rect 34698 31192 34704 31204
rect 34379 31164 34704 31192
rect 34379 31161 34391 31164
rect 34333 31155 34391 31161
rect 34698 31152 34704 31164
rect 34756 31192 34762 31204
rect 35158 31201 35164 31204
rect 35152 31192 35164 31201
rect 34756 31164 35164 31192
rect 34756 31152 34762 31164
rect 35152 31155 35164 31164
rect 35158 31152 35164 31155
rect 35216 31152 35222 31204
rect 31570 31124 31576 31136
rect 31531 31096 31576 31124
rect 31570 31084 31576 31096
rect 31628 31084 31634 31136
rect 31938 31124 31944 31136
rect 31899 31096 31944 31124
rect 31938 31084 31944 31096
rect 31996 31084 32002 31136
rect 1104 31034 38824 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 38824 31034
rect 1104 30960 38824 30982
rect 30374 30880 30380 30932
rect 30432 30920 30438 30932
rect 31573 30923 31631 30929
rect 31573 30920 31585 30923
rect 30432 30892 31585 30920
rect 30432 30880 30438 30892
rect 31573 30889 31585 30892
rect 31619 30920 31631 30923
rect 31938 30920 31944 30932
rect 31619 30892 31944 30920
rect 31619 30889 31631 30892
rect 31573 30883 31631 30889
rect 31938 30880 31944 30892
rect 31996 30880 32002 30932
rect 32585 30923 32643 30929
rect 32585 30889 32597 30923
rect 32631 30920 32643 30923
rect 33042 30920 33048 30932
rect 32631 30892 33048 30920
rect 32631 30889 32643 30892
rect 32585 30883 32643 30889
rect 33042 30880 33048 30892
rect 33100 30880 33106 30932
rect 33321 30923 33379 30929
rect 33321 30889 33333 30923
rect 33367 30920 33379 30923
rect 33594 30920 33600 30932
rect 33367 30892 33600 30920
rect 33367 30889 33379 30892
rect 33321 30883 33379 30889
rect 33594 30880 33600 30892
rect 33652 30920 33658 30932
rect 34238 30920 34244 30932
rect 33652 30892 34244 30920
rect 33652 30880 33658 30892
rect 34238 30880 34244 30892
rect 34296 30880 34302 30932
rect 35158 30880 35164 30932
rect 35216 30920 35222 30932
rect 35805 30923 35863 30929
rect 35805 30920 35817 30923
rect 35216 30892 35817 30920
rect 35216 30880 35222 30892
rect 35805 30889 35817 30892
rect 35851 30889 35863 30923
rect 35805 30883 35863 30889
rect 29816 30855 29874 30861
rect 29816 30821 29828 30855
rect 29862 30852 29874 30855
rect 30098 30852 30104 30864
rect 29862 30824 30104 30852
rect 29862 30821 29874 30824
rect 29816 30815 29874 30821
rect 30098 30812 30104 30824
rect 30156 30812 30162 30864
rect 34606 30812 34612 30864
rect 34664 30861 34670 30864
rect 34664 30855 34728 30861
rect 34664 30821 34682 30855
rect 34716 30821 34728 30855
rect 34664 30815 34728 30821
rect 34664 30812 34670 30815
rect 29362 30744 29368 30796
rect 29420 30784 29426 30796
rect 29549 30787 29607 30793
rect 29549 30784 29561 30787
rect 29420 30756 29561 30784
rect 29420 30744 29426 30756
rect 29549 30753 29561 30756
rect 29595 30753 29607 30787
rect 29549 30747 29607 30753
rect 34425 30787 34483 30793
rect 34425 30753 34437 30787
rect 34471 30784 34483 30787
rect 34514 30784 34520 30796
rect 34471 30756 34520 30784
rect 34471 30753 34483 30756
rect 34425 30747 34483 30753
rect 34514 30744 34520 30756
rect 34572 30744 34578 30796
rect 32674 30716 32680 30728
rect 32635 30688 32680 30716
rect 32674 30676 32680 30688
rect 32732 30676 32738 30728
rect 32861 30719 32919 30725
rect 32861 30685 32873 30719
rect 32907 30716 32919 30719
rect 33134 30716 33140 30728
rect 32907 30688 33140 30716
rect 32907 30685 32919 30688
rect 32861 30679 32919 30685
rect 31662 30608 31668 30660
rect 31720 30648 31726 30660
rect 32122 30648 32128 30660
rect 31720 30620 32128 30648
rect 31720 30608 31726 30620
rect 32122 30608 32128 30620
rect 32180 30648 32186 30660
rect 32876 30648 32904 30679
rect 33134 30676 33140 30688
rect 33192 30676 33198 30728
rect 32180 30620 32904 30648
rect 32180 30608 32186 30620
rect 29457 30583 29515 30589
rect 29457 30549 29469 30583
rect 29503 30580 29515 30583
rect 29546 30580 29552 30592
rect 29503 30552 29552 30580
rect 29503 30549 29515 30552
rect 29457 30543 29515 30549
rect 29546 30540 29552 30552
rect 29604 30580 29610 30592
rect 30834 30580 30840 30592
rect 29604 30552 30840 30580
rect 29604 30540 29610 30552
rect 30834 30540 30840 30552
rect 30892 30580 30898 30592
rect 30929 30583 30987 30589
rect 30929 30580 30941 30583
rect 30892 30552 30941 30580
rect 30892 30540 30898 30552
rect 30929 30549 30941 30552
rect 30975 30549 30987 30583
rect 30929 30543 30987 30549
rect 31754 30540 31760 30592
rect 31812 30580 31818 30592
rect 32217 30583 32275 30589
rect 32217 30580 32229 30583
rect 31812 30552 32229 30580
rect 31812 30540 31818 30552
rect 32217 30549 32229 30552
rect 32263 30549 32275 30583
rect 32217 30543 32275 30549
rect 34333 30583 34391 30589
rect 34333 30549 34345 30583
rect 34379 30580 34391 30583
rect 34606 30580 34612 30592
rect 34379 30552 34612 30580
rect 34379 30549 34391 30552
rect 34333 30543 34391 30549
rect 34606 30540 34612 30552
rect 34664 30540 34670 30592
rect 1104 30490 38824 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 34966 30490
rect 35018 30438 35030 30490
rect 35082 30438 35094 30490
rect 35146 30438 35158 30490
rect 35210 30438 38824 30490
rect 1104 30416 38824 30438
rect 32309 30379 32367 30385
rect 32309 30345 32321 30379
rect 32355 30376 32367 30379
rect 32674 30376 32680 30388
rect 32355 30348 32680 30376
rect 32355 30345 32367 30348
rect 32309 30339 32367 30345
rect 32674 30336 32680 30348
rect 32732 30336 32738 30388
rect 33042 30376 33048 30388
rect 33003 30348 33048 30376
rect 33042 30336 33048 30348
rect 33100 30336 33106 30388
rect 34514 30376 34520 30388
rect 34475 30348 34520 30376
rect 34514 30336 34520 30348
rect 34572 30336 34578 30388
rect 28261 30311 28319 30317
rect 28261 30277 28273 30311
rect 28307 30308 28319 30311
rect 28810 30308 28816 30320
rect 28307 30280 28816 30308
rect 28307 30277 28319 30280
rect 28261 30271 28319 30277
rect 28810 30268 28816 30280
rect 28868 30268 28874 30320
rect 31662 30308 31668 30320
rect 31623 30280 31668 30308
rect 31662 30268 31668 30280
rect 31720 30268 31726 30320
rect 32033 30311 32091 30317
rect 32033 30277 32045 30311
rect 32079 30308 32091 30311
rect 33229 30311 33287 30317
rect 33229 30308 33241 30311
rect 32079 30280 33241 30308
rect 32079 30277 32091 30280
rect 32033 30271 32091 30277
rect 28718 30240 28724 30252
rect 28631 30212 28724 30240
rect 28718 30200 28724 30212
rect 28776 30240 28782 30252
rect 29089 30243 29147 30249
rect 29089 30240 29101 30243
rect 28776 30212 29101 30240
rect 28776 30200 28782 30212
rect 29089 30209 29101 30212
rect 29135 30240 29147 30243
rect 29362 30240 29368 30252
rect 29135 30212 29368 30240
rect 29135 30209 29147 30212
rect 29089 30203 29147 30209
rect 29362 30200 29368 30212
rect 29420 30200 29426 30252
rect 32140 30181 32168 30280
rect 33229 30277 33241 30280
rect 33275 30277 33287 30311
rect 33229 30271 33287 30277
rect 33870 30240 33876 30252
rect 33831 30212 33876 30240
rect 33870 30200 33876 30212
rect 33928 30200 33934 30252
rect 34532 30240 34560 30336
rect 34882 30240 34888 30252
rect 34532 30212 34888 30240
rect 34882 30200 34888 30212
rect 34940 30200 34946 30252
rect 28077 30175 28135 30181
rect 28077 30172 28089 30175
rect 28000 30144 28089 30172
rect 28000 30048 28028 30144
rect 28077 30141 28089 30144
rect 28123 30141 28135 30175
rect 28077 30135 28135 30141
rect 32125 30175 32183 30181
rect 32125 30141 32137 30175
rect 32171 30141 32183 30175
rect 33594 30172 33600 30184
rect 33555 30144 33600 30172
rect 32125 30135 32183 30141
rect 33594 30132 33600 30144
rect 33652 30132 33658 30184
rect 29546 30064 29552 30116
rect 29604 30113 29610 30116
rect 29604 30107 29668 30113
rect 29604 30073 29622 30107
rect 29656 30073 29668 30107
rect 29604 30067 29668 30073
rect 29604 30064 29610 30067
rect 34514 30064 34520 30116
rect 34572 30104 34578 30116
rect 35130 30107 35188 30113
rect 35130 30104 35142 30107
rect 34572 30076 35142 30104
rect 34572 30064 34578 30076
rect 35130 30073 35142 30076
rect 35176 30073 35188 30107
rect 35130 30067 35188 30073
rect 27982 30036 27988 30048
rect 27943 30008 27988 30036
rect 27982 29996 27988 30008
rect 28040 29996 28046 30048
rect 29086 29996 29092 30048
rect 29144 30036 29150 30048
rect 30745 30039 30803 30045
rect 30745 30036 30757 30039
rect 29144 30008 30757 30036
rect 29144 29996 29150 30008
rect 30745 30005 30757 30008
rect 30791 30005 30803 30039
rect 33686 30036 33692 30048
rect 33647 30008 33692 30036
rect 30745 29999 30803 30005
rect 33686 29996 33692 30008
rect 33744 29996 33750 30048
rect 34606 29996 34612 30048
rect 34664 30036 34670 30048
rect 36265 30039 36323 30045
rect 36265 30036 36277 30039
rect 34664 30008 36277 30036
rect 34664 29996 34670 30008
rect 36265 30005 36277 30008
rect 36311 30005 36323 30039
rect 36265 29999 36323 30005
rect 1104 29946 38824 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 38824 29946
rect 1104 29872 38824 29894
rect 30098 29832 30104 29844
rect 30059 29804 30104 29832
rect 30098 29792 30104 29804
rect 30156 29792 30162 29844
rect 33321 29835 33379 29841
rect 33321 29801 33333 29835
rect 33367 29832 33379 29835
rect 33686 29832 33692 29844
rect 33367 29804 33692 29832
rect 33367 29801 33379 29804
rect 33321 29795 33379 29801
rect 33686 29792 33692 29804
rect 33744 29832 33750 29844
rect 34241 29835 34299 29841
rect 34241 29832 34253 29835
rect 33744 29804 34253 29832
rect 33744 29792 33750 29804
rect 34241 29801 34253 29804
rect 34287 29801 34299 29835
rect 34241 29795 34299 29801
rect 34882 29792 34888 29844
rect 34940 29832 34946 29844
rect 35253 29835 35311 29841
rect 35253 29832 35265 29835
rect 34940 29804 35265 29832
rect 34940 29792 34946 29804
rect 35253 29801 35265 29804
rect 35299 29801 35311 29835
rect 35253 29795 35311 29801
rect 35894 29792 35900 29844
rect 35952 29832 35958 29844
rect 35989 29835 36047 29841
rect 35989 29832 36001 29835
rect 35952 29804 36001 29832
rect 35952 29792 35958 29804
rect 35989 29801 36001 29804
rect 36035 29801 36047 29835
rect 35989 29795 36047 29801
rect 28436 29767 28494 29773
rect 28436 29733 28448 29767
rect 28482 29764 28494 29767
rect 29086 29764 29092 29776
rect 28482 29736 29092 29764
rect 28482 29733 28494 29736
rect 28436 29727 28494 29733
rect 29086 29724 29092 29736
rect 29144 29724 29150 29776
rect 30650 29764 30656 29776
rect 30611 29736 30656 29764
rect 30650 29724 30656 29736
rect 30708 29724 30714 29776
rect 34146 29764 34152 29776
rect 34107 29736 34152 29764
rect 34146 29724 34152 29736
rect 34204 29764 34210 29776
rect 34204 29736 34836 29764
rect 34204 29724 34210 29736
rect 28169 29699 28227 29705
rect 28169 29665 28181 29699
rect 28215 29696 28227 29699
rect 28718 29696 28724 29708
rect 28215 29668 28724 29696
rect 28215 29665 28227 29668
rect 28169 29659 28227 29665
rect 28718 29656 28724 29668
rect 28776 29656 28782 29708
rect 30834 29696 30840 29708
rect 30795 29668 30840 29696
rect 30834 29656 30840 29668
rect 30892 29656 30898 29708
rect 31021 29699 31079 29705
rect 31021 29665 31033 29699
rect 31067 29696 31079 29699
rect 32122 29696 32128 29708
rect 31067 29668 32128 29696
rect 31067 29665 31079 29668
rect 31021 29659 31079 29665
rect 32122 29656 32128 29668
rect 32180 29656 32186 29708
rect 34606 29696 34612 29708
rect 34567 29668 34612 29696
rect 34606 29656 34612 29668
rect 34664 29656 34670 29708
rect 34514 29588 34520 29640
rect 34572 29628 34578 29640
rect 34808 29637 34836 29736
rect 35802 29696 35808 29708
rect 35763 29668 35808 29696
rect 35802 29656 35808 29668
rect 35860 29656 35866 29708
rect 34701 29631 34759 29637
rect 34701 29628 34713 29631
rect 34572 29600 34713 29628
rect 34572 29588 34578 29600
rect 34701 29597 34713 29600
rect 34747 29597 34759 29631
rect 34701 29591 34759 29597
rect 34793 29631 34851 29637
rect 34793 29597 34805 29631
rect 34839 29628 34851 29631
rect 35250 29628 35256 29640
rect 34839 29600 35256 29628
rect 34839 29597 34851 29600
rect 34793 29591 34851 29597
rect 34716 29560 34744 29591
rect 35250 29588 35256 29600
rect 35308 29588 35314 29640
rect 35621 29563 35679 29569
rect 35621 29560 35633 29563
rect 34716 29532 35633 29560
rect 35621 29529 35633 29532
rect 35667 29560 35679 29563
rect 36262 29560 36268 29572
rect 35667 29532 36268 29560
rect 35667 29529 35679 29532
rect 35621 29523 35679 29529
rect 36262 29520 36268 29532
rect 36320 29520 36326 29572
rect 27706 29492 27712 29504
rect 27667 29464 27712 29492
rect 27706 29452 27712 29464
rect 27764 29452 27770 29504
rect 28442 29452 28448 29504
rect 28500 29492 28506 29504
rect 29549 29495 29607 29501
rect 29549 29492 29561 29495
rect 28500 29464 29561 29492
rect 28500 29452 28506 29464
rect 29549 29461 29561 29464
rect 29595 29461 29607 29495
rect 29549 29455 29607 29461
rect 30742 29452 30748 29504
rect 30800 29492 30806 29504
rect 32309 29495 32367 29501
rect 32309 29492 32321 29495
rect 30800 29464 32321 29492
rect 30800 29452 30806 29464
rect 32309 29461 32321 29464
rect 32355 29461 32367 29495
rect 32309 29455 32367 29461
rect 33689 29495 33747 29501
rect 33689 29461 33701 29495
rect 33735 29492 33747 29495
rect 33870 29492 33876 29504
rect 33735 29464 33876 29492
rect 33735 29461 33747 29464
rect 33689 29455 33747 29461
rect 33870 29452 33876 29464
rect 33928 29492 33934 29504
rect 36078 29492 36084 29504
rect 33928 29464 36084 29492
rect 33928 29452 33934 29464
rect 36078 29452 36084 29464
rect 36136 29452 36142 29504
rect 1104 29402 38824 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 34966 29402
rect 35018 29350 35030 29402
rect 35082 29350 35094 29402
rect 35146 29350 35158 29402
rect 35210 29350 38824 29402
rect 1104 29328 38824 29350
rect 27982 29248 27988 29300
rect 28040 29288 28046 29300
rect 30009 29291 30067 29297
rect 30009 29288 30021 29291
rect 28040 29260 30021 29288
rect 28040 29248 28046 29260
rect 30009 29257 30021 29260
rect 30055 29257 30067 29291
rect 30009 29251 30067 29257
rect 30650 29248 30656 29300
rect 30708 29288 30714 29300
rect 31021 29291 31079 29297
rect 31021 29288 31033 29291
rect 30708 29260 31033 29288
rect 30708 29248 30714 29260
rect 31021 29257 31033 29260
rect 31067 29257 31079 29291
rect 32122 29288 32128 29300
rect 32083 29260 32128 29288
rect 31021 29251 31079 29257
rect 32122 29248 32128 29260
rect 32180 29248 32186 29300
rect 33597 29291 33655 29297
rect 33597 29257 33609 29291
rect 33643 29288 33655 29291
rect 34606 29288 34612 29300
rect 33643 29260 34612 29288
rect 33643 29257 33655 29260
rect 33597 29251 33655 29257
rect 34606 29248 34612 29260
rect 34664 29248 34670 29300
rect 34701 29291 34759 29297
rect 34701 29257 34713 29291
rect 34747 29288 34759 29291
rect 34790 29288 34796 29300
rect 34747 29260 34796 29288
rect 34747 29257 34759 29260
rect 34701 29251 34759 29257
rect 34790 29248 34796 29260
rect 34848 29248 34854 29300
rect 36262 29288 36268 29300
rect 36223 29260 36268 29288
rect 36262 29248 36268 29260
rect 36320 29248 36326 29300
rect 28718 29220 28724 29232
rect 28679 29192 28724 29220
rect 28718 29180 28724 29192
rect 28776 29180 28782 29232
rect 29086 29220 29092 29232
rect 29047 29192 29092 29220
rect 29086 29180 29092 29192
rect 29144 29220 29150 29232
rect 29822 29220 29828 29232
rect 29144 29192 29828 29220
rect 29144 29180 29150 29192
rect 29822 29180 29828 29192
rect 29880 29180 29886 29232
rect 30834 29180 30840 29232
rect 30892 29220 30898 29232
rect 31389 29223 31447 29229
rect 31389 29220 31401 29223
rect 30892 29192 31401 29220
rect 30892 29180 30898 29192
rect 31389 29189 31401 29192
rect 31435 29189 31447 29223
rect 31389 29183 31447 29189
rect 33134 29180 33140 29232
rect 33192 29220 33198 29232
rect 33873 29223 33931 29229
rect 33873 29220 33885 29223
rect 33192 29192 33885 29220
rect 33192 29180 33198 29192
rect 33873 29189 33885 29192
rect 33919 29189 33931 29223
rect 33873 29183 33931 29189
rect 28261 29155 28319 29161
rect 28261 29121 28273 29155
rect 28307 29152 28319 29155
rect 28442 29152 28448 29164
rect 28307 29124 28448 29152
rect 28307 29121 28319 29124
rect 28261 29115 28319 29121
rect 28442 29112 28448 29124
rect 28500 29112 28506 29164
rect 29549 29155 29607 29161
rect 29549 29121 29561 29155
rect 29595 29152 29607 29155
rect 30653 29155 30711 29161
rect 30653 29152 30665 29155
rect 29595 29124 30665 29152
rect 29595 29121 29607 29124
rect 29549 29115 29607 29121
rect 30653 29121 30665 29124
rect 30699 29152 30711 29155
rect 30742 29152 30748 29164
rect 30699 29124 30748 29152
rect 30699 29121 30711 29124
rect 30653 29115 30711 29121
rect 30742 29112 30748 29124
rect 30800 29112 30806 29164
rect 34330 29152 34336 29164
rect 33704 29124 34336 29152
rect 27706 29044 27712 29096
rect 27764 29084 27770 29096
rect 28077 29087 28135 29093
rect 28077 29084 28089 29087
rect 27764 29056 28089 29084
rect 27764 29044 27770 29056
rect 28077 29053 28089 29056
rect 28123 29084 28135 29087
rect 28902 29084 28908 29096
rect 28123 29056 28908 29084
rect 28123 29053 28135 29056
rect 28077 29047 28135 29053
rect 28902 29044 28908 29056
rect 28960 29044 28966 29096
rect 29917 29087 29975 29093
rect 29917 29053 29929 29087
rect 29963 29084 29975 29087
rect 30466 29084 30472 29096
rect 29963 29056 30472 29084
rect 29963 29053 29975 29056
rect 29917 29047 29975 29053
rect 30466 29044 30472 29056
rect 30524 29084 30530 29096
rect 31662 29084 31668 29096
rect 30524 29056 31668 29084
rect 30524 29044 30530 29056
rect 31662 29044 31668 29056
rect 31720 29044 31726 29096
rect 33704 29093 33732 29124
rect 34330 29112 34336 29124
rect 34388 29112 34394 29164
rect 34808 29152 34836 29248
rect 34885 29155 34943 29161
rect 34885 29152 34897 29155
rect 34808 29124 34897 29152
rect 34885 29121 34897 29124
rect 34931 29121 34943 29155
rect 34885 29115 34943 29121
rect 33689 29087 33747 29093
rect 33689 29053 33701 29087
rect 33735 29053 33747 29087
rect 33689 29047 33747 29053
rect 27525 29019 27583 29025
rect 27525 28985 27537 29019
rect 27571 29016 27583 29019
rect 27985 29019 28043 29025
rect 27985 29016 27997 29019
rect 27571 28988 27997 29016
rect 27571 28985 27583 28988
rect 27525 28979 27583 28985
rect 27985 28985 27997 28988
rect 28031 29016 28043 29019
rect 28166 29016 28172 29028
rect 28031 28988 28172 29016
rect 28031 28985 28043 28988
rect 27985 28979 28043 28985
rect 28166 28976 28172 28988
rect 28224 28976 28230 29028
rect 30374 29016 30380 29028
rect 30287 28988 30380 29016
rect 30374 28976 30380 28988
rect 30432 29016 30438 29028
rect 31570 29016 31576 29028
rect 30432 28988 31576 29016
rect 30432 28976 30438 28988
rect 31570 28976 31576 28988
rect 31628 28976 31634 29028
rect 34974 28976 34980 29028
rect 35032 29016 35038 29028
rect 35130 29019 35188 29025
rect 35130 29016 35142 29019
rect 35032 28988 35142 29016
rect 35032 28976 35038 28988
rect 35130 28985 35142 28988
rect 35176 29016 35188 29019
rect 35802 29016 35808 29028
rect 35176 28988 35808 29016
rect 35176 28985 35188 28988
rect 35130 28979 35188 28985
rect 35802 28976 35808 28988
rect 35860 28976 35866 29028
rect 27614 28948 27620 28960
rect 27575 28920 27620 28948
rect 27614 28908 27620 28920
rect 27672 28908 27678 28960
rect 1104 28858 38824 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 38824 28858
rect 1104 28784 38824 28806
rect 29086 28704 29092 28756
rect 29144 28744 29150 28756
rect 30101 28747 30159 28753
rect 30101 28744 30113 28747
rect 29144 28716 30113 28744
rect 29144 28704 29150 28716
rect 30101 28713 30113 28716
rect 30147 28744 30159 28747
rect 30282 28744 30288 28756
rect 30147 28716 30288 28744
rect 30147 28713 30159 28716
rect 30101 28707 30159 28713
rect 30282 28704 30288 28716
rect 30340 28704 30346 28756
rect 34333 28747 34391 28753
rect 34333 28713 34345 28747
rect 34379 28744 34391 28747
rect 34422 28744 34428 28756
rect 34379 28716 34428 28744
rect 34379 28713 34391 28716
rect 34333 28707 34391 28713
rect 34422 28704 34428 28716
rect 34480 28704 34486 28756
rect 34974 28744 34980 28756
rect 34935 28716 34980 28744
rect 34974 28704 34980 28716
rect 35032 28704 35038 28756
rect 35618 28744 35624 28756
rect 35579 28716 35624 28744
rect 35618 28704 35624 28716
rect 35676 28704 35682 28756
rect 36078 28704 36084 28756
rect 36136 28744 36142 28756
rect 36725 28747 36783 28753
rect 36725 28744 36737 28747
rect 36136 28716 36737 28744
rect 36136 28704 36142 28716
rect 36725 28713 36737 28716
rect 36771 28713 36783 28747
rect 36725 28707 36783 28713
rect 27709 28679 27767 28685
rect 27709 28645 27721 28679
rect 27755 28676 27767 28679
rect 28252 28679 28310 28685
rect 28252 28676 28264 28679
rect 27755 28648 28264 28676
rect 27755 28645 27767 28648
rect 27709 28639 27767 28645
rect 28252 28645 28264 28648
rect 28298 28676 28310 28679
rect 28442 28676 28448 28688
rect 28298 28648 28448 28676
rect 28298 28645 28310 28648
rect 28252 28639 28310 28645
rect 28442 28636 28448 28648
rect 28500 28636 28506 28688
rect 27982 28608 27988 28620
rect 27895 28580 27988 28608
rect 27982 28568 27988 28580
rect 28040 28608 28046 28620
rect 28718 28608 28724 28620
rect 28040 28580 28724 28608
rect 28040 28568 28046 28580
rect 28718 28568 28724 28580
rect 28776 28568 28782 28620
rect 30466 28608 30472 28620
rect 30427 28580 30472 28608
rect 30466 28568 30472 28580
rect 30524 28568 30530 28620
rect 35434 28608 35440 28620
rect 35395 28580 35440 28608
rect 35434 28568 35440 28580
rect 35492 28568 35498 28620
rect 36541 28611 36599 28617
rect 36541 28577 36553 28611
rect 36587 28608 36599 28611
rect 36630 28608 36636 28620
rect 36587 28580 36636 28608
rect 36587 28577 36599 28580
rect 36541 28571 36599 28577
rect 36630 28568 36636 28580
rect 36688 28568 36694 28620
rect 32214 28500 32220 28552
rect 32272 28540 32278 28552
rect 32401 28543 32459 28549
rect 32401 28540 32413 28543
rect 32272 28512 32413 28540
rect 32272 28500 32278 28512
rect 32401 28509 32413 28512
rect 32447 28509 32459 28543
rect 32401 28503 32459 28509
rect 28626 28364 28632 28416
rect 28684 28404 28690 28416
rect 29365 28407 29423 28413
rect 29365 28404 29377 28407
rect 28684 28376 29377 28404
rect 28684 28364 28690 28376
rect 29365 28373 29377 28376
rect 29411 28373 29423 28407
rect 30650 28404 30656 28416
rect 30611 28376 30656 28404
rect 29365 28367 29423 28373
rect 30650 28364 30656 28376
rect 30708 28364 30714 28416
rect 35986 28404 35992 28416
rect 35947 28376 35992 28404
rect 35986 28364 35992 28376
rect 36044 28364 36050 28416
rect 1104 28314 38824 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 34966 28314
rect 35018 28262 35030 28314
rect 35082 28262 35094 28314
rect 35146 28262 35158 28314
rect 35210 28262 38824 28314
rect 1104 28240 38824 28262
rect 27982 28200 27988 28212
rect 27943 28172 27988 28200
rect 27982 28160 27988 28172
rect 28040 28160 28046 28212
rect 28442 28160 28448 28212
rect 28500 28200 28506 28212
rect 28629 28203 28687 28209
rect 28629 28200 28641 28203
rect 28500 28172 28641 28200
rect 28500 28160 28506 28172
rect 28629 28169 28641 28172
rect 28675 28169 28687 28203
rect 28629 28163 28687 28169
rect 28994 28160 29000 28212
rect 29052 28200 29058 28212
rect 29273 28203 29331 28209
rect 29273 28200 29285 28203
rect 29052 28172 29285 28200
rect 29052 28160 29058 28172
rect 29273 28169 29285 28172
rect 29319 28169 29331 28203
rect 29273 28163 29331 28169
rect 30466 28160 30472 28212
rect 30524 28200 30530 28212
rect 30653 28203 30711 28209
rect 30653 28200 30665 28203
rect 30524 28172 30665 28200
rect 30524 28160 30530 28172
rect 30653 28169 30665 28172
rect 30699 28169 30711 28203
rect 32214 28200 32220 28212
rect 32175 28172 32220 28200
rect 30653 28163 30711 28169
rect 32214 28160 32220 28172
rect 32272 28160 32278 28212
rect 32306 28160 32312 28212
rect 32364 28200 32370 28212
rect 32364 28172 32409 28200
rect 32364 28160 32370 28172
rect 35250 28160 35256 28212
rect 35308 28200 35314 28212
rect 35621 28203 35679 28209
rect 35621 28200 35633 28203
rect 35308 28172 35633 28200
rect 35308 28160 35314 28172
rect 35621 28169 35633 28172
rect 35667 28169 35679 28203
rect 35621 28163 35679 28169
rect 30285 28135 30343 28141
rect 30285 28132 30297 28135
rect 29748 28104 30297 28132
rect 28166 28064 28172 28076
rect 28127 28036 28172 28064
rect 28166 28024 28172 28036
rect 28224 28024 28230 28076
rect 28994 28024 29000 28076
rect 29052 28064 29058 28076
rect 29748 28073 29776 28104
rect 30285 28101 30297 28104
rect 30331 28101 30343 28135
rect 30285 28095 30343 28101
rect 29733 28067 29791 28073
rect 29733 28064 29745 28067
rect 29052 28036 29745 28064
rect 29052 28024 29058 28036
rect 29733 28033 29745 28036
rect 29779 28033 29791 28067
rect 29733 28027 29791 28033
rect 29822 28024 29828 28076
rect 29880 28064 29886 28076
rect 31849 28067 31907 28073
rect 29880 28036 29925 28064
rect 29880 28024 29886 28036
rect 31849 28033 31861 28067
rect 31895 28064 31907 28067
rect 32858 28064 32864 28076
rect 31895 28036 32864 28064
rect 31895 28033 31907 28036
rect 31849 28027 31907 28033
rect 32858 28024 32864 28036
rect 32916 28024 32922 28076
rect 29089 27999 29147 28005
rect 29089 27965 29101 27999
rect 29135 27996 29147 27999
rect 29641 27999 29699 28005
rect 29641 27996 29653 27999
rect 29135 27968 29653 27996
rect 29135 27965 29147 27968
rect 29089 27959 29147 27965
rect 29641 27965 29653 27968
rect 29687 27996 29699 27999
rect 30650 27996 30656 28008
rect 29687 27968 30656 27996
rect 29687 27965 29699 27968
rect 29641 27959 29699 27965
rect 30650 27956 30656 27968
rect 30708 27956 30714 28008
rect 32214 27956 32220 28008
rect 32272 27996 32278 28008
rect 32677 27999 32735 28005
rect 32677 27996 32689 27999
rect 32272 27968 32689 27996
rect 32272 27956 32278 27968
rect 32677 27965 32689 27968
rect 32723 27965 32735 27999
rect 32677 27959 32735 27965
rect 35437 27999 35495 28005
rect 35437 27965 35449 27999
rect 35483 27996 35495 27999
rect 36630 27996 36636 28008
rect 35483 27968 35848 27996
rect 36591 27968 36636 27996
rect 35483 27965 35495 27968
rect 35437 27959 35495 27965
rect 31481 27931 31539 27937
rect 31481 27897 31493 27931
rect 31527 27928 31539 27931
rect 31662 27928 31668 27940
rect 31527 27900 31668 27928
rect 31527 27897 31539 27900
rect 31481 27891 31539 27897
rect 31662 27888 31668 27900
rect 31720 27928 31726 27940
rect 32769 27931 32827 27937
rect 32769 27928 32781 27931
rect 31720 27900 32781 27928
rect 31720 27888 31726 27900
rect 32769 27897 32781 27900
rect 32815 27897 32827 27931
rect 32769 27891 32827 27897
rect 35820 27872 35848 27968
rect 36630 27956 36636 27968
rect 36688 27956 36694 28008
rect 35345 27863 35403 27869
rect 35345 27829 35357 27863
rect 35391 27860 35403 27863
rect 35434 27860 35440 27872
rect 35391 27832 35440 27860
rect 35391 27829 35403 27832
rect 35345 27823 35403 27829
rect 35434 27820 35440 27832
rect 35492 27820 35498 27872
rect 35802 27820 35808 27872
rect 35860 27860 35866 27872
rect 35989 27863 36047 27869
rect 35989 27860 36001 27863
rect 35860 27832 36001 27860
rect 35860 27820 35866 27832
rect 35989 27829 36001 27832
rect 36035 27829 36047 27863
rect 35989 27823 36047 27829
rect 1104 27770 38824 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 38824 27770
rect 1104 27696 38824 27718
rect 29822 27616 29828 27668
rect 29880 27656 29886 27668
rect 29917 27659 29975 27665
rect 29917 27656 29929 27659
rect 29880 27628 29929 27656
rect 29880 27616 29886 27628
rect 29917 27625 29929 27628
rect 29963 27625 29975 27659
rect 29917 27619 29975 27625
rect 31662 27616 31668 27668
rect 31720 27656 31726 27668
rect 32125 27659 32183 27665
rect 32125 27656 32137 27659
rect 31720 27628 32137 27656
rect 31720 27616 31726 27628
rect 32125 27625 32137 27628
rect 32171 27625 32183 27659
rect 32125 27619 32183 27625
rect 34140 27591 34198 27597
rect 34140 27557 34152 27591
rect 34186 27588 34198 27591
rect 34238 27588 34244 27600
rect 34186 27560 34244 27588
rect 34186 27557 34198 27560
rect 34140 27551 34198 27557
rect 34238 27548 34244 27560
rect 34296 27548 34302 27600
rect 23106 27520 23112 27532
rect 23067 27492 23112 27520
rect 23106 27480 23112 27492
rect 23164 27480 23170 27532
rect 24302 27480 24308 27532
rect 24360 27520 24366 27532
rect 24397 27523 24455 27529
rect 24397 27520 24409 27523
rect 24360 27492 24409 27520
rect 24360 27480 24366 27492
rect 24397 27489 24409 27492
rect 24443 27520 24455 27523
rect 24949 27523 25007 27529
rect 24949 27520 24961 27523
rect 24443 27492 24961 27520
rect 24443 27489 24455 27492
rect 24397 27483 24455 27489
rect 24949 27489 24961 27492
rect 24995 27489 25007 27523
rect 28902 27520 28908 27532
rect 28863 27492 28908 27520
rect 24949 27483 25007 27489
rect 28902 27480 28908 27492
rect 28960 27480 28966 27532
rect 31846 27480 31852 27532
rect 31904 27520 31910 27532
rect 32493 27523 32551 27529
rect 32493 27520 32505 27523
rect 31904 27492 32505 27520
rect 31904 27480 31910 27492
rect 32493 27489 32505 27492
rect 32539 27489 32551 27523
rect 32493 27483 32551 27489
rect 28445 27455 28503 27461
rect 28445 27421 28457 27455
rect 28491 27452 28503 27455
rect 28994 27452 29000 27464
rect 28491 27424 29000 27452
rect 28491 27421 28503 27424
rect 28445 27415 28503 27421
rect 28994 27412 29000 27424
rect 29052 27412 29058 27464
rect 29089 27455 29147 27461
rect 29089 27421 29101 27455
rect 29135 27421 29147 27455
rect 30098 27452 30104 27464
rect 30059 27424 30104 27452
rect 29089 27415 29147 27421
rect 28077 27387 28135 27393
rect 28077 27353 28089 27387
rect 28123 27384 28135 27387
rect 29104 27384 29132 27415
rect 30098 27412 30104 27424
rect 30156 27412 30162 27464
rect 31294 27412 31300 27464
rect 31352 27452 31358 27464
rect 32582 27452 32588 27464
rect 31352 27424 32588 27452
rect 31352 27412 31358 27424
rect 32582 27412 32588 27424
rect 32640 27412 32646 27464
rect 32677 27455 32735 27461
rect 32677 27421 32689 27455
rect 32723 27421 32735 27455
rect 33870 27452 33876 27464
rect 33831 27424 33876 27452
rect 32677 27415 32735 27421
rect 29546 27384 29552 27396
rect 28123 27356 29552 27384
rect 28123 27353 28135 27356
rect 28077 27347 28135 27353
rect 29546 27344 29552 27356
rect 29604 27344 29610 27396
rect 31941 27387 31999 27393
rect 31941 27353 31953 27387
rect 31987 27384 31999 27387
rect 32030 27384 32036 27396
rect 31987 27356 32036 27384
rect 31987 27353 31999 27356
rect 31941 27347 31999 27353
rect 32030 27344 32036 27356
rect 32088 27384 32094 27396
rect 32692 27384 32720 27415
rect 33870 27412 33876 27424
rect 33928 27412 33934 27464
rect 35710 27412 35716 27464
rect 35768 27452 35774 27464
rect 36357 27455 36415 27461
rect 36357 27452 36369 27455
rect 35768 27424 36369 27452
rect 35768 27412 35774 27424
rect 36357 27421 36369 27424
rect 36403 27421 36415 27455
rect 36357 27415 36415 27421
rect 32088 27356 32720 27384
rect 32088 27344 32094 27356
rect 21910 27316 21916 27328
rect 21871 27288 21916 27316
rect 21910 27276 21916 27288
rect 21968 27276 21974 27328
rect 23290 27316 23296 27328
rect 23251 27288 23296 27316
rect 23290 27276 23296 27288
rect 23348 27276 23354 27328
rect 24581 27319 24639 27325
rect 24581 27285 24593 27319
rect 24627 27316 24639 27319
rect 24762 27316 24768 27328
rect 24627 27288 24768 27316
rect 24627 27285 24639 27288
rect 24581 27279 24639 27285
rect 24762 27276 24768 27288
rect 24820 27276 24826 27328
rect 28537 27319 28595 27325
rect 28537 27285 28549 27319
rect 28583 27316 28595 27319
rect 28810 27316 28816 27328
rect 28583 27288 28816 27316
rect 28583 27285 28595 27288
rect 28537 27279 28595 27285
rect 28810 27276 28816 27288
rect 28868 27276 28874 27328
rect 35250 27316 35256 27328
rect 35211 27288 35256 27316
rect 35250 27276 35256 27288
rect 35308 27276 35314 27328
rect 35526 27276 35532 27328
rect 35584 27316 35590 27328
rect 35805 27319 35863 27325
rect 35805 27316 35817 27319
rect 35584 27288 35817 27316
rect 35584 27276 35590 27288
rect 35805 27285 35817 27288
rect 35851 27285 35863 27319
rect 35805 27279 35863 27285
rect 1104 27226 38824 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 34966 27226
rect 35018 27174 35030 27226
rect 35082 27174 35094 27226
rect 35146 27174 35158 27226
rect 35210 27174 38824 27226
rect 1104 27152 38824 27174
rect 28718 27072 28724 27124
rect 28776 27112 28782 27124
rect 31294 27112 31300 27124
rect 28776 27084 29040 27112
rect 31255 27084 31300 27112
rect 28776 27072 28782 27084
rect 21361 26979 21419 26985
rect 21361 26945 21373 26979
rect 21407 26976 21419 26979
rect 21818 26976 21824 26988
rect 21407 26948 21824 26976
rect 21407 26945 21419 26948
rect 21361 26939 21419 26945
rect 21818 26936 21824 26948
rect 21876 26976 21882 26988
rect 22373 26979 22431 26985
rect 22373 26976 22385 26979
rect 21876 26948 22385 26976
rect 21876 26936 21882 26948
rect 22373 26945 22385 26948
rect 22419 26945 22431 26979
rect 29012 26976 29040 27084
rect 31294 27072 31300 27084
rect 31352 27072 31358 27124
rect 32858 27072 32864 27124
rect 32916 27112 32922 27124
rect 33137 27115 33195 27121
rect 33137 27112 33149 27115
rect 32916 27084 33149 27112
rect 32916 27072 32922 27084
rect 33137 27081 33149 27084
rect 33183 27081 33195 27115
rect 33137 27075 33195 27081
rect 35894 27072 35900 27124
rect 35952 27112 35958 27124
rect 36357 27115 36415 27121
rect 36357 27112 36369 27115
rect 35952 27084 36369 27112
rect 35952 27072 35958 27084
rect 36357 27081 36369 27084
rect 36403 27081 36415 27115
rect 36357 27075 36415 27081
rect 29178 26976 29184 26988
rect 29012 26948 29184 26976
rect 22373 26939 22431 26945
rect 29178 26936 29184 26948
rect 29236 26976 29242 26988
rect 29273 26979 29331 26985
rect 29273 26976 29285 26979
rect 29236 26948 29285 26976
rect 29236 26936 29242 26948
rect 29273 26945 29285 26948
rect 29319 26945 29331 26979
rect 29273 26939 29331 26945
rect 21910 26868 21916 26920
rect 21968 26908 21974 26920
rect 22189 26911 22247 26917
rect 22189 26908 22201 26911
rect 21968 26880 22201 26908
rect 21968 26868 21974 26880
rect 22189 26877 22201 26880
rect 22235 26877 22247 26911
rect 22189 26871 22247 26877
rect 24581 26911 24639 26917
rect 24581 26877 24593 26911
rect 24627 26908 24639 26911
rect 24670 26908 24676 26920
rect 24627 26880 24676 26908
rect 24627 26877 24639 26880
rect 24581 26871 24639 26877
rect 24670 26868 24676 26880
rect 24728 26868 24734 26920
rect 29546 26917 29552 26920
rect 27985 26911 28043 26917
rect 27985 26877 27997 26911
rect 28031 26908 28043 26911
rect 29540 26908 29552 26917
rect 28031 26880 28764 26908
rect 29507 26880 29552 26908
rect 28031 26877 28043 26880
rect 27985 26871 28043 26877
rect 21729 26843 21787 26849
rect 21729 26809 21741 26843
rect 21775 26840 21787 26843
rect 24213 26843 24271 26849
rect 21775 26812 22324 26840
rect 21775 26809 21787 26812
rect 21729 26803 21787 26809
rect 22296 26784 22324 26812
rect 24213 26809 24225 26843
rect 24259 26840 24271 26843
rect 24918 26843 24976 26849
rect 24918 26840 24930 26843
rect 24259 26812 24930 26840
rect 24259 26809 24271 26812
rect 24213 26803 24271 26809
rect 24918 26809 24930 26812
rect 24964 26840 24976 26843
rect 25314 26840 25320 26852
rect 24964 26812 25320 26840
rect 24964 26809 24976 26812
rect 24918 26803 24976 26809
rect 25314 26800 25320 26812
rect 25372 26800 25378 26852
rect 27890 26840 27896 26852
rect 27803 26812 27896 26840
rect 27890 26800 27896 26812
rect 27948 26840 27954 26852
rect 28169 26843 28227 26849
rect 28169 26840 28181 26843
rect 27948 26812 28181 26840
rect 27948 26800 27954 26812
rect 28169 26809 28181 26812
rect 28215 26809 28227 26843
rect 28169 26803 28227 26809
rect 28736 26784 28764 26880
rect 29540 26871 29552 26880
rect 29546 26868 29552 26871
rect 29604 26868 29610 26920
rect 32030 26917 32036 26920
rect 31757 26911 31815 26917
rect 31757 26877 31769 26911
rect 31803 26877 31815 26911
rect 32024 26908 32036 26917
rect 31991 26880 32036 26908
rect 31757 26871 31815 26877
rect 32024 26871 32036 26880
rect 31665 26843 31723 26849
rect 31665 26809 31677 26843
rect 31711 26840 31723 26843
rect 31772 26840 31800 26871
rect 32030 26868 32036 26871
rect 32088 26868 32094 26920
rect 34977 26911 35035 26917
rect 34977 26877 34989 26911
rect 35023 26877 35035 26911
rect 34977 26871 35035 26877
rect 35244 26911 35302 26917
rect 35244 26877 35256 26911
rect 35290 26908 35302 26911
rect 35526 26908 35532 26920
rect 35290 26880 35532 26908
rect 35290 26877 35302 26880
rect 35244 26871 35302 26877
rect 32398 26840 32404 26852
rect 31711 26812 32404 26840
rect 31711 26809 31723 26812
rect 31665 26803 31723 26809
rect 32398 26800 32404 26812
rect 32456 26800 32462 26852
rect 33870 26800 33876 26852
rect 33928 26840 33934 26852
rect 33965 26843 34023 26849
rect 33965 26840 33977 26843
rect 33928 26812 33977 26840
rect 33928 26800 33934 26812
rect 33965 26809 33977 26812
rect 34011 26840 34023 26843
rect 34992 26840 35020 26871
rect 35526 26868 35532 26880
rect 35584 26868 35590 26920
rect 34011 26812 35020 26840
rect 34011 26809 34023 26812
rect 33965 26803 34023 26809
rect 34624 26784 34652 26812
rect 35618 26800 35624 26852
rect 35676 26800 35682 26852
rect 21821 26775 21879 26781
rect 21821 26741 21833 26775
rect 21867 26772 21879 26775
rect 22002 26772 22008 26784
rect 21867 26744 22008 26772
rect 21867 26741 21879 26744
rect 21821 26735 21879 26741
rect 22002 26732 22008 26744
rect 22060 26732 22066 26784
rect 22278 26772 22284 26784
rect 22239 26744 22284 26772
rect 22278 26732 22284 26744
rect 22336 26732 22342 26784
rect 22738 26732 22744 26784
rect 22796 26772 22802 26784
rect 23106 26772 23112 26784
rect 22796 26744 23112 26772
rect 22796 26732 22802 26744
rect 23106 26732 23112 26744
rect 23164 26732 23170 26784
rect 26050 26772 26056 26784
rect 26011 26744 26056 26772
rect 26050 26732 26056 26744
rect 26108 26732 26114 26784
rect 27522 26732 27528 26784
rect 27580 26772 27586 26784
rect 28353 26775 28411 26781
rect 28353 26772 28365 26775
rect 27580 26744 28365 26772
rect 27580 26732 27586 26744
rect 28353 26741 28365 26744
rect 28399 26741 28411 26775
rect 28718 26772 28724 26784
rect 28679 26744 28724 26772
rect 28353 26735 28411 26741
rect 28718 26732 28724 26744
rect 28776 26732 28782 26784
rect 29089 26775 29147 26781
rect 29089 26741 29101 26775
rect 29135 26772 29147 26775
rect 29178 26772 29184 26784
rect 29135 26744 29184 26772
rect 29135 26741 29147 26744
rect 29089 26735 29147 26741
rect 29178 26732 29184 26744
rect 29236 26732 29242 26784
rect 30650 26772 30656 26784
rect 30611 26744 30656 26772
rect 30650 26732 30656 26744
rect 30708 26732 30714 26784
rect 34238 26772 34244 26784
rect 34199 26744 34244 26772
rect 34238 26732 34244 26744
rect 34296 26732 34302 26784
rect 34606 26772 34612 26784
rect 34567 26744 34612 26772
rect 34606 26732 34612 26744
rect 34664 26732 34670 26784
rect 35636 26772 35664 26800
rect 35802 26772 35808 26784
rect 35636 26744 35808 26772
rect 35802 26732 35808 26744
rect 35860 26732 35866 26784
rect 1104 26682 38824 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 38824 26682
rect 1104 26608 38824 26630
rect 21910 26528 21916 26580
rect 21968 26568 21974 26580
rect 22833 26571 22891 26577
rect 22833 26568 22845 26571
rect 21968 26540 22845 26568
rect 21968 26528 21974 26540
rect 22833 26537 22845 26540
rect 22879 26568 22891 26571
rect 23753 26571 23811 26577
rect 23753 26568 23765 26571
rect 22879 26540 23765 26568
rect 22879 26537 22891 26540
rect 22833 26531 22891 26537
rect 23753 26537 23765 26540
rect 23799 26537 23811 26571
rect 27890 26568 27896 26580
rect 27851 26540 27896 26568
rect 23753 26531 23811 26537
rect 21720 26503 21778 26509
rect 21720 26469 21732 26503
rect 21766 26500 21778 26503
rect 22278 26500 22284 26512
rect 21766 26472 22284 26500
rect 21766 26469 21778 26472
rect 21720 26463 21778 26469
rect 22278 26460 22284 26472
rect 22336 26460 22342 26512
rect 23768 26500 23796 26531
rect 27890 26528 27896 26540
rect 27948 26528 27954 26580
rect 29546 26528 29552 26580
rect 29604 26568 29610 26580
rect 30377 26571 30435 26577
rect 30377 26568 30389 26571
rect 29604 26540 30389 26568
rect 29604 26528 29610 26540
rect 30377 26537 30389 26540
rect 30423 26537 30435 26571
rect 30377 26531 30435 26537
rect 33870 26528 33876 26580
rect 33928 26568 33934 26580
rect 34425 26571 34483 26577
rect 34425 26568 34437 26571
rect 33928 26540 34437 26568
rect 33928 26528 33934 26540
rect 34425 26537 34437 26540
rect 34471 26568 34483 26571
rect 35526 26568 35532 26580
rect 34471 26540 35532 26568
rect 34471 26537 34483 26540
rect 34425 26531 34483 26537
rect 35526 26528 35532 26540
rect 35584 26568 35590 26580
rect 36265 26571 36323 26577
rect 36265 26568 36277 26571
rect 35584 26540 36277 26568
rect 35584 26528 35590 26540
rect 36265 26537 36277 26540
rect 36311 26537 36323 26571
rect 36265 26531 36323 26537
rect 24182 26503 24240 26509
rect 24182 26500 24194 26503
rect 23768 26472 24194 26500
rect 24182 26469 24194 26472
rect 24228 26469 24240 26503
rect 27908 26500 27936 26528
rect 29242 26503 29300 26509
rect 29242 26500 29254 26503
rect 24182 26463 24240 26469
rect 26528 26472 26924 26500
rect 27908 26472 29254 26500
rect 26528 26444 26556 26472
rect 23937 26435 23995 26441
rect 23937 26432 23949 26435
rect 21468 26404 23949 26432
rect 20898 26324 20904 26376
rect 20956 26364 20962 26376
rect 21468 26373 21496 26404
rect 23937 26401 23949 26404
rect 23983 26432 23995 26435
rect 24670 26432 24676 26444
rect 23983 26404 24676 26432
rect 23983 26401 23995 26404
rect 23937 26395 23995 26401
rect 24670 26392 24676 26404
rect 24728 26392 24734 26444
rect 26510 26432 26516 26444
rect 26423 26404 26516 26432
rect 26510 26392 26516 26404
rect 26568 26392 26574 26444
rect 26786 26441 26792 26444
rect 26780 26432 26792 26441
rect 26747 26404 26792 26432
rect 26780 26395 26792 26404
rect 26786 26392 26792 26395
rect 26844 26392 26850 26444
rect 26896 26432 26924 26472
rect 29242 26469 29254 26472
rect 29288 26469 29300 26503
rect 29242 26463 29300 26469
rect 29362 26460 29368 26512
rect 29420 26460 29426 26512
rect 31573 26503 31631 26509
rect 31573 26469 31585 26503
rect 31619 26500 31631 26503
rect 32030 26500 32036 26512
rect 31619 26472 32036 26500
rect 31619 26469 31631 26472
rect 31573 26463 31631 26469
rect 32030 26460 32036 26472
rect 32088 26460 32094 26512
rect 32668 26503 32726 26509
rect 32668 26469 32680 26503
rect 32714 26500 32726 26503
rect 32858 26500 32864 26512
rect 32714 26472 32864 26500
rect 32714 26469 32726 26472
rect 32668 26463 32726 26469
rect 32858 26460 32864 26472
rect 32916 26460 32922 26512
rect 35152 26503 35210 26509
rect 35152 26469 35164 26503
rect 35198 26500 35210 26503
rect 35250 26500 35256 26512
rect 35198 26472 35256 26500
rect 35198 26469 35210 26472
rect 35152 26463 35210 26469
rect 35250 26460 35256 26472
rect 35308 26460 35314 26512
rect 28442 26432 28448 26444
rect 26896 26404 28448 26432
rect 28442 26392 28448 26404
rect 28500 26432 28506 26444
rect 28997 26435 29055 26441
rect 28997 26432 29009 26435
rect 28500 26404 29009 26432
rect 28500 26392 28506 26404
rect 28997 26401 29009 26404
rect 29043 26432 29055 26435
rect 29380 26432 29408 26460
rect 29043 26404 29408 26432
rect 29043 26401 29055 26404
rect 28997 26395 29055 26401
rect 21453 26367 21511 26373
rect 21453 26364 21465 26367
rect 20956 26336 21465 26364
rect 20956 26324 20962 26336
rect 21453 26333 21465 26336
rect 21499 26333 21511 26367
rect 32398 26364 32404 26376
rect 32359 26336 32404 26364
rect 21453 26327 21511 26333
rect 32398 26324 32404 26336
rect 32456 26324 32462 26376
rect 34606 26324 34612 26376
rect 34664 26364 34670 26376
rect 34885 26367 34943 26373
rect 34885 26364 34897 26367
rect 34664 26336 34897 26364
rect 34664 26324 34670 26336
rect 34885 26333 34897 26336
rect 34931 26333 34943 26367
rect 34885 26327 34943 26333
rect 25317 26299 25375 26305
rect 25317 26296 25329 26299
rect 24872 26268 25329 26296
rect 21174 26228 21180 26240
rect 21135 26200 21180 26228
rect 21174 26188 21180 26200
rect 21232 26188 21238 26240
rect 24578 26188 24584 26240
rect 24636 26228 24642 26240
rect 24872 26228 24900 26268
rect 25317 26265 25329 26268
rect 25363 26265 25375 26299
rect 28537 26299 28595 26305
rect 28537 26296 28549 26299
rect 25317 26259 25375 26265
rect 27540 26268 28549 26296
rect 24636 26200 24900 26228
rect 24636 26188 24642 26200
rect 27430 26188 27436 26240
rect 27488 26228 27494 26240
rect 27540 26228 27568 26268
rect 28537 26265 28549 26268
rect 28583 26296 28595 26299
rect 28902 26296 28908 26308
rect 28583 26268 28908 26296
rect 28583 26265 28595 26268
rect 28537 26259 28595 26265
rect 28902 26256 28908 26268
rect 28960 26256 28966 26308
rect 31846 26296 31852 26308
rect 31807 26268 31852 26296
rect 31846 26256 31852 26268
rect 31904 26256 31910 26308
rect 33410 26256 33416 26308
rect 33468 26296 33474 26308
rect 33781 26299 33839 26305
rect 33781 26296 33793 26299
rect 33468 26268 33793 26296
rect 33468 26256 33474 26268
rect 33781 26265 33793 26268
rect 33827 26296 33839 26299
rect 34238 26296 34244 26308
rect 33827 26268 34244 26296
rect 33827 26265 33839 26268
rect 33781 26259 33839 26265
rect 34238 26256 34244 26268
rect 34296 26256 34302 26308
rect 34698 26228 34704 26240
rect 27488 26200 27568 26228
rect 34659 26200 34704 26228
rect 27488 26188 27494 26200
rect 34698 26188 34704 26200
rect 34756 26188 34762 26240
rect 1104 26138 38824 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 34966 26138
rect 35018 26086 35030 26138
rect 35082 26086 35094 26138
rect 35146 26086 35158 26138
rect 35210 26086 38824 26138
rect 1104 26064 38824 26086
rect 20441 26027 20499 26033
rect 20441 25993 20453 26027
rect 20487 26024 20499 26027
rect 20809 26027 20867 26033
rect 20809 26024 20821 26027
rect 20487 25996 20821 26024
rect 20487 25993 20499 25996
rect 20441 25987 20499 25993
rect 20809 25993 20821 25996
rect 20855 26024 20867 26027
rect 20898 26024 20904 26036
rect 20855 25996 20904 26024
rect 20855 25993 20867 25996
rect 20809 25987 20867 25993
rect 20898 25984 20904 25996
rect 20956 25984 20962 26036
rect 22278 26024 22284 26036
rect 22191 25996 22284 26024
rect 22278 25984 22284 25996
rect 22336 26024 22342 26036
rect 22833 26027 22891 26033
rect 22833 26024 22845 26027
rect 22336 25996 22845 26024
rect 22336 25984 22342 25996
rect 22833 25993 22845 25996
rect 22879 25993 22891 26027
rect 25314 26024 25320 26036
rect 25275 25996 25320 26024
rect 22833 25987 22891 25993
rect 25314 25984 25320 25996
rect 25372 25984 25378 26036
rect 27890 25984 27896 26036
rect 27948 26024 27954 26036
rect 28629 26027 28687 26033
rect 28629 26024 28641 26027
rect 27948 25996 28641 26024
rect 27948 25984 27954 25996
rect 28629 25993 28641 25996
rect 28675 25993 28687 26027
rect 28629 25987 28687 25993
rect 28994 25984 29000 26036
rect 29052 26024 29058 26036
rect 29457 26027 29515 26033
rect 29457 26024 29469 26027
rect 29052 25996 29469 26024
rect 29052 25984 29058 25996
rect 29457 25993 29469 25996
rect 29503 25993 29515 26027
rect 29457 25987 29515 25993
rect 31757 26027 31815 26033
rect 31757 25993 31769 26027
rect 31803 26024 31815 26027
rect 32030 26024 32036 26036
rect 31803 25996 32036 26024
rect 31803 25993 31815 25996
rect 31757 25987 31815 25993
rect 32030 25984 32036 25996
rect 32088 25984 32094 26036
rect 20916 25897 20944 25984
rect 34790 25916 34796 25968
rect 34848 25956 34854 25968
rect 34885 25959 34943 25965
rect 34885 25956 34897 25959
rect 34848 25928 34897 25956
rect 34848 25916 34854 25928
rect 34885 25925 34897 25928
rect 34931 25956 34943 25959
rect 36078 25956 36084 25968
rect 34931 25928 36084 25956
rect 34931 25925 34943 25928
rect 34885 25919 34943 25925
rect 36078 25916 36084 25928
rect 36136 25916 36142 25968
rect 20901 25891 20959 25897
rect 20901 25857 20913 25891
rect 20947 25857 20959 25891
rect 33870 25888 33876 25900
rect 33831 25860 33876 25888
rect 20901 25851 20959 25857
rect 33870 25848 33876 25860
rect 33928 25848 33934 25900
rect 35250 25848 35256 25900
rect 35308 25888 35314 25900
rect 35437 25891 35495 25897
rect 35437 25888 35449 25891
rect 35308 25860 35449 25888
rect 35308 25848 35314 25860
rect 35437 25857 35449 25860
rect 35483 25888 35495 25891
rect 35897 25891 35955 25897
rect 35897 25888 35909 25891
rect 35483 25860 35909 25888
rect 35483 25857 35495 25860
rect 35437 25851 35495 25857
rect 35897 25857 35909 25860
rect 35943 25888 35955 25891
rect 36265 25891 36323 25897
rect 36265 25888 36277 25891
rect 35943 25860 36277 25888
rect 35943 25857 35955 25860
rect 35897 25851 35955 25857
rect 36265 25857 36277 25860
rect 36311 25857 36323 25891
rect 36265 25851 36323 25857
rect 23477 25823 23535 25829
rect 23477 25789 23489 25823
rect 23523 25820 23535 25823
rect 23937 25823 23995 25829
rect 23937 25820 23949 25823
rect 23523 25792 23949 25820
rect 23523 25789 23535 25792
rect 23477 25783 23535 25789
rect 23937 25789 23949 25792
rect 23983 25820 23995 25823
rect 24026 25820 24032 25832
rect 23983 25792 24032 25820
rect 23983 25789 23995 25792
rect 23937 25783 23995 25789
rect 24026 25780 24032 25792
rect 24084 25820 24090 25832
rect 24670 25820 24676 25832
rect 24084 25792 24676 25820
rect 24084 25780 24090 25792
rect 24670 25780 24676 25792
rect 24728 25820 24734 25832
rect 25961 25823 26019 25829
rect 25961 25820 25973 25823
rect 24728 25792 25973 25820
rect 24728 25780 24734 25792
rect 25961 25789 25973 25792
rect 26007 25820 26019 25823
rect 26329 25823 26387 25829
rect 26329 25820 26341 25823
rect 26007 25792 26341 25820
rect 26007 25789 26019 25792
rect 25961 25783 26019 25789
rect 26329 25789 26341 25792
rect 26375 25820 26387 25823
rect 26421 25823 26479 25829
rect 26421 25820 26433 25823
rect 26375 25792 26433 25820
rect 26375 25789 26387 25792
rect 26329 25783 26387 25789
rect 26421 25789 26433 25792
rect 26467 25820 26479 25823
rect 26510 25820 26516 25832
rect 26467 25792 26516 25820
rect 26467 25789 26479 25792
rect 26421 25783 26479 25789
rect 26510 25780 26516 25792
rect 26568 25780 26574 25832
rect 29270 25820 29276 25832
rect 29231 25792 29276 25820
rect 29270 25780 29276 25792
rect 29328 25780 29334 25832
rect 30374 25820 30380 25832
rect 30335 25792 30380 25820
rect 30374 25780 30380 25792
rect 30432 25780 30438 25832
rect 30650 25829 30656 25832
rect 30644 25820 30656 25829
rect 30484 25792 30656 25820
rect 21174 25761 21180 25764
rect 21168 25752 21180 25761
rect 21087 25724 21180 25752
rect 21168 25715 21180 25724
rect 21232 25752 21238 25764
rect 21542 25752 21548 25764
rect 21232 25724 21548 25752
rect 21174 25712 21180 25715
rect 21232 25712 21238 25724
rect 21542 25712 21548 25724
rect 21600 25712 21606 25764
rect 24204 25755 24262 25761
rect 24204 25721 24216 25755
rect 24250 25752 24262 25755
rect 24578 25752 24584 25764
rect 24250 25724 24584 25752
rect 24250 25721 24262 25724
rect 24204 25715 24262 25721
rect 24578 25712 24584 25724
rect 24636 25712 24642 25764
rect 26050 25712 26056 25764
rect 26108 25752 26114 25764
rect 26666 25755 26724 25761
rect 26666 25752 26678 25755
rect 26108 25724 26678 25752
rect 26108 25712 26114 25724
rect 26666 25721 26678 25724
rect 26712 25721 26724 25755
rect 26666 25715 26724 25721
rect 29917 25755 29975 25761
rect 29917 25721 29929 25755
rect 29963 25752 29975 25755
rect 30282 25752 30288 25764
rect 29963 25724 30288 25752
rect 29963 25721 29975 25724
rect 29917 25715 29975 25721
rect 30282 25712 30288 25724
rect 30340 25752 30346 25764
rect 30484 25752 30512 25792
rect 30644 25783 30656 25792
rect 30650 25780 30656 25783
rect 30708 25780 30714 25832
rect 32398 25820 32404 25832
rect 32311 25792 32404 25820
rect 32398 25780 32404 25792
rect 32456 25820 32462 25832
rect 34606 25820 34612 25832
rect 32456 25792 34612 25820
rect 32456 25780 32462 25792
rect 34606 25780 34612 25792
rect 34664 25780 34670 25832
rect 34698 25780 34704 25832
rect 34756 25820 34762 25832
rect 35345 25823 35403 25829
rect 35345 25820 35357 25823
rect 34756 25792 35357 25820
rect 34756 25780 34762 25792
rect 35345 25789 35357 25792
rect 35391 25789 35403 25823
rect 35345 25783 35403 25789
rect 30340 25724 30512 25752
rect 30340 25712 30346 25724
rect 27798 25684 27804 25696
rect 27759 25656 27804 25684
rect 27798 25644 27804 25656
rect 27856 25644 27862 25696
rect 29089 25687 29147 25693
rect 29089 25653 29101 25687
rect 29135 25684 29147 25687
rect 29178 25684 29184 25696
rect 29135 25656 29184 25684
rect 29135 25653 29147 25656
rect 29089 25647 29147 25653
rect 29178 25644 29184 25656
rect 29236 25684 29242 25696
rect 30193 25687 30251 25693
rect 30193 25684 30205 25687
rect 29236 25656 30205 25684
rect 29236 25644 29242 25656
rect 30193 25653 30205 25656
rect 30239 25684 30251 25687
rect 30374 25684 30380 25696
rect 30239 25656 30380 25684
rect 30239 25653 30251 25656
rect 30193 25647 30251 25653
rect 30374 25644 30380 25656
rect 30432 25684 30438 25696
rect 32122 25684 32128 25696
rect 30432 25656 32128 25684
rect 30432 25644 30438 25656
rect 32122 25644 32128 25656
rect 32180 25684 32186 25696
rect 32416 25693 32444 25780
rect 33137 25755 33195 25761
rect 33137 25721 33149 25755
rect 33183 25752 33195 25755
rect 33597 25755 33655 25761
rect 33597 25752 33609 25755
rect 33183 25724 33609 25752
rect 33183 25721 33195 25724
rect 33137 25715 33195 25721
rect 33597 25721 33609 25724
rect 33643 25752 33655 25755
rect 34333 25755 34391 25761
rect 33643 25724 34284 25752
rect 33643 25721 33655 25724
rect 33597 25715 33655 25721
rect 32401 25687 32459 25693
rect 32401 25684 32413 25687
rect 32180 25656 32413 25684
rect 32180 25644 32186 25656
rect 32401 25653 32413 25656
rect 32447 25653 32459 25687
rect 33226 25684 33232 25696
rect 33187 25656 33232 25684
rect 32401 25647 32459 25653
rect 33226 25644 33232 25656
rect 33284 25644 33290 25696
rect 33686 25684 33692 25696
rect 33647 25656 33692 25684
rect 33686 25644 33692 25656
rect 33744 25644 33750 25696
rect 34256 25684 34284 25724
rect 34333 25721 34345 25755
rect 34379 25752 34391 25755
rect 35253 25755 35311 25761
rect 35253 25752 35265 25755
rect 34379 25724 35265 25752
rect 34379 25721 34391 25724
rect 34333 25715 34391 25721
rect 35253 25721 35265 25724
rect 35299 25752 35311 25755
rect 36449 25755 36507 25761
rect 36449 25752 36461 25755
rect 35299 25724 36461 25752
rect 35299 25721 35311 25724
rect 35253 25715 35311 25721
rect 36449 25721 36461 25724
rect 36495 25721 36507 25755
rect 36449 25715 36507 25721
rect 35158 25684 35164 25696
rect 34256 25656 35164 25684
rect 35158 25644 35164 25656
rect 35216 25644 35222 25696
rect 1104 25594 38824 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 38824 25594
rect 1104 25520 38824 25542
rect 24026 25480 24032 25492
rect 23987 25452 24032 25480
rect 24026 25440 24032 25452
rect 24084 25440 24090 25492
rect 24489 25483 24547 25489
rect 24489 25449 24501 25483
rect 24535 25480 24547 25483
rect 24670 25480 24676 25492
rect 24535 25452 24676 25480
rect 24535 25449 24547 25452
rect 24489 25443 24547 25449
rect 24670 25440 24676 25452
rect 24728 25480 24734 25492
rect 25314 25480 25320 25492
rect 24728 25452 25320 25480
rect 24728 25440 24734 25452
rect 25314 25440 25320 25452
rect 25372 25440 25378 25492
rect 26050 25440 26056 25492
rect 26108 25480 26114 25492
rect 26237 25483 26295 25489
rect 26237 25480 26249 25483
rect 26108 25452 26249 25480
rect 26108 25440 26114 25452
rect 26237 25449 26249 25452
rect 26283 25449 26295 25483
rect 26237 25443 26295 25449
rect 26973 25483 27031 25489
rect 26973 25449 26985 25483
rect 27019 25480 27031 25483
rect 27430 25480 27436 25492
rect 27019 25452 27436 25480
rect 27019 25449 27031 25452
rect 26973 25443 27031 25449
rect 27430 25440 27436 25452
rect 27488 25440 27494 25492
rect 27893 25483 27951 25489
rect 27893 25449 27905 25483
rect 27939 25480 27951 25483
rect 29270 25480 29276 25492
rect 27939 25452 29276 25480
rect 27939 25449 27951 25452
rect 27893 25443 27951 25449
rect 29270 25440 29276 25452
rect 29328 25440 29334 25492
rect 29546 25480 29552 25492
rect 29507 25452 29552 25480
rect 29546 25440 29552 25452
rect 29604 25440 29610 25492
rect 29917 25483 29975 25489
rect 29917 25449 29929 25483
rect 29963 25480 29975 25483
rect 30098 25480 30104 25492
rect 29963 25452 30104 25480
rect 29963 25449 29975 25452
rect 29917 25443 29975 25449
rect 30098 25440 30104 25452
rect 30156 25440 30162 25492
rect 32674 25480 32680 25492
rect 32635 25452 32680 25480
rect 32674 25440 32680 25452
rect 32732 25440 32738 25492
rect 33686 25480 33692 25492
rect 33647 25452 33692 25480
rect 33686 25440 33692 25452
rect 33744 25440 33750 25492
rect 23661 25415 23719 25421
rect 23661 25381 23673 25415
rect 23707 25412 23719 25415
rect 24578 25412 24584 25424
rect 23707 25384 24584 25412
rect 23707 25381 23719 25384
rect 23661 25375 23719 25381
rect 24578 25372 24584 25384
rect 24636 25372 24642 25424
rect 25225 25415 25283 25421
rect 25225 25381 25237 25415
rect 25271 25412 25283 25415
rect 25498 25412 25504 25424
rect 25271 25384 25504 25412
rect 25271 25381 25283 25384
rect 25225 25375 25283 25381
rect 25498 25372 25504 25384
rect 25556 25412 25562 25424
rect 26068 25412 26096 25440
rect 25556 25384 26096 25412
rect 25556 25372 25562 25384
rect 28994 25372 29000 25424
rect 29052 25412 29058 25424
rect 30009 25415 30067 25421
rect 30009 25412 30021 25415
rect 29052 25384 30021 25412
rect 29052 25372 29058 25384
rect 30009 25381 30021 25384
rect 30055 25412 30067 25415
rect 30466 25412 30472 25424
rect 30055 25384 30472 25412
rect 30055 25381 30067 25384
rect 30009 25375 30067 25381
rect 30466 25372 30472 25384
rect 30524 25372 30530 25424
rect 32493 25415 32551 25421
rect 32493 25381 32505 25415
rect 32539 25412 32551 25415
rect 32858 25412 32864 25424
rect 32539 25384 32864 25412
rect 32539 25381 32551 25384
rect 32493 25375 32551 25381
rect 32858 25372 32864 25384
rect 32916 25372 32922 25424
rect 20898 25344 20904 25356
rect 20859 25316 20904 25344
rect 20898 25304 20904 25316
rect 20956 25304 20962 25356
rect 21174 25353 21180 25356
rect 21168 25344 21180 25353
rect 21135 25316 21180 25344
rect 21168 25307 21180 25316
rect 21174 25304 21180 25307
rect 21232 25304 21238 25356
rect 26694 25304 26700 25356
rect 26752 25344 26758 25356
rect 26789 25347 26847 25353
rect 26789 25344 26801 25347
rect 26752 25316 26801 25344
rect 26752 25304 26758 25316
rect 26789 25313 26801 25316
rect 26835 25313 26847 25347
rect 28258 25344 28264 25356
rect 28219 25316 28264 25344
rect 26789 25307 26847 25313
rect 28258 25304 28264 25316
rect 28316 25304 28322 25356
rect 33042 25344 33048 25356
rect 33003 25316 33048 25344
rect 33042 25304 33048 25316
rect 33100 25304 33106 25356
rect 34333 25347 34391 25353
rect 34333 25313 34345 25347
rect 34379 25344 34391 25347
rect 34379 25316 34928 25344
rect 34379 25313 34391 25316
rect 34333 25307 34391 25313
rect 34900 25288 34928 25316
rect 24118 25236 24124 25288
rect 24176 25276 24182 25288
rect 24673 25279 24731 25285
rect 24673 25276 24685 25279
rect 24176 25248 24685 25276
rect 24176 25236 24182 25248
rect 24673 25245 24685 25248
rect 24719 25276 24731 25279
rect 25501 25279 25559 25285
rect 25501 25276 25513 25279
rect 24719 25248 25513 25276
rect 24719 25245 24731 25248
rect 24673 25239 24731 25245
rect 25501 25245 25513 25248
rect 25547 25276 25559 25279
rect 25590 25276 25596 25288
rect 25547 25248 25596 25276
rect 25547 25245 25559 25248
rect 25501 25239 25559 25245
rect 25590 25236 25596 25248
rect 25648 25236 25654 25288
rect 28350 25276 28356 25288
rect 28311 25248 28356 25276
rect 28350 25236 28356 25248
rect 28408 25236 28414 25288
rect 28537 25279 28595 25285
rect 28537 25245 28549 25279
rect 28583 25276 28595 25279
rect 28718 25276 28724 25288
rect 28583 25248 28724 25276
rect 28583 25245 28595 25248
rect 28537 25239 28595 25245
rect 28718 25236 28724 25248
rect 28776 25236 28782 25288
rect 30193 25279 30251 25285
rect 30193 25245 30205 25279
rect 30239 25276 30251 25279
rect 30282 25276 30288 25288
rect 30239 25248 30288 25276
rect 30239 25245 30251 25248
rect 30193 25239 30251 25245
rect 30282 25236 30288 25248
rect 30340 25236 30346 25288
rect 32674 25236 32680 25288
rect 32732 25276 32738 25288
rect 33137 25279 33195 25285
rect 33137 25276 33149 25279
rect 32732 25248 33149 25276
rect 32732 25236 32738 25248
rect 33137 25245 33149 25248
rect 33183 25245 33195 25279
rect 33318 25276 33324 25288
rect 33279 25248 33324 25276
rect 33137 25239 33195 25245
rect 33318 25236 33324 25248
rect 33376 25236 33382 25288
rect 34054 25236 34060 25288
rect 34112 25276 34118 25288
rect 34425 25279 34483 25285
rect 34425 25276 34437 25279
rect 34112 25248 34437 25276
rect 34112 25236 34118 25248
rect 34425 25245 34437 25248
rect 34471 25245 34483 25279
rect 34425 25239 34483 25245
rect 34606 25236 34612 25288
rect 34664 25276 34670 25288
rect 34748 25279 34806 25285
rect 34748 25276 34760 25279
rect 34664 25248 34760 25276
rect 34664 25236 34670 25248
rect 34748 25245 34760 25248
rect 34794 25245 34806 25279
rect 34748 25239 34806 25245
rect 34882 25236 34888 25288
rect 34940 25276 34946 25288
rect 35158 25276 35164 25288
rect 34940 25248 35033 25276
rect 35071 25248 35164 25276
rect 34940 25236 34946 25248
rect 35158 25236 35164 25248
rect 35216 25276 35222 25288
rect 35618 25276 35624 25288
rect 35216 25248 35624 25276
rect 35216 25236 35222 25248
rect 35618 25236 35624 25248
rect 35676 25236 35682 25288
rect 36262 25276 36268 25288
rect 36223 25248 36268 25276
rect 36262 25236 36268 25248
rect 36320 25236 36326 25288
rect 31938 25208 31944 25220
rect 31899 25180 31944 25208
rect 31938 25168 31944 25180
rect 31996 25168 32002 25220
rect 20622 25140 20628 25152
rect 20583 25112 20628 25140
rect 20622 25100 20628 25112
rect 20680 25100 20686 25152
rect 21542 25100 21548 25152
rect 21600 25140 21606 25152
rect 22281 25143 22339 25149
rect 22281 25140 22293 25143
rect 21600 25112 22293 25140
rect 21600 25100 21606 25112
rect 22281 25109 22293 25112
rect 22327 25109 22339 25143
rect 22281 25103 22339 25109
rect 24121 25143 24179 25149
rect 24121 25109 24133 25143
rect 24167 25140 24179 25143
rect 24762 25140 24768 25152
rect 24167 25112 24768 25140
rect 24167 25109 24179 25112
rect 24121 25103 24179 25109
rect 24762 25100 24768 25112
rect 24820 25100 24826 25152
rect 26234 25100 26240 25152
rect 26292 25140 26298 25152
rect 26786 25140 26792 25152
rect 26292 25112 26792 25140
rect 26292 25100 26298 25112
rect 26786 25100 26792 25112
rect 26844 25140 26850 25152
rect 27341 25143 27399 25149
rect 27341 25140 27353 25143
rect 26844 25112 27353 25140
rect 26844 25100 26850 25112
rect 27341 25109 27353 25112
rect 27387 25140 27399 25143
rect 27798 25140 27804 25152
rect 27387 25112 27804 25140
rect 27387 25109 27399 25112
rect 27341 25103 27399 25109
rect 27798 25100 27804 25112
rect 27856 25100 27862 25152
rect 1104 25050 38824 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 34966 25050
rect 35018 24998 35030 25050
rect 35082 24998 35094 25050
rect 35146 24998 35158 25050
rect 35210 24998 38824 25050
rect 1104 24976 38824 24998
rect 20441 24939 20499 24945
rect 20441 24905 20453 24939
rect 20487 24936 20499 24939
rect 20898 24936 20904 24948
rect 20487 24908 20904 24936
rect 20487 24905 20499 24908
rect 20441 24899 20499 24905
rect 20548 24812 20576 24908
rect 20898 24896 20904 24908
rect 20956 24896 20962 24948
rect 24670 24936 24676 24948
rect 24631 24908 24676 24936
rect 24670 24896 24676 24908
rect 24728 24896 24734 24948
rect 26694 24896 26700 24948
rect 26752 24936 26758 24948
rect 27617 24939 27675 24945
rect 27617 24936 27629 24939
rect 26752 24908 27629 24936
rect 26752 24896 26758 24908
rect 27617 24905 27629 24908
rect 27663 24936 27675 24939
rect 27985 24939 28043 24945
rect 27985 24936 27997 24939
rect 27663 24908 27997 24936
rect 27663 24905 27675 24908
rect 27617 24899 27675 24905
rect 27985 24905 27997 24908
rect 28031 24936 28043 24939
rect 28350 24936 28356 24948
rect 28031 24908 28356 24936
rect 28031 24905 28043 24908
rect 27985 24899 28043 24905
rect 28350 24896 28356 24908
rect 28408 24896 28414 24948
rect 29641 24939 29699 24945
rect 29641 24905 29653 24939
rect 29687 24936 29699 24939
rect 30098 24936 30104 24948
rect 29687 24908 30104 24936
rect 29687 24905 29699 24908
rect 29641 24899 29699 24905
rect 30098 24896 30104 24908
rect 30156 24896 30162 24948
rect 31757 24939 31815 24945
rect 31757 24905 31769 24939
rect 31803 24936 31815 24939
rect 34517 24939 34575 24945
rect 34517 24936 34529 24939
rect 31803 24908 34529 24936
rect 31803 24905 31815 24908
rect 31757 24899 31815 24905
rect 24305 24871 24363 24877
rect 24305 24837 24317 24871
rect 24351 24868 24363 24871
rect 24578 24868 24584 24880
rect 24351 24840 24584 24868
rect 24351 24837 24363 24840
rect 24305 24831 24363 24837
rect 24578 24828 24584 24840
rect 24636 24828 24642 24880
rect 30009 24871 30067 24877
rect 30009 24837 30021 24871
rect 30055 24868 30067 24871
rect 30282 24868 30288 24880
rect 30055 24840 30288 24868
rect 30055 24837 30067 24840
rect 30009 24831 30067 24837
rect 30282 24828 30288 24840
rect 30340 24828 30346 24880
rect 20530 24800 20536 24812
rect 20443 24772 20536 24800
rect 20530 24760 20536 24772
rect 20588 24760 20594 24812
rect 25590 24800 25596 24812
rect 25551 24772 25596 24800
rect 25590 24760 25596 24772
rect 25648 24760 25654 24812
rect 26418 24800 26424 24812
rect 26379 24772 26424 24800
rect 26418 24760 26424 24772
rect 26476 24800 26482 24812
rect 27154 24800 27160 24812
rect 26476 24772 27016 24800
rect 27115 24772 27160 24800
rect 26476 24760 26482 24772
rect 23661 24735 23719 24741
rect 23661 24732 23673 24735
rect 23492 24704 23673 24732
rect 20714 24624 20720 24676
rect 20772 24673 20778 24676
rect 20772 24667 20836 24673
rect 20772 24633 20790 24667
rect 20824 24633 20836 24667
rect 20772 24627 20836 24633
rect 20772 24624 20778 24627
rect 23492 24608 23520 24704
rect 23661 24701 23673 24704
rect 23707 24701 23719 24735
rect 23661 24695 23719 24701
rect 24854 24692 24860 24744
rect 24912 24732 24918 24744
rect 26053 24735 26111 24741
rect 26053 24732 26065 24735
rect 24912 24704 26065 24732
rect 24912 24692 24918 24704
rect 26053 24701 26065 24704
rect 26099 24732 26111 24735
rect 26878 24732 26884 24744
rect 26099 24704 26884 24732
rect 26099 24701 26111 24704
rect 26053 24695 26111 24701
rect 26878 24692 26884 24704
rect 26936 24692 26942 24744
rect 26988 24732 27016 24772
rect 27154 24760 27160 24772
rect 27212 24760 27218 24812
rect 31864 24800 31892 24908
rect 34517 24905 34529 24908
rect 34563 24936 34575 24939
rect 34606 24936 34612 24948
rect 34563 24908 34612 24936
rect 34563 24905 34575 24908
rect 34517 24899 34575 24905
rect 34606 24896 34612 24908
rect 34664 24896 34670 24948
rect 34790 24896 34796 24948
rect 34848 24936 34854 24948
rect 34885 24939 34943 24945
rect 34885 24936 34897 24939
rect 34848 24908 34897 24936
rect 34848 24896 34854 24908
rect 34885 24905 34897 24908
rect 34931 24905 34943 24939
rect 34885 24899 34943 24905
rect 33226 24828 33232 24880
rect 33284 24868 33290 24880
rect 33284 24840 34468 24868
rect 33284 24828 33290 24840
rect 32172 24803 32230 24809
rect 32172 24800 32184 24803
rect 31864 24772 32184 24800
rect 32172 24769 32184 24772
rect 32218 24769 32230 24803
rect 32172 24763 32230 24769
rect 32306 24760 32312 24812
rect 32364 24800 32370 24812
rect 32582 24800 32588 24812
rect 32364 24772 32409 24800
rect 32543 24772 32588 24800
rect 32364 24760 32370 24772
rect 32582 24760 32588 24772
rect 32640 24760 32646 24812
rect 34440 24800 34468 24840
rect 35345 24803 35403 24809
rect 35345 24800 35357 24803
rect 34440 24772 35357 24800
rect 35345 24769 35357 24772
rect 35391 24769 35403 24803
rect 35345 24763 35403 24769
rect 35529 24803 35587 24809
rect 35529 24769 35541 24803
rect 35575 24800 35587 24803
rect 35894 24800 35900 24812
rect 35575 24772 35900 24800
rect 35575 24769 35587 24772
rect 35529 24763 35587 24769
rect 27065 24735 27123 24741
rect 27065 24732 27077 24735
rect 26988 24704 27077 24732
rect 27065 24701 27077 24704
rect 27111 24701 27123 24735
rect 27065 24695 27123 24701
rect 30193 24735 30251 24741
rect 30193 24701 30205 24735
rect 30239 24732 30251 24735
rect 30745 24735 30803 24741
rect 30745 24732 30757 24735
rect 30239 24704 30757 24732
rect 30239 24701 30251 24704
rect 30193 24695 30251 24701
rect 30745 24701 30757 24704
rect 30791 24701 30803 24735
rect 31849 24735 31907 24741
rect 31849 24732 31861 24735
rect 30745 24695 30803 24701
rect 31312 24704 31861 24732
rect 26142 24664 26148 24676
rect 25424 24636 26148 24664
rect 25424 24608 25452 24636
rect 26142 24624 26148 24636
rect 26200 24624 26206 24676
rect 28258 24664 28264 24676
rect 26620 24636 28264 24664
rect 20073 24599 20131 24605
rect 20073 24565 20085 24599
rect 20119 24596 20131 24599
rect 20254 24596 20260 24608
rect 20119 24568 20260 24596
rect 20119 24565 20131 24568
rect 20073 24559 20131 24565
rect 20254 24556 20260 24568
rect 20312 24556 20318 24608
rect 21910 24596 21916 24608
rect 21871 24568 21916 24596
rect 21910 24556 21916 24568
rect 21968 24556 21974 24608
rect 23474 24596 23480 24608
rect 23435 24568 23480 24596
rect 23474 24556 23480 24568
rect 23532 24556 23538 24608
rect 23842 24596 23848 24608
rect 23803 24568 23848 24596
rect 23842 24556 23848 24568
rect 23900 24556 23906 24608
rect 25038 24596 25044 24608
rect 24999 24568 25044 24596
rect 25038 24556 25044 24568
rect 25096 24556 25102 24608
rect 25406 24596 25412 24608
rect 25367 24568 25412 24596
rect 25406 24556 25412 24568
rect 25464 24556 25470 24608
rect 25498 24556 25504 24608
rect 25556 24596 25562 24608
rect 26620 24605 26648 24636
rect 28258 24624 28264 24636
rect 28316 24664 28322 24676
rect 28353 24667 28411 24673
rect 28353 24664 28365 24667
rect 28316 24636 28365 24664
rect 28316 24624 28322 24636
rect 28353 24633 28365 24636
rect 28399 24664 28411 24667
rect 30208 24664 30236 24695
rect 28399 24636 30236 24664
rect 28399 24633 28411 24636
rect 28353 24627 28411 24633
rect 30926 24624 30932 24676
rect 30984 24664 30990 24676
rect 31312 24673 31340 24704
rect 31849 24701 31861 24704
rect 31895 24701 31907 24735
rect 35360 24732 35388 24763
rect 35894 24760 35900 24772
rect 35952 24760 35958 24812
rect 36265 24735 36323 24741
rect 36265 24732 36277 24735
rect 35360 24704 36277 24732
rect 31849 24695 31907 24701
rect 36265 24701 36277 24704
rect 36311 24701 36323 24735
rect 36265 24695 36323 24701
rect 31297 24667 31355 24673
rect 31297 24664 31309 24667
rect 30984 24636 31309 24664
rect 30984 24624 30990 24636
rect 31297 24633 31309 24636
rect 31343 24633 31355 24667
rect 31297 24627 31355 24633
rect 34974 24624 34980 24676
rect 35032 24664 35038 24676
rect 35253 24667 35311 24673
rect 35253 24664 35265 24667
rect 35032 24636 35265 24664
rect 35032 24624 35038 24636
rect 35253 24633 35265 24636
rect 35299 24664 35311 24667
rect 35710 24664 35716 24676
rect 35299 24636 35716 24664
rect 35299 24633 35311 24636
rect 35253 24627 35311 24633
rect 35710 24624 35716 24636
rect 35768 24624 35774 24676
rect 26605 24599 26663 24605
rect 25556 24568 25601 24596
rect 25556 24556 25562 24568
rect 26605 24565 26617 24599
rect 26651 24565 26663 24599
rect 26605 24559 26663 24565
rect 26878 24556 26884 24608
rect 26936 24596 26942 24608
rect 26973 24599 27031 24605
rect 26973 24596 26985 24599
rect 26936 24568 26985 24596
rect 26936 24556 26942 24568
rect 26973 24565 26985 24568
rect 27019 24565 27031 24599
rect 28718 24596 28724 24608
rect 28679 24568 28724 24596
rect 26973 24559 27031 24565
rect 28718 24556 28724 24568
rect 28776 24556 28782 24608
rect 30374 24596 30380 24608
rect 30335 24568 30380 24596
rect 30374 24556 30380 24568
rect 30432 24556 30438 24608
rect 32674 24556 32680 24608
rect 32732 24596 32738 24608
rect 33689 24599 33747 24605
rect 33689 24596 33701 24599
rect 32732 24568 33701 24596
rect 32732 24556 32738 24568
rect 33689 24565 33701 24568
rect 33735 24565 33747 24599
rect 33689 24559 33747 24565
rect 1104 24506 38824 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 38824 24506
rect 1104 24432 38824 24454
rect 20530 24392 20536 24404
rect 20491 24364 20536 24392
rect 20530 24352 20536 24364
rect 20588 24352 20594 24404
rect 22738 24392 22744 24404
rect 22699 24364 22744 24392
rect 22738 24352 22744 24364
rect 22796 24352 22802 24404
rect 24302 24392 24308 24404
rect 24263 24364 24308 24392
rect 24302 24352 24308 24364
rect 24360 24352 24366 24404
rect 24673 24395 24731 24401
rect 24673 24361 24685 24395
rect 24719 24392 24731 24395
rect 25038 24392 25044 24404
rect 24719 24364 25044 24392
rect 24719 24361 24731 24364
rect 24673 24355 24731 24361
rect 25038 24352 25044 24364
rect 25096 24352 25102 24404
rect 25406 24392 25412 24404
rect 25367 24364 25412 24392
rect 25406 24352 25412 24364
rect 25464 24352 25470 24404
rect 26142 24352 26148 24404
rect 26200 24392 26206 24404
rect 26789 24395 26847 24401
rect 26789 24392 26801 24395
rect 26200 24364 26801 24392
rect 26200 24352 26206 24364
rect 26789 24361 26801 24364
rect 26835 24392 26847 24395
rect 27154 24392 27160 24404
rect 26835 24364 27160 24392
rect 26835 24361 26847 24364
rect 26789 24355 26847 24361
rect 27154 24352 27160 24364
rect 27212 24352 27218 24404
rect 27525 24395 27583 24401
rect 27525 24361 27537 24395
rect 27571 24392 27583 24395
rect 28718 24392 28724 24404
rect 27571 24364 28724 24392
rect 27571 24361 27583 24364
rect 27525 24355 27583 24361
rect 28718 24352 28724 24364
rect 28776 24352 28782 24404
rect 30374 24352 30380 24404
rect 30432 24392 30438 24404
rect 31941 24395 31999 24401
rect 31941 24392 31953 24395
rect 30432 24364 31953 24392
rect 30432 24352 30438 24364
rect 31941 24361 31953 24364
rect 31987 24392 31999 24395
rect 32306 24392 32312 24404
rect 31987 24364 32312 24392
rect 31987 24361 31999 24364
rect 31941 24355 31999 24361
rect 32306 24352 32312 24364
rect 32364 24392 32370 24404
rect 33042 24392 33048 24404
rect 32364 24364 33048 24392
rect 32364 24352 32370 24364
rect 33042 24352 33048 24364
rect 33100 24352 33106 24404
rect 33318 24352 33324 24404
rect 33376 24392 33382 24404
rect 33413 24395 33471 24401
rect 33413 24392 33425 24395
rect 33376 24364 33425 24392
rect 33376 24352 33382 24364
rect 33413 24361 33425 24364
rect 33459 24361 33471 24395
rect 34974 24392 34980 24404
rect 34935 24364 34980 24392
rect 33413 24355 33471 24361
rect 34974 24352 34980 24364
rect 35032 24352 35038 24404
rect 35342 24392 35348 24404
rect 35303 24364 35348 24392
rect 35342 24352 35348 24364
rect 35400 24352 35406 24404
rect 20254 24284 20260 24336
rect 20312 24324 20318 24336
rect 21174 24324 21180 24336
rect 20312 24296 21180 24324
rect 20312 24284 20318 24296
rect 21174 24284 21180 24296
rect 21232 24324 21238 24336
rect 21637 24327 21695 24333
rect 21637 24324 21649 24327
rect 21232 24296 21649 24324
rect 21232 24284 21238 24296
rect 21637 24293 21649 24296
rect 21683 24324 21695 24327
rect 21910 24324 21916 24336
rect 21683 24296 21916 24324
rect 21683 24293 21695 24296
rect 21637 24287 21695 24293
rect 21910 24284 21916 24296
rect 21968 24284 21974 24336
rect 22094 24284 22100 24336
rect 22152 24324 22158 24336
rect 23106 24324 23112 24336
rect 22152 24296 23112 24324
rect 22152 24284 22158 24296
rect 23106 24284 23112 24296
rect 23164 24284 23170 24336
rect 24762 24324 24768 24336
rect 24723 24296 24768 24324
rect 24762 24284 24768 24296
rect 24820 24284 24826 24336
rect 27985 24327 28043 24333
rect 27985 24293 27997 24327
rect 28031 24324 28043 24327
rect 28258 24324 28264 24336
rect 28031 24296 28264 24324
rect 28031 24293 28043 24296
rect 27985 24287 28043 24293
rect 28258 24284 28264 24296
rect 28316 24324 28322 24336
rect 28626 24324 28632 24336
rect 28316 24296 28632 24324
rect 28316 24284 28322 24296
rect 28626 24284 28632 24296
rect 28684 24284 28690 24336
rect 30466 24324 30472 24336
rect 30427 24296 30472 24324
rect 30466 24284 30472 24296
rect 30524 24284 30530 24336
rect 21542 24256 21548 24268
rect 21503 24228 21548 24256
rect 21542 24216 21548 24228
rect 21600 24216 21606 24268
rect 27341 24259 27399 24265
rect 27341 24225 27353 24259
rect 27387 24256 27399 24259
rect 27522 24256 27528 24268
rect 27387 24228 27528 24256
rect 27387 24225 27399 24228
rect 27341 24219 27399 24225
rect 27522 24216 27528 24228
rect 27580 24216 27586 24268
rect 28442 24256 28448 24268
rect 28403 24228 28448 24256
rect 28442 24216 28448 24228
rect 28500 24216 28506 24268
rect 28644 24256 28672 24284
rect 28712 24259 28770 24265
rect 28712 24256 28724 24259
rect 28644 24228 28724 24256
rect 28712 24225 28724 24228
rect 28758 24225 28770 24259
rect 35710 24256 35716 24268
rect 35671 24228 35716 24256
rect 28712 24219 28770 24225
rect 35710 24216 35716 24228
rect 35768 24216 35774 24268
rect 21818 24188 21824 24200
rect 21779 24160 21824 24188
rect 21818 24148 21824 24160
rect 21876 24148 21882 24200
rect 22830 24148 22836 24200
rect 22888 24188 22894 24200
rect 23201 24191 23259 24197
rect 23201 24188 23213 24191
rect 22888 24160 23213 24188
rect 22888 24148 22894 24160
rect 23201 24157 23213 24160
rect 23247 24157 23259 24191
rect 23201 24151 23259 24157
rect 23385 24191 23443 24197
rect 23385 24157 23397 24191
rect 23431 24188 23443 24191
rect 24949 24191 25007 24197
rect 24949 24188 24961 24191
rect 23431 24160 24961 24188
rect 23431 24157 23443 24160
rect 23385 24151 23443 24157
rect 24949 24157 24961 24160
rect 24995 24188 25007 24191
rect 25406 24188 25412 24200
rect 24995 24160 25412 24188
rect 24995 24157 25007 24160
rect 24949 24151 25007 24157
rect 25406 24148 25412 24160
rect 25464 24148 25470 24200
rect 35802 24188 35808 24200
rect 35763 24160 35808 24188
rect 35802 24148 35808 24160
rect 35860 24148 35866 24200
rect 35989 24191 36047 24197
rect 35989 24157 36001 24191
rect 36035 24188 36047 24191
rect 36262 24188 36268 24200
rect 36035 24160 36268 24188
rect 36035 24157 36047 24160
rect 35989 24151 36047 24157
rect 36262 24148 36268 24160
rect 36320 24148 36326 24200
rect 21177 24055 21235 24061
rect 21177 24021 21189 24055
rect 21223 24052 21235 24055
rect 22830 24052 22836 24064
rect 21223 24024 22836 24052
rect 21223 24021 21235 24024
rect 21177 24015 21235 24021
rect 22830 24012 22836 24024
rect 22888 24012 22894 24064
rect 24118 24052 24124 24064
rect 24079 24024 24124 24052
rect 24118 24012 24124 24024
rect 24176 24012 24182 24064
rect 29822 24052 29828 24064
rect 29783 24024 29828 24052
rect 29822 24012 29828 24024
rect 29880 24012 29886 24064
rect 32674 24052 32680 24064
rect 32635 24024 32680 24052
rect 32674 24012 32680 24024
rect 32732 24012 32738 24064
rect 34054 24052 34060 24064
rect 34015 24024 34060 24052
rect 34054 24012 34060 24024
rect 34112 24012 34118 24064
rect 34517 24055 34575 24061
rect 34517 24021 34529 24055
rect 34563 24052 34575 24055
rect 34606 24052 34612 24064
rect 34563 24024 34612 24052
rect 34563 24021 34575 24024
rect 34517 24015 34575 24021
rect 34606 24012 34612 24024
rect 34664 24012 34670 24064
rect 1104 23962 38824 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 34966 23962
rect 35018 23910 35030 23962
rect 35082 23910 35094 23962
rect 35146 23910 35158 23962
rect 35210 23910 38824 23962
rect 1104 23888 38824 23910
rect 20254 23848 20260 23860
rect 20215 23820 20260 23848
rect 20254 23808 20260 23820
rect 20312 23808 20318 23860
rect 20714 23848 20720 23860
rect 20675 23820 20720 23848
rect 20714 23808 20720 23820
rect 20772 23808 20778 23860
rect 21542 23808 21548 23860
rect 21600 23848 21606 23860
rect 22189 23851 22247 23857
rect 22189 23848 22201 23851
rect 21600 23820 22201 23848
rect 21600 23808 21606 23820
rect 22189 23817 22201 23820
rect 22235 23817 22247 23851
rect 22830 23848 22836 23860
rect 22791 23820 22836 23848
rect 22189 23811 22247 23817
rect 22830 23808 22836 23820
rect 22888 23808 22894 23860
rect 23106 23848 23112 23860
rect 23067 23820 23112 23848
rect 23106 23808 23112 23820
rect 23164 23808 23170 23860
rect 23937 23851 23995 23857
rect 23937 23817 23949 23851
rect 23983 23848 23995 23851
rect 24762 23848 24768 23860
rect 23983 23820 24768 23848
rect 23983 23817 23995 23820
rect 23937 23811 23995 23817
rect 24762 23808 24768 23820
rect 24820 23808 24826 23860
rect 25869 23851 25927 23857
rect 25869 23817 25881 23851
rect 25915 23848 25927 23851
rect 26142 23848 26148 23860
rect 25915 23820 26148 23848
rect 25915 23817 25927 23820
rect 25869 23811 25927 23817
rect 24394 23780 24400 23792
rect 24355 23752 24400 23780
rect 24394 23740 24400 23752
rect 24452 23740 24458 23792
rect 21818 23712 21824 23724
rect 21779 23684 21824 23712
rect 21818 23672 21824 23684
rect 21876 23672 21882 23724
rect 25041 23715 25099 23721
rect 25041 23681 25053 23715
rect 25087 23712 25099 23715
rect 25884 23712 25912 23811
rect 26142 23808 26148 23820
rect 26200 23808 26206 23860
rect 26602 23848 26608 23860
rect 26563 23820 26608 23848
rect 26602 23808 26608 23820
rect 26660 23808 26666 23860
rect 27433 23851 27491 23857
rect 27433 23817 27445 23851
rect 27479 23848 27491 23851
rect 27522 23848 27528 23860
rect 27479 23820 27528 23848
rect 27479 23817 27491 23820
rect 27433 23811 27491 23817
rect 27522 23808 27528 23820
rect 27580 23808 27586 23860
rect 28442 23808 28448 23860
rect 28500 23848 28506 23860
rect 28629 23851 28687 23857
rect 28629 23848 28641 23851
rect 28500 23820 28641 23848
rect 28500 23808 28506 23820
rect 28629 23817 28641 23820
rect 28675 23817 28687 23851
rect 28629 23811 28687 23817
rect 29273 23851 29331 23857
rect 29273 23817 29285 23851
rect 29319 23848 29331 23851
rect 34885 23851 34943 23857
rect 29319 23820 33456 23848
rect 29319 23817 29331 23820
rect 29273 23811 29331 23817
rect 27617 23783 27675 23789
rect 27617 23749 27629 23783
rect 27663 23780 27675 23783
rect 30653 23783 30711 23789
rect 30653 23780 30665 23783
rect 27663 23752 30665 23780
rect 27663 23749 27675 23752
rect 27617 23743 27675 23749
rect 28258 23712 28264 23724
rect 25087 23684 25912 23712
rect 28219 23684 28264 23712
rect 25087 23681 25099 23684
rect 25041 23675 25099 23681
rect 28258 23672 28264 23684
rect 28316 23672 28322 23724
rect 29748 23721 29776 23752
rect 30653 23749 30665 23752
rect 30699 23749 30711 23783
rect 33428 23780 33456 23820
rect 34885 23817 34897 23851
rect 34931 23848 34943 23851
rect 35802 23848 35808 23860
rect 34931 23820 35808 23848
rect 34931 23817 34943 23820
rect 34885 23811 34943 23817
rect 35802 23808 35808 23820
rect 35860 23848 35866 23860
rect 36633 23851 36691 23857
rect 36633 23848 36645 23851
rect 35860 23820 36645 23848
rect 35860 23808 35866 23820
rect 36633 23817 36645 23820
rect 36679 23817 36691 23851
rect 36633 23811 36691 23817
rect 36170 23780 36176 23792
rect 33428 23752 36176 23780
rect 30653 23743 30711 23749
rect 36170 23740 36176 23752
rect 36228 23740 36234 23792
rect 29733 23715 29791 23721
rect 29733 23681 29745 23715
rect 29779 23681 29791 23715
rect 29733 23675 29791 23681
rect 29822 23672 29828 23724
rect 29880 23712 29886 23724
rect 30285 23715 30343 23721
rect 30285 23712 30297 23715
rect 29880 23684 30297 23712
rect 29880 23672 29886 23684
rect 30285 23681 30297 23684
rect 30331 23681 30343 23715
rect 30285 23675 30343 23681
rect 34333 23715 34391 23721
rect 34333 23681 34345 23715
rect 34379 23712 34391 23715
rect 35437 23715 35495 23721
rect 35437 23712 35449 23715
rect 34379 23684 35449 23712
rect 34379 23681 34391 23684
rect 34333 23675 34391 23681
rect 35437 23681 35449 23684
rect 35483 23712 35495 23715
rect 35618 23712 35624 23724
rect 35483 23684 35624 23712
rect 35483 23681 35495 23684
rect 35437 23675 35495 23681
rect 35618 23672 35624 23684
rect 35676 23672 35682 23724
rect 20714 23604 20720 23656
rect 20772 23644 20778 23656
rect 21545 23647 21603 23653
rect 21545 23644 21557 23647
rect 20772 23616 21557 23644
rect 20772 23604 20778 23616
rect 21545 23613 21557 23616
rect 21591 23644 21603 23647
rect 22094 23644 22100 23656
rect 21591 23616 22100 23644
rect 21591 23613 21603 23616
rect 21545 23607 21603 23613
rect 22094 23604 22100 23616
rect 22152 23604 22158 23656
rect 23842 23604 23848 23656
rect 23900 23644 23906 23656
rect 24765 23647 24823 23653
rect 24765 23644 24777 23647
rect 23900 23616 24777 23644
rect 23900 23604 23906 23616
rect 24765 23613 24777 23616
rect 24811 23613 24823 23647
rect 24765 23607 24823 23613
rect 25961 23647 26019 23653
rect 25961 23613 25973 23647
rect 26007 23644 26019 23647
rect 26602 23644 26608 23656
rect 26007 23616 26608 23644
rect 26007 23613 26019 23616
rect 25961 23607 26019 23613
rect 26602 23604 26608 23616
rect 26660 23604 26666 23656
rect 26970 23604 26976 23656
rect 27028 23644 27034 23656
rect 27065 23647 27123 23653
rect 27065 23644 27077 23647
rect 27028 23616 27077 23644
rect 27028 23604 27034 23616
rect 27065 23613 27077 23616
rect 27111 23644 27123 23647
rect 27614 23644 27620 23656
rect 27111 23616 27620 23644
rect 27111 23613 27123 23616
rect 27065 23607 27123 23613
rect 27614 23604 27620 23616
rect 27672 23644 27678 23656
rect 27985 23647 28043 23653
rect 27985 23644 27997 23647
rect 27672 23616 27997 23644
rect 27672 23604 27678 23616
rect 27985 23613 27997 23616
rect 28031 23613 28043 23647
rect 27985 23607 28043 23613
rect 34238 23604 34244 23656
rect 34296 23644 34302 23656
rect 35710 23644 35716 23656
rect 34296 23616 35716 23644
rect 34296 23604 34302 23616
rect 35710 23604 35716 23616
rect 35768 23644 35774 23656
rect 35897 23647 35955 23653
rect 35897 23644 35909 23647
rect 35768 23616 35909 23644
rect 35768 23604 35774 23616
rect 35897 23613 35909 23616
rect 35943 23613 35955 23647
rect 35897 23607 35955 23613
rect 21637 23579 21695 23585
rect 21637 23576 21649 23579
rect 21008 23548 21649 23576
rect 21008 23520 21036 23548
rect 21637 23545 21649 23548
rect 21683 23545 21695 23579
rect 21637 23539 21695 23545
rect 24305 23579 24363 23585
rect 24305 23545 24317 23579
rect 24351 23576 24363 23579
rect 24854 23576 24860 23588
rect 24351 23548 24860 23576
rect 24351 23545 24363 23548
rect 24305 23539 24363 23545
rect 24854 23536 24860 23548
rect 24912 23536 24918 23588
rect 29089 23579 29147 23585
rect 29089 23545 29101 23579
rect 29135 23576 29147 23579
rect 29641 23579 29699 23585
rect 29641 23576 29653 23579
rect 29135 23548 29653 23576
rect 29135 23545 29147 23548
rect 29089 23539 29147 23545
rect 29641 23545 29653 23548
rect 29687 23576 29699 23579
rect 30837 23579 30895 23585
rect 30837 23576 30849 23579
rect 29687 23548 30849 23576
rect 29687 23545 29699 23548
rect 29641 23539 29699 23545
rect 30837 23545 30849 23548
rect 30883 23545 30895 23579
rect 30837 23539 30895 23545
rect 34790 23536 34796 23588
rect 34848 23576 34854 23588
rect 35253 23579 35311 23585
rect 35253 23576 35265 23579
rect 34848 23548 35265 23576
rect 34848 23536 34854 23548
rect 35253 23545 35265 23548
rect 35299 23545 35311 23579
rect 35253 23539 35311 23545
rect 19978 23508 19984 23520
rect 19939 23480 19984 23508
rect 19978 23468 19984 23480
rect 20036 23468 20042 23520
rect 20990 23508 20996 23520
rect 20951 23480 20996 23508
rect 20990 23468 20996 23480
rect 21048 23468 21054 23520
rect 21174 23508 21180 23520
rect 21135 23480 21180 23508
rect 21174 23468 21180 23480
rect 21232 23468 21238 23520
rect 25406 23508 25412 23520
rect 25367 23480 25412 23508
rect 25406 23468 25412 23480
rect 25464 23468 25470 23520
rect 28077 23511 28135 23517
rect 28077 23477 28089 23511
rect 28123 23508 28135 23511
rect 28166 23508 28172 23520
rect 28123 23480 28172 23508
rect 28123 23477 28135 23480
rect 28077 23471 28135 23477
rect 28166 23468 28172 23480
rect 28224 23468 28230 23520
rect 34606 23468 34612 23520
rect 34664 23508 34670 23520
rect 34701 23511 34759 23517
rect 34701 23508 34713 23511
rect 34664 23480 34713 23508
rect 34664 23468 34670 23480
rect 34701 23477 34713 23480
rect 34747 23508 34759 23511
rect 35345 23511 35403 23517
rect 35345 23508 35357 23511
rect 34747 23480 35357 23508
rect 34747 23477 34759 23480
rect 34701 23471 34759 23477
rect 35345 23477 35357 23480
rect 35391 23508 35403 23511
rect 35526 23508 35532 23520
rect 35391 23480 35532 23508
rect 35391 23477 35403 23480
rect 35345 23471 35403 23477
rect 35526 23468 35532 23480
rect 35584 23468 35590 23520
rect 36262 23508 36268 23520
rect 36223 23480 36268 23508
rect 36262 23468 36268 23480
rect 36320 23468 36326 23520
rect 1104 23418 38824 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 38824 23418
rect 1104 23344 38824 23366
rect 19978 23264 19984 23316
rect 20036 23304 20042 23316
rect 20717 23307 20775 23313
rect 20717 23304 20729 23307
rect 20036 23276 20729 23304
rect 20036 23264 20042 23276
rect 20717 23273 20729 23276
rect 20763 23304 20775 23307
rect 21818 23304 21824 23316
rect 20763 23276 21824 23304
rect 20763 23273 20775 23276
rect 20717 23267 20775 23273
rect 21818 23264 21824 23276
rect 21876 23264 21882 23316
rect 22094 23264 22100 23316
rect 22152 23304 22158 23316
rect 22281 23307 22339 23313
rect 22281 23304 22293 23307
rect 22152 23276 22293 23304
rect 22152 23264 22158 23276
rect 22281 23273 22293 23276
rect 22327 23273 22339 23307
rect 23382 23304 23388 23316
rect 23343 23276 23388 23304
rect 22281 23267 22339 23273
rect 23382 23264 23388 23276
rect 23440 23264 23446 23316
rect 23750 23304 23756 23316
rect 23711 23276 23756 23304
rect 23750 23264 23756 23276
rect 23808 23264 23814 23316
rect 23842 23264 23848 23316
rect 23900 23304 23906 23316
rect 24397 23307 24455 23313
rect 24397 23304 24409 23307
rect 23900 23276 24409 23304
rect 23900 23264 23906 23276
rect 24397 23273 24409 23276
rect 24443 23273 24455 23307
rect 24397 23267 24455 23273
rect 24854 23264 24860 23316
rect 24912 23304 24918 23316
rect 25133 23307 25191 23313
rect 25133 23304 25145 23307
rect 24912 23276 25145 23304
rect 24912 23264 24918 23276
rect 25133 23273 25145 23276
rect 25179 23273 25191 23307
rect 26970 23304 26976 23316
rect 26931 23276 26976 23304
rect 25133 23267 25191 23273
rect 26970 23264 26976 23276
rect 27028 23264 27034 23316
rect 28258 23264 28264 23316
rect 28316 23304 28322 23316
rect 28445 23307 28503 23313
rect 28445 23304 28457 23307
rect 28316 23276 28457 23304
rect 28316 23264 28322 23276
rect 28445 23273 28457 23276
rect 28491 23273 28503 23307
rect 28445 23267 28503 23273
rect 34149 23307 34207 23313
rect 34149 23273 34161 23307
rect 34195 23304 34207 23307
rect 34238 23304 34244 23316
rect 34195 23276 34244 23304
rect 34195 23273 34207 23276
rect 34149 23267 34207 23273
rect 34238 23264 34244 23276
rect 34296 23264 34302 23316
rect 35618 23264 35624 23316
rect 35676 23304 35682 23316
rect 36541 23307 36599 23313
rect 36541 23304 36553 23307
rect 35676 23276 36553 23304
rect 35676 23264 35682 23276
rect 36541 23273 36553 23276
rect 36587 23304 36599 23307
rect 36722 23304 36728 23316
rect 36587 23276 36728 23304
rect 36587 23273 36599 23276
rect 36541 23267 36599 23273
rect 36722 23264 36728 23276
rect 36780 23264 36786 23316
rect 28902 23236 28908 23248
rect 27908 23208 28908 23236
rect 27908 23180 27936 23208
rect 28902 23196 28908 23208
rect 28960 23196 28966 23248
rect 20622 23128 20628 23180
rect 20680 23168 20686 23180
rect 20990 23168 20996 23180
rect 20680 23140 20996 23168
rect 20680 23128 20686 23140
rect 20990 23128 20996 23140
rect 21048 23168 21054 23180
rect 21157 23171 21215 23177
rect 21157 23168 21169 23171
rect 21048 23140 21169 23168
rect 21048 23128 21054 23140
rect 21157 23137 21169 23140
rect 21203 23137 21215 23171
rect 21157 23131 21215 23137
rect 22925 23171 22983 23177
rect 22925 23137 22937 23171
rect 22971 23168 22983 23171
rect 23293 23171 23351 23177
rect 23293 23168 23305 23171
rect 22971 23140 23305 23168
rect 22971 23137 22983 23140
rect 22925 23131 22983 23137
rect 23293 23137 23305 23140
rect 23339 23168 23351 23171
rect 24946 23168 24952 23180
rect 23339 23140 24072 23168
rect 24907 23140 24952 23168
rect 23339 23137 23351 23140
rect 23293 23131 23351 23137
rect 24044 23112 24072 23140
rect 24946 23128 24952 23140
rect 25004 23128 25010 23180
rect 27890 23168 27896 23180
rect 27803 23140 27896 23168
rect 27890 23128 27896 23140
rect 27948 23128 27954 23180
rect 28350 23128 28356 23180
rect 28408 23168 28414 23180
rect 29253 23171 29311 23177
rect 29253 23168 29265 23171
rect 28408 23140 29265 23168
rect 28408 23128 28414 23140
rect 29253 23137 29265 23140
rect 29299 23168 29311 23171
rect 29822 23168 29828 23180
rect 29299 23140 29828 23168
rect 29299 23137 29311 23140
rect 29253 23131 29311 23137
rect 29822 23128 29828 23140
rect 29880 23128 29886 23180
rect 35428 23171 35486 23177
rect 35428 23137 35440 23171
rect 35474 23168 35486 23171
rect 35802 23168 35808 23180
rect 35474 23140 35808 23168
rect 35474 23137 35486 23140
rect 35428 23131 35486 23137
rect 35802 23128 35808 23140
rect 35860 23128 35866 23180
rect 20898 23100 20904 23112
rect 20859 23072 20904 23100
rect 20898 23060 20904 23072
rect 20956 23060 20962 23112
rect 23842 23100 23848 23112
rect 23803 23072 23848 23100
rect 23842 23060 23848 23072
rect 23900 23060 23906 23112
rect 24026 23100 24032 23112
rect 23987 23072 24032 23100
rect 24026 23060 24032 23072
rect 24084 23060 24090 23112
rect 24857 23103 24915 23109
rect 24857 23069 24869 23103
rect 24903 23100 24915 23103
rect 25038 23100 25044 23112
rect 24903 23072 25044 23100
rect 24903 23069 24915 23072
rect 24857 23063 24915 23069
rect 25038 23060 25044 23072
rect 25096 23060 25102 23112
rect 28442 23060 28448 23112
rect 28500 23100 28506 23112
rect 28997 23103 29055 23109
rect 28997 23100 29009 23103
rect 28500 23072 29009 23100
rect 28500 23060 28506 23072
rect 28997 23069 29009 23072
rect 29043 23069 29055 23103
rect 28997 23063 29055 23069
rect 35161 23103 35219 23109
rect 35161 23069 35173 23103
rect 35207 23069 35219 23103
rect 35161 23063 35219 23069
rect 27709 23035 27767 23041
rect 27709 23001 27721 23035
rect 27755 23032 27767 23035
rect 28166 23032 28172 23044
rect 27755 23004 28172 23032
rect 27755 23001 27767 23004
rect 27709 22995 27767 23001
rect 28166 22992 28172 23004
rect 28224 22992 28230 23044
rect 28074 22964 28080 22976
rect 28035 22936 28080 22964
rect 28074 22924 28080 22936
rect 28132 22924 28138 22976
rect 28905 22967 28963 22973
rect 28905 22933 28917 22967
rect 28951 22964 28963 22967
rect 29362 22964 29368 22976
rect 28951 22936 29368 22964
rect 28951 22933 28963 22936
rect 28905 22927 28963 22933
rect 29362 22924 29368 22936
rect 29420 22964 29426 22976
rect 30377 22967 30435 22973
rect 30377 22964 30389 22967
rect 29420 22936 30389 22964
rect 29420 22924 29426 22936
rect 30377 22933 30389 22936
rect 30423 22964 30435 22967
rect 30650 22964 30656 22976
rect 30423 22936 30656 22964
rect 30423 22933 30435 22936
rect 30377 22927 30435 22933
rect 30650 22924 30656 22936
rect 30708 22924 30714 22976
rect 34790 22924 34796 22976
rect 34848 22964 34854 22976
rect 34885 22967 34943 22973
rect 34885 22964 34897 22967
rect 34848 22936 34897 22964
rect 34848 22924 34854 22936
rect 34885 22933 34897 22936
rect 34931 22933 34943 22967
rect 35176 22964 35204 23063
rect 35342 22964 35348 22976
rect 35176 22936 35348 22964
rect 34885 22927 34943 22933
rect 35342 22924 35348 22936
rect 35400 22924 35406 22976
rect 1104 22874 38824 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 34966 22874
rect 35018 22822 35030 22874
rect 35082 22822 35094 22874
rect 35146 22822 35158 22874
rect 35210 22822 38824 22874
rect 1104 22800 38824 22822
rect 20898 22760 20904 22772
rect 20859 22732 20904 22760
rect 20898 22720 20904 22732
rect 20956 22720 20962 22772
rect 21542 22760 21548 22772
rect 21503 22732 21548 22760
rect 21542 22720 21548 22732
rect 21600 22720 21606 22772
rect 23842 22720 23848 22772
rect 23900 22760 23906 22772
rect 24673 22763 24731 22769
rect 24673 22760 24685 22763
rect 23900 22732 24685 22760
rect 23900 22720 23906 22732
rect 24673 22729 24685 22732
rect 24719 22729 24731 22763
rect 25406 22760 25412 22772
rect 24673 22723 24731 22729
rect 25056 22732 25412 22760
rect 23661 22695 23719 22701
rect 23661 22661 23673 22695
rect 23707 22692 23719 22695
rect 24946 22692 24952 22704
rect 23707 22664 24952 22692
rect 23707 22661 23719 22664
rect 23661 22655 23719 22661
rect 24946 22652 24952 22664
rect 25004 22652 25010 22704
rect 20257 22627 20315 22633
rect 20257 22593 20269 22627
rect 20303 22624 20315 22627
rect 21818 22624 21824 22636
rect 20303 22596 21824 22624
rect 20303 22593 20315 22596
rect 20257 22587 20315 22593
rect 21818 22584 21824 22596
rect 21876 22624 21882 22636
rect 22097 22627 22155 22633
rect 22097 22624 22109 22627
rect 21876 22596 22109 22624
rect 21876 22584 21882 22596
rect 22097 22593 22109 22596
rect 22143 22593 22155 22627
rect 22097 22587 22155 22593
rect 24026 22584 24032 22636
rect 24084 22624 24090 22636
rect 24305 22627 24363 22633
rect 24305 22624 24317 22627
rect 24084 22596 24317 22624
rect 24084 22584 24090 22596
rect 24305 22593 24317 22596
rect 24351 22624 24363 22627
rect 25056 22624 25084 22732
rect 25406 22720 25412 22732
rect 25464 22720 25470 22772
rect 27890 22760 27896 22772
rect 27851 22732 27896 22760
rect 27890 22720 27896 22732
rect 27948 22720 27954 22772
rect 28350 22760 28356 22772
rect 28311 22732 28356 22760
rect 28350 22720 28356 22732
rect 28408 22720 28414 22772
rect 28442 22720 28448 22772
rect 28500 22760 28506 22772
rect 28626 22760 28632 22772
rect 28500 22732 28632 22760
rect 28500 22720 28506 22732
rect 28626 22720 28632 22732
rect 28684 22760 28690 22772
rect 28997 22763 29055 22769
rect 28997 22760 29009 22763
rect 28684 22732 29009 22760
rect 28684 22720 28690 22732
rect 28997 22729 29009 22732
rect 29043 22729 29055 22763
rect 28997 22723 29055 22729
rect 25866 22624 25872 22636
rect 24351 22596 25084 22624
rect 25240 22596 25872 22624
rect 24351 22593 24363 22596
rect 24305 22587 24363 22593
rect 22005 22559 22063 22565
rect 22005 22556 22017 22559
rect 21376 22528 22017 22556
rect 21376 22432 21404 22528
rect 22005 22525 22017 22528
rect 22051 22525 22063 22559
rect 22005 22519 22063 22525
rect 23477 22559 23535 22565
rect 23477 22525 23489 22559
rect 23523 22556 23535 22559
rect 23658 22556 23664 22568
rect 23523 22528 23664 22556
rect 23523 22525 23535 22528
rect 23477 22519 23535 22525
rect 23658 22516 23664 22528
rect 23716 22556 23722 22568
rect 25240 22565 25268 22596
rect 25866 22584 25872 22596
rect 25924 22584 25930 22636
rect 26234 22584 26240 22636
rect 26292 22624 26298 22636
rect 26421 22627 26479 22633
rect 26421 22624 26433 22627
rect 26292 22596 26433 22624
rect 26292 22584 26298 22596
rect 26421 22593 26433 22596
rect 26467 22624 26479 22627
rect 27433 22627 27491 22633
rect 27433 22624 27445 22627
rect 26467 22596 27445 22624
rect 26467 22593 26479 22596
rect 26421 22587 26479 22593
rect 27433 22593 27445 22596
rect 27479 22624 27491 22627
rect 27522 22624 27528 22636
rect 27479 22596 27528 22624
rect 27479 22593 27491 22596
rect 27433 22587 27491 22593
rect 27522 22584 27528 22596
rect 27580 22584 27586 22636
rect 29012 22624 29040 22723
rect 32950 22720 32956 22772
rect 33008 22760 33014 22772
rect 36262 22760 36268 22772
rect 33008 22732 36268 22760
rect 33008 22720 33014 22732
rect 36262 22720 36268 22732
rect 36320 22760 36326 22772
rect 36725 22763 36783 22769
rect 36725 22760 36737 22763
rect 36320 22732 36737 22760
rect 36320 22720 36326 22732
rect 36725 22729 36737 22732
rect 36771 22729 36783 22763
rect 36725 22723 36783 22729
rect 29273 22627 29331 22633
rect 29273 22624 29285 22627
rect 29012 22596 29285 22624
rect 29273 22593 29285 22596
rect 29319 22593 29331 22627
rect 29273 22587 29331 22593
rect 24121 22559 24179 22565
rect 24121 22556 24133 22559
rect 23716 22528 24133 22556
rect 23716 22516 23722 22528
rect 24121 22525 24133 22528
rect 24167 22525 24179 22559
rect 24121 22519 24179 22525
rect 25225 22559 25283 22565
rect 25225 22525 25237 22559
rect 25271 22525 25283 22559
rect 25225 22519 25283 22525
rect 26970 22516 26976 22568
rect 27028 22556 27034 22568
rect 27341 22559 27399 22565
rect 27341 22556 27353 22559
rect 27028 22528 27353 22556
rect 27028 22516 27034 22528
rect 27341 22525 27353 22528
rect 27387 22525 27399 22559
rect 27341 22519 27399 22525
rect 29362 22516 29368 22568
rect 29420 22556 29426 22568
rect 29529 22559 29587 22565
rect 29529 22556 29541 22559
rect 29420 22528 29541 22556
rect 29420 22516 29426 22528
rect 29529 22525 29541 22528
rect 29575 22525 29587 22559
rect 29529 22519 29587 22525
rect 32122 22516 32128 22568
rect 32180 22556 32186 22568
rect 32217 22559 32275 22565
rect 32217 22556 32229 22559
rect 32180 22528 32229 22556
rect 32180 22516 32186 22528
rect 32217 22525 32229 22528
rect 32263 22525 32275 22559
rect 32217 22519 32275 22525
rect 35158 22516 35164 22568
rect 35216 22556 35222 22568
rect 35342 22556 35348 22568
rect 35216 22528 35348 22556
rect 35216 22516 35222 22528
rect 35342 22516 35348 22528
rect 35400 22516 35406 22568
rect 35618 22565 35624 22568
rect 35612 22556 35624 22565
rect 35579 22528 35624 22556
rect 35612 22519 35624 22528
rect 35618 22516 35624 22519
rect 35676 22516 35682 22568
rect 22557 22491 22615 22497
rect 22557 22488 22569 22491
rect 21928 22460 22569 22488
rect 21928 22432 21956 22460
rect 22557 22457 22569 22460
rect 22603 22457 22615 22491
rect 24029 22491 24087 22497
rect 24029 22488 24041 22491
rect 22557 22451 22615 22457
rect 23124 22460 24041 22488
rect 23124 22432 23152 22460
rect 24029 22457 24041 22460
rect 24075 22457 24087 22491
rect 24029 22451 24087 22457
rect 26789 22491 26847 22497
rect 26789 22457 26801 22491
rect 26835 22488 26847 22491
rect 27154 22488 27160 22500
rect 26835 22460 27160 22488
rect 26835 22457 26847 22460
rect 26789 22451 26847 22457
rect 27154 22448 27160 22460
rect 27212 22488 27218 22500
rect 27249 22491 27307 22497
rect 27249 22488 27261 22491
rect 27212 22460 27261 22488
rect 27212 22448 27218 22460
rect 27249 22457 27261 22460
rect 27295 22457 27307 22491
rect 27249 22451 27307 22457
rect 31757 22491 31815 22497
rect 31757 22457 31769 22491
rect 31803 22488 31815 22491
rect 32462 22491 32520 22497
rect 32462 22488 32474 22491
rect 31803 22460 32474 22488
rect 31803 22457 31815 22460
rect 31757 22451 31815 22457
rect 32462 22457 32474 22460
rect 32508 22488 32520 22491
rect 32950 22488 32956 22500
rect 32508 22460 32956 22488
rect 32508 22457 32520 22460
rect 32462 22451 32520 22457
rect 32950 22448 32956 22460
rect 33008 22448 33014 22500
rect 34333 22491 34391 22497
rect 34333 22457 34345 22491
rect 34379 22488 34391 22491
rect 34379 22460 35296 22488
rect 34379 22457 34391 22460
rect 34333 22451 34391 22457
rect 20622 22420 20628 22432
rect 20583 22392 20628 22420
rect 20622 22380 20628 22392
rect 20680 22380 20686 22432
rect 21358 22420 21364 22432
rect 21319 22392 21364 22420
rect 21358 22380 21364 22392
rect 21416 22380 21422 22432
rect 21910 22420 21916 22432
rect 21871 22392 21916 22420
rect 21910 22380 21916 22392
rect 21968 22380 21974 22432
rect 23106 22420 23112 22432
rect 23067 22392 23112 22420
rect 23106 22380 23112 22392
rect 23164 22380 23170 22432
rect 23750 22380 23756 22432
rect 23808 22420 23814 22432
rect 25041 22423 25099 22429
rect 25041 22420 25053 22423
rect 23808 22392 25053 22420
rect 23808 22380 23814 22392
rect 25041 22389 25053 22392
rect 25087 22389 25099 22423
rect 26878 22420 26884 22432
rect 26839 22392 26884 22420
rect 25041 22383 25099 22389
rect 26878 22380 26884 22392
rect 26936 22380 26942 22432
rect 30466 22380 30472 22432
rect 30524 22420 30530 22432
rect 30653 22423 30711 22429
rect 30653 22420 30665 22423
rect 30524 22392 30665 22420
rect 30524 22380 30530 22392
rect 30653 22389 30665 22392
rect 30699 22389 30711 22423
rect 32122 22420 32128 22432
rect 32083 22392 32128 22420
rect 30653 22383 30711 22389
rect 32122 22380 32128 22392
rect 32180 22380 32186 22432
rect 33594 22420 33600 22432
rect 33555 22392 33600 22420
rect 33594 22380 33600 22392
rect 33652 22380 33658 22432
rect 34238 22380 34244 22432
rect 34296 22420 34302 22432
rect 34609 22423 34667 22429
rect 34609 22420 34621 22423
rect 34296 22392 34621 22420
rect 34296 22380 34302 22392
rect 34609 22389 34621 22392
rect 34655 22420 34667 22423
rect 35158 22420 35164 22432
rect 34655 22392 35164 22420
rect 34655 22389 34667 22392
rect 34609 22383 34667 22389
rect 35158 22380 35164 22392
rect 35216 22380 35222 22432
rect 35268 22420 35296 22460
rect 35802 22420 35808 22432
rect 35268 22392 35808 22420
rect 35802 22380 35808 22392
rect 35860 22380 35866 22432
rect 1104 22330 38824 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 38824 22330
rect 1104 22256 38824 22278
rect 20622 22176 20628 22228
rect 20680 22216 20686 22228
rect 22281 22219 22339 22225
rect 22281 22216 22293 22219
rect 20680 22188 22293 22216
rect 20680 22176 20686 22188
rect 22281 22185 22293 22188
rect 22327 22185 22339 22219
rect 22281 22179 22339 22185
rect 23106 22176 23112 22228
rect 23164 22216 23170 22228
rect 23385 22219 23443 22225
rect 23385 22216 23397 22219
rect 23164 22188 23397 22216
rect 23164 22176 23170 22188
rect 23385 22185 23397 22188
rect 23431 22185 23443 22219
rect 24026 22216 24032 22228
rect 23385 22179 23443 22185
rect 23584 22188 24032 22216
rect 21818 22108 21824 22160
rect 21876 22148 21882 22160
rect 23293 22151 23351 22157
rect 21876 22120 22048 22148
rect 21876 22108 21882 22120
rect 20714 22040 20720 22092
rect 20772 22080 20778 22092
rect 21157 22083 21215 22089
rect 21157 22080 21169 22083
rect 20772 22052 21169 22080
rect 20772 22040 20778 22052
rect 21157 22049 21169 22052
rect 21203 22080 21215 22083
rect 21910 22080 21916 22092
rect 21203 22052 21916 22080
rect 21203 22049 21215 22052
rect 21157 22043 21215 22049
rect 21910 22040 21916 22052
rect 21968 22040 21974 22092
rect 22020 22080 22048 22120
rect 23293 22117 23305 22151
rect 23339 22148 23351 22151
rect 23584 22148 23612 22188
rect 24026 22176 24032 22188
rect 24084 22176 24090 22228
rect 24946 22216 24952 22228
rect 24907 22188 24952 22216
rect 24946 22176 24952 22188
rect 25004 22176 25010 22228
rect 27251 22219 27309 22225
rect 27251 22185 27263 22219
rect 27297 22216 27309 22219
rect 27430 22216 27436 22228
rect 27297 22188 27436 22216
rect 27297 22185 27309 22188
rect 27251 22179 27309 22185
rect 27430 22176 27436 22188
rect 27488 22176 27494 22228
rect 34330 22176 34336 22228
rect 34388 22216 34394 22228
rect 34698 22216 34704 22228
rect 34388 22188 34704 22216
rect 34388 22176 34394 22188
rect 34698 22176 34704 22188
rect 34756 22216 34762 22228
rect 34795 22219 34853 22225
rect 34795 22216 34807 22219
rect 34756 22188 34807 22216
rect 34756 22176 34762 22188
rect 34795 22185 34807 22188
rect 34841 22185 34853 22219
rect 34795 22179 34853 22185
rect 35526 22176 35532 22228
rect 35584 22216 35590 22228
rect 35710 22216 35716 22228
rect 35584 22188 35716 22216
rect 35584 22176 35590 22188
rect 35710 22176 35716 22188
rect 35768 22176 35774 22228
rect 36722 22216 36728 22228
rect 36683 22188 36728 22216
rect 36722 22176 36728 22188
rect 36780 22176 36786 22228
rect 23750 22148 23756 22160
rect 23339 22120 23612 22148
rect 23663 22120 23756 22148
rect 23339 22117 23351 22120
rect 23293 22111 23351 22117
rect 23750 22108 23756 22120
rect 23808 22148 23814 22160
rect 24762 22148 24768 22160
rect 23808 22120 24768 22148
rect 23808 22108 23814 22120
rect 24762 22108 24768 22120
rect 24820 22108 24826 22160
rect 23198 22080 23204 22092
rect 22020 22052 23204 22080
rect 23198 22040 23204 22052
rect 23256 22080 23262 22092
rect 25314 22080 25320 22092
rect 23256 22052 23980 22080
rect 25275 22052 25320 22080
rect 23256 22040 23262 22052
rect 20898 22012 20904 22024
rect 20859 21984 20904 22012
rect 20898 21972 20904 21984
rect 20956 21972 20962 22024
rect 23952 22021 23980 22052
rect 25314 22040 25320 22052
rect 25372 22080 25378 22092
rect 25774 22080 25780 22092
rect 25372 22052 25780 22080
rect 25372 22040 25378 22052
rect 25774 22040 25780 22052
rect 25832 22040 25838 22092
rect 27154 22040 27160 22092
rect 27212 22080 27218 22092
rect 27212 22052 27568 22080
rect 27212 22040 27218 22052
rect 23845 22015 23903 22021
rect 23845 21981 23857 22015
rect 23891 21981 23903 22015
rect 23845 21975 23903 21981
rect 23937 22015 23995 22021
rect 23937 21981 23949 22015
rect 23983 22012 23995 22015
rect 24210 22012 24216 22024
rect 23983 21984 24216 22012
rect 23983 21981 23995 21984
rect 23937 21975 23995 21981
rect 23860 21876 23888 21975
rect 24210 21972 24216 21984
rect 24268 22012 24274 22024
rect 24397 22015 24455 22021
rect 24397 22012 24409 22015
rect 24268 21984 24409 22012
rect 24268 21972 24274 21984
rect 24397 21981 24409 21984
rect 24443 21981 24455 22015
rect 26786 22012 26792 22024
rect 26747 21984 26792 22012
rect 24397 21975 24455 21981
rect 24412 21944 24440 21975
rect 26786 21972 26792 21984
rect 26844 21972 26850 22024
rect 27246 22012 27252 22024
rect 27207 21984 27252 22012
rect 27246 21972 27252 21984
rect 27304 21972 27310 22024
rect 27540 22021 27568 22052
rect 29546 22040 29552 22092
rect 29604 22080 29610 22092
rect 30101 22083 30159 22089
rect 30101 22080 30113 22083
rect 29604 22052 30113 22080
rect 29604 22040 29610 22052
rect 30101 22049 30113 22052
rect 30147 22049 30159 22083
rect 30101 22043 30159 22049
rect 31754 22040 31760 22092
rect 31812 22080 31818 22092
rect 32493 22083 32551 22089
rect 32493 22080 32505 22083
rect 31812 22052 32505 22080
rect 31812 22040 31818 22052
rect 32493 22049 32505 22052
rect 32539 22049 32551 22083
rect 32493 22043 32551 22049
rect 33873 22083 33931 22089
rect 33873 22049 33885 22083
rect 33919 22080 33931 22083
rect 34422 22080 34428 22092
rect 33919 22052 34428 22080
rect 33919 22049 33931 22052
rect 33873 22043 33931 22049
rect 34422 22040 34428 22052
rect 34480 22080 34486 22092
rect 35069 22083 35127 22089
rect 35069 22080 35081 22083
rect 34480 22052 35081 22080
rect 34480 22040 34486 22052
rect 35069 22049 35081 22052
rect 35115 22049 35127 22083
rect 35069 22043 35127 22049
rect 35802 22040 35808 22092
rect 35860 22080 35866 22092
rect 36262 22080 36268 22092
rect 35860 22052 36268 22080
rect 35860 22040 35866 22052
rect 36262 22040 36268 22052
rect 36320 22040 36326 22092
rect 27525 22015 27583 22021
rect 27525 21981 27537 22015
rect 27571 22012 27583 22015
rect 27706 22012 27712 22024
rect 27571 21984 27712 22012
rect 27571 21981 27583 21984
rect 27525 21975 27583 21981
rect 27706 21972 27712 21984
rect 27764 21972 27770 22024
rect 28166 21972 28172 22024
rect 28224 22012 28230 22024
rect 28629 22015 28687 22021
rect 28629 22012 28641 22015
rect 28224 21984 28641 22012
rect 28224 21972 28230 21984
rect 28629 21981 28641 21984
rect 28675 22012 28687 22015
rect 29181 22015 29239 22021
rect 29181 22012 29193 22015
rect 28675 21984 29193 22012
rect 28675 21981 28687 21984
rect 28629 21975 28687 21981
rect 29181 21981 29193 21984
rect 29227 22012 29239 22015
rect 30006 22012 30012 22024
rect 29227 21984 30012 22012
rect 29227 21981 29239 21984
rect 29181 21975 29239 21981
rect 30006 21972 30012 21984
rect 30064 21972 30070 22024
rect 30193 22015 30251 22021
rect 30193 21981 30205 22015
rect 30239 22012 30251 22015
rect 30282 22012 30288 22024
rect 30239 21984 30288 22012
rect 30239 21981 30251 21984
rect 30193 21975 30251 21981
rect 30282 21972 30288 21984
rect 30340 21972 30346 22024
rect 30377 22015 30435 22021
rect 30377 21981 30389 22015
rect 30423 22012 30435 22015
rect 30650 22012 30656 22024
rect 30423 21984 30656 22012
rect 30423 21981 30435 21984
rect 30377 21975 30435 21981
rect 30650 21972 30656 21984
rect 30708 21972 30714 22024
rect 31941 22015 31999 22021
rect 31941 21981 31953 22015
rect 31987 22012 31999 22015
rect 32582 22012 32588 22024
rect 31987 21984 32588 22012
rect 31987 21981 31999 21984
rect 31941 21975 31999 21981
rect 32582 21972 32588 21984
rect 32640 21972 32646 22024
rect 32677 22015 32735 22021
rect 32677 21981 32689 22015
rect 32723 21981 32735 22015
rect 34333 22015 34391 22021
rect 34333 22012 34345 22015
rect 32677 21975 32735 21981
rect 34072 21984 34345 22012
rect 25501 21947 25559 21953
rect 25501 21944 25513 21947
rect 24412 21916 25513 21944
rect 25501 21913 25513 21916
rect 25547 21913 25559 21947
rect 25501 21907 25559 21913
rect 29270 21904 29276 21956
rect 29328 21944 29334 21956
rect 30745 21947 30803 21953
rect 30745 21944 30757 21947
rect 29328 21916 30757 21944
rect 29328 21904 29334 21916
rect 30745 21913 30757 21916
rect 30791 21944 30803 21947
rect 30926 21944 30932 21956
rect 30791 21916 30932 21944
rect 30791 21913 30803 21916
rect 30745 21907 30803 21913
rect 30926 21904 30932 21916
rect 30984 21904 30990 21956
rect 32306 21904 32312 21956
rect 32364 21944 32370 21956
rect 32692 21944 32720 21975
rect 34072 21956 34100 21984
rect 34333 21981 34345 21984
rect 34379 21981 34391 22015
rect 34790 22012 34796 22024
rect 34751 21984 34796 22012
rect 34333 21975 34391 21981
rect 34790 21972 34796 21984
rect 34848 21972 34854 22024
rect 35894 21972 35900 22024
rect 35952 22012 35958 22024
rect 36173 22015 36231 22021
rect 36173 22012 36185 22015
rect 35952 21984 36185 22012
rect 35952 21972 35958 21984
rect 36173 21981 36185 21984
rect 36219 21981 36231 22015
rect 36173 21975 36231 21981
rect 34054 21944 34060 21956
rect 32364 21916 32720 21944
rect 33428 21916 34060 21944
rect 32364 21904 32370 21916
rect 24670 21876 24676 21888
rect 23860 21848 24676 21876
rect 24670 21836 24676 21848
rect 24728 21836 24734 21888
rect 26329 21879 26387 21885
rect 26329 21845 26341 21879
rect 26375 21876 26387 21879
rect 26510 21876 26516 21888
rect 26375 21848 26516 21876
rect 26375 21845 26387 21848
rect 26329 21839 26387 21845
rect 26510 21836 26516 21848
rect 26568 21836 26574 21888
rect 29546 21876 29552 21888
rect 29507 21848 29552 21876
rect 29546 21836 29552 21848
rect 29604 21836 29610 21888
rect 29730 21876 29736 21888
rect 29691 21848 29736 21876
rect 29730 21836 29736 21848
rect 29788 21836 29794 21888
rect 32125 21879 32183 21885
rect 32125 21845 32137 21879
rect 32171 21876 32183 21879
rect 32950 21876 32956 21888
rect 32171 21848 32956 21876
rect 32171 21845 32183 21848
rect 32125 21839 32183 21845
rect 32950 21836 32956 21848
rect 33008 21836 33014 21888
rect 33134 21836 33140 21888
rect 33192 21876 33198 21888
rect 33428 21885 33456 21916
rect 34054 21904 34060 21916
rect 34112 21904 34118 21956
rect 33413 21879 33471 21885
rect 33413 21876 33425 21879
rect 33192 21848 33425 21876
rect 33192 21836 33198 21848
rect 33413 21845 33425 21848
rect 33459 21845 33471 21879
rect 33413 21839 33471 21845
rect 33870 21836 33876 21888
rect 33928 21876 33934 21888
rect 34149 21879 34207 21885
rect 34149 21876 34161 21879
rect 33928 21848 34161 21876
rect 33928 21836 33934 21848
rect 34149 21845 34161 21848
rect 34195 21876 34207 21879
rect 34790 21876 34796 21888
rect 34195 21848 34796 21876
rect 34195 21845 34207 21848
rect 34149 21839 34207 21845
rect 34790 21836 34796 21848
rect 34848 21836 34854 21888
rect 1104 21786 38824 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 34966 21786
rect 35018 21734 35030 21786
rect 35082 21734 35094 21786
rect 35146 21734 35158 21786
rect 35210 21734 38824 21786
rect 1104 21712 38824 21734
rect 20898 21672 20904 21684
rect 20859 21644 20904 21672
rect 20898 21632 20904 21644
rect 20956 21632 20962 21684
rect 21910 21632 21916 21684
rect 21968 21672 21974 21684
rect 22373 21675 22431 21681
rect 22373 21672 22385 21675
rect 21968 21644 22385 21672
rect 21968 21632 21974 21644
rect 22373 21641 22385 21644
rect 22419 21641 22431 21675
rect 23658 21672 23664 21684
rect 23619 21644 23664 21672
rect 22373 21635 22431 21641
rect 23658 21632 23664 21644
rect 23716 21632 23722 21684
rect 24762 21632 24768 21684
rect 24820 21672 24826 21684
rect 25041 21675 25099 21681
rect 25041 21672 25053 21675
rect 24820 21644 25053 21672
rect 24820 21632 24826 21644
rect 25041 21641 25053 21644
rect 25087 21641 25099 21675
rect 25041 21635 25099 21641
rect 25314 21632 25320 21684
rect 25372 21672 25378 21684
rect 25685 21675 25743 21681
rect 25685 21672 25697 21675
rect 25372 21644 25697 21672
rect 25372 21632 25378 21644
rect 25685 21641 25697 21644
rect 25731 21641 25743 21675
rect 27614 21672 27620 21684
rect 27575 21644 27620 21672
rect 25685 21635 25743 21641
rect 27614 21632 27620 21644
rect 27672 21632 27678 21684
rect 28074 21632 28080 21684
rect 28132 21672 28138 21684
rect 28629 21675 28687 21681
rect 28629 21672 28641 21675
rect 28132 21644 28641 21672
rect 28132 21632 28138 21644
rect 28629 21641 28641 21644
rect 28675 21672 28687 21675
rect 29546 21672 29552 21684
rect 28675 21644 29552 21672
rect 28675 21641 28687 21644
rect 28629 21635 28687 21641
rect 29546 21632 29552 21644
rect 29604 21632 29610 21684
rect 31754 21632 31760 21684
rect 31812 21672 31818 21684
rect 34330 21672 34336 21684
rect 31812 21644 31857 21672
rect 34291 21644 34336 21672
rect 31812 21632 31818 21644
rect 34330 21632 34336 21644
rect 34388 21632 34394 21684
rect 36262 21672 36268 21684
rect 36223 21644 36268 21672
rect 36262 21632 36268 21644
rect 36320 21632 36326 21684
rect 20533 21539 20591 21545
rect 20533 21505 20545 21539
rect 20579 21536 20591 21539
rect 20916 21536 20944 21632
rect 20993 21539 21051 21545
rect 20993 21536 21005 21539
rect 20579 21508 21005 21536
rect 20579 21505 20591 21508
rect 20533 21499 20591 21505
rect 20993 21505 21005 21508
rect 21039 21505 21051 21539
rect 24210 21536 24216 21548
rect 24171 21508 24216 21536
rect 20993 21499 21051 21505
rect 24210 21496 24216 21508
rect 24268 21496 24274 21548
rect 29270 21536 29276 21548
rect 29231 21508 29276 21536
rect 29270 21496 29276 21508
rect 29328 21496 29334 21548
rect 29546 21496 29552 21548
rect 29604 21536 29610 21548
rect 29733 21539 29791 21545
rect 29733 21536 29745 21539
rect 29604 21508 29745 21536
rect 29604 21496 29610 21508
rect 29733 21505 29745 21508
rect 29779 21505 29791 21539
rect 30006 21536 30012 21548
rect 29967 21508 30012 21536
rect 29733 21499 29791 21505
rect 30006 21496 30012 21508
rect 30064 21496 30070 21548
rect 32122 21496 32128 21548
rect 32180 21536 32186 21548
rect 32217 21539 32275 21545
rect 32217 21536 32229 21539
rect 32180 21508 32229 21536
rect 32180 21496 32186 21508
rect 32217 21505 32229 21508
rect 32263 21505 32275 21539
rect 32217 21499 32275 21505
rect 26237 21471 26295 21477
rect 26237 21437 26249 21471
rect 26283 21468 26295 21471
rect 26326 21468 26332 21480
rect 26283 21440 26332 21468
rect 26283 21437 26295 21440
rect 26237 21431 26295 21437
rect 26326 21428 26332 21440
rect 26384 21428 26390 21480
rect 31938 21428 31944 21480
rect 31996 21468 32002 21480
rect 32484 21471 32542 21477
rect 32484 21468 32496 21471
rect 31996 21440 32496 21468
rect 31996 21428 32002 21440
rect 32484 21437 32496 21440
rect 32530 21468 32542 21471
rect 33226 21468 33232 21480
rect 32530 21440 33232 21468
rect 32530 21437 32542 21440
rect 32484 21431 32542 21437
rect 33226 21428 33232 21440
rect 33284 21468 33290 21480
rect 33594 21468 33600 21480
rect 33284 21440 33600 21468
rect 33284 21428 33290 21440
rect 33594 21428 33600 21440
rect 33652 21428 33658 21480
rect 34238 21428 34244 21480
rect 34296 21468 34302 21480
rect 34882 21468 34888 21480
rect 34296 21440 34888 21468
rect 34296 21428 34302 21440
rect 34882 21428 34888 21440
rect 34940 21428 34946 21480
rect 35618 21428 35624 21480
rect 35676 21468 35682 21480
rect 36170 21468 36176 21480
rect 35676 21440 36176 21468
rect 35676 21428 35682 21440
rect 36170 21428 36176 21440
rect 36228 21428 36234 21480
rect 20165 21403 20223 21409
rect 20165 21369 20177 21403
rect 20211 21400 20223 21403
rect 21260 21403 21318 21409
rect 21260 21400 21272 21403
rect 20211 21372 21272 21400
rect 20211 21369 20223 21372
rect 20165 21363 20223 21369
rect 21260 21369 21272 21372
rect 21306 21400 21318 21403
rect 21358 21400 21364 21412
rect 21306 21372 21364 21400
rect 21306 21369 21318 21372
rect 21260 21363 21318 21369
rect 21358 21360 21364 21372
rect 21416 21400 21422 21412
rect 22278 21400 22284 21412
rect 21416 21372 22284 21400
rect 21416 21360 21422 21372
rect 22278 21360 22284 21372
rect 22336 21360 22342 21412
rect 23109 21403 23167 21409
rect 23109 21369 23121 21403
rect 23155 21400 23167 21403
rect 23934 21400 23940 21412
rect 23155 21372 23940 21400
rect 23155 21369 23167 21372
rect 23109 21363 23167 21369
rect 23934 21360 23940 21372
rect 23992 21400 23998 21412
rect 24029 21403 24087 21409
rect 24029 21400 24041 21403
rect 23992 21372 24041 21400
rect 23992 21360 23998 21372
rect 24029 21369 24041 21372
rect 24075 21400 24087 21403
rect 24762 21400 24768 21412
rect 24075 21372 24768 21400
rect 24075 21369 24087 21372
rect 24029 21363 24087 21369
rect 24762 21360 24768 21372
rect 24820 21360 24826 21412
rect 26510 21409 26516 21412
rect 26504 21400 26516 21409
rect 26471 21372 26516 21400
rect 26504 21363 26516 21372
rect 26510 21360 26516 21363
rect 26568 21360 26574 21412
rect 27246 21360 27252 21412
rect 27304 21400 27310 21412
rect 28169 21403 28227 21409
rect 28169 21400 28181 21403
rect 27304 21372 28181 21400
rect 27304 21360 27310 21372
rect 28169 21369 28181 21372
rect 28215 21369 28227 21403
rect 32122 21400 32128 21412
rect 32035 21372 32128 21400
rect 28169 21363 28227 21369
rect 32122 21360 32128 21372
rect 32180 21400 32186 21412
rect 34256 21400 34284 21428
rect 32180 21372 34284 21400
rect 35152 21403 35210 21409
rect 32180 21360 32186 21372
rect 35152 21369 35164 21403
rect 35198 21400 35210 21403
rect 35342 21400 35348 21412
rect 35198 21372 35348 21400
rect 35198 21369 35210 21372
rect 35152 21363 35210 21369
rect 35342 21360 35348 21372
rect 35400 21400 35406 21412
rect 36817 21403 36875 21409
rect 36817 21400 36829 21403
rect 35400 21372 36829 21400
rect 35400 21360 35406 21372
rect 36817 21369 36829 21372
rect 36863 21369 36875 21403
rect 36817 21363 36875 21369
rect 23477 21335 23535 21341
rect 23477 21301 23489 21335
rect 23523 21332 23535 21335
rect 23658 21332 23664 21344
rect 23523 21304 23664 21332
rect 23523 21301 23535 21304
rect 23477 21295 23535 21301
rect 23658 21292 23664 21304
rect 23716 21332 23722 21344
rect 24118 21332 24124 21344
rect 23716 21304 24124 21332
rect 23716 21292 23722 21304
rect 24118 21292 24124 21304
rect 24176 21292 24182 21344
rect 24670 21332 24676 21344
rect 24631 21304 24676 21332
rect 24670 21292 24676 21304
rect 24728 21292 24734 21344
rect 25222 21332 25228 21344
rect 25183 21304 25228 21332
rect 25222 21292 25228 21304
rect 25280 21292 25286 21344
rect 26050 21332 26056 21344
rect 26011 21304 26056 21332
rect 26050 21292 26056 21304
rect 26108 21292 26114 21344
rect 29086 21332 29092 21344
rect 28999 21304 29092 21332
rect 29086 21292 29092 21304
rect 29144 21332 29150 21344
rect 29735 21335 29793 21341
rect 29735 21332 29747 21335
rect 29144 21304 29747 21332
rect 29144 21292 29150 21304
rect 29735 21301 29747 21304
rect 29781 21332 29793 21335
rect 29822 21332 29828 21344
rect 29781 21304 29828 21332
rect 29781 21301 29793 21304
rect 29735 21295 29793 21301
rect 29822 21292 29828 21304
rect 29880 21292 29886 21344
rect 30374 21292 30380 21344
rect 30432 21332 30438 21344
rect 31113 21335 31171 21341
rect 31113 21332 31125 21335
rect 30432 21304 31125 21332
rect 30432 21292 30438 21304
rect 31113 21301 31125 21304
rect 31159 21301 31171 21335
rect 31113 21295 31171 21301
rect 32306 21292 32312 21344
rect 32364 21332 32370 21344
rect 33597 21335 33655 21341
rect 33597 21332 33609 21335
rect 32364 21304 33609 21332
rect 32364 21292 32370 21304
rect 33597 21301 33609 21304
rect 33643 21301 33655 21335
rect 37366 21332 37372 21344
rect 37327 21304 37372 21332
rect 33597 21295 33655 21301
rect 37366 21292 37372 21304
rect 37424 21292 37430 21344
rect 1104 21242 38824 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 38824 21242
rect 1104 21168 38824 21190
rect 20714 21128 20720 21140
rect 20675 21100 20720 21128
rect 20714 21088 20720 21100
rect 20772 21088 20778 21140
rect 22278 21128 22284 21140
rect 22239 21100 22284 21128
rect 22278 21088 22284 21100
rect 22336 21088 22342 21140
rect 23198 21128 23204 21140
rect 23159 21100 23204 21128
rect 23198 21088 23204 21100
rect 23256 21088 23262 21140
rect 24762 21128 24768 21140
rect 24723 21100 24768 21128
rect 24762 21088 24768 21100
rect 24820 21088 24826 21140
rect 25961 21131 26019 21137
rect 25961 21097 25973 21131
rect 26007 21128 26019 21131
rect 26786 21128 26792 21140
rect 26007 21100 26792 21128
rect 26007 21097 26019 21100
rect 25961 21091 26019 21097
rect 26786 21088 26792 21100
rect 26844 21088 26850 21140
rect 26878 21088 26884 21140
rect 26936 21128 26942 21140
rect 26973 21131 27031 21137
rect 26973 21128 26985 21131
rect 26936 21100 26985 21128
rect 26936 21088 26942 21100
rect 26973 21097 26985 21100
rect 27019 21097 27031 21131
rect 26973 21091 27031 21097
rect 27617 21131 27675 21137
rect 27617 21097 27629 21131
rect 27663 21128 27675 21131
rect 27706 21128 27712 21140
rect 27663 21100 27712 21128
rect 27663 21097 27675 21100
rect 27617 21091 27675 21097
rect 27706 21088 27712 21100
rect 27764 21088 27770 21140
rect 28994 21088 29000 21140
rect 29052 21128 29058 21140
rect 29733 21131 29791 21137
rect 29733 21128 29745 21131
rect 29052 21100 29745 21128
rect 29052 21088 29058 21100
rect 29733 21097 29745 21100
rect 29779 21097 29791 21131
rect 30650 21128 30656 21140
rect 30611 21100 30656 21128
rect 29733 21091 29791 21097
rect 30650 21088 30656 21100
rect 30708 21088 30714 21140
rect 31938 21128 31944 21140
rect 31899 21100 31944 21128
rect 31938 21088 31944 21100
rect 31996 21088 32002 21140
rect 32766 21128 32772 21140
rect 32048 21100 32772 21128
rect 21168 21063 21226 21069
rect 21168 21029 21180 21063
rect 21214 21060 21226 21063
rect 21358 21060 21364 21072
rect 21214 21032 21364 21060
rect 21214 21029 21226 21032
rect 21168 21023 21226 21029
rect 21358 21020 21364 21032
rect 21416 21020 21422 21072
rect 23474 21020 23480 21072
rect 23532 21060 23538 21072
rect 23658 21069 23664 21072
rect 23652 21060 23664 21069
rect 23532 21032 23664 21060
rect 23532 21020 23538 21032
rect 23652 21023 23664 21032
rect 23658 21020 23664 21023
rect 23716 21020 23722 21072
rect 26142 21020 26148 21072
rect 26200 21060 26206 21072
rect 26326 21060 26332 21072
rect 26200 21032 26332 21060
rect 26200 21020 26206 21032
rect 26326 21020 26332 21032
rect 26384 21060 26390 21072
rect 26384 21032 28396 21060
rect 26384 21020 26390 21032
rect 20898 20992 20904 21004
rect 20859 20964 20904 20992
rect 20898 20952 20904 20964
rect 20956 20952 20962 21004
rect 25222 20952 25228 21004
rect 25280 20992 25286 21004
rect 26694 20992 26700 21004
rect 25280 20964 26700 20992
rect 25280 20952 25286 20964
rect 26694 20952 26700 20964
rect 26752 20992 26758 21004
rect 28368 21001 28396 21032
rect 29822 21020 29828 21072
rect 29880 21060 29886 21072
rect 32048 21060 32076 21100
rect 32766 21088 32772 21100
rect 32824 21128 32830 21140
rect 32955 21131 33013 21137
rect 32955 21128 32967 21131
rect 32824 21100 32967 21128
rect 32824 21088 32830 21100
rect 32955 21097 32967 21100
rect 33001 21128 33013 21131
rect 34238 21128 34244 21140
rect 33001 21100 34244 21128
rect 33001 21097 33013 21100
rect 32955 21091 33013 21097
rect 34238 21088 34244 21100
rect 34296 21088 34302 21140
rect 34333 21131 34391 21137
rect 34333 21097 34345 21131
rect 34379 21128 34391 21131
rect 34422 21128 34428 21140
rect 34379 21100 34428 21128
rect 34379 21097 34391 21100
rect 34333 21091 34391 21097
rect 34422 21088 34428 21100
rect 34480 21128 34486 21140
rect 34606 21128 34612 21140
rect 34480 21100 34612 21128
rect 34480 21088 34486 21100
rect 34606 21088 34612 21100
rect 34664 21088 34670 21140
rect 34882 21128 34888 21140
rect 34843 21100 34888 21128
rect 34882 21088 34888 21100
rect 34940 21088 34946 21140
rect 35342 21128 35348 21140
rect 35303 21100 35348 21128
rect 35342 21088 35348 21100
rect 35400 21088 35406 21140
rect 35802 21128 35808 21140
rect 35763 21100 35808 21128
rect 35802 21088 35808 21100
rect 35860 21088 35866 21140
rect 29880 21032 32076 21060
rect 29880 21020 29886 21032
rect 26881 20995 26939 21001
rect 26881 20992 26893 20995
rect 26752 20964 26893 20992
rect 26752 20952 26758 20964
rect 26881 20961 26893 20964
rect 26927 20961 26939 20995
rect 26881 20955 26939 20961
rect 28353 20995 28411 21001
rect 28353 20961 28365 20995
rect 28399 20992 28411 20995
rect 28442 20992 28448 21004
rect 28399 20964 28448 20992
rect 28399 20961 28411 20964
rect 28353 20955 28411 20961
rect 28442 20952 28448 20964
rect 28500 20952 28506 21004
rect 28626 21001 28632 21004
rect 28620 20992 28632 21001
rect 28587 20964 28632 20992
rect 28620 20955 28632 20964
rect 28626 20952 28632 20955
rect 28684 20952 28690 21004
rect 30926 20952 30932 21004
rect 30984 20992 30990 21004
rect 33134 20992 33140 21004
rect 30984 20964 33140 20992
rect 30984 20952 30990 20964
rect 32416 20936 32444 20964
rect 33134 20952 33140 20964
rect 33192 20952 33198 21004
rect 23290 20884 23296 20936
rect 23348 20924 23354 20936
rect 23385 20927 23443 20933
rect 23385 20924 23397 20927
rect 23348 20896 23397 20924
rect 23348 20884 23354 20896
rect 23385 20893 23397 20896
rect 23431 20893 23443 20927
rect 27154 20924 27160 20936
rect 27115 20896 27160 20924
rect 23385 20887 23443 20893
rect 27154 20884 27160 20896
rect 27212 20884 27218 20936
rect 30282 20884 30288 20936
rect 30340 20924 30346 20936
rect 30837 20927 30895 20933
rect 30837 20924 30849 20927
rect 30340 20896 30849 20924
rect 30340 20884 30346 20896
rect 30837 20893 30849 20896
rect 30883 20893 30895 20927
rect 32306 20924 32312 20936
rect 32267 20896 32312 20924
rect 30837 20887 30895 20893
rect 32306 20884 32312 20896
rect 32364 20884 32370 20936
rect 32398 20884 32404 20936
rect 32456 20924 32462 20936
rect 32493 20927 32551 20933
rect 32493 20924 32505 20927
rect 32456 20896 32505 20924
rect 32456 20884 32462 20896
rect 32493 20893 32505 20896
rect 32539 20893 32551 20927
rect 32950 20924 32956 20936
rect 32911 20896 32956 20924
rect 32493 20887 32551 20893
rect 32950 20884 32956 20896
rect 33008 20884 33014 20936
rect 33229 20927 33287 20933
rect 33229 20893 33241 20927
rect 33275 20924 33287 20927
rect 33318 20924 33324 20936
rect 33275 20896 33324 20924
rect 33275 20893 33287 20896
rect 33229 20887 33287 20893
rect 33318 20884 33324 20896
rect 33376 20884 33382 20936
rect 35710 20884 35716 20936
rect 35768 20924 35774 20936
rect 35897 20927 35955 20933
rect 35897 20924 35909 20927
rect 35768 20896 35909 20924
rect 35768 20884 35774 20896
rect 35897 20893 35909 20896
rect 35943 20893 35955 20927
rect 35897 20887 35955 20893
rect 36081 20927 36139 20933
rect 36081 20893 36093 20927
rect 36127 20924 36139 20927
rect 36262 20924 36268 20936
rect 36127 20896 36268 20924
rect 36127 20893 36139 20896
rect 36081 20887 36139 20893
rect 36262 20884 36268 20896
rect 36320 20884 36326 20936
rect 26513 20859 26571 20865
rect 26513 20825 26525 20859
rect 26559 20856 26571 20859
rect 27246 20856 27252 20868
rect 26559 20828 27252 20856
rect 26559 20825 26571 20828
rect 26513 20819 26571 20825
rect 27246 20816 27252 20828
rect 27304 20816 27310 20868
rect 35437 20859 35495 20865
rect 35437 20825 35449 20859
rect 35483 20856 35495 20859
rect 37458 20856 37464 20868
rect 35483 20828 37464 20856
rect 35483 20825 35495 20828
rect 35437 20819 35495 20825
rect 36096 20800 36124 20828
rect 37458 20816 37464 20828
rect 37516 20816 37522 20868
rect 29638 20748 29644 20800
rect 29696 20788 29702 20800
rect 30285 20791 30343 20797
rect 30285 20788 30297 20791
rect 29696 20760 30297 20788
rect 29696 20748 29702 20760
rect 30285 20757 30297 20760
rect 30331 20788 30343 20791
rect 30374 20788 30380 20800
rect 30331 20760 30380 20788
rect 30331 20757 30343 20760
rect 30285 20751 30343 20757
rect 30374 20748 30380 20760
rect 30432 20748 30438 20800
rect 36078 20748 36084 20800
rect 36136 20748 36142 20800
rect 1104 20698 38824 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 34966 20698
rect 35018 20646 35030 20698
rect 35082 20646 35094 20698
rect 35146 20646 35158 20698
rect 35210 20646 38824 20698
rect 1104 20624 38824 20646
rect 20898 20584 20904 20596
rect 20859 20556 20904 20584
rect 20898 20544 20904 20556
rect 20956 20544 20962 20596
rect 21358 20584 21364 20596
rect 21319 20556 21364 20584
rect 21358 20544 21364 20556
rect 21416 20544 21422 20596
rect 22741 20587 22799 20593
rect 22741 20553 22753 20587
rect 22787 20584 22799 20587
rect 23382 20584 23388 20596
rect 22787 20556 23388 20584
rect 22787 20553 22799 20556
rect 22741 20547 22799 20553
rect 23382 20544 23388 20556
rect 23440 20544 23446 20596
rect 25685 20587 25743 20593
rect 25685 20553 25697 20587
rect 25731 20584 25743 20587
rect 25866 20584 25872 20596
rect 25731 20556 25872 20584
rect 25731 20553 25743 20556
rect 25685 20547 25743 20553
rect 25866 20544 25872 20556
rect 25924 20584 25930 20596
rect 27154 20584 27160 20596
rect 25924 20556 27160 20584
rect 25924 20544 25930 20556
rect 27154 20544 27160 20556
rect 27212 20584 27218 20596
rect 27525 20587 27583 20593
rect 27525 20584 27537 20587
rect 27212 20556 27537 20584
rect 27212 20544 27218 20556
rect 27525 20553 27537 20556
rect 27571 20553 27583 20587
rect 32582 20584 32588 20596
rect 32543 20556 32588 20584
rect 27525 20547 27583 20553
rect 32582 20544 32588 20556
rect 32640 20544 32646 20596
rect 33134 20544 33140 20596
rect 33192 20584 33198 20596
rect 33597 20587 33655 20593
rect 33597 20584 33609 20587
rect 33192 20556 33609 20584
rect 33192 20544 33198 20556
rect 33597 20553 33609 20556
rect 33643 20553 33655 20587
rect 34606 20584 34612 20596
rect 34567 20556 34612 20584
rect 33597 20547 33655 20553
rect 34606 20544 34612 20556
rect 34664 20544 34670 20596
rect 35894 20584 35900 20596
rect 35855 20556 35900 20584
rect 35894 20544 35900 20556
rect 35952 20544 35958 20596
rect 36262 20584 36268 20596
rect 36223 20556 36268 20584
rect 36262 20544 36268 20556
rect 36320 20544 36326 20596
rect 20916 20516 20944 20544
rect 22462 20516 22468 20528
rect 20916 20488 22468 20516
rect 22462 20476 22468 20488
rect 22520 20476 22526 20528
rect 29362 20516 29368 20528
rect 29323 20488 29368 20516
rect 29362 20476 29368 20488
rect 29420 20476 29426 20528
rect 30377 20519 30435 20525
rect 30377 20516 30389 20519
rect 29840 20488 30389 20516
rect 26053 20451 26111 20457
rect 26053 20417 26065 20451
rect 26099 20448 26111 20451
rect 26142 20448 26148 20460
rect 26099 20420 26148 20448
rect 26099 20417 26111 20420
rect 26053 20411 26111 20417
rect 23934 20389 23940 20392
rect 23661 20383 23719 20389
rect 23661 20349 23673 20383
rect 23707 20349 23719 20383
rect 23928 20380 23940 20389
rect 23895 20352 23940 20380
rect 23661 20343 23719 20349
rect 23928 20343 23940 20352
rect 23109 20315 23167 20321
rect 23109 20281 23121 20315
rect 23155 20312 23167 20315
rect 23290 20312 23296 20324
rect 23155 20284 23296 20312
rect 23155 20281 23167 20284
rect 23109 20275 23167 20281
rect 23290 20272 23296 20284
rect 23348 20312 23354 20324
rect 23477 20315 23535 20321
rect 23477 20312 23489 20315
rect 23348 20284 23489 20312
rect 23348 20272 23354 20284
rect 23477 20281 23489 20284
rect 23523 20312 23535 20315
rect 23676 20312 23704 20343
rect 23934 20340 23940 20343
rect 23992 20340 23998 20392
rect 26068 20312 26096 20411
rect 26142 20408 26148 20420
rect 26200 20408 26206 20460
rect 29730 20408 29736 20460
rect 29788 20448 29794 20460
rect 29840 20457 29868 20488
rect 30377 20485 30389 20488
rect 30423 20485 30435 20519
rect 30377 20479 30435 20485
rect 32493 20519 32551 20525
rect 32493 20485 32505 20519
rect 32539 20516 32551 20519
rect 32766 20516 32772 20528
rect 32539 20488 32772 20516
rect 32539 20485 32551 20488
rect 32493 20479 32551 20485
rect 32600 20460 32628 20488
rect 32766 20476 32772 20488
rect 32824 20476 32830 20528
rect 34885 20519 34943 20525
rect 34885 20485 34897 20519
rect 34931 20516 34943 20519
rect 35710 20516 35716 20528
rect 34931 20488 35716 20516
rect 34931 20485 34943 20488
rect 34885 20479 34943 20485
rect 35710 20476 35716 20488
rect 35768 20516 35774 20528
rect 36633 20519 36691 20525
rect 36633 20516 36645 20519
rect 35768 20488 36645 20516
rect 35768 20476 35774 20488
rect 36633 20485 36645 20488
rect 36679 20485 36691 20519
rect 36633 20479 36691 20485
rect 29825 20451 29883 20457
rect 29825 20448 29837 20451
rect 29788 20420 29837 20448
rect 29788 20408 29794 20420
rect 29825 20417 29837 20420
rect 29871 20417 29883 20451
rect 30006 20448 30012 20460
rect 29919 20420 30012 20448
rect 29825 20411 29883 20417
rect 30006 20408 30012 20420
rect 30064 20448 30070 20460
rect 30466 20448 30472 20460
rect 30064 20420 30472 20448
rect 30064 20408 30070 20420
rect 30466 20408 30472 20420
rect 30524 20408 30530 20460
rect 31573 20451 31631 20457
rect 31573 20417 31585 20451
rect 31619 20448 31631 20451
rect 31662 20448 31668 20460
rect 31619 20420 31668 20448
rect 31619 20417 31631 20420
rect 31573 20411 31631 20417
rect 31662 20408 31668 20420
rect 31720 20408 31726 20460
rect 32582 20408 32588 20460
rect 32640 20408 32646 20460
rect 33226 20448 33232 20460
rect 33187 20420 33232 20448
rect 33226 20408 33232 20420
rect 33284 20408 33290 20460
rect 35342 20408 35348 20460
rect 35400 20448 35406 20460
rect 35437 20451 35495 20457
rect 35437 20448 35449 20451
rect 35400 20420 35449 20448
rect 35400 20408 35406 20420
rect 35437 20417 35449 20420
rect 35483 20417 35495 20451
rect 35437 20411 35495 20417
rect 26234 20340 26240 20392
rect 26292 20380 26298 20392
rect 26401 20383 26459 20389
rect 26401 20380 26413 20383
rect 26292 20352 26413 20380
rect 26292 20340 26298 20352
rect 26401 20349 26413 20352
rect 26447 20349 26459 20383
rect 26401 20343 26459 20349
rect 23523 20284 26096 20312
rect 29089 20315 29147 20321
rect 23523 20281 23535 20284
rect 23477 20275 23535 20281
rect 29089 20281 29101 20315
rect 29135 20312 29147 20315
rect 29733 20315 29791 20321
rect 29733 20312 29745 20315
rect 29135 20284 29745 20312
rect 29135 20281 29147 20284
rect 29089 20275 29147 20281
rect 29733 20281 29745 20284
rect 29779 20312 29791 20315
rect 30282 20312 30288 20324
rect 29779 20284 30288 20312
rect 29779 20281 29791 20284
rect 29733 20275 29791 20281
rect 30282 20272 30288 20284
rect 30340 20272 30346 20324
rect 32125 20315 32183 20321
rect 32125 20281 32137 20315
rect 32171 20312 32183 20315
rect 33318 20312 33324 20324
rect 32171 20284 33324 20312
rect 32171 20281 32183 20284
rect 32125 20275 32183 20281
rect 32968 20256 32996 20284
rect 33318 20272 33324 20284
rect 33376 20272 33382 20324
rect 34606 20272 34612 20324
rect 34664 20312 34670 20324
rect 35345 20315 35403 20321
rect 35345 20312 35357 20315
rect 34664 20284 35357 20312
rect 34664 20272 34670 20284
rect 35345 20281 35357 20284
rect 35391 20281 35403 20315
rect 35345 20275 35403 20281
rect 25038 20244 25044 20256
rect 24999 20216 25044 20244
rect 25038 20204 25044 20216
rect 25096 20204 25102 20256
rect 28442 20244 28448 20256
rect 28355 20216 28448 20244
rect 28442 20204 28448 20216
rect 28500 20244 28506 20256
rect 28810 20244 28816 20256
rect 28500 20216 28816 20244
rect 28500 20204 28506 20216
rect 28810 20204 28816 20216
rect 28868 20204 28874 20256
rect 32950 20244 32956 20256
rect 32911 20216 32956 20244
rect 32950 20204 32956 20216
rect 33008 20204 33014 20256
rect 33042 20204 33048 20256
rect 33100 20244 33106 20256
rect 34333 20247 34391 20253
rect 34333 20244 34345 20247
rect 33100 20216 34345 20244
rect 33100 20204 33106 20216
rect 34333 20213 34345 20216
rect 34379 20244 34391 20247
rect 34422 20244 34428 20256
rect 34379 20216 34428 20244
rect 34379 20213 34391 20216
rect 34333 20207 34391 20213
rect 34422 20204 34428 20216
rect 34480 20244 34486 20256
rect 35253 20247 35311 20253
rect 35253 20244 35265 20247
rect 34480 20216 35265 20244
rect 34480 20204 34486 20216
rect 35253 20213 35265 20216
rect 35299 20213 35311 20247
rect 35253 20207 35311 20213
rect 1104 20154 38824 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 38824 20154
rect 1104 20080 38824 20102
rect 23750 20000 23756 20052
rect 23808 20040 23814 20052
rect 23845 20043 23903 20049
rect 23845 20040 23857 20043
rect 23808 20012 23857 20040
rect 23808 20000 23814 20012
rect 23845 20009 23857 20012
rect 23891 20009 23903 20043
rect 23845 20003 23903 20009
rect 23934 20000 23940 20052
rect 23992 20040 23998 20052
rect 24397 20043 24455 20049
rect 24397 20040 24409 20043
rect 23992 20012 24409 20040
rect 23992 20000 23998 20012
rect 24397 20009 24409 20012
rect 24443 20009 24455 20043
rect 26234 20040 26240 20052
rect 26195 20012 26240 20040
rect 24397 20003 24455 20009
rect 26234 20000 26240 20012
rect 26292 20000 26298 20052
rect 26694 20040 26700 20052
rect 26655 20012 26700 20040
rect 26694 20000 26700 20012
rect 26752 20000 26758 20052
rect 26878 20000 26884 20052
rect 26936 20040 26942 20052
rect 27065 20043 27123 20049
rect 27065 20040 27077 20043
rect 26936 20012 27077 20040
rect 26936 20000 26942 20012
rect 27065 20009 27077 20012
rect 27111 20009 27123 20043
rect 27065 20003 27123 20009
rect 28445 20043 28503 20049
rect 28445 20009 28457 20043
rect 28491 20040 28503 20043
rect 28626 20040 28632 20052
rect 28491 20012 28632 20040
rect 28491 20009 28503 20012
rect 28445 20003 28503 20009
rect 28626 20000 28632 20012
rect 28684 20000 28690 20052
rect 29457 20043 29515 20049
rect 29457 20009 29469 20043
rect 29503 20040 29515 20043
rect 30006 20040 30012 20052
rect 29503 20012 30012 20040
rect 29503 20009 29515 20012
rect 29457 20003 29515 20009
rect 30006 20000 30012 20012
rect 30064 20000 30070 20052
rect 33042 20040 33048 20052
rect 33003 20012 33048 20040
rect 33042 20000 33048 20012
rect 33100 20000 33106 20052
rect 33226 20000 33232 20052
rect 33284 20040 33290 20052
rect 33321 20043 33379 20049
rect 33321 20040 33333 20043
rect 33284 20012 33333 20040
rect 33284 20000 33290 20012
rect 33321 20009 33333 20012
rect 33367 20009 33379 20043
rect 33321 20003 33379 20009
rect 35342 20000 35348 20052
rect 35400 20040 35406 20052
rect 36081 20043 36139 20049
rect 36081 20040 36093 20043
rect 35400 20012 36093 20040
rect 35400 20000 35406 20012
rect 36081 20009 36093 20012
rect 36127 20009 36139 20043
rect 36081 20003 36139 20009
rect 22738 19913 22744 19916
rect 22732 19904 22744 19913
rect 22699 19876 22744 19904
rect 22732 19867 22744 19876
rect 22738 19864 22744 19867
rect 22796 19864 22802 19916
rect 34968 19907 35026 19913
rect 34968 19873 34980 19907
rect 35014 19904 35026 19907
rect 35526 19904 35532 19916
rect 35014 19876 35532 19904
rect 35014 19873 35026 19876
rect 34968 19867 35026 19873
rect 35526 19864 35532 19876
rect 35584 19864 35590 19916
rect 22462 19836 22468 19848
rect 22423 19808 22468 19836
rect 22462 19796 22468 19808
rect 22520 19796 22526 19848
rect 33689 19839 33747 19845
rect 33689 19805 33701 19839
rect 33735 19836 33747 19839
rect 34606 19836 34612 19848
rect 33735 19808 34612 19836
rect 33735 19805 33747 19808
rect 33689 19799 33747 19805
rect 34606 19796 34612 19808
rect 34664 19796 34670 19848
rect 34701 19839 34759 19845
rect 34701 19805 34713 19839
rect 34747 19805 34759 19839
rect 34701 19799 34759 19805
rect 29825 19703 29883 19709
rect 29825 19669 29837 19703
rect 29871 19700 29883 19703
rect 30006 19700 30012 19712
rect 29871 19672 30012 19700
rect 29871 19669 29883 19672
rect 29825 19663 29883 19669
rect 30006 19660 30012 19672
rect 30064 19660 30070 19712
rect 32677 19703 32735 19709
rect 32677 19669 32689 19703
rect 32723 19700 32735 19703
rect 33042 19700 33048 19712
rect 32723 19672 33048 19700
rect 32723 19669 32735 19672
rect 32677 19663 32735 19669
rect 33042 19660 33048 19672
rect 33100 19660 33106 19712
rect 34606 19700 34612 19712
rect 34567 19672 34612 19700
rect 34606 19660 34612 19672
rect 34664 19660 34670 19712
rect 34716 19700 34744 19799
rect 35342 19700 35348 19712
rect 34716 19672 35348 19700
rect 35342 19660 35348 19672
rect 35400 19660 35406 19712
rect 1104 19610 38824 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 34966 19610
rect 35018 19558 35030 19610
rect 35082 19558 35094 19610
rect 35146 19558 35158 19610
rect 35210 19558 38824 19610
rect 1104 19536 38824 19558
rect 22738 19456 22744 19508
rect 22796 19496 22802 19508
rect 22833 19499 22891 19505
rect 22833 19496 22845 19499
rect 22796 19468 22845 19496
rect 22796 19456 22802 19468
rect 22833 19465 22845 19468
rect 22879 19465 22891 19499
rect 33870 19496 33876 19508
rect 33831 19468 33876 19496
rect 22833 19459 22891 19465
rect 33870 19456 33876 19468
rect 33928 19456 33934 19508
rect 34422 19456 34428 19508
rect 34480 19496 34486 19508
rect 34885 19499 34943 19505
rect 34885 19496 34897 19499
rect 34480 19468 34897 19496
rect 34480 19456 34486 19468
rect 34885 19465 34897 19468
rect 34931 19465 34943 19499
rect 34885 19459 34943 19465
rect 22462 19388 22468 19440
rect 22520 19428 22526 19440
rect 22557 19431 22615 19437
rect 22557 19428 22569 19431
rect 22520 19400 22569 19428
rect 22520 19388 22526 19400
rect 22557 19397 22569 19400
rect 22603 19428 22615 19431
rect 23290 19428 23296 19440
rect 22603 19400 23296 19428
rect 22603 19397 22615 19400
rect 22557 19391 22615 19397
rect 23290 19388 23296 19400
rect 23348 19388 23354 19440
rect 34333 19431 34391 19437
rect 34333 19397 34345 19431
rect 34379 19428 34391 19431
rect 34379 19400 35572 19428
rect 34379 19397 34391 19400
rect 34333 19391 34391 19397
rect 35544 19372 35572 19400
rect 34606 19320 34612 19372
rect 34664 19360 34670 19372
rect 35158 19360 35164 19372
rect 34664 19332 35164 19360
rect 34664 19320 34670 19332
rect 35158 19320 35164 19332
rect 35216 19360 35222 19372
rect 35345 19363 35403 19369
rect 35345 19360 35357 19363
rect 35216 19332 35357 19360
rect 35216 19320 35222 19332
rect 35345 19329 35357 19332
rect 35391 19329 35403 19363
rect 35526 19360 35532 19372
rect 35439 19332 35532 19360
rect 35345 19323 35403 19329
rect 35526 19320 35532 19332
rect 35584 19360 35590 19372
rect 35584 19332 35940 19360
rect 35584 19320 35590 19332
rect 29733 19295 29791 19301
rect 29733 19292 29745 19295
rect 29564 19264 29745 19292
rect 28810 19116 28816 19168
rect 28868 19156 28874 19168
rect 29564 19165 29592 19264
rect 29733 19261 29745 19264
rect 29779 19261 29791 19295
rect 33689 19295 33747 19301
rect 33689 19292 33701 19295
rect 29733 19255 29791 19261
rect 33520 19264 33701 19292
rect 30006 19233 30012 19236
rect 30000 19224 30012 19233
rect 29967 19196 30012 19224
rect 30000 19187 30012 19196
rect 30006 19184 30012 19187
rect 30064 19184 30070 19236
rect 33520 19168 33548 19264
rect 33689 19261 33701 19264
rect 33735 19261 33747 19295
rect 33689 19255 33747 19261
rect 34698 19184 34704 19236
rect 34756 19224 34762 19236
rect 35253 19227 35311 19233
rect 35253 19224 35265 19227
rect 34756 19196 35265 19224
rect 34756 19184 34762 19196
rect 35253 19193 35265 19196
rect 35299 19193 35311 19227
rect 35253 19187 35311 19193
rect 29549 19159 29607 19165
rect 29549 19156 29561 19159
rect 28868 19128 29561 19156
rect 28868 19116 28874 19128
rect 29549 19125 29561 19128
rect 29595 19125 29607 19159
rect 29549 19119 29607 19125
rect 31018 19116 31024 19168
rect 31076 19156 31082 19168
rect 31113 19159 31171 19165
rect 31113 19156 31125 19159
rect 31076 19128 31125 19156
rect 31076 19116 31082 19128
rect 31113 19125 31125 19128
rect 31159 19125 31171 19159
rect 31113 19119 31171 19125
rect 32398 19116 32404 19168
rect 32456 19156 32462 19168
rect 32493 19159 32551 19165
rect 32493 19156 32505 19159
rect 32456 19128 32505 19156
rect 32456 19116 32462 19128
rect 32493 19125 32505 19128
rect 32539 19125 32551 19159
rect 33502 19156 33508 19168
rect 33463 19128 33508 19156
rect 32493 19119 32551 19125
rect 33502 19116 33508 19128
rect 33560 19116 33566 19168
rect 34330 19116 34336 19168
rect 34388 19156 34394 19168
rect 34609 19159 34667 19165
rect 34609 19156 34621 19159
rect 34388 19128 34621 19156
rect 34388 19116 34394 19128
rect 34609 19125 34621 19128
rect 34655 19156 34667 19159
rect 35342 19156 35348 19168
rect 34655 19128 35348 19156
rect 34655 19125 34667 19128
rect 34609 19119 34667 19125
rect 35342 19116 35348 19128
rect 35400 19116 35406 19168
rect 35912 19156 35940 19332
rect 36449 19295 36507 19301
rect 36449 19261 36461 19295
rect 36495 19292 36507 19295
rect 37182 19292 37188 19304
rect 36495 19264 37188 19292
rect 36495 19261 36507 19264
rect 36449 19255 36507 19261
rect 37182 19252 37188 19264
rect 37240 19252 37246 19304
rect 36633 19227 36691 19233
rect 36633 19224 36645 19227
rect 36280 19196 36645 19224
rect 36280 19168 36308 19196
rect 36633 19193 36645 19196
rect 36679 19193 36691 19227
rect 36633 19187 36691 19193
rect 35986 19156 35992 19168
rect 35912 19128 35992 19156
rect 35986 19116 35992 19128
rect 36044 19116 36050 19168
rect 36262 19156 36268 19168
rect 36223 19128 36268 19156
rect 36262 19116 36268 19128
rect 36320 19116 36326 19168
rect 36814 19156 36820 19168
rect 36775 19128 36820 19156
rect 36814 19116 36820 19128
rect 36872 19116 36878 19168
rect 1104 19066 38824 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 38824 19066
rect 1104 18992 38824 19014
rect 25866 18952 25872 18964
rect 25827 18924 25872 18952
rect 25866 18912 25872 18924
rect 25924 18912 25930 18964
rect 34698 18912 34704 18964
rect 34756 18952 34762 18964
rect 34885 18955 34943 18961
rect 34885 18952 34897 18955
rect 34756 18924 34897 18952
rect 34756 18912 34762 18924
rect 34885 18921 34897 18924
rect 34931 18921 34943 18955
rect 35158 18952 35164 18964
rect 35119 18924 35164 18952
rect 34885 18915 34943 18921
rect 35158 18912 35164 18924
rect 35216 18912 35222 18964
rect 28258 18844 28264 18896
rect 28316 18884 28322 18896
rect 28721 18887 28779 18893
rect 28721 18884 28733 18887
rect 28316 18856 28733 18884
rect 28316 18844 28322 18856
rect 28721 18853 28733 18856
rect 28767 18884 28779 18887
rect 29914 18884 29920 18896
rect 28767 18856 29920 18884
rect 28767 18853 28779 18856
rect 28721 18847 28779 18853
rect 29914 18844 29920 18856
rect 29972 18844 29978 18896
rect 28166 18776 28172 18828
rect 28224 18816 28230 18828
rect 29069 18819 29127 18825
rect 29069 18816 29081 18819
rect 28224 18788 29081 18816
rect 28224 18776 28230 18788
rect 29069 18785 29081 18788
rect 29115 18785 29127 18819
rect 29069 18779 29127 18785
rect 32677 18819 32735 18825
rect 32677 18785 32689 18819
rect 32723 18816 32735 18819
rect 32766 18816 32772 18828
rect 32723 18788 32772 18816
rect 32723 18785 32735 18788
rect 32677 18779 32735 18785
rect 32766 18776 32772 18788
rect 32824 18776 32830 18828
rect 32950 18825 32956 18828
rect 32944 18816 32956 18825
rect 32911 18788 32956 18816
rect 32944 18779 32956 18788
rect 32950 18776 32956 18779
rect 33008 18776 33014 18828
rect 34238 18776 34244 18828
rect 34296 18816 34302 18828
rect 35529 18819 35587 18825
rect 35529 18816 35541 18819
rect 34296 18788 35541 18816
rect 34296 18776 34302 18788
rect 35529 18785 35541 18788
rect 35575 18785 35587 18819
rect 35529 18779 35587 18785
rect 28810 18748 28816 18760
rect 28771 18720 28816 18748
rect 28810 18708 28816 18720
rect 28868 18708 28874 18760
rect 34422 18708 34428 18760
rect 34480 18748 34486 18760
rect 35621 18751 35679 18757
rect 35621 18748 35633 18751
rect 34480 18720 35633 18748
rect 34480 18708 34486 18720
rect 35621 18717 35633 18720
rect 35667 18717 35679 18751
rect 35621 18711 35679 18717
rect 35636 18680 35664 18711
rect 35710 18708 35716 18760
rect 35768 18748 35774 18760
rect 36173 18751 36231 18757
rect 36173 18748 36185 18751
rect 35768 18720 36185 18748
rect 35768 18708 35774 18720
rect 36173 18717 36185 18720
rect 36219 18717 36231 18751
rect 36173 18711 36231 18717
rect 36814 18680 36820 18692
rect 35636 18652 36820 18680
rect 36814 18640 36820 18652
rect 36872 18640 36878 18692
rect 28994 18572 29000 18624
rect 29052 18612 29058 18624
rect 30006 18612 30012 18624
rect 29052 18584 30012 18612
rect 29052 18572 29058 18584
rect 30006 18572 30012 18584
rect 30064 18612 30070 18624
rect 30193 18615 30251 18621
rect 30193 18612 30205 18615
rect 30064 18584 30205 18612
rect 30064 18572 30070 18584
rect 30193 18581 30205 18584
rect 30239 18581 30251 18615
rect 31018 18612 31024 18624
rect 30979 18584 31024 18612
rect 30193 18575 30251 18581
rect 31018 18572 31024 18584
rect 31076 18572 31082 18624
rect 34054 18612 34060 18624
rect 34015 18584 34060 18612
rect 34054 18572 34060 18584
rect 34112 18572 34118 18624
rect 1104 18522 38824 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 34966 18522
rect 35018 18470 35030 18522
rect 35082 18470 35094 18522
rect 35146 18470 35158 18522
rect 35210 18470 38824 18522
rect 1104 18448 38824 18470
rect 25685 18411 25743 18417
rect 25685 18377 25697 18411
rect 25731 18408 25743 18411
rect 26142 18408 26148 18420
rect 25731 18380 26148 18408
rect 25731 18377 25743 18380
rect 25685 18371 25743 18377
rect 24486 18232 24492 18284
rect 24544 18272 24550 18284
rect 25792 18281 25820 18380
rect 26142 18368 26148 18380
rect 26200 18368 26206 18420
rect 35986 18368 35992 18420
rect 36044 18408 36050 18420
rect 36265 18411 36323 18417
rect 36265 18408 36277 18411
rect 36044 18380 36277 18408
rect 36044 18368 36050 18380
rect 36265 18377 36277 18380
rect 36311 18377 36323 18411
rect 36814 18408 36820 18420
rect 36775 18380 36820 18408
rect 36265 18371 36323 18377
rect 36814 18368 36820 18380
rect 36872 18368 36878 18420
rect 29089 18343 29147 18349
rect 29089 18309 29101 18343
rect 29135 18340 29147 18343
rect 30745 18343 30803 18349
rect 30745 18340 30757 18343
rect 29135 18312 30757 18340
rect 29135 18309 29147 18312
rect 29089 18303 29147 18309
rect 30745 18309 30757 18312
rect 30791 18340 30803 18343
rect 33873 18343 33931 18349
rect 30791 18312 30972 18340
rect 30791 18309 30803 18312
rect 30745 18303 30803 18309
rect 25777 18275 25835 18281
rect 25777 18272 25789 18275
rect 24544 18244 25789 18272
rect 24544 18232 24550 18244
rect 25777 18241 25789 18244
rect 25823 18241 25835 18275
rect 29914 18272 29920 18284
rect 29875 18244 29920 18272
rect 25777 18235 25835 18241
rect 29914 18232 29920 18244
rect 29972 18232 29978 18284
rect 30944 18281 30972 18312
rect 33873 18309 33885 18343
rect 33919 18340 33931 18343
rect 34606 18340 34612 18352
rect 33919 18312 34612 18340
rect 33919 18309 33931 18312
rect 33873 18303 33931 18309
rect 34606 18300 34612 18312
rect 34664 18300 34670 18352
rect 30929 18275 30987 18281
rect 30929 18241 30941 18275
rect 30975 18241 30987 18275
rect 30929 18235 30987 18241
rect 18874 18204 18880 18216
rect 18835 18176 18880 18204
rect 18874 18164 18880 18176
rect 18932 18164 18938 18216
rect 25866 18164 25872 18216
rect 25924 18204 25930 18216
rect 26033 18207 26091 18213
rect 26033 18204 26045 18207
rect 25924 18176 26045 18204
rect 25924 18164 25930 18176
rect 26033 18173 26045 18176
rect 26079 18173 26091 18207
rect 28534 18204 28540 18216
rect 28447 18176 28540 18204
rect 26033 18167 26091 18173
rect 28534 18164 28540 18176
rect 28592 18204 28598 18216
rect 29730 18204 29736 18216
rect 28592 18176 29736 18204
rect 28592 18164 28598 18176
rect 29730 18164 29736 18176
rect 29788 18164 29794 18216
rect 30944 18204 30972 18235
rect 32766 18204 32772 18216
rect 30944 18176 32772 18204
rect 32766 18164 32772 18176
rect 32824 18204 32830 18216
rect 32861 18207 32919 18213
rect 32861 18204 32873 18207
rect 32824 18176 32873 18204
rect 32824 18164 32830 18176
rect 32861 18173 32873 18176
rect 32907 18204 32919 18207
rect 33686 18204 33692 18216
rect 32907 18176 33364 18204
rect 33647 18176 33692 18204
rect 32907 18173 32919 18176
rect 32861 18167 32919 18173
rect 18690 18136 18696 18148
rect 18651 18108 18696 18136
rect 18690 18096 18696 18108
rect 18748 18136 18754 18148
rect 19122 18139 19180 18145
rect 19122 18136 19134 18139
rect 18748 18108 19134 18136
rect 18748 18096 18754 18108
rect 19122 18105 19134 18108
rect 19168 18105 19180 18139
rect 19122 18099 19180 18105
rect 28074 18096 28080 18148
rect 28132 18136 28138 18148
rect 28810 18136 28816 18148
rect 28132 18108 28816 18136
rect 28132 18096 28138 18108
rect 28810 18096 28816 18108
rect 28868 18136 28874 18148
rect 29089 18139 29147 18145
rect 29089 18136 29101 18139
rect 28868 18108 29101 18136
rect 28868 18096 28874 18108
rect 29089 18105 29101 18108
rect 29135 18105 29147 18139
rect 29089 18099 29147 18105
rect 29641 18139 29699 18145
rect 29641 18105 29653 18139
rect 29687 18136 29699 18139
rect 29687 18108 30328 18136
rect 29687 18105 29699 18108
rect 29641 18099 29699 18105
rect 30300 18080 30328 18108
rect 31018 18096 31024 18148
rect 31076 18136 31082 18148
rect 31196 18139 31254 18145
rect 31196 18136 31208 18139
rect 31076 18108 31208 18136
rect 31076 18096 31082 18108
rect 31196 18105 31208 18108
rect 31242 18136 31254 18139
rect 31662 18136 31668 18148
rect 31242 18108 31668 18136
rect 31242 18105 31254 18108
rect 31196 18099 31254 18105
rect 31662 18096 31668 18108
rect 31720 18096 31726 18148
rect 32950 18136 32956 18148
rect 32324 18108 32956 18136
rect 32324 18080 32352 18108
rect 32950 18096 32956 18108
rect 33008 18136 33014 18148
rect 33229 18139 33287 18145
rect 33229 18136 33241 18139
rect 33008 18108 33241 18136
rect 33008 18096 33014 18108
rect 33229 18105 33241 18108
rect 33275 18105 33287 18139
rect 33336 18136 33364 18176
rect 33686 18164 33692 18176
rect 33744 18164 33750 18216
rect 34885 18207 34943 18213
rect 34885 18173 34897 18207
rect 34931 18173 34943 18207
rect 34885 18167 34943 18173
rect 34330 18136 34336 18148
rect 33336 18108 34336 18136
rect 33229 18099 33287 18105
rect 34330 18096 34336 18108
rect 34388 18136 34394 18148
rect 34609 18139 34667 18145
rect 34609 18136 34621 18139
rect 34388 18108 34621 18136
rect 34388 18096 34394 18108
rect 34609 18105 34621 18108
rect 34655 18136 34667 18139
rect 34900 18136 34928 18167
rect 34655 18108 34928 18136
rect 34655 18105 34667 18108
rect 34609 18099 34667 18105
rect 35066 18096 35072 18148
rect 35124 18145 35130 18148
rect 35124 18139 35188 18145
rect 35124 18105 35142 18139
rect 35176 18105 35188 18139
rect 35124 18099 35188 18105
rect 35124 18096 35130 18099
rect 20254 18068 20260 18080
rect 20215 18040 20260 18068
rect 20254 18028 20260 18040
rect 20312 18028 20318 18080
rect 27154 18068 27160 18080
rect 27115 18040 27160 18068
rect 27154 18028 27160 18040
rect 27212 18028 27218 18080
rect 28166 18068 28172 18080
rect 28127 18040 28172 18068
rect 28166 18028 28172 18040
rect 28224 18028 28230 18080
rect 29270 18068 29276 18080
rect 29231 18040 29276 18068
rect 29270 18028 29276 18040
rect 29328 18028 29334 18080
rect 30282 18068 30288 18080
rect 30243 18040 30288 18068
rect 30282 18028 30288 18040
rect 30340 18028 30346 18080
rect 32306 18068 32312 18080
rect 32267 18040 32312 18068
rect 32306 18028 32312 18040
rect 32364 18028 32370 18080
rect 33134 18028 33140 18080
rect 33192 18068 33198 18080
rect 34238 18068 34244 18080
rect 33192 18040 34244 18068
rect 33192 18028 33198 18040
rect 34238 18028 34244 18040
rect 34296 18028 34302 18080
rect 1104 17978 38824 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 38824 17978
rect 1104 17904 38824 17926
rect 29546 17864 29552 17876
rect 29459 17836 29552 17864
rect 29546 17824 29552 17836
rect 29604 17864 29610 17876
rect 30193 17867 30251 17873
rect 30193 17864 30205 17867
rect 29604 17836 30205 17864
rect 29604 17824 29610 17836
rect 30193 17833 30205 17836
rect 30239 17864 30251 17867
rect 30282 17864 30288 17876
rect 30239 17836 30288 17864
rect 30239 17833 30251 17836
rect 30193 17827 30251 17833
rect 30282 17824 30288 17836
rect 30340 17824 30346 17876
rect 31113 17867 31171 17873
rect 31113 17833 31125 17867
rect 31159 17864 31171 17867
rect 33134 17864 33140 17876
rect 31159 17836 33140 17864
rect 31159 17833 31171 17836
rect 31113 17827 31171 17833
rect 33134 17824 33140 17836
rect 33192 17864 33198 17876
rect 33229 17867 33287 17873
rect 33229 17864 33241 17867
rect 33192 17836 33241 17864
rect 33192 17824 33198 17836
rect 33229 17833 33241 17836
rect 33275 17833 33287 17867
rect 33229 17827 33287 17833
rect 33686 17824 33692 17876
rect 33744 17864 33750 17876
rect 33873 17867 33931 17873
rect 33873 17864 33885 17867
rect 33744 17836 33885 17864
rect 33744 17824 33750 17836
rect 33873 17833 33885 17836
rect 33919 17833 33931 17867
rect 33873 17827 33931 17833
rect 34333 17867 34391 17873
rect 34333 17833 34345 17867
rect 34379 17864 34391 17867
rect 35066 17864 35072 17876
rect 34379 17836 35072 17864
rect 34379 17833 34391 17836
rect 34333 17827 34391 17833
rect 35066 17824 35072 17836
rect 35124 17864 35130 17876
rect 35710 17864 35716 17876
rect 35124 17836 35716 17864
rect 35124 17824 35130 17836
rect 35710 17824 35716 17836
rect 35768 17864 35774 17876
rect 35805 17867 35863 17873
rect 35805 17864 35817 17867
rect 35768 17836 35817 17864
rect 35768 17824 35774 17836
rect 35805 17833 35817 17836
rect 35851 17833 35863 17867
rect 35805 17827 35863 17833
rect 28436 17799 28494 17805
rect 28436 17765 28448 17799
rect 28482 17796 28494 17799
rect 28534 17796 28540 17808
rect 28482 17768 28540 17796
rect 28482 17765 28494 17768
rect 28436 17759 28494 17765
rect 28534 17756 28540 17768
rect 28592 17756 28598 17808
rect 11606 17737 11612 17740
rect 11600 17728 11612 17737
rect 11567 17700 11612 17728
rect 11600 17691 11612 17700
rect 11606 17688 11612 17691
rect 11664 17688 11670 17740
rect 21720 17731 21778 17737
rect 21720 17697 21732 17731
rect 21766 17728 21778 17731
rect 22646 17728 22652 17740
rect 21766 17700 22652 17728
rect 21766 17697 21778 17700
rect 21720 17691 21778 17697
rect 22646 17688 22652 17700
rect 22704 17688 22710 17740
rect 23106 17688 23112 17740
rect 23164 17728 23170 17740
rect 24193 17731 24251 17737
rect 24193 17728 24205 17731
rect 23164 17700 24205 17728
rect 23164 17688 23170 17700
rect 24193 17697 24205 17700
rect 24239 17697 24251 17731
rect 30926 17728 30932 17740
rect 30887 17700 30932 17728
rect 24193 17691 24251 17697
rect 30926 17688 30932 17700
rect 30984 17688 30990 17740
rect 33594 17688 33600 17740
rect 33652 17728 33658 17740
rect 34054 17728 34060 17740
rect 33652 17700 34060 17728
rect 33652 17688 33658 17700
rect 34054 17688 34060 17700
rect 34112 17728 34118 17740
rect 34681 17731 34739 17737
rect 34681 17728 34693 17731
rect 34112 17700 34693 17728
rect 34112 17688 34118 17700
rect 34681 17697 34693 17700
rect 34727 17697 34739 17731
rect 34681 17691 34739 17697
rect 11330 17660 11336 17672
rect 11291 17632 11336 17660
rect 11330 17620 11336 17632
rect 11388 17620 11394 17672
rect 21450 17660 21456 17672
rect 21411 17632 21456 17660
rect 21450 17620 21456 17632
rect 21508 17620 21514 17672
rect 23937 17663 23995 17669
rect 23937 17629 23949 17663
rect 23983 17629 23995 17663
rect 23937 17623 23995 17629
rect 8018 17524 8024 17536
rect 7979 17496 8024 17524
rect 8018 17484 8024 17496
rect 8076 17484 8082 17536
rect 10870 17524 10876 17536
rect 10831 17496 10876 17524
rect 10870 17484 10876 17496
rect 10928 17484 10934 17536
rect 12713 17527 12771 17533
rect 12713 17493 12725 17527
rect 12759 17524 12771 17527
rect 12802 17524 12808 17536
rect 12759 17496 12808 17524
rect 12759 17493 12771 17496
rect 12713 17487 12771 17493
rect 12802 17484 12808 17496
rect 12860 17484 12866 17536
rect 13262 17524 13268 17536
rect 13223 17496 13268 17524
rect 13262 17484 13268 17496
rect 13320 17484 13326 17536
rect 18874 17524 18880 17536
rect 18835 17496 18880 17524
rect 18874 17484 18880 17496
rect 18932 17484 18938 17536
rect 22833 17527 22891 17533
rect 22833 17493 22845 17527
rect 22879 17524 22891 17527
rect 23661 17527 23719 17533
rect 23661 17524 23673 17527
rect 22879 17496 23673 17524
rect 22879 17493 22891 17496
rect 22833 17487 22891 17493
rect 23661 17493 23673 17496
rect 23707 17524 23719 17527
rect 23750 17524 23756 17536
rect 23707 17496 23756 17524
rect 23707 17493 23719 17496
rect 23661 17487 23719 17493
rect 23750 17484 23756 17496
rect 23808 17484 23814 17536
rect 23952 17524 23980 17623
rect 28074 17620 28080 17672
rect 28132 17660 28138 17672
rect 28169 17663 28227 17669
rect 28169 17660 28181 17663
rect 28132 17632 28181 17660
rect 28132 17620 28138 17632
rect 28169 17629 28181 17632
rect 28215 17629 28227 17663
rect 33318 17660 33324 17672
rect 33279 17632 33324 17660
rect 28169 17623 28227 17629
rect 33318 17620 33324 17632
rect 33376 17620 33382 17672
rect 33413 17663 33471 17669
rect 33413 17629 33425 17663
rect 33459 17629 33471 17663
rect 33413 17623 33471 17629
rect 32769 17595 32827 17601
rect 32769 17561 32781 17595
rect 32815 17592 32827 17595
rect 33428 17592 33456 17623
rect 34330 17620 34336 17672
rect 34388 17660 34394 17672
rect 34425 17663 34483 17669
rect 34425 17660 34437 17663
rect 34388 17632 34437 17660
rect 34388 17620 34394 17632
rect 34425 17629 34437 17632
rect 34471 17629 34483 17663
rect 34425 17623 34483 17629
rect 34054 17592 34060 17604
rect 32815 17564 34060 17592
rect 32815 17561 32827 17564
rect 32769 17555 32827 17561
rect 34054 17552 34060 17564
rect 34112 17552 34118 17604
rect 24302 17524 24308 17536
rect 23952 17496 24308 17524
rect 24302 17484 24308 17496
rect 24360 17484 24366 17536
rect 25314 17524 25320 17536
rect 25275 17496 25320 17524
rect 25314 17484 25320 17496
rect 25372 17484 25378 17536
rect 27709 17527 27767 17533
rect 27709 17493 27721 17527
rect 27755 17524 27767 17527
rect 27982 17524 27988 17536
rect 27755 17496 27988 17524
rect 27755 17493 27767 17496
rect 27709 17487 27767 17493
rect 27982 17484 27988 17496
rect 28040 17524 28046 17536
rect 28902 17524 28908 17536
rect 28040 17496 28908 17524
rect 28040 17484 28046 17496
rect 28902 17484 28908 17496
rect 28960 17484 28966 17536
rect 30374 17484 30380 17536
rect 30432 17524 30438 17536
rect 31846 17524 31852 17536
rect 30432 17496 31852 17524
rect 30432 17484 30438 17496
rect 31846 17484 31852 17496
rect 31904 17484 31910 17536
rect 32858 17524 32864 17536
rect 32819 17496 32864 17524
rect 32858 17484 32864 17496
rect 32916 17484 32922 17536
rect 1104 17434 38824 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 34966 17434
rect 35018 17382 35030 17434
rect 35082 17382 35094 17434
rect 35146 17382 35158 17434
rect 35210 17382 38824 17434
rect 1104 17360 38824 17382
rect 11330 17280 11336 17332
rect 11388 17320 11394 17332
rect 11793 17323 11851 17329
rect 11793 17320 11805 17323
rect 11388 17292 11805 17320
rect 11388 17280 11394 17292
rect 11793 17289 11805 17292
rect 11839 17320 11851 17323
rect 11882 17320 11888 17332
rect 11839 17292 11888 17320
rect 11839 17289 11851 17292
rect 11793 17283 11851 17289
rect 11882 17280 11888 17292
rect 11940 17280 11946 17332
rect 22646 17320 22652 17332
rect 22607 17292 22652 17320
rect 22646 17280 22652 17292
rect 22704 17280 22710 17332
rect 23106 17320 23112 17332
rect 23067 17292 23112 17320
rect 23106 17280 23112 17292
rect 23164 17320 23170 17332
rect 24578 17320 24584 17332
rect 23164 17292 24584 17320
rect 23164 17280 23170 17292
rect 24578 17280 24584 17292
rect 24636 17320 24642 17332
rect 25041 17323 25099 17329
rect 25041 17320 25053 17323
rect 24636 17292 25053 17320
rect 24636 17280 24642 17292
rect 25041 17289 25053 17292
rect 25087 17289 25099 17323
rect 25041 17283 25099 17289
rect 30926 17280 30932 17332
rect 30984 17320 30990 17332
rect 31205 17323 31263 17329
rect 31205 17320 31217 17323
rect 30984 17292 31217 17320
rect 30984 17280 30990 17292
rect 31205 17289 31217 17292
rect 31251 17320 31263 17323
rect 31757 17323 31815 17329
rect 31757 17320 31769 17323
rect 31251 17292 31769 17320
rect 31251 17289 31263 17292
rect 31205 17283 31263 17289
rect 31757 17289 31769 17292
rect 31803 17289 31815 17323
rect 31757 17283 31815 17289
rect 32953 17323 33011 17329
rect 32953 17289 32965 17323
rect 32999 17320 33011 17323
rect 33318 17320 33324 17332
rect 32999 17292 33324 17320
rect 32999 17289 33011 17292
rect 32953 17283 33011 17289
rect 27525 17255 27583 17261
rect 27525 17221 27537 17255
rect 27571 17252 27583 17255
rect 28166 17252 28172 17264
rect 27571 17224 28172 17252
rect 27571 17221 27583 17224
rect 27525 17215 27583 17221
rect 28166 17212 28172 17224
rect 28224 17212 28230 17264
rect 10870 17144 10876 17196
rect 10928 17184 10934 17196
rect 11425 17187 11483 17193
rect 11425 17184 11437 17187
rect 10928 17156 11437 17184
rect 10928 17144 10934 17156
rect 11425 17153 11437 17156
rect 11471 17184 11483 17187
rect 13081 17187 13139 17193
rect 13081 17184 13093 17187
rect 11471 17156 13093 17184
rect 11471 17153 11483 17156
rect 11425 17147 11483 17153
rect 13081 17153 13093 17156
rect 13127 17184 13139 17187
rect 13262 17184 13268 17196
rect 13127 17156 13268 17184
rect 13127 17153 13139 17156
rect 13081 17147 13139 17153
rect 13262 17144 13268 17156
rect 13320 17144 13326 17196
rect 27157 17187 27215 17193
rect 27157 17153 27169 17187
rect 27203 17184 27215 17187
rect 28258 17184 28264 17196
rect 27203 17156 28264 17184
rect 27203 17153 27215 17156
rect 27157 17147 27215 17153
rect 28258 17144 28264 17156
rect 28316 17144 28322 17196
rect 31846 17144 31852 17196
rect 31904 17184 31910 17196
rect 32401 17187 32459 17193
rect 32401 17184 32413 17187
rect 31904 17156 32413 17184
rect 31904 17144 31910 17156
rect 32401 17153 32413 17156
rect 32447 17184 32459 17187
rect 32766 17184 32772 17196
rect 32447 17156 32772 17184
rect 32447 17153 32459 17156
rect 32401 17147 32459 17153
rect 32766 17144 32772 17156
rect 32824 17144 32830 17196
rect 7929 17119 7987 17125
rect 7929 17116 7941 17119
rect 7760 17088 7941 17116
rect 7098 16940 7104 16992
rect 7156 16980 7162 16992
rect 7760 16989 7788 17088
rect 7929 17085 7941 17088
rect 7975 17085 7987 17119
rect 7929 17079 7987 17085
rect 8018 17076 8024 17128
rect 8076 17116 8082 17128
rect 8185 17119 8243 17125
rect 8185 17116 8197 17119
rect 8076 17088 8197 17116
rect 8076 17076 8082 17088
rect 8185 17085 8197 17088
rect 8231 17085 8243 17119
rect 8185 17079 8243 17085
rect 10689 17119 10747 17125
rect 10689 17085 10701 17119
rect 10735 17116 10747 17119
rect 11241 17119 11299 17125
rect 11241 17116 11253 17119
rect 10735 17088 11253 17116
rect 10735 17085 10747 17088
rect 10689 17079 10747 17085
rect 11241 17085 11253 17088
rect 11287 17116 11299 17119
rect 11514 17116 11520 17128
rect 11287 17088 11520 17116
rect 11287 17085 11299 17088
rect 11241 17079 11299 17085
rect 11514 17076 11520 17088
rect 11572 17076 11578 17128
rect 11606 17076 11612 17128
rect 11664 17116 11670 17128
rect 12253 17119 12311 17125
rect 12253 17116 12265 17119
rect 11664 17088 12265 17116
rect 11664 17076 11670 17088
rect 12253 17085 12265 17088
rect 12299 17116 12311 17119
rect 12897 17119 12955 17125
rect 12897 17116 12909 17119
rect 12299 17088 12909 17116
rect 12299 17085 12311 17088
rect 12253 17079 12311 17085
rect 12897 17085 12909 17088
rect 12943 17116 12955 17119
rect 13538 17116 13544 17128
rect 12943 17088 13544 17116
rect 12943 17085 12955 17088
rect 12897 17079 12955 17085
rect 13538 17076 13544 17088
rect 13596 17076 13602 17128
rect 20625 17119 20683 17125
rect 20625 17085 20637 17119
rect 20671 17116 20683 17119
rect 20717 17119 20775 17125
rect 20717 17116 20729 17119
rect 20671 17088 20729 17116
rect 20671 17085 20683 17088
rect 20625 17079 20683 17085
rect 20717 17085 20729 17088
rect 20763 17116 20775 17119
rect 21450 17116 21456 17128
rect 20763 17088 21456 17116
rect 20763 17085 20775 17088
rect 20717 17079 20775 17085
rect 21450 17076 21456 17088
rect 21508 17076 21514 17128
rect 23477 17119 23535 17125
rect 23477 17085 23489 17119
rect 23523 17116 23535 17119
rect 23661 17119 23719 17125
rect 23661 17116 23673 17119
rect 23523 17088 23673 17116
rect 23523 17085 23535 17088
rect 23477 17079 23535 17085
rect 23661 17085 23673 17088
rect 23707 17085 23719 17119
rect 23661 17079 23719 17085
rect 20254 17048 20260 17060
rect 20167 17020 20260 17048
rect 20254 17008 20260 17020
rect 20312 17048 20318 17060
rect 20984 17051 21042 17057
rect 20984 17048 20996 17051
rect 20312 17020 20996 17048
rect 20312 17008 20318 17020
rect 20984 17017 20996 17020
rect 21030 17048 21042 17051
rect 22186 17048 22192 17060
rect 21030 17020 22192 17048
rect 21030 17017 21042 17020
rect 20984 17011 21042 17017
rect 22186 17008 22192 17020
rect 22244 17008 22250 17060
rect 23676 17048 23704 17079
rect 23750 17076 23756 17128
rect 23808 17116 23814 17128
rect 23917 17119 23975 17125
rect 23917 17116 23929 17119
rect 23808 17088 23929 17116
rect 23808 17076 23814 17088
rect 23917 17085 23929 17088
rect 23963 17085 23975 17119
rect 27982 17116 27988 17128
rect 27943 17088 27988 17116
rect 23917 17079 23975 17085
rect 27982 17076 27988 17088
rect 28040 17076 28046 17128
rect 28077 17119 28135 17125
rect 28077 17085 28089 17119
rect 28123 17116 28135 17119
rect 28166 17116 28172 17128
rect 28123 17088 28172 17116
rect 28123 17085 28135 17088
rect 28077 17079 28135 17085
rect 28166 17076 28172 17088
rect 28224 17076 28230 17128
rect 29546 17125 29552 17128
rect 28905 17119 28963 17125
rect 28905 17085 28917 17119
rect 28951 17116 28963 17119
rect 29273 17119 29331 17125
rect 29273 17116 29285 17119
rect 28951 17088 29285 17116
rect 28951 17085 28963 17088
rect 28905 17079 28963 17085
rect 29273 17085 29285 17088
rect 29319 17085 29331 17119
rect 29540 17116 29552 17125
rect 29507 17088 29552 17116
rect 29273 17079 29331 17085
rect 29540 17079 29552 17088
rect 29546 17076 29552 17079
rect 29604 17076 29610 17128
rect 31110 17076 31116 17128
rect 31168 17116 31174 17128
rect 32968 17116 32996 17283
rect 33318 17280 33324 17292
rect 33376 17280 33382 17332
rect 33594 17320 33600 17332
rect 33555 17292 33600 17320
rect 33594 17280 33600 17292
rect 33652 17280 33658 17332
rect 33873 17323 33931 17329
rect 33873 17289 33885 17323
rect 33919 17320 33931 17323
rect 34422 17320 34428 17332
rect 33919 17292 34428 17320
rect 33919 17289 33931 17292
rect 33873 17283 33931 17289
rect 34422 17280 34428 17292
rect 34480 17280 34486 17332
rect 37090 17320 37096 17332
rect 37051 17292 37096 17320
rect 37090 17280 37096 17292
rect 37148 17280 37154 17332
rect 34330 17144 34336 17196
rect 34388 17184 34394 17196
rect 34425 17187 34483 17193
rect 34425 17184 34437 17187
rect 34388 17156 34437 17184
rect 34388 17144 34394 17156
rect 34425 17153 34437 17156
rect 34471 17153 34483 17187
rect 34425 17147 34483 17153
rect 34606 17144 34612 17196
rect 34664 17184 34670 17196
rect 35437 17187 35495 17193
rect 35437 17184 35449 17187
rect 34664 17156 35449 17184
rect 34664 17144 34670 17156
rect 35437 17153 35449 17156
rect 35483 17184 35495 17187
rect 35618 17184 35624 17196
rect 35483 17156 35624 17184
rect 35483 17153 35495 17156
rect 35437 17147 35495 17153
rect 35618 17144 35624 17156
rect 35676 17144 35682 17196
rect 31168 17088 32996 17116
rect 33689 17119 33747 17125
rect 31168 17076 31174 17088
rect 33689 17085 33701 17119
rect 33735 17116 33747 17119
rect 33778 17116 33784 17128
rect 33735 17088 33784 17116
rect 33735 17085 33747 17088
rect 33689 17079 33747 17085
rect 33778 17076 33784 17088
rect 33836 17116 33842 17128
rect 33836 17088 34928 17116
rect 33836 17076 33842 17088
rect 24486 17048 24492 17060
rect 23676 17020 24492 17048
rect 24486 17008 24492 17020
rect 24544 17008 24550 17060
rect 31573 17051 31631 17057
rect 31573 17048 31585 17051
rect 27632 17020 31585 17048
rect 7745 16983 7803 16989
rect 7745 16980 7757 16983
rect 7156 16952 7757 16980
rect 7156 16940 7162 16952
rect 7745 16949 7757 16952
rect 7791 16949 7803 16983
rect 7745 16943 7803 16949
rect 8294 16940 8300 16992
rect 8352 16980 8358 16992
rect 9309 16983 9367 16989
rect 9309 16980 9321 16983
rect 8352 16952 9321 16980
rect 8352 16940 8358 16952
rect 9309 16949 9321 16952
rect 9355 16949 9367 16983
rect 9309 16943 9367 16949
rect 10686 16940 10692 16992
rect 10744 16980 10750 16992
rect 10781 16983 10839 16989
rect 10781 16980 10793 16983
rect 10744 16952 10793 16980
rect 10744 16940 10750 16952
rect 10781 16949 10793 16952
rect 10827 16949 10839 16983
rect 11146 16980 11152 16992
rect 11107 16952 11152 16980
rect 10781 16943 10839 16949
rect 11146 16940 11152 16952
rect 11204 16940 11210 16992
rect 12434 16980 12440 16992
rect 12395 16952 12440 16980
rect 12434 16940 12440 16952
rect 12492 16940 12498 16992
rect 12802 16980 12808 16992
rect 12763 16952 12808 16980
rect 12802 16940 12808 16952
rect 12860 16940 12866 16992
rect 22094 16940 22100 16992
rect 22152 16980 22158 16992
rect 27632 16989 27660 17020
rect 31573 17017 31585 17020
rect 31619 17048 31631 17051
rect 32217 17051 32275 17057
rect 32217 17048 32229 17051
rect 31619 17020 32229 17048
rect 31619 17017 31631 17020
rect 31573 17011 31631 17017
rect 32217 17017 32229 17020
rect 32263 17017 32275 17051
rect 32217 17011 32275 17017
rect 27617 16983 27675 16989
rect 22152 16952 22197 16980
rect 22152 16940 22158 16952
rect 27617 16949 27629 16983
rect 27663 16949 27675 16983
rect 27617 16943 27675 16949
rect 28074 16940 28080 16992
rect 28132 16980 28138 16992
rect 28350 16980 28356 16992
rect 28132 16952 28356 16980
rect 28132 16940 28138 16952
rect 28350 16940 28356 16952
rect 28408 16980 28414 16992
rect 28629 16983 28687 16989
rect 28629 16980 28641 16983
rect 28408 16952 28641 16980
rect 28408 16940 28414 16952
rect 28629 16949 28641 16952
rect 28675 16980 28687 16983
rect 28905 16983 28963 16989
rect 28905 16980 28917 16983
rect 28675 16952 28917 16980
rect 28675 16949 28687 16952
rect 28629 16943 28687 16949
rect 28905 16949 28917 16952
rect 28951 16980 28963 16983
rect 28997 16983 29055 16989
rect 28997 16980 29009 16983
rect 28951 16952 29009 16980
rect 28951 16949 28963 16952
rect 28905 16943 28963 16949
rect 28997 16949 29009 16952
rect 29043 16949 29055 16983
rect 30650 16980 30656 16992
rect 30611 16952 30656 16980
rect 28997 16943 29055 16949
rect 30650 16940 30656 16952
rect 30708 16940 30714 16992
rect 32122 16980 32128 16992
rect 32083 16952 32128 16980
rect 32122 16940 32128 16952
rect 32180 16940 32186 16992
rect 34900 16989 34928 17088
rect 34974 17076 34980 17128
rect 35032 17116 35038 17128
rect 35253 17119 35311 17125
rect 35253 17116 35265 17119
rect 35032 17088 35265 17116
rect 35032 17076 35038 17088
rect 35253 17085 35265 17088
rect 35299 17116 35311 17119
rect 35897 17119 35955 17125
rect 35897 17116 35909 17119
rect 35299 17088 35909 17116
rect 35299 17085 35311 17088
rect 35253 17079 35311 17085
rect 35897 17085 35909 17088
rect 35943 17085 35955 17119
rect 35897 17079 35955 17085
rect 36449 17119 36507 17125
rect 36449 17085 36461 17119
rect 36495 17116 36507 17119
rect 37090 17116 37096 17128
rect 36495 17088 37096 17116
rect 36495 17085 36507 17088
rect 36449 17079 36507 17085
rect 37090 17076 37096 17088
rect 37148 17076 37154 17128
rect 34885 16983 34943 16989
rect 34885 16949 34897 16983
rect 34931 16949 34943 16983
rect 35342 16980 35348 16992
rect 35303 16952 35348 16980
rect 34885 16943 34943 16949
rect 35342 16940 35348 16952
rect 35400 16940 35406 16992
rect 36446 16940 36452 16992
rect 36504 16980 36510 16992
rect 36633 16983 36691 16989
rect 36633 16980 36645 16983
rect 36504 16952 36645 16980
rect 36504 16940 36510 16952
rect 36633 16949 36645 16952
rect 36679 16949 36691 16983
rect 36633 16943 36691 16949
rect 1104 16890 38824 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 38824 16890
rect 1104 16816 38824 16838
rect 7285 16779 7343 16785
rect 7285 16745 7297 16779
rect 7331 16776 7343 16779
rect 7466 16776 7472 16788
rect 7331 16748 7472 16776
rect 7331 16745 7343 16748
rect 7285 16739 7343 16745
rect 7466 16736 7472 16748
rect 7524 16776 7530 16788
rect 8294 16776 8300 16788
rect 7524 16748 8300 16776
rect 7524 16736 7530 16748
rect 8294 16736 8300 16748
rect 8352 16736 8358 16788
rect 11606 16736 11612 16788
rect 11664 16776 11670 16788
rect 12713 16779 12771 16785
rect 12713 16776 12725 16779
rect 11664 16748 12725 16776
rect 11664 16736 11670 16748
rect 12713 16745 12725 16748
rect 12759 16745 12771 16779
rect 12713 16739 12771 16745
rect 22646 16736 22652 16788
rect 22704 16776 22710 16788
rect 23109 16779 23167 16785
rect 23109 16776 23121 16779
rect 22704 16748 23121 16776
rect 22704 16736 22710 16748
rect 23109 16745 23121 16748
rect 23155 16745 23167 16779
rect 23109 16739 23167 16745
rect 7760 16680 7972 16708
rect 7760 16652 7788 16680
rect 7742 16640 7748 16652
rect 7703 16612 7748 16640
rect 7742 16600 7748 16612
rect 7800 16600 7806 16652
rect 7944 16640 7972 16680
rect 8018 16668 8024 16720
rect 8076 16708 8082 16720
rect 9401 16711 9459 16717
rect 9401 16708 9413 16711
rect 8076 16680 9413 16708
rect 8076 16668 8082 16680
rect 9401 16677 9413 16680
rect 9447 16708 9459 16711
rect 10045 16711 10103 16717
rect 10045 16708 10057 16711
rect 9447 16680 10057 16708
rect 9447 16677 9459 16680
rect 9401 16671 9459 16677
rect 10045 16677 10057 16680
rect 10091 16677 10103 16711
rect 10045 16671 10103 16677
rect 10873 16711 10931 16717
rect 10873 16677 10885 16711
rect 10919 16708 10931 16711
rect 11146 16708 11152 16720
rect 10919 16680 11152 16708
rect 10919 16677 10931 16680
rect 10873 16671 10931 16677
rect 8202 16640 8208 16652
rect 7944 16612 8064 16640
rect 8163 16612 8208 16640
rect 8036 16572 8064 16612
rect 8202 16600 8208 16612
rect 8260 16600 8266 16652
rect 10060 16640 10088 16671
rect 11146 16668 11152 16680
rect 11204 16708 11210 16720
rect 12526 16708 12532 16720
rect 11204 16680 12532 16708
rect 11204 16668 11210 16680
rect 12526 16668 12532 16680
rect 12584 16668 12590 16720
rect 21996 16711 22054 16717
rect 21996 16677 22008 16711
rect 22042 16708 22054 16711
rect 22094 16708 22100 16720
rect 22042 16680 22100 16708
rect 22042 16677 22054 16680
rect 21996 16671 22054 16677
rect 22094 16668 22100 16680
rect 22152 16668 22158 16720
rect 23124 16708 23152 16739
rect 23474 16736 23480 16788
rect 23532 16776 23538 16788
rect 24213 16779 24271 16785
rect 24213 16776 24225 16779
rect 23532 16748 24225 16776
rect 23532 16736 23538 16748
rect 24213 16745 24225 16748
rect 24259 16745 24271 16779
rect 24213 16739 24271 16745
rect 28261 16779 28319 16785
rect 28261 16745 28273 16779
rect 28307 16776 28319 16779
rect 29730 16776 29736 16788
rect 28307 16748 29736 16776
rect 28307 16745 28319 16748
rect 28261 16739 28319 16745
rect 29730 16736 29736 16748
rect 29788 16736 29794 16788
rect 30374 16776 30380 16788
rect 30335 16748 30380 16776
rect 30374 16736 30380 16748
rect 30432 16736 30438 16788
rect 31110 16776 31116 16788
rect 31071 16748 31116 16776
rect 31110 16736 31116 16748
rect 31168 16736 31174 16788
rect 31849 16779 31907 16785
rect 31849 16745 31861 16779
rect 31895 16776 31907 16779
rect 32122 16776 32128 16788
rect 31895 16748 32128 16776
rect 31895 16745 31907 16748
rect 31849 16739 31907 16745
rect 32122 16736 32128 16748
rect 32180 16736 32186 16788
rect 33134 16776 33140 16788
rect 33095 16748 33140 16776
rect 33134 16736 33140 16748
rect 33192 16736 33198 16788
rect 33778 16776 33784 16788
rect 33739 16748 33784 16776
rect 33778 16736 33784 16748
rect 33836 16736 33842 16788
rect 33962 16736 33968 16788
rect 34020 16776 34026 16788
rect 34241 16779 34299 16785
rect 34241 16776 34253 16779
rect 34020 16748 34253 16776
rect 34020 16736 34026 16748
rect 34241 16745 34253 16748
rect 34287 16776 34299 16779
rect 35342 16776 35348 16788
rect 34287 16748 35348 16776
rect 34287 16745 34299 16748
rect 34241 16739 34299 16745
rect 35342 16736 35348 16748
rect 35400 16736 35406 16788
rect 35618 16776 35624 16788
rect 35579 16748 35624 16776
rect 35618 16736 35624 16748
rect 35676 16736 35682 16788
rect 23658 16708 23664 16720
rect 23124 16680 23664 16708
rect 23658 16668 23664 16680
rect 23716 16668 23722 16720
rect 23750 16668 23756 16720
rect 23808 16708 23814 16720
rect 24302 16708 24308 16720
rect 23808 16680 24308 16708
rect 23808 16668 23814 16680
rect 24302 16668 24308 16680
rect 24360 16708 24366 16720
rect 24581 16711 24639 16717
rect 24581 16708 24593 16711
rect 24360 16680 24593 16708
rect 24360 16668 24366 16680
rect 24581 16677 24593 16680
rect 24627 16677 24639 16711
rect 24581 16671 24639 16677
rect 31754 16668 31760 16720
rect 31812 16708 31818 16720
rect 32214 16708 32220 16720
rect 31812 16680 32220 16708
rect 31812 16668 31818 16680
rect 32214 16668 32220 16680
rect 32272 16708 32278 16720
rect 32585 16711 32643 16717
rect 32585 16708 32597 16711
rect 32272 16680 32597 16708
rect 32272 16668 32278 16680
rect 32585 16677 32597 16680
rect 32631 16677 32643 16711
rect 34054 16708 34060 16720
rect 34015 16680 34060 16708
rect 32585 16671 32643 16677
rect 34054 16668 34060 16680
rect 34112 16708 34118 16720
rect 34112 16680 34836 16708
rect 34112 16668 34118 16680
rect 10060 16612 11100 16640
rect 8481 16575 8539 16581
rect 8481 16572 8493 16575
rect 8036 16544 8493 16572
rect 8481 16541 8493 16544
rect 8527 16541 8539 16575
rect 10134 16572 10140 16584
rect 10095 16544 10140 16572
rect 8481 16535 8539 16541
rect 8496 16504 8524 16535
rect 10134 16532 10140 16544
rect 10192 16532 10198 16584
rect 10321 16575 10379 16581
rect 10321 16541 10333 16575
rect 10367 16572 10379 16575
rect 10870 16572 10876 16584
rect 10367 16544 10876 16572
rect 10367 16541 10379 16544
rect 10321 16535 10379 16541
rect 9122 16504 9128 16516
rect 8496 16476 9128 16504
rect 9122 16464 9128 16476
rect 9180 16504 9186 16516
rect 10336 16504 10364 16535
rect 10870 16532 10876 16544
rect 10928 16532 10934 16584
rect 11072 16572 11100 16612
rect 11238 16600 11244 16652
rect 11296 16640 11302 16652
rect 11589 16643 11647 16649
rect 11589 16640 11601 16643
rect 11296 16612 11601 16640
rect 11296 16600 11302 16612
rect 11589 16609 11601 16612
rect 11635 16640 11647 16643
rect 12802 16640 12808 16652
rect 11635 16612 12808 16640
rect 11635 16609 11647 16612
rect 11589 16603 11647 16609
rect 12802 16600 12808 16612
rect 12860 16640 12866 16652
rect 13265 16643 13323 16649
rect 13265 16640 13277 16643
rect 12860 16612 13277 16640
rect 12860 16600 12866 16612
rect 13265 16609 13277 16612
rect 13311 16609 13323 16643
rect 23676 16640 23704 16668
rect 24673 16643 24731 16649
rect 24673 16640 24685 16643
rect 23676 16612 24685 16640
rect 13265 16603 13323 16609
rect 24673 16609 24685 16612
rect 24719 16609 24731 16643
rect 24673 16603 24731 16609
rect 24854 16600 24860 16652
rect 24912 16640 24918 16652
rect 25225 16643 25283 16649
rect 25225 16640 25237 16643
rect 24912 16612 25237 16640
rect 24912 16600 24918 16612
rect 25225 16609 25237 16612
rect 25271 16640 25283 16643
rect 25314 16640 25320 16652
rect 25271 16612 25320 16640
rect 25271 16609 25283 16612
rect 25225 16603 25283 16609
rect 25314 16600 25320 16612
rect 25372 16600 25378 16652
rect 26510 16640 26516 16652
rect 26471 16612 26516 16640
rect 26510 16600 26516 16612
rect 26568 16640 26574 16652
rect 28626 16649 28632 16652
rect 27065 16643 27123 16649
rect 27065 16640 27077 16643
rect 26568 16612 27077 16640
rect 26568 16600 26574 16612
rect 27065 16609 27077 16612
rect 27111 16609 27123 16643
rect 27065 16603 27123 16609
rect 28620 16603 28632 16649
rect 28684 16640 28690 16652
rect 30926 16640 30932 16652
rect 28684 16612 28720 16640
rect 30887 16612 30932 16640
rect 28626 16600 28632 16603
rect 28684 16600 28690 16612
rect 30926 16600 30932 16612
rect 30984 16600 30990 16652
rect 31846 16600 31852 16652
rect 31904 16640 31910 16652
rect 32306 16640 32312 16652
rect 31904 16612 32312 16640
rect 31904 16600 31910 16612
rect 32306 16600 32312 16612
rect 32364 16640 32370 16652
rect 32493 16643 32551 16649
rect 32493 16640 32505 16643
rect 32364 16612 32505 16640
rect 32364 16600 32370 16612
rect 32493 16609 32505 16612
rect 32539 16609 32551 16643
rect 32493 16603 32551 16609
rect 32766 16600 32772 16652
rect 32824 16640 32830 16652
rect 34606 16640 34612 16652
rect 32824 16612 33088 16640
rect 34567 16612 34612 16640
rect 32824 16600 32830 16612
rect 11146 16572 11152 16584
rect 11072 16544 11152 16572
rect 11146 16532 11152 16544
rect 11204 16532 11210 16584
rect 11330 16572 11336 16584
rect 11291 16544 11336 16572
rect 11330 16532 11336 16544
rect 11388 16532 11394 16584
rect 21729 16575 21787 16581
rect 21729 16572 21741 16575
rect 21468 16544 21741 16572
rect 9180 16476 10364 16504
rect 9180 16464 9186 16476
rect 21468 16448 21496 16544
rect 21729 16541 21741 16544
rect 21775 16541 21787 16575
rect 21729 16535 21787 16541
rect 24210 16532 24216 16584
rect 24268 16572 24274 16584
rect 24765 16575 24823 16581
rect 24765 16572 24777 16575
rect 24268 16544 24777 16572
rect 24268 16532 24274 16544
rect 24765 16541 24777 16544
rect 24811 16572 24823 16575
rect 27433 16575 27491 16581
rect 27433 16572 27445 16575
rect 24811 16544 27445 16572
rect 24811 16541 24823 16544
rect 24765 16535 24823 16541
rect 27433 16541 27445 16544
rect 27479 16572 27491 16575
rect 27522 16572 27528 16584
rect 27479 16544 27528 16572
rect 27479 16541 27491 16544
rect 27433 16535 27491 16541
rect 27522 16532 27528 16544
rect 27580 16532 27586 16584
rect 28350 16572 28356 16584
rect 28311 16544 28356 16572
rect 28350 16532 28356 16544
rect 28408 16532 28414 16584
rect 32677 16575 32735 16581
rect 32677 16541 32689 16575
rect 32723 16572 32735 16575
rect 32858 16572 32864 16584
rect 32723 16544 32864 16572
rect 32723 16541 32735 16544
rect 32677 16535 32735 16541
rect 32858 16532 32864 16544
rect 32916 16532 32922 16584
rect 33060 16572 33088 16612
rect 34606 16600 34612 16612
rect 34664 16600 34670 16652
rect 33870 16572 33876 16584
rect 33060 16544 33876 16572
rect 33870 16532 33876 16544
rect 33928 16532 33934 16584
rect 34330 16532 34336 16584
rect 34388 16572 34394 16584
rect 34808 16581 34836 16680
rect 35802 16640 35808 16652
rect 35763 16612 35808 16640
rect 35802 16600 35808 16612
rect 35860 16600 35866 16652
rect 34701 16575 34759 16581
rect 34701 16572 34713 16575
rect 34388 16544 34713 16572
rect 34388 16532 34394 16544
rect 34701 16541 34713 16544
rect 34747 16541 34759 16575
rect 34701 16535 34759 16541
rect 34793 16575 34851 16581
rect 34793 16541 34805 16575
rect 34839 16572 34851 16575
rect 35618 16572 35624 16584
rect 34839 16544 35624 16572
rect 34839 16541 34851 16544
rect 34793 16535 34851 16541
rect 35618 16532 35624 16544
rect 35676 16532 35682 16584
rect 24029 16507 24087 16513
rect 24029 16473 24041 16507
rect 24075 16504 24087 16507
rect 24486 16504 24492 16516
rect 24075 16476 24492 16504
rect 24075 16473 24087 16476
rect 24029 16467 24087 16473
rect 24486 16464 24492 16476
rect 24544 16464 24550 16516
rect 7834 16436 7840 16448
rect 7795 16408 7840 16436
rect 7834 16396 7840 16408
rect 7892 16396 7898 16448
rect 9674 16436 9680 16448
rect 9635 16408 9680 16436
rect 9674 16396 9680 16408
rect 9732 16396 9738 16448
rect 21450 16436 21456 16448
rect 21411 16408 21456 16436
rect 21450 16396 21456 16408
rect 21508 16396 21514 16448
rect 26694 16436 26700 16448
rect 26655 16408 26700 16436
rect 26694 16396 26700 16408
rect 26752 16396 26758 16448
rect 35989 16439 36047 16445
rect 35989 16405 36001 16439
rect 36035 16436 36047 16439
rect 36170 16436 36176 16448
rect 36035 16408 36176 16436
rect 36035 16405 36047 16408
rect 35989 16399 36047 16405
rect 36170 16396 36176 16408
rect 36228 16396 36234 16448
rect 1104 16346 38824 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 34966 16346
rect 35018 16294 35030 16346
rect 35082 16294 35094 16346
rect 35146 16294 35158 16346
rect 35210 16294 38824 16346
rect 1104 16272 38824 16294
rect 7098 16232 7104 16244
rect 7059 16204 7104 16232
rect 7098 16192 7104 16204
rect 7156 16192 7162 16244
rect 11146 16232 11152 16244
rect 11107 16204 11152 16232
rect 11146 16192 11152 16204
rect 11204 16192 11210 16244
rect 23658 16192 23664 16244
rect 23716 16232 23722 16244
rect 23937 16235 23995 16241
rect 23937 16232 23949 16235
rect 23716 16204 23949 16232
rect 23716 16192 23722 16204
rect 23937 16201 23949 16204
rect 23983 16201 23995 16235
rect 23937 16195 23995 16201
rect 24762 16192 24768 16244
rect 24820 16232 24826 16244
rect 24820 16204 25912 16232
rect 24820 16192 24826 16204
rect 7116 16096 7144 16192
rect 25884 16173 25912 16204
rect 28626 16192 28632 16244
rect 28684 16232 28690 16244
rect 28721 16235 28779 16241
rect 28721 16232 28733 16235
rect 28684 16204 28733 16232
rect 28684 16192 28690 16204
rect 28721 16201 28733 16204
rect 28767 16201 28779 16235
rect 28721 16195 28779 16201
rect 29270 16192 29276 16244
rect 29328 16232 29334 16244
rect 29549 16235 29607 16241
rect 29549 16232 29561 16235
rect 29328 16204 29561 16232
rect 29328 16192 29334 16204
rect 29549 16201 29561 16204
rect 29595 16201 29607 16235
rect 31846 16232 31852 16244
rect 31807 16204 31852 16232
rect 29549 16195 29607 16201
rect 25869 16167 25927 16173
rect 25869 16133 25881 16167
rect 25915 16164 25927 16167
rect 25915 16136 26924 16164
rect 25915 16133 25927 16136
rect 25869 16127 25927 16133
rect 7193 16099 7251 16105
rect 7193 16096 7205 16099
rect 7116 16068 7205 16096
rect 7193 16065 7205 16068
rect 7239 16065 7251 16099
rect 7193 16059 7251 16065
rect 22186 16056 22192 16108
rect 22244 16096 22250 16108
rect 22465 16099 22523 16105
rect 22465 16096 22477 16099
rect 22244 16068 22477 16096
rect 22244 16056 22250 16068
rect 22465 16065 22477 16068
rect 22511 16065 22523 16099
rect 22465 16059 22523 16065
rect 22649 16099 22707 16105
rect 22649 16065 22661 16099
rect 22695 16096 22707 16099
rect 23017 16099 23075 16105
rect 23017 16096 23029 16099
rect 22695 16068 23029 16096
rect 22695 16065 22707 16068
rect 22649 16059 22707 16065
rect 23017 16065 23029 16068
rect 23063 16096 23075 16099
rect 23385 16099 23443 16105
rect 23385 16096 23397 16099
rect 23063 16068 23397 16096
rect 23063 16065 23075 16068
rect 23017 16059 23075 16065
rect 23385 16065 23397 16068
rect 23431 16096 23443 16099
rect 24210 16096 24216 16108
rect 23431 16068 24216 16096
rect 23431 16065 23443 16068
rect 23385 16059 23443 16065
rect 24210 16056 24216 16068
rect 24268 16056 24274 16108
rect 7466 16037 7472 16040
rect 7460 15991 7472 16037
rect 7524 16028 7530 16040
rect 9677 16031 9735 16037
rect 7524 16000 7560 16028
rect 7466 15988 7472 15991
rect 7524 15988 7530 16000
rect 9677 15997 9689 16031
rect 9723 16028 9735 16031
rect 9769 16031 9827 16037
rect 9769 16028 9781 16031
rect 9723 16000 9781 16028
rect 9723 15997 9735 16000
rect 9677 15991 9735 15997
rect 9769 15997 9781 16000
rect 9815 16028 9827 16031
rect 11330 16028 11336 16040
rect 9815 16000 11336 16028
rect 9815 15997 9827 16000
rect 9769 15991 9827 15997
rect 11330 15988 11336 16000
rect 11388 16028 11394 16040
rect 11701 16031 11759 16037
rect 11701 16028 11713 16031
rect 11388 16000 11713 16028
rect 11388 15988 11394 16000
rect 11701 15997 11713 16000
rect 11747 16028 11759 16031
rect 11882 16028 11888 16040
rect 11747 16000 11888 16028
rect 11747 15997 11759 16000
rect 11701 15991 11759 15997
rect 11882 15988 11888 16000
rect 11940 16028 11946 16040
rect 12161 16031 12219 16037
rect 12161 16028 12173 16031
rect 11940 16000 12173 16028
rect 11940 15988 11946 16000
rect 12161 15997 12173 16000
rect 12207 16028 12219 16031
rect 12437 16031 12495 16037
rect 12437 16028 12449 16031
rect 12207 16000 12449 16028
rect 12207 15997 12219 16000
rect 12161 15991 12219 15997
rect 12437 15997 12449 16000
rect 12483 15997 12495 16031
rect 12437 15991 12495 15997
rect 12526 15988 12532 16040
rect 12584 16028 12590 16040
rect 12693 16031 12751 16037
rect 12693 16028 12705 16031
rect 12584 16000 12705 16028
rect 12584 15988 12590 16000
rect 12693 15997 12705 16000
rect 12739 15997 12751 16031
rect 12693 15991 12751 15997
rect 21453 16031 21511 16037
rect 21453 15997 21465 16031
rect 21499 16028 21511 16031
rect 22094 16028 22100 16040
rect 21499 16000 22100 16028
rect 21499 15997 21511 16000
rect 21453 15991 21511 15997
rect 22094 15988 22100 16000
rect 22152 16028 22158 16040
rect 22373 16031 22431 16037
rect 22373 16028 22385 16031
rect 22152 16000 22385 16028
rect 22152 15988 22158 16000
rect 22373 15997 22385 16000
rect 22419 15997 22431 16031
rect 22373 15991 22431 15997
rect 24397 16031 24455 16037
rect 24397 15997 24409 16031
rect 24443 16028 24455 16031
rect 24486 16028 24492 16040
rect 24443 16000 24492 16028
rect 24443 15997 24455 16000
rect 24397 15991 24455 15997
rect 24486 15988 24492 16000
rect 24544 15988 24550 16040
rect 26896 16037 26924 16136
rect 27522 16096 27528 16108
rect 27483 16068 27528 16096
rect 27522 16056 27528 16068
rect 27580 16056 27586 16108
rect 26881 16031 26939 16037
rect 26881 15997 26893 16031
rect 26927 16028 26939 16031
rect 27433 16031 27491 16037
rect 27433 16028 27445 16031
rect 26927 16000 27445 16028
rect 26927 15997 26939 16000
rect 26881 15991 26939 15997
rect 27433 15997 27445 16000
rect 27479 15997 27491 16031
rect 29564 16028 29592 16195
rect 31846 16192 31852 16204
rect 31904 16192 31910 16244
rect 32214 16232 32220 16244
rect 32175 16204 32220 16232
rect 32214 16192 32220 16204
rect 32272 16192 32278 16244
rect 32769 16235 32827 16241
rect 32769 16201 32781 16235
rect 32815 16232 32827 16235
rect 33042 16232 33048 16244
rect 32815 16204 33048 16232
rect 32815 16201 32827 16204
rect 32769 16195 32827 16201
rect 33042 16192 33048 16204
rect 33100 16192 33106 16244
rect 33873 16235 33931 16241
rect 33873 16201 33885 16235
rect 33919 16232 33931 16235
rect 34330 16232 34336 16244
rect 33919 16204 34336 16232
rect 33919 16201 33931 16204
rect 33873 16195 33931 16201
rect 34330 16192 34336 16204
rect 34388 16192 34394 16244
rect 34606 16232 34612 16244
rect 34567 16204 34612 16232
rect 34606 16192 34612 16204
rect 34664 16192 34670 16244
rect 35618 16232 35624 16244
rect 35579 16204 35624 16232
rect 35618 16192 35624 16204
rect 35676 16192 35682 16244
rect 35894 16192 35900 16244
rect 35952 16232 35958 16244
rect 35989 16235 36047 16241
rect 35989 16232 36001 16235
rect 35952 16204 36001 16232
rect 35952 16192 35958 16204
rect 35989 16201 36001 16204
rect 36035 16201 36047 16235
rect 35989 16195 36047 16201
rect 30101 16167 30159 16173
rect 30101 16133 30113 16167
rect 30147 16164 30159 16167
rect 30926 16164 30932 16176
rect 30147 16136 30932 16164
rect 30147 16133 30159 16136
rect 30101 16127 30159 16133
rect 30926 16124 30932 16136
rect 30984 16164 30990 16176
rect 31113 16167 31171 16173
rect 31113 16164 31125 16167
rect 30984 16136 31125 16164
rect 30984 16124 30990 16136
rect 31113 16133 31125 16136
rect 31159 16133 31171 16167
rect 31113 16127 31171 16133
rect 33229 16167 33287 16173
rect 33229 16133 33241 16167
rect 33275 16164 33287 16167
rect 33962 16164 33968 16176
rect 33275 16136 33968 16164
rect 33275 16133 33287 16136
rect 33229 16127 33287 16133
rect 30374 16056 30380 16108
rect 30432 16096 30438 16108
rect 30653 16099 30711 16105
rect 30653 16096 30665 16099
rect 30432 16068 30665 16096
rect 30432 16056 30438 16068
rect 30653 16065 30665 16068
rect 30699 16065 30711 16099
rect 30653 16059 30711 16065
rect 30469 16031 30527 16037
rect 30469 16028 30481 16031
rect 29564 16000 30481 16028
rect 27433 15991 27491 15997
rect 30469 15997 30481 16000
rect 30515 15997 30527 16031
rect 30469 15991 30527 15997
rect 32585 16031 32643 16037
rect 32585 15997 32597 16031
rect 32631 16028 32643 16031
rect 33244 16028 33272 16127
rect 33962 16124 33968 16136
rect 34020 16124 34026 16176
rect 35345 16167 35403 16173
rect 35345 16133 35357 16167
rect 35391 16164 35403 16167
rect 35526 16164 35532 16176
rect 35391 16136 35532 16164
rect 35391 16133 35403 16136
rect 35345 16127 35403 16133
rect 35452 16037 35480 16136
rect 35526 16124 35532 16136
rect 35584 16124 35590 16176
rect 32631 16000 33272 16028
rect 33689 16031 33747 16037
rect 32631 15997 32643 16000
rect 32585 15991 32643 15997
rect 33689 15997 33701 16031
rect 33735 15997 33747 16031
rect 33689 15991 33747 15997
rect 35437 16031 35495 16037
rect 35437 15997 35449 16031
rect 35483 15997 35495 16031
rect 35437 15991 35495 15997
rect 9309 15963 9367 15969
rect 9309 15929 9321 15963
rect 9355 15960 9367 15963
rect 9490 15960 9496 15972
rect 9355 15932 9496 15960
rect 9355 15929 9367 15932
rect 9309 15923 9367 15929
rect 9490 15920 9496 15932
rect 9548 15960 9554 15972
rect 10036 15963 10094 15969
rect 10036 15960 10048 15963
rect 9548 15932 10048 15960
rect 9548 15920 9554 15932
rect 10036 15929 10048 15932
rect 10082 15960 10094 15963
rect 10134 15960 10140 15972
rect 10082 15932 10140 15960
rect 10082 15929 10094 15932
rect 10036 15923 10094 15929
rect 10134 15920 10140 15932
rect 10192 15920 10198 15972
rect 24670 15920 24676 15972
rect 24728 15969 24734 15972
rect 24728 15963 24792 15969
rect 24728 15929 24746 15963
rect 24780 15929 24792 15963
rect 27341 15963 27399 15969
rect 27341 15960 27353 15963
rect 24728 15923 24792 15929
rect 26436 15932 27353 15960
rect 24728 15920 24734 15923
rect 8570 15892 8576 15904
rect 8531 15864 8576 15892
rect 8570 15852 8576 15864
rect 8628 15852 8634 15904
rect 13814 15892 13820 15904
rect 13775 15864 13820 15892
rect 13814 15852 13820 15864
rect 13872 15852 13878 15904
rect 20898 15852 20904 15904
rect 20956 15892 20962 15904
rect 21450 15892 21456 15904
rect 20956 15864 21456 15892
rect 20956 15852 20962 15864
rect 21450 15852 21456 15864
rect 21508 15892 21514 15904
rect 21729 15895 21787 15901
rect 21729 15892 21741 15895
rect 21508 15864 21741 15892
rect 21508 15852 21514 15864
rect 21729 15861 21741 15864
rect 21775 15861 21787 15895
rect 21729 15855 21787 15861
rect 22005 15895 22063 15901
rect 22005 15861 22017 15895
rect 22051 15892 22063 15895
rect 22738 15892 22744 15904
rect 22051 15864 22744 15892
rect 22051 15861 22063 15864
rect 22005 15855 22063 15861
rect 22738 15852 22744 15864
rect 22796 15852 22802 15904
rect 26234 15852 26240 15904
rect 26292 15892 26298 15904
rect 26436 15901 26464 15932
rect 27341 15929 27353 15932
rect 27387 15929 27399 15963
rect 30561 15963 30619 15969
rect 30561 15960 30573 15963
rect 27341 15923 27399 15929
rect 29932 15932 30573 15960
rect 26421 15895 26479 15901
rect 26421 15892 26433 15895
rect 26292 15864 26433 15892
rect 26292 15852 26298 15864
rect 26421 15861 26433 15864
rect 26467 15861 26479 15895
rect 26421 15855 26479 15861
rect 26878 15852 26884 15904
rect 26936 15892 26942 15904
rect 26973 15895 27031 15901
rect 26973 15892 26985 15895
rect 26936 15864 26985 15892
rect 26936 15852 26942 15864
rect 26973 15861 26985 15864
rect 27019 15861 27031 15895
rect 26973 15855 27031 15861
rect 28350 15852 28356 15904
rect 28408 15892 28414 15904
rect 28445 15895 28503 15901
rect 28445 15892 28457 15895
rect 28408 15864 28457 15892
rect 28408 15852 28414 15864
rect 28445 15861 28457 15864
rect 28491 15892 28503 15895
rect 29178 15892 29184 15904
rect 28491 15864 29184 15892
rect 28491 15861 28503 15864
rect 28445 15855 28503 15861
rect 29178 15852 29184 15864
rect 29236 15852 29242 15904
rect 29822 15852 29828 15904
rect 29880 15892 29886 15904
rect 29932 15901 29960 15932
rect 30561 15929 30573 15932
rect 30607 15929 30619 15963
rect 30561 15923 30619 15929
rect 29917 15895 29975 15901
rect 29917 15892 29929 15895
rect 29880 15864 29929 15892
rect 29880 15852 29886 15864
rect 29917 15861 29929 15864
rect 29963 15861 29975 15895
rect 29917 15855 29975 15861
rect 33597 15895 33655 15901
rect 33597 15861 33609 15895
rect 33643 15892 33655 15895
rect 33704 15892 33732 15991
rect 34422 15892 34428 15904
rect 33643 15864 34428 15892
rect 33643 15861 33655 15864
rect 33597 15855 33655 15861
rect 34422 15852 34428 15864
rect 34480 15852 34486 15904
rect 1104 15802 38824 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 38824 15802
rect 1104 15728 38824 15750
rect 8294 15688 8300 15700
rect 8255 15660 8300 15688
rect 8294 15648 8300 15660
rect 8352 15648 8358 15700
rect 9122 15688 9128 15700
rect 9083 15660 9128 15688
rect 9122 15648 9128 15660
rect 9180 15648 9186 15700
rect 9490 15688 9496 15700
rect 9451 15660 9496 15688
rect 9490 15648 9496 15660
rect 9548 15648 9554 15700
rect 10042 15688 10048 15700
rect 10003 15660 10048 15688
rect 10042 15648 10048 15660
rect 10100 15648 10106 15700
rect 11238 15688 11244 15700
rect 11199 15660 11244 15688
rect 11238 15648 11244 15660
rect 11296 15648 11302 15700
rect 12526 15648 12532 15700
rect 12584 15688 12590 15700
rect 12713 15691 12771 15697
rect 12713 15688 12725 15691
rect 12584 15660 12725 15688
rect 12584 15648 12590 15660
rect 12713 15657 12725 15660
rect 12759 15688 12771 15691
rect 13265 15691 13323 15697
rect 13265 15688 13277 15691
rect 12759 15660 13277 15688
rect 12759 15657 12771 15660
rect 12713 15651 12771 15657
rect 13265 15657 13277 15660
rect 13311 15657 13323 15691
rect 13265 15651 13323 15657
rect 22094 15648 22100 15700
rect 22152 15688 22158 15700
rect 22373 15691 22431 15697
rect 22373 15688 22385 15691
rect 22152 15660 22385 15688
rect 22152 15648 22158 15660
rect 22373 15657 22385 15660
rect 22419 15657 22431 15691
rect 22373 15651 22431 15657
rect 22738 15648 22744 15700
rect 22796 15688 22802 15700
rect 23293 15691 23351 15697
rect 23293 15688 23305 15691
rect 22796 15660 23305 15688
rect 22796 15648 22802 15660
rect 23293 15657 23305 15660
rect 23339 15657 23351 15691
rect 24302 15688 24308 15700
rect 24263 15660 24308 15688
rect 23293 15651 23351 15657
rect 24302 15648 24308 15660
rect 24360 15648 24366 15700
rect 24578 15648 24584 15700
rect 24636 15688 24642 15700
rect 24857 15691 24915 15697
rect 24857 15688 24869 15691
rect 24636 15660 24869 15688
rect 24636 15648 24642 15660
rect 24857 15657 24869 15660
rect 24903 15657 24915 15691
rect 30558 15688 30564 15700
rect 30519 15660 30564 15688
rect 24857 15651 24915 15657
rect 30558 15648 30564 15660
rect 30616 15648 30622 15700
rect 34241 15691 34299 15697
rect 34241 15657 34253 15691
rect 34287 15688 34299 15691
rect 34606 15688 34612 15700
rect 34287 15660 34612 15688
rect 34287 15657 34299 15660
rect 34241 15651 34299 15657
rect 34606 15648 34612 15660
rect 34664 15648 34670 15700
rect 6273 15623 6331 15629
rect 6273 15589 6285 15623
rect 6319 15620 6331 15623
rect 6610 15623 6668 15629
rect 6610 15620 6622 15623
rect 6319 15592 6622 15620
rect 6319 15589 6331 15592
rect 6273 15583 6331 15589
rect 6610 15589 6622 15592
rect 6656 15620 6668 15623
rect 8202 15620 8208 15632
rect 6656 15592 8208 15620
rect 6656 15589 6668 15592
rect 6610 15583 6668 15589
rect 8202 15580 8208 15592
rect 8260 15620 8266 15632
rect 8570 15620 8576 15632
rect 8260 15592 8576 15620
rect 8260 15580 8266 15592
rect 8570 15580 8576 15592
rect 8628 15620 8634 15632
rect 11606 15629 11612 15632
rect 8665 15623 8723 15629
rect 8665 15620 8677 15623
rect 8628 15592 8677 15620
rect 8628 15580 8634 15592
rect 8665 15589 8677 15592
rect 8711 15589 8723 15623
rect 11600 15620 11612 15629
rect 11567 15592 11612 15620
rect 8665 15583 8723 15589
rect 11600 15583 11612 15592
rect 11606 15580 11612 15583
rect 11664 15580 11670 15632
rect 23201 15623 23259 15629
rect 23201 15589 23213 15623
rect 23247 15620 23259 15623
rect 23382 15620 23388 15632
rect 23247 15592 23388 15620
rect 23247 15589 23259 15592
rect 23201 15583 23259 15589
rect 23382 15580 23388 15592
rect 23440 15580 23446 15632
rect 32861 15623 32919 15629
rect 32861 15589 32873 15623
rect 32907 15620 32919 15623
rect 32950 15620 32956 15632
rect 32907 15592 32956 15620
rect 32907 15589 32919 15592
rect 32861 15583 32919 15589
rect 32950 15580 32956 15592
rect 33008 15580 33014 15632
rect 7098 15552 7104 15564
rect 6380 15524 7104 15552
rect 6380 15496 6408 15524
rect 7098 15512 7104 15524
rect 7156 15512 7162 15564
rect 11330 15552 11336 15564
rect 11291 15524 11336 15552
rect 11330 15512 11336 15524
rect 11388 15512 11394 15564
rect 22097 15555 22155 15561
rect 22097 15521 22109 15555
rect 22143 15552 22155 15555
rect 22186 15552 22192 15564
rect 22143 15524 22192 15552
rect 22143 15521 22155 15524
rect 22097 15515 22155 15521
rect 22186 15512 22192 15524
rect 22244 15512 22250 15564
rect 23474 15512 23480 15564
rect 23532 15552 23538 15564
rect 24670 15552 24676 15564
rect 23532 15524 24676 15552
rect 23532 15512 23538 15524
rect 24670 15512 24676 15524
rect 24728 15552 24734 15564
rect 24765 15555 24823 15561
rect 24765 15552 24777 15555
rect 24728 15524 24777 15552
rect 24728 15512 24734 15524
rect 24765 15521 24777 15524
rect 24811 15521 24823 15555
rect 26878 15552 26884 15564
rect 26791 15524 26884 15552
rect 24765 15515 24823 15521
rect 26878 15512 26884 15524
rect 26936 15552 26942 15564
rect 27522 15552 27528 15564
rect 26936 15524 27528 15552
rect 26936 15512 26942 15524
rect 27522 15512 27528 15524
rect 27580 15512 27586 15564
rect 29178 15552 29184 15564
rect 29139 15524 29184 15552
rect 29178 15512 29184 15524
rect 29236 15512 29242 15564
rect 29454 15561 29460 15564
rect 29448 15552 29460 15561
rect 29415 15524 29460 15552
rect 29448 15515 29460 15524
rect 29454 15512 29460 15515
rect 29512 15512 29518 15564
rect 34054 15552 34060 15564
rect 34015 15524 34060 15552
rect 34054 15512 34060 15524
rect 34112 15512 34118 15564
rect 34606 15512 34612 15564
rect 34664 15552 34670 15564
rect 35529 15555 35587 15561
rect 35529 15552 35541 15555
rect 34664 15524 35541 15552
rect 34664 15512 34670 15524
rect 35529 15521 35541 15524
rect 35575 15521 35587 15555
rect 35529 15515 35587 15521
rect 6362 15484 6368 15496
rect 6323 15456 6368 15484
rect 6362 15444 6368 15456
rect 6420 15444 6426 15496
rect 9674 15444 9680 15496
rect 9732 15484 9738 15496
rect 10137 15487 10195 15493
rect 10137 15484 10149 15487
rect 9732 15456 10149 15484
rect 9732 15444 9738 15456
rect 10137 15453 10149 15456
rect 10183 15453 10195 15487
rect 10137 15447 10195 15453
rect 10226 15444 10232 15496
rect 10284 15484 10290 15496
rect 10284 15456 10329 15484
rect 10284 15444 10290 15456
rect 22922 15444 22928 15496
rect 22980 15484 22986 15496
rect 23385 15487 23443 15493
rect 23385 15484 23397 15487
rect 22980 15456 23397 15484
rect 22980 15444 22986 15456
rect 23385 15453 23397 15456
rect 23431 15453 23443 15487
rect 23385 15447 23443 15453
rect 24210 15444 24216 15496
rect 24268 15484 24274 15496
rect 24949 15487 25007 15493
rect 24949 15484 24961 15487
rect 24268 15456 24961 15484
rect 24268 15444 24274 15456
rect 24949 15453 24961 15456
rect 24995 15484 25007 15487
rect 25409 15487 25467 15493
rect 25409 15484 25421 15487
rect 24995 15456 25421 15484
rect 24995 15453 25007 15456
rect 24949 15447 25007 15453
rect 25409 15453 25421 15456
rect 25455 15484 25467 15487
rect 25958 15484 25964 15496
rect 25455 15456 25964 15484
rect 25455 15453 25467 15456
rect 25409 15447 25467 15453
rect 25958 15444 25964 15456
rect 26016 15444 26022 15496
rect 26418 15444 26424 15496
rect 26476 15484 26482 15496
rect 26973 15487 27031 15493
rect 26973 15484 26985 15487
rect 26476 15456 26985 15484
rect 26476 15444 26482 15456
rect 26973 15453 26985 15456
rect 27019 15453 27031 15487
rect 26973 15447 27031 15453
rect 27065 15487 27123 15493
rect 27065 15453 27077 15487
rect 27111 15453 27123 15487
rect 27065 15447 27123 15453
rect 22830 15416 22836 15428
rect 22791 15388 22836 15416
rect 22830 15376 22836 15388
rect 22888 15376 22894 15428
rect 23937 15419 23995 15425
rect 23937 15385 23949 15419
rect 23983 15416 23995 15419
rect 24762 15416 24768 15428
rect 23983 15388 24768 15416
rect 23983 15385 23995 15388
rect 23937 15379 23995 15385
rect 24762 15376 24768 15388
rect 24820 15376 24826 15428
rect 26786 15416 26792 15428
rect 26344 15388 26792 15416
rect 26344 15360 26372 15388
rect 26786 15376 26792 15388
rect 26844 15416 26850 15428
rect 27080 15416 27108 15447
rect 32398 15444 32404 15496
rect 32456 15484 32462 15496
rect 32953 15487 33011 15493
rect 32953 15484 32965 15487
rect 32456 15456 32965 15484
rect 32456 15444 32462 15456
rect 32953 15453 32965 15456
rect 32999 15453 33011 15487
rect 32953 15447 33011 15453
rect 33045 15487 33103 15493
rect 33045 15453 33057 15487
rect 33091 15453 33103 15487
rect 35618 15484 35624 15496
rect 35579 15456 35624 15484
rect 33045 15447 33103 15453
rect 26844 15388 27108 15416
rect 31941 15419 31999 15425
rect 26844 15376 26850 15388
rect 31941 15385 31953 15419
rect 31987 15416 31999 15419
rect 32858 15416 32864 15428
rect 31987 15388 32864 15416
rect 31987 15385 31999 15388
rect 31941 15379 31999 15385
rect 32858 15376 32864 15388
rect 32916 15416 32922 15428
rect 33060 15416 33088 15447
rect 35618 15444 35624 15456
rect 35676 15444 35682 15496
rect 35805 15487 35863 15493
rect 35805 15453 35817 15487
rect 35851 15484 35863 15487
rect 35851 15456 36032 15484
rect 35851 15453 35863 15456
rect 35805 15447 35863 15453
rect 32916 15388 33088 15416
rect 34977 15419 35035 15425
rect 32916 15376 32922 15388
rect 34977 15385 34989 15419
rect 35023 15416 35035 15419
rect 35342 15416 35348 15428
rect 35023 15388 35348 15416
rect 35023 15385 35035 15388
rect 34977 15379 35035 15385
rect 35342 15376 35348 15388
rect 35400 15376 35406 15428
rect 36004 15360 36032 15456
rect 5258 15348 5264 15360
rect 5219 15320 5264 15348
rect 5258 15308 5264 15320
rect 5316 15308 5322 15360
rect 7742 15348 7748 15360
rect 7703 15320 7748 15348
rect 7742 15308 7748 15320
rect 7800 15308 7806 15360
rect 9490 15308 9496 15360
rect 9548 15348 9554 15360
rect 9677 15351 9735 15357
rect 9677 15348 9689 15351
rect 9548 15320 9689 15348
rect 9548 15308 9554 15320
rect 9677 15317 9689 15320
rect 9723 15317 9735 15351
rect 19242 15348 19248 15360
rect 19203 15320 19248 15348
rect 9677 15311 9735 15317
rect 19242 15308 19248 15320
rect 19300 15308 19306 15360
rect 24394 15348 24400 15360
rect 24355 15320 24400 15348
rect 24394 15308 24400 15320
rect 24452 15308 24458 15360
rect 26326 15348 26332 15360
rect 26287 15320 26332 15348
rect 26326 15308 26332 15320
rect 26384 15308 26390 15360
rect 26510 15348 26516 15360
rect 26471 15320 26516 15348
rect 26510 15308 26516 15320
rect 26568 15308 26574 15360
rect 27522 15308 27528 15360
rect 27580 15348 27586 15360
rect 27617 15351 27675 15357
rect 27617 15348 27629 15351
rect 27580 15320 27629 15348
rect 27580 15308 27586 15320
rect 27617 15317 27629 15320
rect 27663 15317 27675 15351
rect 27617 15311 27675 15317
rect 32401 15351 32459 15357
rect 32401 15317 32413 15351
rect 32447 15348 32459 15351
rect 32493 15351 32551 15357
rect 32493 15348 32505 15351
rect 32447 15320 32505 15348
rect 32447 15317 32459 15320
rect 32401 15311 32459 15317
rect 32493 15317 32505 15320
rect 32539 15348 32551 15351
rect 33042 15348 33048 15360
rect 32539 15320 33048 15348
rect 32539 15317 32551 15320
rect 32493 15311 32551 15317
rect 33042 15308 33048 15320
rect 33100 15308 33106 15360
rect 33410 15308 33416 15360
rect 33468 15348 33474 15360
rect 33505 15351 33563 15357
rect 33505 15348 33517 15351
rect 33468 15320 33517 15348
rect 33468 15308 33474 15320
rect 33505 15317 33517 15320
rect 33551 15317 33563 15351
rect 33962 15348 33968 15360
rect 33923 15320 33968 15348
rect 33505 15311 33563 15317
rect 33962 15308 33968 15320
rect 34020 15308 34026 15360
rect 35161 15351 35219 15357
rect 35161 15317 35173 15351
rect 35207 15348 35219 15351
rect 35250 15348 35256 15360
rect 35207 15320 35256 15348
rect 35207 15317 35219 15320
rect 35161 15311 35219 15317
rect 35250 15308 35256 15320
rect 35308 15308 35314 15360
rect 35986 15308 35992 15360
rect 36044 15348 36050 15360
rect 36170 15348 36176 15360
rect 36044 15320 36176 15348
rect 36044 15308 36050 15320
rect 36170 15308 36176 15320
rect 36228 15308 36234 15360
rect 1104 15258 38824 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 34966 15258
rect 35018 15206 35030 15258
rect 35082 15206 35094 15258
rect 35146 15206 35158 15258
rect 35210 15206 38824 15258
rect 1104 15184 38824 15206
rect 9401 15147 9459 15153
rect 9401 15113 9413 15147
rect 9447 15144 9459 15147
rect 9582 15144 9588 15156
rect 9447 15116 9588 15144
rect 9447 15113 9459 15116
rect 9401 15107 9459 15113
rect 9582 15104 9588 15116
rect 9640 15104 9646 15156
rect 11330 15144 11336 15156
rect 11291 15116 11336 15144
rect 11330 15104 11336 15116
rect 11388 15104 11394 15156
rect 11606 15104 11612 15156
rect 11664 15144 11670 15156
rect 11701 15147 11759 15153
rect 11701 15144 11713 15147
rect 11664 15116 11713 15144
rect 11664 15104 11670 15116
rect 11701 15113 11713 15116
rect 11747 15113 11759 15147
rect 11701 15107 11759 15113
rect 18874 15104 18880 15156
rect 18932 15144 18938 15156
rect 18969 15147 19027 15153
rect 18969 15144 18981 15147
rect 18932 15116 18981 15144
rect 18932 15104 18938 15116
rect 18969 15113 18981 15116
rect 19015 15113 19027 15147
rect 18969 15107 19027 15113
rect 5258 14968 5264 15020
rect 5316 15008 5322 15020
rect 5810 15008 5816 15020
rect 5316 14980 5816 15008
rect 5316 14968 5322 14980
rect 5810 14968 5816 14980
rect 5868 14968 5874 15020
rect 9858 14968 9864 15020
rect 9916 15008 9922 15020
rect 10226 15008 10232 15020
rect 9916 14980 10232 15008
rect 9916 14968 9922 14980
rect 10226 14968 10232 14980
rect 10284 15008 10290 15020
rect 10781 15011 10839 15017
rect 10781 15008 10793 15011
rect 10284 14980 10793 15008
rect 10284 14968 10290 14980
rect 10781 14977 10793 14980
rect 10827 14977 10839 15011
rect 10781 14971 10839 14977
rect 17954 14968 17960 15020
rect 18012 15008 18018 15020
rect 18984 15008 19012 15107
rect 22738 15104 22744 15156
rect 22796 15144 22802 15156
rect 22833 15147 22891 15153
rect 22833 15144 22845 15147
rect 22796 15116 22845 15144
rect 22796 15104 22802 15116
rect 22833 15113 22845 15116
rect 22879 15113 22891 15147
rect 23474 15144 23480 15156
rect 23435 15116 23480 15144
rect 22833 15107 22891 15113
rect 23474 15104 23480 15116
rect 23532 15104 23538 15156
rect 24029 15147 24087 15153
rect 24029 15113 24041 15147
rect 24075 15144 24087 15147
rect 24486 15144 24492 15156
rect 24075 15116 24492 15144
rect 24075 15113 24087 15116
rect 24029 15107 24087 15113
rect 24486 15104 24492 15116
rect 24544 15104 24550 15156
rect 26418 15104 26424 15156
rect 26476 15144 26482 15156
rect 26513 15147 26571 15153
rect 26513 15144 26525 15147
rect 26476 15116 26525 15144
rect 26476 15104 26482 15116
rect 26513 15113 26525 15116
rect 26559 15113 26571 15147
rect 27614 15144 27620 15156
rect 27575 15116 27620 15144
rect 26513 15107 26571 15113
rect 27614 15104 27620 15116
rect 27672 15104 27678 15156
rect 29178 15104 29184 15156
rect 29236 15144 29242 15156
rect 29457 15147 29515 15153
rect 29457 15144 29469 15147
rect 29236 15116 29469 15144
rect 29236 15104 29242 15116
rect 29457 15113 29469 15116
rect 29503 15144 29515 15147
rect 30285 15147 30343 15153
rect 30285 15144 30297 15147
rect 29503 15116 30297 15144
rect 29503 15113 29515 15116
rect 29457 15107 29515 15113
rect 30285 15113 30297 15116
rect 30331 15113 30343 15147
rect 30285 15107 30343 15113
rect 22557 15079 22615 15085
rect 22557 15045 22569 15079
rect 22603 15076 22615 15079
rect 23382 15076 23388 15088
rect 22603 15048 23388 15076
rect 22603 15045 22615 15048
rect 22557 15039 22615 15045
rect 23382 15036 23388 15048
rect 23440 15036 23446 15088
rect 24302 15076 24308 15088
rect 24263 15048 24308 15076
rect 24302 15036 24308 15048
rect 24360 15076 24366 15088
rect 24360 15048 24532 15076
rect 24360 15036 24366 15048
rect 24504 15017 24532 15048
rect 19153 15011 19211 15017
rect 19153 15008 19165 15011
rect 18012 14980 19165 15008
rect 18012 14968 18018 14980
rect 19153 14977 19165 14980
rect 19199 14977 19211 15011
rect 19153 14971 19211 14977
rect 24489 15011 24547 15017
rect 24489 14977 24501 15011
rect 24535 14977 24547 15011
rect 30300 15008 30328 15107
rect 34422 15104 34428 15156
rect 34480 15144 34486 15156
rect 34885 15147 34943 15153
rect 34885 15144 34897 15147
rect 34480 15116 34897 15144
rect 34480 15104 34486 15116
rect 34885 15113 34897 15116
rect 34931 15113 34943 15147
rect 37090 15144 37096 15156
rect 37051 15116 37096 15144
rect 34885 15107 34943 15113
rect 37090 15104 37096 15116
rect 37148 15104 37154 15156
rect 32953 15079 33011 15085
rect 32953 15045 32965 15079
rect 32999 15076 33011 15079
rect 34054 15076 34060 15088
rect 32999 15048 34060 15076
rect 32999 15045 33011 15048
rect 32953 15039 33011 15045
rect 34054 15036 34060 15048
rect 34112 15036 34118 15088
rect 30469 15011 30527 15017
rect 30469 15008 30481 15011
rect 30300 14980 30481 15008
rect 24489 14971 24547 14977
rect 30469 14977 30481 14980
rect 30515 14977 30527 15011
rect 33410 15008 33416 15020
rect 33371 14980 33416 15008
rect 30469 14971 30527 14977
rect 6362 14900 6368 14952
rect 6420 14940 6426 14952
rect 6457 14943 6515 14949
rect 6457 14940 6469 14943
rect 6420 14912 6469 14940
rect 6420 14900 6426 14912
rect 6457 14909 6469 14912
rect 6503 14940 6515 14943
rect 6825 14943 6883 14949
rect 6825 14940 6837 14943
rect 6503 14912 6837 14940
rect 6503 14909 6515 14912
rect 6457 14903 6515 14909
rect 6825 14909 6837 14912
rect 6871 14909 6883 14943
rect 6825 14903 6883 14909
rect 9769 14943 9827 14949
rect 9769 14909 9781 14943
rect 9815 14940 9827 14943
rect 10597 14943 10655 14949
rect 10597 14940 10609 14943
rect 9815 14912 10609 14940
rect 9815 14909 9827 14912
rect 9769 14903 9827 14909
rect 10597 14909 10609 14912
rect 10643 14940 10655 14943
rect 10686 14940 10692 14952
rect 10643 14912 10692 14940
rect 10643 14909 10655 14912
rect 10597 14903 10655 14909
rect 10686 14900 10692 14912
rect 10744 14900 10750 14952
rect 19242 14900 19248 14952
rect 19300 14940 19306 14952
rect 24762 14949 24768 14952
rect 19409 14943 19467 14949
rect 19409 14940 19421 14943
rect 19300 14912 19421 14940
rect 19300 14900 19306 14912
rect 19409 14909 19421 14912
rect 19455 14909 19467 14943
rect 24756 14940 24768 14949
rect 24723 14912 24768 14940
rect 19409 14903 19467 14909
rect 24756 14903 24768 14912
rect 24762 14900 24768 14903
rect 24820 14900 24826 14952
rect 26510 14900 26516 14952
rect 26568 14940 26574 14952
rect 26973 14943 27031 14949
rect 26973 14940 26985 14943
rect 26568 14912 26985 14940
rect 26568 14900 26574 14912
rect 26973 14909 26985 14912
rect 27019 14940 27031 14943
rect 27893 14943 27951 14949
rect 27893 14940 27905 14943
rect 27019 14912 27905 14940
rect 27019 14909 27031 14912
rect 26973 14903 27031 14909
rect 27893 14909 27905 14912
rect 27939 14909 27951 14943
rect 27893 14903 27951 14909
rect 29089 14943 29147 14949
rect 29089 14909 29101 14943
rect 29135 14940 29147 14943
rect 29454 14940 29460 14952
rect 29135 14912 29460 14940
rect 29135 14909 29147 14912
rect 29089 14903 29147 14909
rect 29454 14900 29460 14912
rect 29512 14940 29518 14952
rect 30282 14940 30288 14952
rect 29512 14912 30288 14940
rect 29512 14900 29518 14912
rect 30282 14900 30288 14912
rect 30340 14900 30346 14952
rect 30484 14940 30512 14971
rect 33410 14968 33416 14980
rect 33468 14968 33474 15020
rect 33597 15011 33655 15017
rect 33597 14977 33609 15011
rect 33643 15008 33655 15011
rect 33962 15008 33968 15020
rect 33643 14980 33968 15008
rect 33643 14977 33655 14980
rect 33597 14971 33655 14977
rect 33962 14968 33968 14980
rect 34020 15008 34026 15020
rect 35526 15008 35532 15020
rect 34020 14980 35532 15008
rect 34020 14968 34026 14980
rect 35526 14968 35532 14980
rect 35584 14968 35590 15020
rect 32122 14940 32128 14952
rect 30484 14912 32128 14940
rect 32122 14900 32128 14912
rect 32180 14900 32186 14952
rect 33134 14900 33140 14952
rect 33192 14940 33198 14952
rect 33321 14943 33379 14949
rect 33321 14940 33333 14943
rect 33192 14912 33333 14940
rect 33192 14900 33198 14912
rect 33321 14909 33333 14912
rect 33367 14909 33379 14943
rect 35250 14940 35256 14952
rect 35211 14912 35256 14940
rect 33321 14903 33379 14909
rect 35250 14900 35256 14912
rect 35308 14940 35314 14952
rect 36265 14943 36323 14949
rect 36265 14940 36277 14943
rect 35308 14912 36277 14940
rect 35308 14900 35314 14912
rect 36265 14909 36277 14912
rect 36311 14909 36323 14943
rect 36265 14903 36323 14909
rect 36449 14943 36507 14949
rect 36449 14909 36461 14943
rect 36495 14940 36507 14943
rect 37090 14940 37096 14952
rect 36495 14912 37096 14940
rect 36495 14909 36507 14912
rect 36449 14903 36507 14909
rect 37090 14900 37096 14912
rect 37148 14900 37154 14952
rect 5077 14875 5135 14881
rect 5077 14841 5089 14875
rect 5123 14872 5135 14875
rect 5629 14875 5687 14881
rect 5629 14872 5641 14875
rect 5123 14844 5641 14872
rect 5123 14841 5135 14844
rect 5077 14835 5135 14841
rect 5629 14841 5641 14844
rect 5675 14872 5687 14875
rect 7092 14875 7150 14881
rect 7092 14872 7104 14875
rect 5675 14844 7104 14872
rect 5675 14841 5687 14844
rect 5629 14835 5687 14841
rect 7092 14841 7104 14844
rect 7138 14872 7150 14875
rect 7742 14872 7748 14884
rect 7138 14844 7748 14872
rect 7138 14841 7150 14844
rect 7092 14835 7150 14841
rect 7742 14832 7748 14844
rect 7800 14832 7806 14884
rect 7834 14832 7840 14884
rect 7892 14872 7898 14884
rect 8941 14875 8999 14881
rect 8941 14872 8953 14875
rect 7892 14844 8953 14872
rect 7892 14832 7898 14844
rect 8941 14841 8953 14844
rect 8987 14872 8999 14875
rect 9858 14872 9864 14884
rect 8987 14844 9864 14872
rect 8987 14841 8999 14844
rect 8941 14835 8999 14841
rect 9858 14832 9864 14844
rect 9916 14832 9922 14884
rect 10137 14875 10195 14881
rect 10137 14841 10149 14875
rect 10183 14872 10195 14875
rect 10183 14844 10732 14872
rect 10183 14841 10195 14844
rect 10137 14835 10195 14841
rect 5166 14804 5172 14816
rect 5127 14776 5172 14804
rect 5166 14764 5172 14776
rect 5224 14764 5230 14816
rect 5534 14804 5540 14816
rect 5495 14776 5540 14804
rect 5534 14764 5540 14776
rect 5592 14764 5598 14816
rect 5718 14764 5724 14816
rect 5776 14804 5782 14816
rect 6181 14807 6239 14813
rect 6181 14804 6193 14807
rect 5776 14776 6193 14804
rect 5776 14764 5782 14776
rect 6181 14773 6193 14776
rect 6227 14804 6239 14807
rect 6457 14807 6515 14813
rect 6457 14804 6469 14807
rect 6227 14776 6469 14804
rect 6227 14773 6239 14776
rect 6181 14767 6239 14773
rect 6457 14773 6469 14776
rect 6503 14804 6515 14807
rect 6549 14807 6607 14813
rect 6549 14804 6561 14807
rect 6503 14776 6561 14804
rect 6503 14773 6515 14776
rect 6457 14767 6515 14773
rect 6549 14773 6561 14776
rect 6595 14773 6607 14807
rect 6549 14767 6607 14773
rect 6638 14764 6644 14816
rect 6696 14804 6702 14816
rect 8205 14807 8263 14813
rect 8205 14804 8217 14807
rect 6696 14776 8217 14804
rect 6696 14764 6702 14776
rect 8205 14773 8217 14776
rect 8251 14773 8263 14807
rect 10226 14804 10232 14816
rect 10187 14776 10232 14804
rect 8205 14767 8263 14773
rect 10226 14764 10232 14776
rect 10284 14764 10290 14816
rect 10704 14813 10732 14844
rect 26786 14832 26792 14884
rect 26844 14872 26850 14884
rect 28261 14875 28319 14881
rect 28261 14872 28273 14875
rect 26844 14844 28273 14872
rect 26844 14832 26850 14844
rect 28261 14841 28273 14844
rect 28307 14872 28319 14875
rect 28442 14872 28448 14884
rect 28307 14844 28448 14872
rect 28307 14841 28319 14844
rect 28261 14835 28319 14841
rect 28442 14832 28448 14844
rect 28500 14832 28506 14884
rect 30742 14881 30748 14884
rect 30009 14875 30067 14881
rect 30009 14841 30021 14875
rect 30055 14872 30067 14875
rect 30736 14872 30748 14881
rect 30055 14844 30748 14872
rect 30055 14841 30067 14844
rect 30009 14835 30067 14841
rect 30736 14835 30748 14844
rect 30742 14832 30748 14835
rect 30800 14832 30806 14884
rect 10689 14807 10747 14813
rect 10689 14773 10701 14807
rect 10735 14804 10747 14807
rect 10778 14804 10784 14816
rect 10735 14776 10784 14804
rect 10735 14773 10747 14776
rect 10689 14767 10747 14773
rect 10778 14764 10784 14776
rect 10836 14764 10842 14816
rect 20530 14804 20536 14816
rect 20491 14776 20536 14804
rect 20530 14764 20536 14776
rect 20588 14764 20594 14816
rect 25866 14804 25872 14816
rect 25827 14776 25872 14804
rect 25866 14764 25872 14776
rect 25924 14804 25930 14816
rect 26234 14804 26240 14816
rect 25924 14776 26240 14804
rect 25924 14764 25930 14776
rect 26234 14764 26240 14776
rect 26292 14764 26298 14816
rect 27062 14764 27068 14816
rect 27120 14804 27126 14816
rect 27157 14807 27215 14813
rect 27157 14804 27169 14807
rect 27120 14776 27169 14804
rect 27120 14764 27126 14776
rect 27157 14773 27169 14776
rect 27203 14773 27215 14807
rect 31846 14804 31852 14816
rect 31807 14776 31852 14804
rect 27157 14767 27215 14773
rect 31846 14764 31852 14776
rect 31904 14764 31910 14816
rect 32398 14764 32404 14816
rect 32456 14804 32462 14816
rect 32493 14807 32551 14813
rect 32493 14804 32505 14807
rect 32456 14776 32505 14804
rect 32456 14764 32462 14776
rect 32493 14773 32505 14776
rect 32539 14773 32551 14807
rect 32493 14767 32551 14773
rect 32950 14764 32956 14816
rect 33008 14804 33014 14816
rect 33594 14804 33600 14816
rect 33008 14776 33600 14804
rect 33008 14764 33014 14776
rect 33594 14764 33600 14776
rect 33652 14804 33658 14816
rect 33965 14807 34023 14813
rect 33965 14804 33977 14807
rect 33652 14776 33977 14804
rect 33652 14764 33658 14776
rect 33965 14773 33977 14776
rect 34011 14773 34023 14807
rect 34606 14804 34612 14816
rect 34567 14776 34612 14804
rect 33965 14767 34023 14773
rect 34606 14764 34612 14776
rect 34664 14764 34670 14816
rect 35250 14764 35256 14816
rect 35308 14804 35314 14816
rect 35345 14807 35403 14813
rect 35345 14804 35357 14807
rect 35308 14776 35357 14804
rect 35308 14764 35314 14776
rect 35345 14773 35357 14776
rect 35391 14773 35403 14807
rect 35345 14767 35403 14773
rect 35618 14764 35624 14816
rect 35676 14804 35682 14816
rect 35897 14807 35955 14813
rect 35897 14804 35909 14807
rect 35676 14776 35909 14804
rect 35676 14764 35682 14776
rect 35897 14773 35909 14776
rect 35943 14773 35955 14807
rect 36630 14804 36636 14816
rect 36591 14776 36636 14804
rect 35897 14767 35955 14773
rect 36630 14764 36636 14776
rect 36688 14764 36694 14816
rect 1104 14714 38824 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 38824 14714
rect 1104 14640 38824 14662
rect 7742 14600 7748 14612
rect 7703 14572 7748 14600
rect 7742 14560 7748 14572
rect 7800 14560 7806 14612
rect 9953 14603 10011 14609
rect 9953 14569 9965 14603
rect 9999 14600 10011 14603
rect 10042 14600 10048 14612
rect 9999 14572 10048 14600
rect 9999 14569 10011 14572
rect 9953 14563 10011 14569
rect 10042 14560 10048 14572
rect 10100 14560 10106 14612
rect 19242 14560 19248 14612
rect 19300 14600 19306 14612
rect 19337 14603 19395 14609
rect 19337 14600 19349 14603
rect 19300 14572 19349 14600
rect 19300 14560 19306 14572
rect 19337 14569 19349 14572
rect 19383 14569 19395 14603
rect 22922 14600 22928 14612
rect 22883 14572 22928 14600
rect 19337 14563 19395 14569
rect 22922 14560 22928 14572
rect 22980 14560 22986 14612
rect 23753 14603 23811 14609
rect 23753 14569 23765 14603
rect 23799 14600 23811 14603
rect 24302 14600 24308 14612
rect 23799 14572 24308 14600
rect 23799 14569 23811 14572
rect 23753 14563 23811 14569
rect 24302 14560 24308 14572
rect 24360 14560 24366 14612
rect 26694 14560 26700 14612
rect 26752 14600 26758 14612
rect 27157 14603 27215 14609
rect 27157 14600 27169 14603
rect 26752 14572 27169 14600
rect 26752 14560 26758 14572
rect 27157 14569 27169 14572
rect 27203 14600 27215 14603
rect 28074 14600 28080 14612
rect 27203 14572 28080 14600
rect 27203 14569 27215 14572
rect 27157 14563 27215 14569
rect 28074 14560 28080 14572
rect 28132 14560 28138 14612
rect 28442 14600 28448 14612
rect 28403 14572 28448 14600
rect 28442 14560 28448 14572
rect 28500 14560 28506 14612
rect 29822 14600 29828 14612
rect 29783 14572 29828 14600
rect 29822 14560 29828 14572
rect 29880 14560 29886 14612
rect 30282 14600 30288 14612
rect 30243 14572 30288 14600
rect 30282 14560 30288 14572
rect 30340 14560 30346 14612
rect 32953 14603 33011 14609
rect 32953 14569 32965 14603
rect 32999 14600 33011 14603
rect 33410 14600 33416 14612
rect 32999 14572 33416 14600
rect 32999 14569 33011 14572
rect 32953 14563 33011 14569
rect 33410 14560 33416 14572
rect 33468 14560 33474 14612
rect 34054 14600 34060 14612
rect 34015 14572 34060 14600
rect 34054 14560 34060 14572
rect 34112 14560 34118 14612
rect 35526 14560 35532 14612
rect 35584 14600 35590 14612
rect 36446 14600 36452 14612
rect 35584 14572 36452 14600
rect 35584 14560 35590 14572
rect 36446 14560 36452 14572
rect 36504 14560 36510 14612
rect 8754 14532 8760 14544
rect 8496 14504 8760 14532
rect 5261 14467 5319 14473
rect 5261 14433 5273 14467
rect 5307 14464 5319 14467
rect 5534 14464 5540 14476
rect 5307 14436 5540 14464
rect 5307 14433 5319 14436
rect 5261 14427 5319 14433
rect 5534 14424 5540 14436
rect 5592 14464 5598 14476
rect 6080 14467 6138 14473
rect 6080 14464 6092 14467
rect 5592 14436 6092 14464
rect 5592 14424 5598 14436
rect 6080 14433 6092 14436
rect 6126 14464 6138 14467
rect 6638 14464 6644 14476
rect 6126 14436 6644 14464
rect 6126 14433 6138 14436
rect 6080 14427 6138 14433
rect 6638 14424 6644 14436
rect 6696 14424 6702 14476
rect 8496 14473 8524 14504
rect 8754 14492 8760 14504
rect 8812 14532 8818 14544
rect 9490 14532 9496 14544
rect 8812 14504 9496 14532
rect 8812 14492 8818 14504
rect 9490 14492 9496 14504
rect 9548 14492 9554 14544
rect 9858 14492 9864 14544
rect 9916 14532 9922 14544
rect 10597 14535 10655 14541
rect 10597 14532 10609 14535
rect 9916 14504 10609 14532
rect 9916 14492 9922 14504
rect 10597 14501 10609 14504
rect 10643 14501 10655 14535
rect 10597 14495 10655 14501
rect 16853 14535 16911 14541
rect 16853 14501 16865 14535
rect 16899 14532 16911 14535
rect 16942 14532 16948 14544
rect 16899 14504 16948 14532
rect 16899 14501 16911 14504
rect 16853 14495 16911 14501
rect 16942 14492 16948 14504
rect 17000 14492 17006 14544
rect 30190 14532 30196 14544
rect 30151 14504 30196 14532
rect 30190 14492 30196 14504
rect 30248 14492 30254 14544
rect 31846 14492 31852 14544
rect 31904 14532 31910 14544
rect 31941 14535 31999 14541
rect 31941 14532 31953 14535
rect 31904 14504 31953 14532
rect 31904 14492 31910 14504
rect 31941 14501 31953 14504
rect 31987 14532 31999 14535
rect 32858 14532 32864 14544
rect 31987 14504 32864 14532
rect 31987 14501 31999 14504
rect 31941 14495 31999 14501
rect 32858 14492 32864 14504
rect 32916 14532 32922 14544
rect 32916 14504 33640 14532
rect 32916 14492 32922 14504
rect 8481 14467 8539 14473
rect 8481 14433 8493 14467
rect 8527 14433 8539 14467
rect 8481 14427 8539 14433
rect 9214 14424 9220 14476
rect 9272 14464 9278 14476
rect 10045 14467 10103 14473
rect 10045 14464 10057 14467
rect 9272 14436 10057 14464
rect 9272 14424 9278 14436
rect 10045 14433 10057 14436
rect 10091 14464 10103 14467
rect 10226 14464 10232 14476
rect 10091 14436 10232 14464
rect 10091 14433 10103 14436
rect 10045 14427 10103 14433
rect 10226 14424 10232 14436
rect 10284 14424 10290 14476
rect 11054 14424 11060 14476
rect 11112 14464 11118 14476
rect 11149 14467 11207 14473
rect 11149 14464 11161 14467
rect 11112 14436 11161 14464
rect 11112 14424 11118 14436
rect 11149 14433 11161 14436
rect 11195 14433 11207 14467
rect 11149 14427 11207 14433
rect 16301 14467 16359 14473
rect 16301 14433 16313 14467
rect 16347 14464 16359 14467
rect 16761 14467 16819 14473
rect 16761 14464 16773 14467
rect 16347 14436 16773 14464
rect 16347 14433 16359 14436
rect 16301 14427 16359 14433
rect 16761 14433 16773 14436
rect 16807 14464 16819 14467
rect 18046 14464 18052 14476
rect 16807 14436 18052 14464
rect 16807 14433 16819 14436
rect 16761 14427 16819 14433
rect 18046 14424 18052 14436
rect 18104 14464 18110 14476
rect 18213 14467 18271 14473
rect 18213 14464 18225 14467
rect 18104 14436 18225 14464
rect 18104 14424 18110 14436
rect 18213 14433 18225 14436
rect 18259 14433 18271 14467
rect 18213 14427 18271 14433
rect 23566 14424 23572 14476
rect 23624 14464 23630 14476
rect 24121 14467 24179 14473
rect 24121 14464 24133 14467
rect 23624 14436 24133 14464
rect 23624 14424 23630 14436
rect 24121 14433 24133 14436
rect 24167 14433 24179 14467
rect 27062 14464 27068 14476
rect 27023 14436 27068 14464
rect 24121 14427 24179 14433
rect 27062 14424 27068 14436
rect 27120 14424 27126 14476
rect 32582 14424 32588 14476
rect 32640 14464 32646 14476
rect 33321 14467 33379 14473
rect 33321 14464 33333 14467
rect 32640 14436 33333 14464
rect 32640 14424 32646 14436
rect 33321 14433 33333 14436
rect 33367 14433 33379 14467
rect 33321 14427 33379 14433
rect 5718 14356 5724 14408
rect 5776 14396 5782 14408
rect 5813 14399 5871 14405
rect 5813 14396 5825 14399
rect 5776 14368 5825 14396
rect 5776 14356 5782 14368
rect 5813 14365 5825 14368
rect 5859 14365 5871 14399
rect 5813 14359 5871 14365
rect 17037 14399 17095 14405
rect 17037 14365 17049 14399
rect 17083 14365 17095 14399
rect 17954 14396 17960 14408
rect 17915 14368 17960 14396
rect 17037 14359 17095 14365
rect 16574 14288 16580 14340
rect 16632 14328 16638 14340
rect 17052 14328 17080 14359
rect 17954 14356 17960 14368
rect 18012 14356 18018 14408
rect 27341 14399 27399 14405
rect 27341 14365 27353 14399
rect 27387 14396 27399 14399
rect 27522 14396 27528 14408
rect 27387 14368 27528 14396
rect 27387 14365 27399 14368
rect 27341 14359 27399 14365
rect 27522 14356 27528 14368
rect 27580 14356 27586 14408
rect 29914 14356 29920 14408
rect 29972 14396 29978 14408
rect 30466 14396 30472 14408
rect 29972 14368 30472 14396
rect 29972 14356 29978 14368
rect 30466 14356 30472 14368
rect 30524 14356 30530 14408
rect 33612 14405 33640 14504
rect 34606 14424 34612 14476
rect 34664 14464 34670 14476
rect 34773 14467 34831 14473
rect 34773 14464 34785 14467
rect 34664 14436 34785 14464
rect 34664 14424 34670 14436
rect 34773 14433 34785 14436
rect 34819 14433 34831 14467
rect 34773 14427 34831 14433
rect 33413 14399 33471 14405
rect 33413 14365 33425 14399
rect 33459 14365 33471 14399
rect 33413 14359 33471 14365
rect 33597 14399 33655 14405
rect 33597 14365 33609 14399
rect 33643 14396 33655 14399
rect 33686 14396 33692 14408
rect 33643 14368 33692 14396
rect 33643 14365 33655 14368
rect 33597 14359 33655 14365
rect 16632 14300 17908 14328
rect 16632 14288 16638 14300
rect 6822 14220 6828 14272
rect 6880 14260 6886 14272
rect 7193 14263 7251 14269
rect 7193 14260 7205 14263
rect 6880 14232 7205 14260
rect 6880 14220 6886 14232
rect 7193 14229 7205 14232
rect 7239 14229 7251 14263
rect 7193 14223 7251 14229
rect 8665 14263 8723 14269
rect 8665 14229 8677 14263
rect 8711 14260 8723 14263
rect 9490 14260 9496 14272
rect 8711 14232 9496 14260
rect 8711 14229 8723 14232
rect 8665 14223 8723 14229
rect 9490 14220 9496 14232
rect 9548 14220 9554 14272
rect 9950 14220 9956 14272
rect 10008 14260 10014 14272
rect 10229 14263 10287 14269
rect 10229 14260 10241 14263
rect 10008 14232 10241 14260
rect 10008 14220 10014 14232
rect 10229 14229 10241 14232
rect 10275 14229 10287 14263
rect 10229 14223 10287 14229
rect 11238 14220 11244 14272
rect 11296 14260 11302 14272
rect 11333 14263 11391 14269
rect 11333 14260 11345 14263
rect 11296 14232 11345 14260
rect 11296 14220 11302 14232
rect 11333 14229 11345 14232
rect 11379 14229 11391 14263
rect 11333 14223 11391 14229
rect 15565 14263 15623 14269
rect 15565 14229 15577 14263
rect 15611 14260 15623 14263
rect 15746 14260 15752 14272
rect 15611 14232 15752 14260
rect 15611 14229 15623 14232
rect 15565 14223 15623 14229
rect 15746 14220 15752 14232
rect 15804 14220 15810 14272
rect 16390 14260 16396 14272
rect 16351 14232 16396 14260
rect 16390 14220 16396 14232
rect 16448 14220 16454 14272
rect 17880 14269 17908 14300
rect 17865 14263 17923 14269
rect 17865 14229 17877 14263
rect 17911 14260 17923 14263
rect 18966 14260 18972 14272
rect 17911 14232 18972 14260
rect 17911 14229 17923 14232
rect 17865 14223 17923 14229
rect 18966 14220 18972 14232
rect 19024 14220 19030 14272
rect 25406 14260 25412 14272
rect 25367 14232 25412 14260
rect 25406 14220 25412 14232
rect 25464 14220 25470 14272
rect 26326 14260 26332 14272
rect 26287 14232 26332 14260
rect 26326 14220 26332 14232
rect 26384 14220 26390 14272
rect 26694 14260 26700 14272
rect 26655 14232 26700 14260
rect 26694 14220 26700 14232
rect 26752 14220 26758 14272
rect 27614 14220 27620 14272
rect 27672 14260 27678 14272
rect 27709 14263 27767 14269
rect 27709 14260 27721 14263
rect 27672 14232 27721 14260
rect 27672 14220 27678 14232
rect 27709 14229 27721 14232
rect 27755 14229 27767 14263
rect 27709 14223 27767 14229
rect 27798 14220 27804 14272
rect 27856 14260 27862 14272
rect 28077 14263 28135 14269
rect 28077 14260 28089 14263
rect 27856 14232 28089 14260
rect 27856 14220 27862 14232
rect 28077 14229 28089 14232
rect 28123 14229 28135 14263
rect 28077 14223 28135 14229
rect 32493 14263 32551 14269
rect 32493 14229 32505 14263
rect 32539 14260 32551 14263
rect 32582 14260 32588 14272
rect 32539 14232 32588 14260
rect 32539 14229 32551 14232
rect 32493 14223 32551 14229
rect 32582 14220 32588 14232
rect 32640 14220 32646 14272
rect 32861 14263 32919 14269
rect 32861 14229 32873 14263
rect 32907 14260 32919 14263
rect 32950 14260 32956 14272
rect 32907 14232 32956 14260
rect 32907 14229 32919 14232
rect 32861 14223 32919 14229
rect 32950 14220 32956 14232
rect 33008 14260 33014 14272
rect 33428 14260 33456 14359
rect 33686 14356 33692 14368
rect 33744 14356 33750 14408
rect 34422 14356 34428 14408
rect 34480 14396 34486 14408
rect 34517 14399 34575 14405
rect 34517 14396 34529 14399
rect 34480 14368 34529 14396
rect 34480 14356 34486 14368
rect 34517 14365 34529 14368
rect 34563 14365 34575 14399
rect 34517 14359 34575 14365
rect 35897 14263 35955 14269
rect 35897 14260 35909 14263
rect 33008 14232 35909 14260
rect 33008 14220 33014 14232
rect 35897 14229 35909 14232
rect 35943 14229 35955 14263
rect 35897 14223 35955 14229
rect 1104 14170 38824 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 34966 14170
rect 35018 14118 35030 14170
rect 35082 14118 35094 14170
rect 35146 14118 35158 14170
rect 35210 14118 38824 14170
rect 1104 14096 38824 14118
rect 6638 14056 6644 14068
rect 6599 14028 6644 14056
rect 6638 14016 6644 14028
rect 6696 14016 6702 14068
rect 8754 14056 8760 14068
rect 8715 14028 8760 14056
rect 8754 14016 8760 14028
rect 8812 14016 8818 14068
rect 9214 14056 9220 14068
rect 9175 14028 9220 14056
rect 9214 14016 9220 14028
rect 9272 14016 9278 14068
rect 9490 14056 9496 14068
rect 9451 14028 9496 14056
rect 9490 14016 9496 14028
rect 9548 14016 9554 14068
rect 9950 14056 9956 14068
rect 9911 14028 9956 14056
rect 9950 14016 9956 14028
rect 10008 14016 10014 14068
rect 17865 14059 17923 14065
rect 17865 14025 17877 14059
rect 17911 14056 17923 14059
rect 17954 14056 17960 14068
rect 17911 14028 17960 14056
rect 17911 14025 17923 14028
rect 17865 14019 17923 14025
rect 17954 14016 17960 14028
rect 18012 14016 18018 14068
rect 27062 14016 27068 14068
rect 27120 14056 27126 14068
rect 28445 14059 28503 14065
rect 28445 14056 28457 14059
rect 27120 14028 28457 14056
rect 27120 14016 27126 14028
rect 28445 14025 28457 14028
rect 28491 14025 28503 14059
rect 28445 14019 28503 14025
rect 29917 14059 29975 14065
rect 29917 14025 29929 14059
rect 29963 14056 29975 14059
rect 30282 14056 30288 14068
rect 29963 14028 30288 14056
rect 29963 14025 29975 14028
rect 29917 14019 29975 14025
rect 30282 14016 30288 14028
rect 30340 14016 30346 14068
rect 30466 14016 30472 14068
rect 30524 14056 30530 14068
rect 30653 14059 30711 14065
rect 30653 14056 30665 14059
rect 30524 14028 30665 14056
rect 30524 14016 30530 14028
rect 30653 14025 30665 14028
rect 30699 14056 30711 14059
rect 31846 14056 31852 14068
rect 30699 14028 31852 14056
rect 30699 14025 30711 14028
rect 30653 14019 30711 14025
rect 31846 14016 31852 14028
rect 31904 14016 31910 14068
rect 32122 14056 32128 14068
rect 32083 14028 32128 14056
rect 32122 14016 32128 14028
rect 32180 14016 32186 14068
rect 32490 14016 32496 14068
rect 32548 14056 32554 14068
rect 33689 14059 33747 14065
rect 33689 14056 33701 14059
rect 32548 14028 33701 14056
rect 32548 14016 32554 14028
rect 33689 14025 33701 14028
rect 33735 14025 33747 14059
rect 33689 14019 33747 14025
rect 34606 14016 34612 14068
rect 34664 14056 34670 14068
rect 36725 14059 36783 14065
rect 36725 14056 36737 14059
rect 34664 14028 36737 14056
rect 34664 14016 34670 14028
rect 36725 14025 36737 14028
rect 36771 14025 36783 14059
rect 36725 14019 36783 14025
rect 5166 13988 5172 14000
rect 5127 13960 5172 13988
rect 5166 13948 5172 13960
rect 5224 13948 5230 14000
rect 4709 13923 4767 13929
rect 4709 13889 4721 13923
rect 4755 13920 4767 13923
rect 5810 13920 5816 13932
rect 4755 13892 5816 13920
rect 4755 13889 4767 13892
rect 4709 13883 4767 13889
rect 5810 13880 5816 13892
rect 5868 13920 5874 13932
rect 6546 13920 6552 13932
rect 5868 13892 6552 13920
rect 5868 13880 5874 13892
rect 6546 13880 6552 13892
rect 6604 13880 6610 13932
rect 7374 13920 7380 13932
rect 7335 13892 7380 13920
rect 7374 13880 7380 13892
rect 7432 13880 7438 13932
rect 7561 13923 7619 13929
rect 7561 13889 7573 13923
rect 7607 13920 7619 13923
rect 7742 13920 7748 13932
rect 7607 13892 7748 13920
rect 7607 13889 7619 13892
rect 7561 13883 7619 13889
rect 7742 13880 7748 13892
rect 7800 13880 7806 13932
rect 9968 13920 9996 14016
rect 10318 13948 10324 14000
rect 10376 13988 10382 14000
rect 11057 13991 11115 13997
rect 11057 13988 11069 13991
rect 10376 13960 11069 13988
rect 10376 13948 10382 13960
rect 10612 13929 10640 13960
rect 11057 13957 11069 13960
rect 11103 13957 11115 13991
rect 11057 13951 11115 13957
rect 25409 13991 25467 13997
rect 25409 13957 25421 13991
rect 25455 13988 25467 13991
rect 28074 13988 28080 14000
rect 25455 13960 26372 13988
rect 28035 13960 28080 13988
rect 25455 13957 25467 13960
rect 25409 13951 25467 13957
rect 26344 13932 26372 13960
rect 28074 13948 28080 13960
rect 28132 13948 28138 14000
rect 30190 13988 30196 14000
rect 30151 13960 30196 13988
rect 30190 13948 30196 13960
rect 30248 13948 30254 14000
rect 10505 13923 10563 13929
rect 10505 13920 10517 13923
rect 9968 13892 10517 13920
rect 10505 13889 10517 13892
rect 10551 13889 10563 13923
rect 10505 13883 10563 13889
rect 10597 13923 10655 13929
rect 10597 13889 10609 13923
rect 10643 13920 10655 13923
rect 18785 13923 18843 13929
rect 10643 13892 10677 13920
rect 10643 13889 10655 13892
rect 10597 13883 10655 13889
rect 18785 13889 18797 13923
rect 18831 13920 18843 13923
rect 18966 13920 18972 13932
rect 18831 13892 18972 13920
rect 18831 13889 18843 13892
rect 18785 13883 18843 13889
rect 18966 13880 18972 13892
rect 19024 13880 19030 13932
rect 19058 13880 19064 13932
rect 19116 13920 19122 13932
rect 19153 13923 19211 13929
rect 19153 13920 19165 13923
rect 19116 13892 19165 13920
rect 19116 13880 19122 13892
rect 19153 13889 19165 13892
rect 19199 13920 19211 13923
rect 23109 13923 23167 13929
rect 19199 13892 19840 13920
rect 19199 13889 19211 13892
rect 19153 13883 19211 13889
rect 5077 13855 5135 13861
rect 5077 13821 5089 13855
rect 5123 13852 5135 13855
rect 7392 13852 7420 13880
rect 7929 13855 7987 13861
rect 7929 13852 7941 13855
rect 5123 13824 5580 13852
rect 7392 13824 7941 13852
rect 5123 13821 5135 13824
rect 5077 13815 5135 13821
rect 5552 13784 5580 13824
rect 7929 13821 7941 13824
rect 7975 13821 7987 13855
rect 7929 13815 7987 13821
rect 8297 13855 8355 13861
rect 8297 13821 8309 13855
rect 8343 13821 8355 13855
rect 8297 13815 8355 13821
rect 5629 13787 5687 13793
rect 5629 13784 5641 13787
rect 5552 13756 5641 13784
rect 5629 13753 5641 13756
rect 5675 13784 5687 13787
rect 5994 13784 6000 13796
rect 5675 13756 6000 13784
rect 5675 13753 5687 13756
rect 5629 13747 5687 13753
rect 5994 13744 6000 13756
rect 6052 13784 6058 13796
rect 6822 13784 6828 13796
rect 6052 13756 6828 13784
rect 6052 13744 6058 13756
rect 6822 13744 6828 13756
rect 6880 13744 6886 13796
rect 7282 13784 7288 13796
rect 7243 13756 7288 13784
rect 7282 13744 7288 13756
rect 7340 13784 7346 13796
rect 8312 13784 8340 13815
rect 9490 13812 9496 13864
rect 9548 13852 9554 13864
rect 9548 13824 9628 13852
rect 9548 13812 9554 13824
rect 7340 13756 8340 13784
rect 9600 13784 9628 13824
rect 11054 13812 11060 13864
rect 11112 13852 11118 13864
rect 15746 13861 15752 13864
rect 11425 13855 11483 13861
rect 11425 13852 11437 13855
rect 11112 13824 11437 13852
rect 11112 13812 11118 13824
rect 11425 13821 11437 13824
rect 11471 13821 11483 13855
rect 15473 13855 15531 13861
rect 15473 13852 15485 13855
rect 11425 13815 11483 13821
rect 15304 13824 15485 13852
rect 10413 13787 10471 13793
rect 10413 13784 10425 13787
rect 9600 13756 10425 13784
rect 7340 13744 7346 13756
rect 10413 13753 10425 13756
rect 10459 13753 10471 13787
rect 10413 13747 10471 13753
rect 5534 13716 5540 13728
rect 5495 13688 5540 13716
rect 5534 13676 5540 13688
rect 5592 13676 5598 13728
rect 5718 13676 5724 13728
rect 5776 13716 5782 13728
rect 6181 13719 6239 13725
rect 6181 13716 6193 13719
rect 5776 13688 6193 13716
rect 5776 13676 5782 13688
rect 6181 13685 6193 13688
rect 6227 13685 6239 13719
rect 6181 13679 6239 13685
rect 6917 13719 6975 13725
rect 6917 13685 6929 13719
rect 6963 13716 6975 13719
rect 8202 13716 8208 13728
rect 6963 13688 8208 13716
rect 6963 13685 6975 13688
rect 6917 13679 6975 13685
rect 8202 13676 8208 13688
rect 8260 13676 8266 13728
rect 10042 13716 10048 13728
rect 10003 13688 10048 13716
rect 10042 13676 10048 13688
rect 10100 13676 10106 13728
rect 15194 13676 15200 13728
rect 15252 13716 15258 13728
rect 15304 13725 15332 13824
rect 15473 13821 15485 13824
rect 15519 13821 15531 13855
rect 15740 13852 15752 13861
rect 15707 13824 15752 13852
rect 15473 13815 15531 13821
rect 15740 13815 15752 13824
rect 15746 13812 15752 13815
rect 15804 13812 15810 13864
rect 17497 13855 17555 13861
rect 17497 13821 17509 13855
rect 17543 13852 17555 13855
rect 18046 13852 18052 13864
rect 17543 13824 18052 13852
rect 17543 13821 17555 13824
rect 17497 13815 17555 13821
rect 18046 13812 18052 13824
rect 18104 13812 18110 13864
rect 18598 13852 18604 13864
rect 18511 13824 18604 13852
rect 18598 13812 18604 13824
rect 18656 13852 18662 13864
rect 19242 13852 19248 13864
rect 18656 13824 19248 13852
rect 18656 13812 18662 13824
rect 19242 13812 19248 13824
rect 19300 13812 19306 13864
rect 19705 13855 19763 13861
rect 19705 13821 19717 13855
rect 19751 13821 19763 13855
rect 19812 13852 19840 13892
rect 23109 13889 23121 13923
rect 23155 13920 23167 13923
rect 25958 13920 25964 13932
rect 23155 13892 23796 13920
rect 25919 13892 25964 13920
rect 23155 13889 23167 13892
rect 23109 13883 23167 13889
rect 19972 13855 20030 13861
rect 19972 13852 19984 13855
rect 19812 13824 19984 13852
rect 19705 13815 19763 13821
rect 19972 13821 19984 13824
rect 20018 13852 20030 13855
rect 20530 13852 20536 13864
rect 20018 13824 20536 13852
rect 20018 13821 20030 13824
rect 19972 13815 20030 13821
rect 18509 13787 18567 13793
rect 18509 13753 18521 13787
rect 18555 13784 18567 13787
rect 19058 13784 19064 13796
rect 18555 13756 19064 13784
rect 18555 13753 18567 13756
rect 18509 13747 18567 13753
rect 19058 13744 19064 13756
rect 19116 13744 19122 13796
rect 15289 13719 15347 13725
rect 15289 13716 15301 13719
rect 15252 13688 15301 13716
rect 15252 13676 15258 13688
rect 15289 13685 15301 13688
rect 15335 13685 15347 13719
rect 15289 13679 15347 13685
rect 16853 13719 16911 13725
rect 16853 13685 16865 13719
rect 16899 13716 16911 13719
rect 16942 13716 16948 13728
rect 16899 13688 16948 13716
rect 16899 13685 16911 13688
rect 16853 13679 16911 13685
rect 16942 13676 16948 13688
rect 17000 13676 17006 13728
rect 18138 13716 18144 13728
rect 18099 13688 18144 13716
rect 18138 13676 18144 13688
rect 18196 13676 18202 13728
rect 19613 13719 19671 13725
rect 19613 13685 19625 13719
rect 19659 13716 19671 13719
rect 19720 13716 19748 13815
rect 20530 13812 20536 13824
rect 20588 13812 20594 13864
rect 23477 13855 23535 13861
rect 23477 13821 23489 13855
rect 23523 13852 23535 13855
rect 23566 13852 23572 13864
rect 23523 13824 23572 13852
rect 23523 13821 23535 13824
rect 23477 13815 23535 13821
rect 23566 13812 23572 13824
rect 23624 13812 23630 13864
rect 23661 13855 23719 13861
rect 23661 13821 23673 13855
rect 23707 13821 23719 13855
rect 23768 13852 23796 13892
rect 25958 13880 25964 13892
rect 26016 13880 26022 13932
rect 26326 13880 26332 13932
rect 26384 13920 26390 13932
rect 26697 13923 26755 13929
rect 26697 13920 26709 13923
rect 26384 13892 26709 13920
rect 26384 13880 26390 13892
rect 26697 13889 26709 13892
rect 26743 13889 26755 13923
rect 26697 13883 26755 13889
rect 26786 13880 26792 13932
rect 26844 13920 26850 13932
rect 27617 13923 27675 13929
rect 27617 13920 27629 13923
rect 26844 13892 27629 13920
rect 26844 13880 26850 13892
rect 27617 13889 27629 13892
rect 27663 13889 27675 13923
rect 32140 13920 32168 14016
rect 32309 13923 32367 13929
rect 32309 13920 32321 13923
rect 32140 13892 32321 13920
rect 27617 13883 27675 13889
rect 32309 13889 32321 13892
rect 32355 13889 32367 13923
rect 32309 13883 32367 13889
rect 23917 13855 23975 13861
rect 23917 13852 23929 13855
rect 23768 13824 23929 13852
rect 23661 13815 23719 13821
rect 23917 13821 23929 13824
rect 23963 13852 23975 13855
rect 25866 13852 25872 13864
rect 23963 13824 25872 13852
rect 23963 13821 23975 13824
rect 23917 13815 23975 13821
rect 23676 13784 23704 13815
rect 25866 13812 25872 13824
rect 25924 13812 25930 13864
rect 26602 13812 26608 13864
rect 26660 13852 26666 13864
rect 27525 13855 27583 13861
rect 27525 13852 27537 13855
rect 26660 13824 27537 13852
rect 26660 13812 26666 13824
rect 27525 13821 27537 13824
rect 27571 13852 27583 13855
rect 28813 13855 28871 13861
rect 28813 13852 28825 13855
rect 27571 13824 28825 13852
rect 27571 13821 27583 13824
rect 27525 13815 27583 13821
rect 28813 13821 28825 13824
rect 28859 13821 28871 13855
rect 32324 13852 32352 13883
rect 34422 13852 34428 13864
rect 32324 13824 34428 13852
rect 28813 13815 28871 13821
rect 34422 13812 34428 13824
rect 34480 13852 34486 13864
rect 34517 13855 34575 13861
rect 34517 13852 34529 13855
rect 34480 13824 34529 13852
rect 34480 13812 34486 13824
rect 34517 13821 34529 13824
rect 34563 13852 34575 13855
rect 35161 13855 35219 13861
rect 35161 13852 35173 13855
rect 34563 13824 35173 13852
rect 34563 13821 34575 13824
rect 34517 13815 34575 13821
rect 35161 13821 35173 13824
rect 35207 13852 35219 13855
rect 35345 13855 35403 13861
rect 35345 13852 35357 13855
rect 35207 13824 35357 13852
rect 35207 13821 35219 13824
rect 35161 13815 35219 13821
rect 35345 13821 35357 13824
rect 35391 13821 35403 13855
rect 35345 13815 35403 13821
rect 24210 13784 24216 13796
rect 23676 13756 24216 13784
rect 24210 13744 24216 13756
rect 24268 13744 24274 13796
rect 27433 13787 27491 13793
rect 25056 13756 25912 13784
rect 20898 13716 20904 13728
rect 19659 13688 20904 13716
rect 19659 13685 19671 13688
rect 19613 13679 19671 13685
rect 20898 13676 20904 13688
rect 20956 13676 20962 13728
rect 21082 13716 21088 13728
rect 21043 13688 21088 13716
rect 21082 13676 21088 13688
rect 21140 13676 21146 13728
rect 24302 13676 24308 13728
rect 24360 13716 24366 13728
rect 25056 13725 25084 13756
rect 25884 13728 25912 13756
rect 26620 13756 27200 13784
rect 25041 13719 25099 13725
rect 25041 13716 25053 13719
rect 24360 13688 25053 13716
rect 24360 13676 24366 13688
rect 25041 13685 25053 13688
rect 25087 13685 25099 13719
rect 25774 13716 25780 13728
rect 25735 13688 25780 13716
rect 25041 13679 25099 13685
rect 25774 13676 25780 13688
rect 25832 13676 25838 13728
rect 25866 13676 25872 13728
rect 25924 13716 25930 13728
rect 26234 13716 26240 13728
rect 25924 13688 25969 13716
rect 26195 13688 26240 13716
rect 25924 13676 25930 13688
rect 26234 13676 26240 13688
rect 26292 13676 26298 13728
rect 26510 13676 26516 13728
rect 26568 13716 26574 13728
rect 26620 13725 26648 13756
rect 26605 13719 26663 13725
rect 26605 13716 26617 13719
rect 26568 13688 26617 13716
rect 26568 13676 26574 13688
rect 26605 13685 26617 13688
rect 26651 13685 26663 13719
rect 27062 13716 27068 13728
rect 27023 13688 27068 13716
rect 26605 13679 26663 13685
rect 27062 13676 27068 13688
rect 27120 13676 27126 13728
rect 27172 13716 27200 13756
rect 27433 13753 27445 13787
rect 27479 13784 27491 13787
rect 27798 13784 27804 13796
rect 27479 13756 27804 13784
rect 27479 13753 27491 13756
rect 27433 13747 27491 13753
rect 27798 13744 27804 13756
rect 27856 13744 27862 13796
rect 32582 13793 32588 13796
rect 32576 13784 32588 13793
rect 32543 13756 32588 13784
rect 32576 13747 32588 13756
rect 32582 13744 32588 13747
rect 32640 13744 32646 13796
rect 35618 13793 35624 13796
rect 35612 13784 35624 13793
rect 35579 13756 35624 13784
rect 35612 13747 35624 13756
rect 35618 13744 35624 13747
rect 35676 13744 35682 13796
rect 27522 13716 27528 13728
rect 27172 13688 27528 13716
rect 27522 13676 27528 13688
rect 27580 13676 27586 13728
rect 1104 13626 38824 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 38824 13626
rect 1104 13552 38824 13574
rect 5261 13515 5319 13521
rect 5261 13481 5273 13515
rect 5307 13512 5319 13515
rect 5534 13512 5540 13524
rect 5307 13484 5540 13512
rect 5307 13481 5319 13484
rect 5261 13475 5319 13481
rect 5534 13472 5540 13484
rect 5592 13512 5598 13524
rect 7098 13512 7104 13524
rect 5592 13484 7104 13512
rect 5592 13472 5598 13484
rect 7098 13472 7104 13484
rect 7156 13512 7162 13524
rect 7653 13515 7711 13521
rect 7653 13512 7665 13515
rect 7156 13484 7665 13512
rect 7156 13472 7162 13484
rect 7653 13481 7665 13484
rect 7699 13481 7711 13515
rect 18046 13512 18052 13524
rect 18007 13484 18052 13512
rect 7653 13475 7711 13481
rect 18046 13472 18052 13484
rect 18104 13472 18110 13524
rect 18598 13512 18604 13524
rect 18559 13484 18604 13512
rect 18598 13472 18604 13484
rect 18656 13472 18662 13524
rect 19058 13512 19064 13524
rect 19019 13484 19064 13512
rect 19058 13472 19064 13484
rect 19116 13472 19122 13524
rect 25501 13515 25559 13521
rect 25501 13481 25513 13515
rect 25547 13512 25559 13515
rect 25866 13512 25872 13524
rect 25547 13484 25872 13512
rect 25547 13481 25559 13484
rect 25501 13475 25559 13481
rect 25866 13472 25872 13484
rect 25924 13472 25930 13524
rect 26237 13515 26295 13521
rect 26237 13481 26249 13515
rect 26283 13481 26295 13515
rect 26602 13512 26608 13524
rect 26563 13484 26608 13512
rect 26237 13475 26295 13481
rect 5994 13453 6000 13456
rect 5988 13444 6000 13453
rect 5955 13416 6000 13444
rect 5988 13407 6000 13416
rect 5994 13404 6000 13407
rect 6052 13404 6058 13456
rect 19705 13447 19763 13453
rect 19705 13413 19717 13447
rect 19751 13444 19763 13447
rect 20070 13444 20076 13456
rect 19751 13416 20076 13444
rect 19751 13413 19763 13416
rect 19705 13407 19763 13413
rect 20070 13404 20076 13416
rect 20128 13444 20134 13456
rect 21082 13444 21088 13456
rect 20128 13416 21088 13444
rect 20128 13404 20134 13416
rect 21082 13404 21088 13416
rect 21140 13453 21146 13456
rect 21140 13447 21204 13453
rect 21140 13413 21158 13447
rect 21192 13413 21204 13447
rect 24210 13444 24216 13456
rect 21140 13407 21204 13413
rect 23492 13416 24216 13444
rect 21140 13404 21146 13407
rect 8202 13376 8208 13388
rect 8163 13348 8208 13376
rect 8202 13336 8208 13348
rect 8260 13336 8266 13388
rect 9861 13379 9919 13385
rect 9861 13345 9873 13379
rect 9907 13376 9919 13379
rect 9950 13376 9956 13388
rect 9907 13348 9956 13376
rect 9907 13345 9919 13348
rect 9861 13339 9919 13345
rect 9950 13336 9956 13348
rect 10008 13336 10014 13388
rect 11698 13376 11704 13388
rect 11659 13348 11704 13376
rect 11698 13336 11704 13348
rect 11756 13336 11762 13388
rect 11793 13379 11851 13385
rect 11793 13345 11805 13379
rect 11839 13376 11851 13379
rect 12342 13376 12348 13388
rect 11839 13348 12348 13376
rect 11839 13345 11851 13348
rect 11793 13339 11851 13345
rect 12342 13336 12348 13348
rect 12400 13336 12406 13388
rect 16942 13385 16948 13388
rect 16485 13379 16543 13385
rect 16485 13345 16497 13379
rect 16531 13376 16543 13379
rect 16936 13376 16948 13385
rect 16531 13348 16948 13376
rect 16531 13345 16543 13348
rect 16485 13339 16543 13345
rect 16936 13339 16948 13348
rect 17000 13376 17006 13388
rect 17770 13376 17776 13388
rect 17000 13348 17776 13376
rect 16942 13336 16948 13339
rect 17000 13336 17006 13348
rect 17770 13336 17776 13348
rect 17828 13336 17834 13388
rect 19613 13379 19671 13385
rect 19613 13345 19625 13379
rect 19659 13376 19671 13379
rect 20622 13376 20628 13388
rect 19659 13348 20628 13376
rect 19659 13345 19671 13348
rect 19613 13339 19671 13345
rect 20622 13336 20628 13348
rect 20680 13336 20686 13388
rect 23492 13385 23520 13416
rect 24210 13404 24216 13416
rect 24268 13404 24274 13456
rect 26252 13444 26280 13475
rect 26602 13472 26608 13484
rect 26660 13472 26666 13524
rect 27709 13515 27767 13521
rect 27709 13481 27721 13515
rect 27755 13512 27767 13515
rect 27798 13512 27804 13524
rect 27755 13484 27804 13512
rect 27755 13481 27767 13484
rect 27709 13475 27767 13481
rect 27798 13472 27804 13484
rect 27856 13472 27862 13524
rect 32401 13515 32459 13521
rect 32401 13481 32413 13515
rect 32447 13512 32459 13515
rect 32582 13512 32588 13524
rect 32447 13484 32588 13512
rect 32447 13481 32459 13484
rect 32401 13475 32459 13481
rect 32582 13472 32588 13484
rect 32640 13512 32646 13524
rect 34057 13515 34115 13521
rect 34057 13512 34069 13515
rect 32640 13484 34069 13512
rect 32640 13472 32646 13484
rect 34057 13481 34069 13484
rect 34103 13481 34115 13515
rect 34606 13512 34612 13524
rect 34567 13484 34612 13512
rect 34057 13475 34115 13481
rect 34606 13472 34612 13484
rect 34664 13472 34670 13524
rect 35069 13515 35127 13521
rect 35069 13481 35081 13515
rect 35115 13512 35127 13515
rect 35618 13512 35624 13524
rect 35115 13484 35624 13512
rect 35115 13481 35127 13484
rect 35069 13475 35127 13481
rect 35618 13472 35624 13484
rect 35676 13512 35682 13524
rect 36541 13515 36599 13521
rect 36541 13512 36553 13515
rect 35676 13484 36553 13512
rect 35676 13472 35682 13484
rect 36541 13481 36553 13484
rect 36587 13481 36599 13515
rect 36541 13475 36599 13481
rect 26786 13444 26792 13456
rect 26252 13416 26792 13444
rect 26786 13404 26792 13416
rect 26844 13404 26850 13456
rect 32950 13453 32956 13456
rect 32944 13444 32956 13453
rect 32911 13416 32956 13444
rect 32944 13407 32956 13416
rect 32950 13404 32956 13407
rect 33008 13404 33014 13456
rect 35342 13404 35348 13456
rect 35400 13404 35406 13456
rect 23477 13379 23535 13385
rect 23477 13345 23489 13379
rect 23523 13345 23535 13379
rect 23477 13339 23535 13345
rect 23744 13379 23802 13385
rect 23744 13345 23756 13379
rect 23790 13376 23802 13379
rect 24302 13376 24308 13388
rect 23790 13348 24308 13376
rect 23790 13345 23802 13348
rect 23744 13339 23802 13345
rect 24302 13336 24308 13348
rect 24360 13336 24366 13388
rect 25866 13336 25872 13388
rect 25924 13376 25930 13388
rect 26053 13379 26111 13385
rect 26053 13376 26065 13379
rect 25924 13348 26065 13376
rect 25924 13336 25930 13348
rect 26053 13345 26065 13348
rect 26099 13345 26111 13379
rect 26970 13376 26976 13388
rect 26931 13348 26976 13376
rect 26053 13339 26111 13345
rect 26970 13336 26976 13348
rect 27028 13336 27034 13388
rect 28074 13376 28080 13388
rect 28035 13348 28080 13376
rect 28074 13336 28080 13348
rect 28132 13336 28138 13388
rect 29917 13379 29975 13385
rect 29917 13345 29929 13379
rect 29963 13376 29975 13379
rect 30558 13376 30564 13388
rect 29963 13348 30564 13376
rect 29963 13345 29975 13348
rect 29917 13339 29975 13345
rect 30558 13336 30564 13348
rect 30616 13336 30622 13388
rect 32122 13336 32128 13388
rect 32180 13376 32186 13388
rect 32677 13379 32735 13385
rect 32677 13376 32689 13379
rect 32180 13348 32689 13376
rect 32180 13336 32186 13348
rect 32677 13345 32689 13348
rect 32723 13345 32735 13379
rect 35360 13376 35388 13404
rect 35428 13379 35486 13385
rect 35428 13376 35440 13379
rect 35360 13348 35440 13376
rect 32677 13339 32735 13345
rect 35428 13345 35440 13348
rect 35474 13376 35486 13379
rect 36814 13376 36820 13388
rect 35474 13348 36820 13376
rect 35474 13345 35486 13348
rect 35428 13339 35486 13345
rect 36814 13336 36820 13348
rect 36872 13336 36878 13388
rect 5718 13308 5724 13320
rect 5679 13280 5724 13308
rect 5718 13268 5724 13280
rect 5776 13268 5782 13320
rect 11974 13308 11980 13320
rect 11935 13280 11980 13308
rect 11974 13268 11980 13280
rect 12032 13268 12038 13320
rect 15194 13268 15200 13320
rect 15252 13308 15258 13320
rect 16669 13311 16727 13317
rect 16669 13308 16681 13311
rect 15252 13280 16681 13308
rect 15252 13268 15258 13280
rect 16669 13277 16681 13280
rect 16715 13277 16727 13311
rect 16669 13271 16727 13277
rect 16025 13243 16083 13249
rect 16025 13240 16037 13243
rect 14476 13212 16037 13240
rect 14476 13184 14504 13212
rect 16025 13209 16037 13212
rect 16071 13240 16083 13243
rect 16298 13240 16304 13252
rect 16071 13212 16304 13240
rect 16071 13209 16083 13212
rect 16025 13203 16083 13209
rect 16298 13200 16304 13212
rect 16356 13240 16362 13252
rect 16574 13240 16580 13252
rect 16356 13212 16580 13240
rect 16356 13200 16362 13212
rect 16574 13200 16580 13212
rect 16632 13200 16638 13252
rect 7742 13132 7748 13184
rect 7800 13172 7806 13184
rect 8021 13175 8079 13181
rect 8021 13172 8033 13175
rect 7800 13144 8033 13172
rect 7800 13132 7806 13144
rect 8021 13141 8033 13144
rect 8067 13141 8079 13175
rect 8386 13172 8392 13184
rect 8347 13144 8392 13172
rect 8021 13135 8079 13141
rect 8386 13132 8392 13144
rect 8444 13132 8450 13184
rect 10045 13175 10103 13181
rect 10045 13141 10057 13175
rect 10091 13172 10103 13175
rect 10318 13172 10324 13184
rect 10091 13144 10324 13172
rect 10091 13141 10103 13144
rect 10045 13135 10103 13141
rect 10318 13132 10324 13144
rect 10376 13132 10382 13184
rect 10686 13172 10692 13184
rect 10647 13144 10692 13172
rect 10686 13132 10692 13144
rect 10744 13132 10750 13184
rect 11333 13175 11391 13181
rect 11333 13141 11345 13175
rect 11379 13172 11391 13175
rect 12250 13172 12256 13184
rect 11379 13144 12256 13172
rect 11379 13141 11391 13144
rect 11333 13135 11391 13141
rect 12250 13132 12256 13144
rect 12308 13132 12314 13184
rect 14001 13175 14059 13181
rect 14001 13141 14013 13175
rect 14047 13172 14059 13175
rect 14458 13172 14464 13184
rect 14047 13144 14464 13172
rect 14047 13141 14059 13144
rect 14001 13135 14059 13141
rect 14458 13132 14464 13144
rect 14516 13132 14522 13184
rect 15562 13172 15568 13184
rect 15523 13144 15568 13172
rect 15562 13132 15568 13144
rect 15620 13132 15626 13184
rect 16684 13172 16712 13271
rect 18966 13268 18972 13320
rect 19024 13308 19030 13320
rect 19886 13308 19892 13320
rect 19024 13280 19892 13308
rect 19024 13268 19030 13280
rect 19886 13268 19892 13280
rect 19944 13268 19950 13320
rect 20898 13308 20904 13320
rect 20859 13280 20904 13308
rect 20898 13268 20904 13280
rect 20956 13268 20962 13320
rect 26786 13268 26792 13320
rect 26844 13308 26850 13320
rect 27065 13311 27123 13317
rect 27065 13308 27077 13311
rect 26844 13280 27077 13308
rect 26844 13268 26850 13280
rect 27065 13277 27077 13280
rect 27111 13277 27123 13311
rect 27065 13271 27123 13277
rect 27157 13311 27215 13317
rect 27157 13277 27169 13311
rect 27203 13277 27215 13311
rect 28166 13308 28172 13320
rect 28127 13280 28172 13308
rect 27157 13271 27215 13277
rect 25958 13200 25964 13252
rect 26016 13240 26022 13252
rect 27172 13240 27200 13271
rect 28166 13268 28172 13280
rect 28224 13268 28230 13320
rect 28353 13311 28411 13317
rect 28353 13277 28365 13311
rect 28399 13308 28411 13311
rect 28721 13311 28779 13317
rect 28721 13308 28733 13311
rect 28399 13280 28733 13308
rect 28399 13277 28411 13280
rect 28353 13271 28411 13277
rect 28721 13277 28733 13280
rect 28767 13277 28779 13311
rect 28721 13271 28779 13277
rect 26016 13212 27200 13240
rect 26016 13200 26022 13212
rect 17862 13172 17868 13184
rect 16684 13144 17868 13172
rect 17862 13132 17868 13144
rect 17920 13132 17926 13184
rect 19242 13172 19248 13184
rect 19203 13144 19248 13172
rect 19242 13132 19248 13144
rect 19300 13132 19306 13184
rect 22278 13172 22284 13184
rect 22239 13144 22284 13172
rect 22278 13132 22284 13144
rect 22336 13132 22342 13184
rect 24854 13172 24860 13184
rect 24815 13144 24860 13172
rect 24854 13132 24860 13144
rect 24912 13172 24918 13184
rect 25774 13172 25780 13184
rect 24912 13144 25780 13172
rect 24912 13132 24918 13144
rect 25774 13132 25780 13144
rect 25832 13132 25838 13184
rect 27172 13172 27200 13212
rect 28258 13172 28264 13184
rect 27172 13144 28264 13172
rect 28258 13132 28264 13144
rect 28316 13172 28322 13184
rect 28368 13172 28396 13271
rect 34422 13268 34428 13320
rect 34480 13308 34486 13320
rect 35161 13311 35219 13317
rect 35161 13308 35173 13311
rect 34480 13280 35173 13308
rect 34480 13268 34486 13280
rect 35161 13277 35173 13280
rect 35207 13277 35219 13311
rect 35161 13271 35219 13277
rect 29362 13172 29368 13184
rect 28316 13144 28396 13172
rect 29323 13144 29368 13172
rect 28316 13132 28322 13144
rect 29362 13132 29368 13144
rect 29420 13132 29426 13184
rect 29638 13172 29644 13184
rect 29599 13144 29644 13172
rect 29638 13132 29644 13144
rect 29696 13132 29702 13184
rect 30101 13175 30159 13181
rect 30101 13141 30113 13175
rect 30147 13172 30159 13175
rect 30190 13172 30196 13184
rect 30147 13144 30196 13172
rect 30147 13141 30159 13144
rect 30101 13135 30159 13141
rect 30190 13132 30196 13144
rect 30248 13132 30254 13184
rect 30558 13172 30564 13184
rect 30519 13144 30564 13172
rect 30558 13132 30564 13144
rect 30616 13132 30622 13184
rect 1104 13082 38824 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 34966 13082
rect 35018 13030 35030 13082
rect 35082 13030 35094 13082
rect 35146 13030 35158 13082
rect 35210 13030 38824 13082
rect 1104 13008 38824 13030
rect 5994 12928 6000 12980
rect 6052 12968 6058 12980
rect 6089 12971 6147 12977
rect 6089 12968 6101 12971
rect 6052 12940 6101 12968
rect 6052 12928 6058 12940
rect 6089 12937 6101 12940
rect 6135 12937 6147 12971
rect 6089 12931 6147 12937
rect 8202 12928 8208 12980
rect 8260 12968 8266 12980
rect 8757 12971 8815 12977
rect 8757 12968 8769 12971
rect 8260 12940 8769 12968
rect 8260 12928 8266 12940
rect 8757 12937 8769 12940
rect 8803 12937 8815 12971
rect 8757 12931 8815 12937
rect 10042 12928 10048 12980
rect 10100 12968 10106 12980
rect 10413 12971 10471 12977
rect 10413 12968 10425 12971
rect 10100 12940 10425 12968
rect 10100 12928 10106 12940
rect 10413 12937 10425 12940
rect 10459 12937 10471 12971
rect 11698 12968 11704 12980
rect 11659 12940 11704 12968
rect 10413 12931 10471 12937
rect 7098 12773 7104 12776
rect 6825 12767 6883 12773
rect 6825 12764 6837 12767
rect 6748 12736 6837 12764
rect 6748 12640 6776 12736
rect 6825 12733 6837 12736
rect 6871 12733 6883 12767
rect 7092 12764 7104 12773
rect 7059 12736 7104 12764
rect 6825 12727 6883 12733
rect 7092 12727 7104 12736
rect 7098 12724 7104 12727
rect 7156 12724 7162 12776
rect 9309 12767 9367 12773
rect 9309 12733 9321 12767
rect 9355 12733 9367 12767
rect 9309 12727 9367 12733
rect 7834 12656 7840 12708
rect 7892 12696 7898 12708
rect 9125 12699 9183 12705
rect 9125 12696 9137 12699
rect 7892 12668 9137 12696
rect 7892 12656 7898 12668
rect 9125 12665 9137 12668
rect 9171 12696 9183 12699
rect 9324 12696 9352 12727
rect 9171 12668 9352 12696
rect 10428 12696 10456 12931
rect 11698 12928 11704 12940
rect 11756 12968 11762 12980
rect 12621 12971 12679 12977
rect 12621 12968 12633 12971
rect 11756 12940 12633 12968
rect 11756 12928 11762 12940
rect 12621 12937 12633 12940
rect 12667 12937 12679 12971
rect 17770 12968 17776 12980
rect 17731 12940 17776 12968
rect 12621 12931 12679 12937
rect 17770 12928 17776 12940
rect 17828 12928 17834 12980
rect 18138 12928 18144 12980
rect 18196 12968 18202 12980
rect 18417 12971 18475 12977
rect 18417 12968 18429 12971
rect 18196 12940 18429 12968
rect 18196 12928 18202 12940
rect 18417 12937 18429 12940
rect 18463 12968 18475 12971
rect 20070 12968 20076 12980
rect 18463 12940 19472 12968
rect 20031 12940 20076 12968
rect 18463 12937 18475 12940
rect 18417 12931 18475 12937
rect 17497 12903 17555 12909
rect 17497 12869 17509 12903
rect 17543 12900 17555 12903
rect 17862 12900 17868 12912
rect 17543 12872 17868 12900
rect 17543 12869 17555 12872
rect 17497 12863 17555 12869
rect 17862 12860 17868 12872
rect 17920 12860 17926 12912
rect 10778 12792 10784 12844
rect 10836 12832 10842 12844
rect 11238 12832 11244 12844
rect 10836 12804 11244 12832
rect 10836 12792 10842 12804
rect 11238 12792 11244 12804
rect 11296 12792 11302 12844
rect 14458 12832 14464 12844
rect 14419 12804 14464 12832
rect 14458 12792 14464 12804
rect 14516 12792 14522 12844
rect 19444 12841 19472 12940
rect 20070 12928 20076 12940
rect 20128 12928 20134 12980
rect 24302 12968 24308 12980
rect 24263 12940 24308 12968
rect 24302 12928 24308 12940
rect 24360 12928 24366 12980
rect 25038 12928 25044 12980
rect 25096 12968 25102 12980
rect 25133 12971 25191 12977
rect 25133 12968 25145 12971
rect 25096 12940 25145 12968
rect 25096 12928 25102 12940
rect 25133 12937 25145 12940
rect 25179 12968 25191 12971
rect 25406 12968 25412 12980
rect 25179 12940 25412 12968
rect 25179 12937 25191 12940
rect 25133 12931 25191 12937
rect 25406 12928 25412 12940
rect 25464 12928 25470 12980
rect 25501 12971 25559 12977
rect 25501 12937 25513 12971
rect 25547 12968 25559 12971
rect 25958 12968 25964 12980
rect 25547 12940 25964 12968
rect 25547 12937 25559 12940
rect 25501 12931 25559 12937
rect 25958 12928 25964 12940
rect 26016 12928 26022 12980
rect 27430 12968 27436 12980
rect 27391 12940 27436 12968
rect 27430 12928 27436 12940
rect 27488 12928 27494 12980
rect 28166 12928 28172 12980
rect 28224 12968 28230 12980
rect 28721 12971 28779 12977
rect 28721 12968 28733 12971
rect 28224 12940 28733 12968
rect 28224 12928 28230 12940
rect 28721 12937 28733 12940
rect 28767 12968 28779 12971
rect 28810 12968 28816 12980
rect 28767 12940 28816 12968
rect 28767 12937 28779 12940
rect 28721 12931 28779 12937
rect 28810 12928 28816 12940
rect 28868 12928 28874 12980
rect 30558 12928 30564 12980
rect 30616 12968 30622 12980
rect 31205 12971 31263 12977
rect 31205 12968 31217 12971
rect 30616 12940 31217 12968
rect 30616 12928 30622 12940
rect 31205 12937 31217 12940
rect 31251 12937 31263 12971
rect 31570 12968 31576 12980
rect 31531 12940 31576 12968
rect 31205 12931 31263 12937
rect 31570 12928 31576 12940
rect 31628 12928 31634 12980
rect 32122 12968 32128 12980
rect 32083 12940 32128 12968
rect 32122 12928 32128 12940
rect 32180 12928 32186 12980
rect 33594 12968 33600 12980
rect 33555 12940 33600 12968
rect 33594 12928 33600 12940
rect 33652 12928 33658 12980
rect 34422 12928 34428 12980
rect 34480 12968 34486 12980
rect 34609 12971 34667 12977
rect 34609 12968 34621 12971
rect 34480 12940 34621 12968
rect 34480 12928 34486 12940
rect 34609 12937 34621 12940
rect 34655 12968 34667 12971
rect 35161 12971 35219 12977
rect 35161 12968 35173 12971
rect 34655 12940 35173 12968
rect 34655 12937 34667 12940
rect 34609 12931 34667 12937
rect 35161 12937 35173 12940
rect 35207 12937 35219 12971
rect 36814 12968 36820 12980
rect 36775 12940 36820 12968
rect 35161 12931 35219 12937
rect 23474 12860 23480 12912
rect 23532 12900 23538 12912
rect 23937 12903 23995 12909
rect 23937 12900 23949 12903
rect 23532 12872 23949 12900
rect 23532 12860 23538 12872
rect 23937 12869 23949 12872
rect 23983 12900 23995 12903
rect 24210 12900 24216 12912
rect 23983 12872 24216 12900
rect 23983 12869 23995 12872
rect 23937 12863 23995 12869
rect 24210 12860 24216 12872
rect 24268 12860 24274 12912
rect 26970 12860 26976 12912
rect 27028 12900 27034 12912
rect 27890 12900 27896 12912
rect 27028 12872 27896 12900
rect 27028 12860 27034 12872
rect 27890 12860 27896 12872
rect 27948 12900 27954 12912
rect 28353 12903 28411 12909
rect 28353 12900 28365 12903
rect 27948 12872 28365 12900
rect 27948 12860 27954 12872
rect 28353 12869 28365 12872
rect 28399 12869 28411 12903
rect 28353 12863 28411 12869
rect 28994 12860 29000 12912
rect 29052 12900 29058 12912
rect 30285 12903 30343 12909
rect 30285 12900 30297 12903
rect 29052 12872 30297 12900
rect 29052 12860 29058 12872
rect 19429 12835 19487 12841
rect 19429 12801 19441 12835
rect 19475 12801 19487 12835
rect 19429 12795 19487 12801
rect 19518 12792 19524 12844
rect 19576 12832 19582 12844
rect 19576 12804 19621 12832
rect 19576 12792 19582 12804
rect 29362 12792 29368 12844
rect 29420 12832 29426 12844
rect 29730 12832 29736 12844
rect 29420 12804 29736 12832
rect 29420 12792 29426 12804
rect 29730 12792 29736 12804
rect 29788 12792 29794 12844
rect 29840 12841 29868 12872
rect 30285 12869 30297 12872
rect 30331 12900 30343 12903
rect 30374 12900 30380 12912
rect 30331 12872 30380 12900
rect 30331 12869 30343 12872
rect 30285 12863 30343 12869
rect 30374 12860 30380 12872
rect 30432 12860 30438 12912
rect 29825 12835 29883 12841
rect 29825 12801 29837 12835
rect 29871 12801 29883 12835
rect 32140 12832 32168 12928
rect 32217 12835 32275 12841
rect 32217 12832 32229 12835
rect 32140 12804 32229 12832
rect 29825 12795 29883 12801
rect 32217 12801 32229 12804
rect 32263 12801 32275 12835
rect 35176 12832 35204 12931
rect 36814 12928 36820 12940
rect 36872 12928 36878 12980
rect 35437 12835 35495 12841
rect 35437 12832 35449 12835
rect 35176 12804 35449 12832
rect 32217 12795 32275 12801
rect 35437 12801 35449 12804
rect 35483 12801 35495 12835
rect 35437 12795 35495 12801
rect 10686 12724 10692 12776
rect 10744 12764 10750 12776
rect 10965 12767 11023 12773
rect 10965 12764 10977 12767
rect 10744 12736 10977 12764
rect 10744 12724 10750 12736
rect 10965 12733 10977 12736
rect 11011 12733 11023 12767
rect 10965 12727 11023 12733
rect 12437 12767 12495 12773
rect 12437 12733 12449 12767
rect 12483 12764 12495 12767
rect 12989 12767 13047 12773
rect 12989 12764 13001 12767
rect 12483 12736 13001 12764
rect 12483 12733 12495 12736
rect 12437 12727 12495 12733
rect 12989 12733 13001 12736
rect 13035 12733 13047 12767
rect 12989 12727 13047 12733
rect 11057 12699 11115 12705
rect 11057 12696 11069 12699
rect 10428 12668 11069 12696
rect 9171 12665 9183 12668
rect 9125 12659 9183 12665
rect 11057 12665 11069 12668
rect 11103 12696 11115 12699
rect 12452 12696 12480 12727
rect 15194 12724 15200 12776
rect 15252 12764 15258 12776
rect 15473 12767 15531 12773
rect 15473 12764 15485 12767
rect 15252 12736 15485 12764
rect 15252 12724 15258 12736
rect 15473 12733 15485 12736
rect 15519 12733 15531 12767
rect 15473 12727 15531 12733
rect 19242 12724 19248 12776
rect 19300 12764 19306 12776
rect 19337 12767 19395 12773
rect 19337 12764 19349 12767
rect 19300 12736 19349 12764
rect 19300 12724 19306 12736
rect 19337 12733 19349 12736
rect 19383 12733 19395 12767
rect 19337 12727 19395 12733
rect 20533 12767 20591 12773
rect 20533 12733 20545 12767
rect 20579 12733 20591 12767
rect 20533 12727 20591 12733
rect 11103 12668 12480 12696
rect 13817 12699 13875 12705
rect 11103 12665 11115 12668
rect 11057 12659 11115 12665
rect 13817 12665 13829 12699
rect 13863 12696 13875 12699
rect 14369 12699 14427 12705
rect 14369 12696 14381 12699
rect 13863 12668 14381 12696
rect 13863 12665 13875 12668
rect 13817 12659 13875 12665
rect 14369 12665 14381 12668
rect 14415 12696 14427 12699
rect 15562 12696 15568 12708
rect 14415 12668 15568 12696
rect 14415 12665 14427 12668
rect 14369 12659 14427 12665
rect 15562 12656 15568 12668
rect 15620 12696 15626 12708
rect 15740 12699 15798 12705
rect 15740 12696 15752 12699
rect 15620 12668 15752 12696
rect 15620 12656 15626 12668
rect 15740 12665 15752 12668
rect 15786 12696 15798 12699
rect 16482 12696 16488 12708
rect 15786 12668 16488 12696
rect 15786 12665 15798 12668
rect 15740 12659 15798 12665
rect 16482 12656 16488 12668
rect 16540 12656 16546 12708
rect 18877 12699 18935 12705
rect 18877 12665 18889 12699
rect 18923 12696 18935 12699
rect 20070 12696 20076 12708
rect 18923 12668 20076 12696
rect 18923 12665 18935 12668
rect 18877 12659 18935 12665
rect 20070 12656 20076 12668
rect 20128 12656 20134 12708
rect 5718 12588 5724 12640
rect 5776 12628 5782 12640
rect 5813 12631 5871 12637
rect 5813 12628 5825 12631
rect 5776 12600 5825 12628
rect 5776 12588 5782 12600
rect 5813 12597 5825 12600
rect 5859 12628 5871 12631
rect 6641 12631 6699 12637
rect 6641 12628 6653 12631
rect 5859 12600 6653 12628
rect 5859 12597 5871 12600
rect 5813 12591 5871 12597
rect 6641 12597 6653 12600
rect 6687 12628 6699 12631
rect 6730 12628 6736 12640
rect 6687 12600 6736 12628
rect 6687 12597 6699 12600
rect 6641 12591 6699 12597
rect 6730 12588 6736 12600
rect 6788 12588 6794 12640
rect 6914 12588 6920 12640
rect 6972 12628 6978 12640
rect 8205 12631 8263 12637
rect 8205 12628 8217 12631
rect 6972 12600 8217 12628
rect 6972 12588 6978 12600
rect 8205 12597 8217 12600
rect 8251 12597 8263 12631
rect 8205 12591 8263 12597
rect 9493 12631 9551 12637
rect 9493 12597 9505 12631
rect 9539 12628 9551 12631
rect 9582 12628 9588 12640
rect 9539 12600 9588 12628
rect 9539 12597 9551 12600
rect 9493 12591 9551 12597
rect 9582 12588 9588 12600
rect 9640 12588 9646 12640
rect 9950 12628 9956 12640
rect 9911 12600 9956 12628
rect 9950 12588 9956 12600
rect 10008 12588 10014 12640
rect 10597 12631 10655 12637
rect 10597 12597 10609 12631
rect 10643 12628 10655 12631
rect 10962 12628 10968 12640
rect 10643 12600 10968 12628
rect 10643 12597 10655 12600
rect 10597 12591 10655 12597
rect 10962 12588 10968 12600
rect 11020 12588 11026 12640
rect 12069 12631 12127 12637
rect 12069 12597 12081 12631
rect 12115 12628 12127 12631
rect 12342 12628 12348 12640
rect 12115 12600 12348 12628
rect 12115 12597 12127 12600
rect 12069 12591 12127 12597
rect 12342 12588 12348 12600
rect 12400 12588 12406 12640
rect 13906 12628 13912 12640
rect 13867 12600 13912 12628
rect 13906 12588 13912 12600
rect 13964 12588 13970 12640
rect 14274 12628 14280 12640
rect 14235 12600 14280 12628
rect 14274 12588 14280 12600
rect 14332 12588 14338 12640
rect 15194 12588 15200 12640
rect 15252 12628 15258 12640
rect 15289 12631 15347 12637
rect 15289 12628 15301 12631
rect 15252 12600 15301 12628
rect 15252 12588 15258 12600
rect 15289 12597 15301 12600
rect 15335 12597 15347 12631
rect 16850 12628 16856 12640
rect 16811 12600 16856 12628
rect 15289 12591 15347 12597
rect 16850 12588 16856 12600
rect 16908 12588 16914 12640
rect 18966 12628 18972 12640
rect 18927 12600 18972 12628
rect 18966 12588 18972 12600
rect 19024 12588 19030 12640
rect 20441 12631 20499 12637
rect 20441 12597 20453 12631
rect 20487 12628 20499 12631
rect 20548 12628 20576 12727
rect 20622 12724 20628 12776
rect 20680 12764 20686 12776
rect 20800 12767 20858 12773
rect 20800 12764 20812 12767
rect 20680 12736 20812 12764
rect 20680 12724 20686 12736
rect 20800 12733 20812 12736
rect 20846 12764 20858 12767
rect 22278 12764 22284 12776
rect 20846 12736 22284 12764
rect 20846 12733 20858 12736
rect 20800 12727 20858 12733
rect 22278 12724 22284 12736
rect 22336 12724 22342 12776
rect 25406 12724 25412 12776
rect 25464 12764 25470 12776
rect 25961 12767 26019 12773
rect 25961 12764 25973 12767
rect 25464 12736 25973 12764
rect 25464 12724 25470 12736
rect 25961 12733 25973 12736
rect 26007 12733 26019 12767
rect 25961 12727 26019 12733
rect 26786 12724 26792 12776
rect 26844 12764 26850 12776
rect 27985 12767 28043 12773
rect 27985 12764 27997 12767
rect 26844 12736 27997 12764
rect 26844 12724 26850 12736
rect 27985 12733 27997 12736
rect 28031 12733 28043 12767
rect 29638 12764 29644 12776
rect 29599 12736 29644 12764
rect 27985 12727 28043 12733
rect 29638 12724 29644 12736
rect 29696 12724 29702 12776
rect 30837 12767 30895 12773
rect 30837 12733 30849 12767
rect 30883 12764 30895 12767
rect 31570 12764 31576 12776
rect 30883 12736 31576 12764
rect 30883 12733 30895 12736
rect 30837 12727 30895 12733
rect 31570 12724 31576 12736
rect 31628 12724 31634 12776
rect 34333 12767 34391 12773
rect 34333 12733 34345 12767
rect 34379 12764 34391 12767
rect 35342 12764 35348 12776
rect 34379 12736 35348 12764
rect 34379 12733 34391 12736
rect 34333 12727 34391 12733
rect 35342 12724 35348 12736
rect 35400 12724 35406 12776
rect 25866 12696 25872 12708
rect 25827 12668 25872 12696
rect 25866 12656 25872 12668
rect 25924 12656 25930 12708
rect 31021 12699 31079 12705
rect 31021 12665 31033 12699
rect 31067 12665 31079 12699
rect 31021 12659 31079 12665
rect 20898 12628 20904 12640
rect 20487 12600 20904 12628
rect 20487 12597 20499 12600
rect 20441 12591 20499 12597
rect 20898 12588 20904 12600
rect 20956 12588 20962 12640
rect 21910 12628 21916 12640
rect 21871 12600 21916 12628
rect 21910 12588 21916 12600
rect 21968 12588 21974 12640
rect 29270 12628 29276 12640
rect 29231 12600 29276 12628
rect 29270 12588 29276 12600
rect 29328 12588 29334 12640
rect 30374 12588 30380 12640
rect 30432 12628 30438 12640
rect 30653 12631 30711 12637
rect 30653 12628 30665 12631
rect 30432 12600 30665 12628
rect 30432 12588 30438 12600
rect 30653 12597 30665 12600
rect 30699 12628 30711 12631
rect 31036 12628 31064 12659
rect 32398 12656 32404 12708
rect 32456 12705 32462 12708
rect 35710 12705 35716 12708
rect 32456 12699 32520 12705
rect 32456 12665 32474 12699
rect 32508 12665 32520 12699
rect 32456 12659 32520 12665
rect 35704 12659 35716 12705
rect 35768 12696 35774 12708
rect 35768 12668 35804 12696
rect 32456 12656 32462 12659
rect 35710 12656 35716 12659
rect 35768 12656 35774 12668
rect 30699 12600 31064 12628
rect 30699 12597 30711 12600
rect 30653 12591 30711 12597
rect 1104 12538 38824 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 38824 12538
rect 1104 12464 38824 12486
rect 9677 12427 9735 12433
rect 9677 12393 9689 12427
rect 9723 12424 9735 12427
rect 9950 12424 9956 12436
rect 9723 12396 9956 12424
rect 9723 12393 9735 12396
rect 9677 12387 9735 12393
rect 9950 12384 9956 12396
rect 10008 12424 10014 12436
rect 10594 12424 10600 12436
rect 10008 12396 10600 12424
rect 10008 12384 10014 12396
rect 10594 12384 10600 12396
rect 10652 12384 10658 12436
rect 10778 12424 10784 12436
rect 10739 12396 10784 12424
rect 10778 12384 10784 12396
rect 10836 12384 10842 12436
rect 14001 12427 14059 12433
rect 14001 12393 14013 12427
rect 14047 12424 14059 12427
rect 14274 12424 14280 12436
rect 14047 12396 14280 12424
rect 14047 12393 14059 12396
rect 14001 12387 14059 12393
rect 14274 12384 14280 12396
rect 14332 12384 14338 12436
rect 16574 12384 16580 12436
rect 16632 12424 16638 12436
rect 16761 12427 16819 12433
rect 16761 12424 16773 12427
rect 16632 12396 16773 12424
rect 16632 12384 16638 12396
rect 16761 12393 16773 12396
rect 16807 12393 16819 12427
rect 18322 12424 18328 12436
rect 18283 12396 18328 12424
rect 16761 12387 16819 12393
rect 18322 12384 18328 12396
rect 18380 12384 18386 12436
rect 19334 12384 19340 12436
rect 19392 12424 19398 12436
rect 19613 12427 19671 12433
rect 19613 12424 19625 12427
rect 19392 12396 19625 12424
rect 19392 12384 19398 12396
rect 19613 12393 19625 12396
rect 19659 12393 19671 12427
rect 20622 12424 20628 12436
rect 20583 12396 20628 12424
rect 19613 12387 19671 12393
rect 20622 12384 20628 12396
rect 20680 12384 20686 12436
rect 25958 12384 25964 12436
rect 26016 12424 26022 12436
rect 26237 12427 26295 12433
rect 26237 12424 26249 12427
rect 26016 12396 26249 12424
rect 26016 12384 26022 12396
rect 26237 12393 26249 12396
rect 26283 12393 26295 12427
rect 27890 12424 27896 12436
rect 27851 12396 27896 12424
rect 26237 12387 26295 12393
rect 27890 12384 27896 12396
rect 27948 12384 27954 12436
rect 28074 12384 28080 12436
rect 28132 12424 28138 12436
rect 28445 12427 28503 12433
rect 28445 12424 28457 12427
rect 28132 12396 28457 12424
rect 28132 12384 28138 12396
rect 28445 12393 28457 12396
rect 28491 12393 28503 12427
rect 30374 12424 30380 12436
rect 30335 12396 30380 12424
rect 28445 12387 28503 12393
rect 6908 12359 6966 12365
rect 6908 12325 6920 12359
rect 6954 12356 6966 12359
rect 7006 12356 7012 12368
rect 6954 12328 7012 12356
rect 6954 12325 6966 12328
rect 6908 12319 6966 12325
rect 7006 12316 7012 12328
rect 7064 12316 7070 12368
rect 8386 12316 8392 12368
rect 8444 12356 8450 12368
rect 10137 12359 10195 12365
rect 10137 12356 10149 12359
rect 8444 12328 10149 12356
rect 8444 12316 8450 12328
rect 10137 12325 10149 12328
rect 10183 12325 10195 12359
rect 10137 12319 10195 12325
rect 6641 12291 6699 12297
rect 6641 12257 6653 12291
rect 6687 12288 6699 12291
rect 6730 12288 6736 12300
rect 6687 12260 6736 12288
rect 6687 12257 6699 12260
rect 6641 12251 6699 12257
rect 6730 12248 6736 12260
rect 6788 12248 6794 12300
rect 9674 12248 9680 12300
rect 9732 12288 9738 12300
rect 10042 12288 10048 12300
rect 9732 12260 10048 12288
rect 9732 12248 9738 12260
rect 10042 12248 10048 12260
rect 10100 12248 10106 12300
rect 11425 12291 11483 12297
rect 11425 12257 11437 12291
rect 11471 12288 11483 12291
rect 11793 12291 11851 12297
rect 11793 12288 11805 12291
rect 11471 12260 11805 12288
rect 11471 12257 11483 12260
rect 11425 12251 11483 12257
rect 11793 12257 11805 12260
rect 11839 12288 11851 12291
rect 11974 12288 11980 12300
rect 11839 12260 11980 12288
rect 11839 12257 11851 12260
rect 11793 12251 11851 12257
rect 11974 12248 11980 12260
rect 12032 12288 12038 12300
rect 12152 12291 12210 12297
rect 12152 12288 12164 12291
rect 12032 12260 12164 12288
rect 12032 12248 12038 12260
rect 12152 12257 12164 12260
rect 12198 12288 12210 12291
rect 12434 12288 12440 12300
rect 12198 12260 12440 12288
rect 12198 12257 12210 12260
rect 12152 12251 12210 12257
rect 12434 12248 12440 12260
rect 12492 12248 12498 12300
rect 14826 12248 14832 12300
rect 14884 12288 14890 12300
rect 15637 12291 15695 12297
rect 15637 12288 15649 12291
rect 14884 12260 15649 12288
rect 14884 12248 14890 12260
rect 15637 12257 15649 12260
rect 15683 12288 15695 12291
rect 16206 12288 16212 12300
rect 15683 12260 16212 12288
rect 15683 12257 15695 12260
rect 15637 12251 15695 12257
rect 16206 12248 16212 12260
rect 16264 12248 16270 12300
rect 18230 12288 18236 12300
rect 18191 12260 18236 12288
rect 18230 12248 18236 12260
rect 18288 12248 18294 12300
rect 19337 12291 19395 12297
rect 19337 12257 19349 12291
rect 19383 12288 19395 12291
rect 20640 12288 20668 12384
rect 26786 12365 26792 12368
rect 26780 12356 26792 12365
rect 26747 12328 26792 12356
rect 26780 12319 26792 12328
rect 26786 12316 26792 12319
rect 26844 12316 26850 12368
rect 28460 12356 28488 12387
rect 30374 12384 30380 12396
rect 30432 12384 30438 12436
rect 32398 12424 32404 12436
rect 32359 12396 32404 12424
rect 32398 12384 32404 12396
rect 32456 12384 32462 12436
rect 32950 12384 32956 12436
rect 33008 12424 33014 12436
rect 33137 12427 33195 12433
rect 33137 12424 33149 12427
rect 33008 12396 33149 12424
rect 33008 12384 33014 12396
rect 33137 12393 33149 12396
rect 33183 12393 33195 12427
rect 35250 12424 35256 12436
rect 35211 12396 35256 12424
rect 33137 12387 33195 12393
rect 35250 12384 35256 12396
rect 35308 12384 35314 12436
rect 35342 12384 35348 12436
rect 35400 12424 35406 12436
rect 35621 12427 35679 12433
rect 35621 12424 35633 12427
rect 35400 12396 35633 12424
rect 35400 12384 35406 12396
rect 35621 12393 35633 12396
rect 35667 12393 35679 12427
rect 35621 12387 35679 12393
rect 29086 12356 29092 12368
rect 28460 12328 29092 12356
rect 29086 12316 29092 12328
rect 29144 12356 29150 12368
rect 29242 12359 29300 12365
rect 29242 12356 29254 12359
rect 29144 12328 29254 12356
rect 29144 12316 29150 12328
rect 29242 12325 29254 12328
rect 29288 12325 29300 12359
rect 29242 12319 29300 12325
rect 32122 12316 32128 12368
rect 32180 12356 32186 12368
rect 32677 12359 32735 12365
rect 32677 12356 32689 12359
rect 32180 12328 32689 12356
rect 32180 12316 32186 12328
rect 32677 12325 32689 12328
rect 32723 12325 32735 12359
rect 32677 12319 32735 12325
rect 19383 12260 20668 12288
rect 19383 12257 19395 12260
rect 19337 12251 19395 12257
rect 23658 12248 23664 12300
rect 23716 12288 23722 12300
rect 24009 12291 24067 12297
rect 24009 12288 24021 12291
rect 23716 12260 24021 12288
rect 23716 12248 23722 12260
rect 24009 12257 24021 12260
rect 24055 12288 24067 12291
rect 24762 12288 24768 12300
rect 24055 12260 24768 12288
rect 24055 12257 24067 12260
rect 24009 12251 24067 12257
rect 24762 12248 24768 12260
rect 24820 12248 24826 12300
rect 28994 12248 29000 12300
rect 29052 12288 29058 12300
rect 32140 12288 32168 12316
rect 29052 12260 32168 12288
rect 29052 12248 29058 12260
rect 10318 12220 10324 12232
rect 10231 12192 10324 12220
rect 10318 12180 10324 12192
rect 10376 12220 10382 12232
rect 11238 12220 11244 12232
rect 10376 12192 11244 12220
rect 10376 12180 10382 12192
rect 11238 12180 11244 12192
rect 11296 12180 11302 12232
rect 11330 12180 11336 12232
rect 11388 12220 11394 12232
rect 11882 12220 11888 12232
rect 11388 12192 11888 12220
rect 11388 12180 11394 12192
rect 11882 12180 11888 12192
rect 11940 12180 11946 12232
rect 15194 12180 15200 12232
rect 15252 12220 15258 12232
rect 15381 12223 15439 12229
rect 15381 12220 15393 12223
rect 15252 12192 15393 12220
rect 15252 12180 15258 12192
rect 15381 12189 15393 12192
rect 15427 12189 15439 12223
rect 15381 12183 15439 12189
rect 18138 12180 18144 12232
rect 18196 12220 18202 12232
rect 18417 12223 18475 12229
rect 18417 12220 18429 12223
rect 18196 12192 18429 12220
rect 18196 12180 18202 12192
rect 18417 12189 18429 12192
rect 18463 12220 18475 12223
rect 18877 12223 18935 12229
rect 18877 12220 18889 12223
rect 18463 12192 18889 12220
rect 18463 12189 18475 12192
rect 18417 12183 18475 12189
rect 18877 12189 18889 12192
rect 18923 12220 18935 12223
rect 19426 12220 19432 12232
rect 18923 12192 19432 12220
rect 18923 12189 18935 12192
rect 18877 12183 18935 12189
rect 19426 12180 19432 12192
rect 19484 12180 19490 12232
rect 23474 12180 23480 12232
rect 23532 12220 23538 12232
rect 23753 12223 23811 12229
rect 23753 12220 23765 12223
rect 23532 12192 23765 12220
rect 23532 12180 23538 12192
rect 23753 12189 23765 12192
rect 23799 12189 23811 12223
rect 23753 12183 23811 12189
rect 25682 12180 25688 12232
rect 25740 12220 25746 12232
rect 26513 12223 26571 12229
rect 26513 12220 26525 12223
rect 25740 12192 26525 12220
rect 25740 12180 25746 12192
rect 26513 12189 26525 12192
rect 26559 12189 26571 12223
rect 35710 12220 35716 12232
rect 35623 12192 35716 12220
rect 26513 12183 26571 12189
rect 35710 12180 35716 12192
rect 35768 12180 35774 12232
rect 35897 12223 35955 12229
rect 35897 12189 35909 12223
rect 35943 12220 35955 12223
rect 35986 12220 35992 12232
rect 35943 12192 35992 12220
rect 35943 12189 35955 12192
rect 35897 12183 35955 12189
rect 35986 12180 35992 12192
rect 36044 12180 36050 12232
rect 35728 12152 35756 12180
rect 35728 12124 36400 12152
rect 8018 12084 8024 12096
rect 7979 12056 8024 12084
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 13262 12084 13268 12096
rect 13223 12056 13268 12084
rect 13262 12044 13268 12056
rect 13320 12044 13326 12096
rect 17862 12084 17868 12096
rect 17823 12056 17868 12084
rect 17862 12044 17868 12056
rect 17920 12044 17926 12096
rect 19886 12044 19892 12096
rect 19944 12084 19950 12096
rect 19981 12087 20039 12093
rect 19981 12084 19993 12087
rect 19944 12056 19993 12084
rect 19944 12044 19950 12056
rect 19981 12053 19993 12056
rect 20027 12053 20039 12087
rect 19981 12047 20039 12053
rect 20898 12044 20904 12096
rect 20956 12084 20962 12096
rect 21085 12087 21143 12093
rect 21085 12084 21097 12087
rect 20956 12056 21097 12084
rect 20956 12044 20962 12056
rect 21085 12053 21097 12056
rect 21131 12053 21143 12087
rect 25130 12084 25136 12096
rect 25091 12056 25136 12084
rect 21085 12047 21143 12053
rect 25130 12044 25136 12056
rect 25188 12044 25194 12096
rect 25314 12044 25320 12096
rect 25372 12084 25378 12096
rect 25685 12087 25743 12093
rect 25685 12084 25697 12087
rect 25372 12056 25697 12084
rect 25372 12044 25378 12056
rect 25685 12053 25697 12056
rect 25731 12053 25743 12087
rect 28810 12084 28816 12096
rect 28771 12056 28816 12084
rect 25685 12047 25743 12053
rect 28810 12044 28816 12056
rect 28868 12044 28874 12096
rect 36372 12093 36400 12124
rect 36357 12087 36415 12093
rect 36357 12053 36369 12087
rect 36403 12084 36415 12087
rect 36814 12084 36820 12096
rect 36403 12056 36820 12084
rect 36403 12053 36415 12056
rect 36357 12047 36415 12053
rect 36814 12044 36820 12056
rect 36872 12044 36878 12096
rect 1104 11994 38824 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 34966 11994
rect 35018 11942 35030 11994
rect 35082 11942 35094 11994
rect 35146 11942 35158 11994
rect 35210 11942 38824 11994
rect 1104 11920 38824 11942
rect 5905 11883 5963 11889
rect 5905 11849 5917 11883
rect 5951 11880 5963 11883
rect 7006 11880 7012 11892
rect 5951 11852 7012 11880
rect 5951 11849 5963 11852
rect 5905 11843 5963 11849
rect 7006 11840 7012 11852
rect 7064 11880 7070 11892
rect 8205 11883 8263 11889
rect 8205 11880 8217 11883
rect 7064 11852 8217 11880
rect 7064 11840 7070 11852
rect 8205 11849 8217 11852
rect 8251 11849 8263 11883
rect 8205 11843 8263 11849
rect 8386 11840 8392 11892
rect 8444 11880 8450 11892
rect 8757 11883 8815 11889
rect 8757 11880 8769 11883
rect 8444 11852 8769 11880
rect 8444 11840 8450 11852
rect 8757 11849 8769 11852
rect 8803 11849 8815 11883
rect 11238 11880 11244 11892
rect 11199 11852 11244 11880
rect 8757 11843 8815 11849
rect 11238 11840 11244 11852
rect 11296 11840 11302 11892
rect 11882 11880 11888 11892
rect 11843 11852 11888 11880
rect 11882 11840 11888 11852
rect 11940 11880 11946 11892
rect 12161 11883 12219 11889
rect 12161 11880 12173 11883
rect 11940 11852 12173 11880
rect 11940 11840 11946 11852
rect 12161 11849 12173 11852
rect 12207 11849 12219 11883
rect 14826 11880 14832 11892
rect 14787 11852 14832 11880
rect 12161 11843 12219 11849
rect 12176 11744 12204 11843
rect 14826 11840 14832 11852
rect 14884 11840 14890 11892
rect 16574 11840 16580 11892
rect 16632 11880 16638 11892
rect 17773 11883 17831 11889
rect 17773 11880 17785 11883
rect 16632 11852 17785 11880
rect 16632 11840 16638 11852
rect 17773 11849 17785 11852
rect 17819 11880 17831 11883
rect 18230 11880 18236 11892
rect 17819 11852 18236 11880
rect 17819 11849 17831 11852
rect 17773 11843 17831 11849
rect 18230 11840 18236 11852
rect 18288 11840 18294 11892
rect 18322 11840 18328 11892
rect 18380 11880 18386 11892
rect 18601 11883 18659 11889
rect 18601 11880 18613 11883
rect 18380 11852 18613 11880
rect 18380 11840 18386 11852
rect 18601 11849 18613 11852
rect 18647 11849 18659 11883
rect 18601 11843 18659 11849
rect 20898 11840 20904 11892
rect 20956 11880 20962 11892
rect 23474 11880 23480 11892
rect 20956 11852 23480 11880
rect 20956 11840 20962 11852
rect 23474 11840 23480 11852
rect 23532 11840 23538 11892
rect 25314 11880 25320 11892
rect 25275 11852 25320 11880
rect 25314 11840 25320 11852
rect 25372 11840 25378 11892
rect 26786 11840 26792 11892
rect 26844 11880 26850 11892
rect 27065 11883 27123 11889
rect 27065 11880 27077 11883
rect 26844 11852 27077 11880
rect 26844 11840 26850 11852
rect 27065 11849 27077 11852
rect 27111 11880 27123 11883
rect 27617 11883 27675 11889
rect 27617 11880 27629 11883
rect 27111 11852 27629 11880
rect 27111 11849 27123 11852
rect 27065 11843 27123 11849
rect 27617 11849 27629 11852
rect 27663 11849 27675 11883
rect 28258 11880 28264 11892
rect 28219 11852 28264 11880
rect 27617 11843 27675 11849
rect 28258 11840 28264 11852
rect 28316 11840 28322 11892
rect 28718 11880 28724 11892
rect 28679 11852 28724 11880
rect 28718 11840 28724 11852
rect 28776 11840 28782 11892
rect 28994 11840 29000 11892
rect 29052 11880 29058 11892
rect 29052 11852 29097 11880
rect 29052 11840 29058 11852
rect 35342 11840 35348 11892
rect 35400 11880 35406 11892
rect 35621 11883 35679 11889
rect 35621 11880 35633 11883
rect 35400 11852 35633 11880
rect 35400 11840 35406 11852
rect 35621 11849 35633 11852
rect 35667 11849 35679 11883
rect 35986 11880 35992 11892
rect 35947 11852 35992 11880
rect 35621 11843 35679 11849
rect 35986 11840 35992 11852
rect 36044 11840 36050 11892
rect 16298 11772 16304 11824
rect 16356 11812 16362 11824
rect 16356 11784 16528 11812
rect 16356 11772 16362 11784
rect 16500 11753 16528 11784
rect 12437 11747 12495 11753
rect 12437 11744 12449 11747
rect 12176 11716 12449 11744
rect 12437 11713 12449 11716
rect 12483 11713 12495 11747
rect 12437 11707 12495 11713
rect 16485 11747 16543 11753
rect 16485 11713 16497 11747
rect 16531 11744 16543 11747
rect 16666 11744 16672 11756
rect 16531 11716 16672 11744
rect 16531 11713 16543 11716
rect 16485 11707 16543 11713
rect 16666 11704 16672 11716
rect 16724 11744 16730 11756
rect 17313 11747 17371 11753
rect 17313 11744 17325 11747
rect 16724 11716 17325 11744
rect 16724 11704 16730 11716
rect 17313 11713 17325 11716
rect 17359 11713 17371 11747
rect 20901 11747 20959 11753
rect 20901 11744 20913 11747
rect 17313 11707 17371 11713
rect 19904 11716 20913 11744
rect 6549 11679 6607 11685
rect 6549 11645 6561 11679
rect 6595 11676 6607 11679
rect 6822 11676 6828 11688
rect 6595 11648 6828 11676
rect 6595 11645 6607 11648
rect 6549 11639 6607 11645
rect 6822 11636 6828 11648
rect 6880 11636 6886 11688
rect 7926 11636 7932 11688
rect 7984 11676 7990 11688
rect 9217 11679 9275 11685
rect 9217 11676 9229 11679
rect 7984 11648 9229 11676
rect 7984 11636 7990 11648
rect 9217 11645 9229 11648
rect 9263 11676 9275 11679
rect 9309 11679 9367 11685
rect 9309 11676 9321 11679
rect 9263 11648 9321 11676
rect 9263 11645 9275 11648
rect 9217 11639 9275 11645
rect 9309 11645 9321 11648
rect 9355 11645 9367 11679
rect 9309 11639 9367 11645
rect 13814 11636 13820 11688
rect 13872 11676 13878 11688
rect 14921 11679 14979 11685
rect 14921 11676 14933 11679
rect 13872 11648 14933 11676
rect 13872 11636 13878 11648
rect 14921 11645 14933 11648
rect 14967 11645 14979 11679
rect 14921 11639 14979 11645
rect 16206 11636 16212 11688
rect 16264 11676 16270 11688
rect 16301 11679 16359 11685
rect 16301 11676 16313 11679
rect 16264 11648 16313 11676
rect 16264 11636 16270 11648
rect 16301 11645 16313 11648
rect 16347 11676 16359 11679
rect 16347 11648 16896 11676
rect 16347 11645 16359 11648
rect 16301 11639 16359 11645
rect 6273 11611 6331 11617
rect 6273 11577 6285 11611
rect 6319 11608 6331 11611
rect 6638 11608 6644 11620
rect 6319 11580 6644 11608
rect 6319 11577 6331 11580
rect 6273 11571 6331 11577
rect 6638 11568 6644 11580
rect 6696 11608 6702 11620
rect 6914 11608 6920 11620
rect 6696 11580 6920 11608
rect 6696 11568 6702 11580
rect 6914 11568 6920 11580
rect 6972 11608 6978 11620
rect 7070 11611 7128 11617
rect 7070 11608 7082 11611
rect 6972 11580 7082 11608
rect 6972 11568 6978 11580
rect 7070 11577 7082 11580
rect 7116 11577 7128 11611
rect 7070 11571 7128 11577
rect 9398 11568 9404 11620
rect 9456 11608 9462 11620
rect 9554 11611 9612 11617
rect 9554 11608 9566 11611
rect 9456 11580 9566 11608
rect 9456 11568 9462 11580
rect 9554 11577 9566 11580
rect 9600 11577 9612 11611
rect 9554 11571 9612 11577
rect 12704 11611 12762 11617
rect 12704 11577 12716 11611
rect 12750 11608 12762 11611
rect 13262 11608 13268 11620
rect 12750 11580 13268 11608
rect 12750 11577 12762 11580
rect 12704 11571 12762 11577
rect 13262 11568 13268 11580
rect 13320 11568 13326 11620
rect 16393 11611 16451 11617
rect 16393 11608 16405 11611
rect 15764 11580 16405 11608
rect 15764 11552 15792 11580
rect 16393 11577 16405 11580
rect 16439 11577 16451 11611
rect 16393 11571 16451 11577
rect 16868 11552 16896 11648
rect 17862 11636 17868 11688
rect 17920 11676 17926 11688
rect 18049 11679 18107 11685
rect 18049 11676 18061 11679
rect 17920 11648 18061 11676
rect 17920 11636 17926 11648
rect 18049 11645 18061 11648
rect 18095 11645 18107 11679
rect 18049 11639 18107 11645
rect 19904 11620 19932 11716
rect 20901 11713 20913 11716
rect 20947 11713 20959 11747
rect 25332 11744 25360 11840
rect 29012 11744 29040 11840
rect 29273 11747 29331 11753
rect 29273 11744 29285 11747
rect 25332 11716 25820 11744
rect 29012 11716 29285 11744
rect 20901 11707 20959 11713
rect 20254 11676 20260 11688
rect 20167 11648 20260 11676
rect 20254 11636 20260 11648
rect 20312 11676 20318 11688
rect 20809 11679 20867 11685
rect 20809 11676 20821 11679
rect 20312 11648 20821 11676
rect 20312 11636 20318 11648
rect 20809 11645 20821 11648
rect 20855 11676 20867 11679
rect 21174 11676 21180 11688
rect 20855 11648 21180 11676
rect 20855 11645 20867 11648
rect 20809 11639 20867 11645
rect 21174 11636 21180 11648
rect 21232 11676 21238 11688
rect 21910 11676 21916 11688
rect 21232 11648 21916 11676
rect 21232 11636 21238 11648
rect 21910 11636 21916 11648
rect 21968 11636 21974 11688
rect 23474 11676 23480 11688
rect 23435 11648 23480 11676
rect 23474 11636 23480 11648
rect 23532 11676 23538 11688
rect 23944 11679 24002 11685
rect 23944 11676 23956 11679
rect 23532 11648 23956 11676
rect 23532 11636 23538 11648
rect 23944 11645 23956 11648
rect 23990 11645 24002 11679
rect 25682 11676 25688 11688
rect 25643 11648 25688 11676
rect 23944 11639 24002 11645
rect 25682 11636 25688 11648
rect 25740 11636 25746 11688
rect 25792 11676 25820 11716
rect 29273 11713 29285 11716
rect 29319 11713 29331 11747
rect 29273 11707 29331 11713
rect 35345 11747 35403 11753
rect 35345 11713 35357 11747
rect 35391 11744 35403 11747
rect 35710 11744 35716 11756
rect 35391 11716 35716 11744
rect 35391 11713 35403 11716
rect 35345 11707 35403 11713
rect 35710 11704 35716 11716
rect 35768 11704 35774 11756
rect 25941 11679 25999 11685
rect 25941 11676 25953 11679
rect 25792 11648 25953 11676
rect 25941 11645 25953 11648
rect 25987 11645 25999 11679
rect 25941 11639 25999 11645
rect 28077 11679 28135 11685
rect 28077 11645 28089 11679
rect 28123 11676 28135 11679
rect 28718 11676 28724 11688
rect 28123 11648 28724 11676
rect 28123 11645 28135 11648
rect 28077 11639 28135 11645
rect 28718 11636 28724 11648
rect 28776 11636 28782 11688
rect 19886 11608 19892 11620
rect 19847 11580 19892 11608
rect 19886 11568 19892 11580
rect 19944 11568 19950 11620
rect 23109 11611 23167 11617
rect 23109 11577 23121 11611
rect 23155 11608 23167 11611
rect 24204 11611 24262 11617
rect 24204 11608 24216 11611
rect 23155 11580 24216 11608
rect 23155 11577 23167 11580
rect 23109 11571 23167 11577
rect 24204 11577 24216 11580
rect 24250 11608 24262 11611
rect 25130 11608 25136 11620
rect 24250 11580 25136 11608
rect 24250 11577 24262 11580
rect 24204 11571 24262 11577
rect 25130 11568 25136 11580
rect 25188 11568 25194 11620
rect 28810 11568 28816 11620
rect 28868 11608 28874 11620
rect 29518 11611 29576 11617
rect 29518 11608 29530 11611
rect 28868 11580 29530 11608
rect 28868 11568 28874 11580
rect 29518 11577 29530 11580
rect 29564 11577 29576 11611
rect 29518 11571 29576 11577
rect 10686 11540 10692 11552
rect 10647 11512 10692 11540
rect 10686 11500 10692 11512
rect 10744 11500 10750 11552
rect 13817 11543 13875 11549
rect 13817 11509 13829 11543
rect 13863 11540 13875 11543
rect 13906 11540 13912 11552
rect 13863 11512 13912 11540
rect 13863 11509 13875 11512
rect 13817 11503 13875 11509
rect 13906 11500 13912 11512
rect 13964 11500 13970 11552
rect 15194 11500 15200 11552
rect 15252 11540 15258 11552
rect 15381 11543 15439 11549
rect 15381 11540 15393 11543
rect 15252 11512 15393 11540
rect 15252 11500 15258 11512
rect 15381 11509 15393 11512
rect 15427 11509 15439 11543
rect 15746 11540 15752 11552
rect 15707 11512 15752 11540
rect 15381 11503 15439 11509
rect 15746 11500 15752 11512
rect 15804 11500 15810 11552
rect 15930 11540 15936 11552
rect 15891 11512 15936 11540
rect 15930 11500 15936 11512
rect 15988 11500 15994 11552
rect 16850 11500 16856 11552
rect 16908 11540 16914 11552
rect 16945 11543 17003 11549
rect 16945 11540 16957 11543
rect 16908 11512 16957 11540
rect 16908 11500 16914 11512
rect 16945 11509 16957 11512
rect 16991 11509 17003 11543
rect 18230 11540 18236 11552
rect 18191 11512 18236 11540
rect 16945 11503 17003 11509
rect 18230 11500 18236 11512
rect 18288 11500 18294 11552
rect 20346 11540 20352 11552
rect 20307 11512 20352 11540
rect 20346 11500 20352 11512
rect 20404 11500 20410 11552
rect 20438 11500 20444 11552
rect 20496 11540 20502 11552
rect 20717 11543 20775 11549
rect 20717 11540 20729 11543
rect 20496 11512 20729 11540
rect 20496 11500 20502 11512
rect 20717 11509 20729 11512
rect 20763 11509 20775 11543
rect 20717 11503 20775 11509
rect 20806 11500 20812 11552
rect 20864 11540 20870 11552
rect 21358 11540 21364 11552
rect 20864 11512 21364 11540
rect 20864 11500 20870 11512
rect 21358 11500 21364 11512
rect 21416 11500 21422 11552
rect 29086 11500 29092 11552
rect 29144 11540 29150 11552
rect 30653 11543 30711 11549
rect 30653 11540 30665 11543
rect 29144 11512 30665 11540
rect 29144 11500 29150 11512
rect 30653 11509 30665 11512
rect 30699 11509 30711 11543
rect 30653 11503 30711 11509
rect 1104 11450 38824 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 38824 11450
rect 1104 11376 38824 11398
rect 8481 11339 8539 11345
rect 8481 11305 8493 11339
rect 8527 11336 8539 11339
rect 8754 11336 8760 11348
rect 8527 11308 8760 11336
rect 8527 11305 8539 11308
rect 8481 11299 8539 11305
rect 8754 11296 8760 11308
rect 8812 11336 8818 11348
rect 9398 11336 9404 11348
rect 8812 11308 9404 11336
rect 8812 11296 8818 11308
rect 9398 11296 9404 11308
rect 9456 11296 9462 11348
rect 10042 11296 10048 11348
rect 10100 11336 10106 11348
rect 10505 11339 10563 11345
rect 10505 11336 10517 11339
rect 10100 11308 10517 11336
rect 10100 11296 10106 11308
rect 10505 11305 10517 11308
rect 10551 11305 10563 11339
rect 12434 11336 12440 11348
rect 12395 11308 12440 11336
rect 10505 11299 10563 11305
rect 12434 11296 12440 11308
rect 12492 11296 12498 11348
rect 13081 11339 13139 11345
rect 13081 11305 13093 11339
rect 13127 11336 13139 11339
rect 13262 11336 13268 11348
rect 13127 11308 13268 11336
rect 13127 11305 13139 11308
rect 13081 11299 13139 11305
rect 13262 11296 13268 11308
rect 13320 11296 13326 11348
rect 16850 11336 16856 11348
rect 16811 11308 16856 11336
rect 16850 11296 16856 11308
rect 16908 11296 16914 11348
rect 17862 11296 17868 11348
rect 17920 11336 17926 11348
rect 18049 11339 18107 11345
rect 18049 11336 18061 11339
rect 17920 11308 18061 11336
rect 17920 11296 17926 11308
rect 18049 11305 18061 11308
rect 18095 11305 18107 11339
rect 18049 11299 18107 11305
rect 19337 11339 19395 11345
rect 19337 11305 19349 11339
rect 19383 11336 19395 11339
rect 20346 11336 20352 11348
rect 19383 11308 20352 11336
rect 19383 11305 19395 11308
rect 19337 11299 19395 11305
rect 19720 11280 19748 11308
rect 20346 11296 20352 11308
rect 20404 11296 20410 11348
rect 20438 11296 20444 11348
rect 20496 11336 20502 11348
rect 22281 11339 22339 11345
rect 22281 11336 22293 11339
rect 20496 11308 22293 11336
rect 20496 11296 20502 11308
rect 22281 11305 22293 11308
rect 22327 11305 22339 11339
rect 23658 11336 23664 11348
rect 23619 11308 23664 11336
rect 22281 11299 22339 11305
rect 23658 11296 23664 11308
rect 23716 11296 23722 11348
rect 24394 11336 24400 11348
rect 24355 11308 24400 11336
rect 24394 11296 24400 11308
rect 24452 11296 24458 11348
rect 24765 11339 24823 11345
rect 24765 11305 24777 11339
rect 24811 11336 24823 11339
rect 24854 11336 24860 11348
rect 24811 11308 24860 11336
rect 24811 11305 24823 11308
rect 24765 11299 24823 11305
rect 24854 11296 24860 11308
rect 24912 11336 24918 11348
rect 25314 11336 25320 11348
rect 24912 11308 25320 11336
rect 24912 11296 24918 11308
rect 25314 11296 25320 11308
rect 25372 11296 25378 11348
rect 28537 11339 28595 11345
rect 28537 11305 28549 11339
rect 28583 11336 28595 11339
rect 28810 11336 28816 11348
rect 28583 11308 28816 11336
rect 28583 11305 28595 11308
rect 28537 11299 28595 11305
rect 28810 11296 28816 11308
rect 28868 11296 28874 11348
rect 28994 11296 29000 11348
rect 29052 11336 29058 11348
rect 29273 11339 29331 11345
rect 29273 11336 29285 11339
rect 29052 11308 29285 11336
rect 29052 11296 29058 11308
rect 29273 11305 29285 11308
rect 29319 11336 29331 11339
rect 29362 11336 29368 11348
rect 29319 11308 29368 11336
rect 29319 11305 29331 11308
rect 29273 11299 29331 11305
rect 29362 11296 29368 11308
rect 29420 11296 29426 11348
rect 30098 11336 30104 11348
rect 30059 11308 30104 11336
rect 30098 11296 30104 11308
rect 30156 11296 30162 11348
rect 31754 11296 31760 11348
rect 31812 11336 31818 11348
rect 32309 11339 32367 11345
rect 32309 11336 32321 11339
rect 31812 11308 32321 11336
rect 31812 11296 31818 11308
rect 32309 11305 32321 11308
rect 32355 11305 32367 11339
rect 32309 11299 32367 11305
rect 6914 11228 6920 11280
rect 6972 11268 6978 11280
rect 7368 11271 7426 11277
rect 7368 11268 7380 11271
rect 6972 11240 7380 11268
rect 6972 11228 6978 11240
rect 7368 11237 7380 11240
rect 7414 11268 7426 11271
rect 8018 11268 8024 11280
rect 7414 11240 8024 11268
rect 7414 11237 7426 11240
rect 7368 11231 7426 11237
rect 8018 11228 8024 11240
rect 8076 11228 8082 11280
rect 10686 11228 10692 11280
rect 10744 11268 10750 11280
rect 11302 11271 11360 11277
rect 11302 11268 11314 11271
rect 10744 11240 11314 11268
rect 10744 11228 10750 11240
rect 11302 11237 11314 11240
rect 11348 11237 11360 11271
rect 11302 11231 11360 11237
rect 19702 11228 19708 11280
rect 19760 11228 19766 11280
rect 21174 11277 21180 11280
rect 21168 11268 21180 11277
rect 21135 11240 21180 11268
rect 21168 11231 21180 11240
rect 21174 11228 21180 11231
rect 21232 11228 21238 11280
rect 23474 11228 23480 11280
rect 23532 11268 23538 11280
rect 24029 11271 24087 11277
rect 24029 11268 24041 11271
rect 23532 11240 24041 11268
rect 23532 11228 23538 11240
rect 24029 11237 24041 11240
rect 24075 11268 24087 11271
rect 27424 11271 27482 11277
rect 24075 11240 25728 11268
rect 24075 11237 24087 11240
rect 24029 11231 24087 11237
rect 25700 11212 25728 11240
rect 27424 11237 27436 11271
rect 27470 11268 27482 11271
rect 27890 11268 27896 11280
rect 27470 11240 27896 11268
rect 27470 11237 27482 11240
rect 27424 11231 27482 11237
rect 27890 11228 27896 11240
rect 27948 11228 27954 11280
rect 7101 11203 7159 11209
rect 7101 11169 7113 11203
rect 7147 11200 7159 11203
rect 7926 11200 7932 11212
rect 7147 11172 7932 11200
rect 7147 11169 7159 11172
rect 7101 11163 7159 11169
rect 6822 11132 6828 11144
rect 6735 11104 6828 11132
rect 6822 11092 6828 11104
rect 6880 11132 6886 11144
rect 7116 11132 7144 11163
rect 7926 11160 7932 11172
rect 7984 11160 7990 11212
rect 9950 11200 9956 11212
rect 9911 11172 9956 11200
rect 9950 11160 9956 11172
rect 10008 11160 10014 11212
rect 11057 11203 11115 11209
rect 11057 11169 11069 11203
rect 11103 11200 11115 11203
rect 11882 11200 11888 11212
rect 11103 11172 11888 11200
rect 11103 11169 11115 11172
rect 11057 11163 11115 11169
rect 11882 11160 11888 11172
rect 11940 11160 11946 11212
rect 13538 11200 13544 11212
rect 13499 11172 13544 11200
rect 13538 11160 13544 11172
rect 13596 11160 13602 11212
rect 15746 11209 15752 11212
rect 15740 11200 15752 11209
rect 15707 11172 15752 11200
rect 15740 11163 15752 11172
rect 15746 11160 15752 11163
rect 15804 11160 15810 11212
rect 18693 11203 18751 11209
rect 18693 11169 18705 11203
rect 18739 11200 18751 11203
rect 18966 11200 18972 11212
rect 18739 11172 18972 11200
rect 18739 11169 18751 11172
rect 18693 11163 18751 11169
rect 18966 11160 18972 11172
rect 19024 11160 19030 11212
rect 24486 11160 24492 11212
rect 24544 11200 24550 11212
rect 24857 11203 24915 11209
rect 24857 11200 24869 11203
rect 24544 11172 24869 11200
rect 24544 11160 24550 11172
rect 24857 11169 24869 11172
rect 24903 11200 24915 11203
rect 25130 11200 25136 11212
rect 24903 11172 25136 11200
rect 24903 11169 24915 11172
rect 24857 11163 24915 11169
rect 25130 11160 25136 11172
rect 25188 11160 25194 11212
rect 25682 11160 25688 11212
rect 25740 11200 25746 11212
rect 25777 11203 25835 11209
rect 25777 11200 25789 11203
rect 25740 11172 25789 11200
rect 25740 11160 25746 11172
rect 25777 11169 25789 11172
rect 25823 11200 25835 11203
rect 26789 11203 26847 11209
rect 26789 11200 26801 11203
rect 25823 11172 26801 11200
rect 25823 11169 25835 11172
rect 25777 11163 25835 11169
rect 26789 11169 26801 11172
rect 26835 11200 26847 11203
rect 27157 11203 27215 11209
rect 27157 11200 27169 11203
rect 26835 11172 27169 11200
rect 26835 11169 26847 11172
rect 26789 11163 26847 11169
rect 27157 11169 27169 11172
rect 27203 11200 27215 11203
rect 27246 11200 27252 11212
rect 27203 11172 27252 11200
rect 27203 11169 27215 11172
rect 27157 11163 27215 11169
rect 27246 11160 27252 11172
rect 27304 11160 27310 11212
rect 30006 11200 30012 11212
rect 29967 11172 30012 11200
rect 30006 11160 30012 11172
rect 30064 11160 30070 11212
rect 32122 11200 32128 11212
rect 32083 11172 32128 11200
rect 32122 11160 32128 11172
rect 32180 11160 32186 11212
rect 6880 11104 7144 11132
rect 6880 11092 6886 11104
rect 15194 11092 15200 11144
rect 15252 11132 15258 11144
rect 15473 11135 15531 11141
rect 15473 11132 15485 11135
rect 15252 11104 15485 11132
rect 15252 11092 15258 11104
rect 15473 11101 15485 11104
rect 15519 11101 15531 11135
rect 20898 11132 20904 11144
rect 20859 11104 20904 11132
rect 15473 11095 15531 11101
rect 20898 11092 20904 11104
rect 20956 11092 20962 11144
rect 25041 11135 25099 11141
rect 25041 11101 25053 11135
rect 25087 11132 25099 11135
rect 25222 11132 25228 11144
rect 25087 11104 25228 11132
rect 25087 11101 25099 11104
rect 25041 11095 25099 11101
rect 25222 11092 25228 11104
rect 25280 11132 25286 11144
rect 25958 11132 25964 11144
rect 25280 11104 25964 11132
rect 25280 11092 25286 11104
rect 25958 11092 25964 11104
rect 26016 11092 26022 11144
rect 28994 11092 29000 11144
rect 29052 11132 29058 11144
rect 30190 11132 30196 11144
rect 29052 11104 30196 11132
rect 29052 11092 29058 11104
rect 30190 11092 30196 11104
rect 30248 11092 30254 11144
rect 10137 11067 10195 11073
rect 10137 11033 10149 11067
rect 10183 11064 10195 11067
rect 10962 11064 10968 11076
rect 10183 11036 10968 11064
rect 10183 11033 10195 11036
rect 10137 11027 10195 11033
rect 10962 11024 10968 11036
rect 11020 11024 11026 11076
rect 12526 11024 12532 11076
rect 12584 11064 12590 11076
rect 13725 11067 13783 11073
rect 13725 11064 13737 11067
rect 12584 11036 13737 11064
rect 12584 11024 12590 11036
rect 13725 11033 13737 11036
rect 13771 11033 13783 11067
rect 13725 11027 13783 11033
rect 18782 11024 18788 11076
rect 18840 11064 18846 11076
rect 18877 11067 18935 11073
rect 18877 11064 18889 11067
rect 18840 11036 18889 11064
rect 18840 11024 18846 11036
rect 18877 11033 18889 11036
rect 18923 11033 18935 11067
rect 20346 11064 20352 11076
rect 20307 11036 20352 11064
rect 18877 11027 18935 11033
rect 20346 11024 20352 11036
rect 20404 11024 20410 11076
rect 29641 11067 29699 11073
rect 29641 11033 29653 11067
rect 29687 11064 29699 11067
rect 32122 11064 32128 11076
rect 29687 11036 32128 11064
rect 29687 11033 29699 11036
rect 29641 11027 29699 11033
rect 32122 11024 32128 11036
rect 32180 11024 32186 11076
rect 18138 10956 18144 11008
rect 18196 10996 18202 11008
rect 18417 10999 18475 11005
rect 18417 10996 18429 10999
rect 18196 10968 18429 10996
rect 18196 10956 18202 10968
rect 18417 10965 18429 10968
rect 18463 10965 18475 10999
rect 19610 10996 19616 11008
rect 19571 10968 19616 10996
rect 18417 10959 18475 10965
rect 19610 10956 19616 10968
rect 19668 10956 19674 11008
rect 19978 10996 19984 11008
rect 19939 10968 19984 10996
rect 19978 10956 19984 10968
rect 20036 10956 20042 11008
rect 35526 10996 35532 11008
rect 35487 10968 35532 10996
rect 35526 10956 35532 10968
rect 35584 10956 35590 11008
rect 1104 10906 38824 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 34966 10906
rect 35018 10854 35030 10906
rect 35082 10854 35094 10906
rect 35146 10854 35158 10906
rect 35210 10854 38824 10906
rect 1104 10832 38824 10854
rect 6638 10792 6644 10804
rect 6599 10764 6644 10792
rect 6638 10752 6644 10764
rect 6696 10792 6702 10804
rect 7926 10792 7932 10804
rect 6696 10764 7328 10792
rect 7887 10764 7932 10792
rect 6696 10752 6702 10764
rect 6273 10727 6331 10733
rect 6273 10693 6285 10727
rect 6319 10724 6331 10727
rect 6914 10724 6920 10736
rect 6319 10696 6920 10724
rect 6319 10693 6331 10696
rect 6273 10687 6331 10693
rect 6914 10684 6920 10696
rect 6972 10684 6978 10736
rect 7300 10665 7328 10764
rect 7926 10752 7932 10764
rect 7984 10752 7990 10804
rect 8294 10792 8300 10804
rect 8255 10764 8300 10792
rect 8294 10752 8300 10764
rect 8352 10792 8358 10804
rect 9950 10792 9956 10804
rect 8352 10764 8892 10792
rect 9911 10764 9956 10792
rect 8352 10752 8358 10764
rect 7285 10659 7343 10665
rect 7285 10625 7297 10659
rect 7331 10625 7343 10659
rect 7285 10619 7343 10625
rect 7374 10616 7380 10668
rect 7432 10656 7438 10668
rect 8864 10665 8892 10764
rect 9950 10752 9956 10764
rect 10008 10752 10014 10804
rect 10505 10795 10563 10801
rect 10505 10761 10517 10795
rect 10551 10792 10563 10795
rect 10686 10792 10692 10804
rect 10551 10764 10692 10792
rect 10551 10761 10563 10764
rect 10505 10755 10563 10761
rect 10686 10752 10692 10764
rect 10744 10752 10750 10804
rect 10965 10795 11023 10801
rect 10965 10761 10977 10795
rect 11011 10792 11023 10795
rect 11054 10792 11060 10804
rect 11011 10764 11060 10792
rect 11011 10761 11023 10764
rect 10965 10755 11023 10761
rect 11054 10752 11060 10764
rect 11112 10752 11118 10804
rect 11698 10792 11704 10804
rect 11611 10764 11704 10792
rect 11698 10752 11704 10764
rect 11756 10792 11762 10804
rect 11882 10792 11888 10804
rect 11756 10764 11888 10792
rect 11756 10752 11762 10764
rect 11882 10752 11888 10764
rect 11940 10752 11946 10804
rect 13538 10792 13544 10804
rect 13499 10764 13544 10792
rect 13538 10752 13544 10764
rect 13596 10752 13602 10804
rect 15746 10752 15752 10804
rect 15804 10792 15810 10804
rect 16853 10795 16911 10801
rect 16853 10792 16865 10795
rect 15804 10764 16865 10792
rect 15804 10752 15810 10764
rect 16853 10761 16865 10764
rect 16899 10761 16911 10795
rect 18966 10792 18972 10804
rect 18927 10764 18972 10792
rect 16853 10755 16911 10761
rect 18966 10752 18972 10764
rect 19024 10752 19030 10804
rect 20254 10792 20260 10804
rect 20215 10764 20260 10792
rect 20254 10752 20260 10764
rect 20312 10752 20318 10804
rect 24486 10792 24492 10804
rect 24447 10764 24492 10792
rect 24486 10752 24492 10764
rect 24544 10752 24550 10804
rect 24854 10792 24860 10804
rect 24815 10764 24860 10792
rect 24854 10752 24860 10764
rect 24912 10752 24918 10804
rect 25222 10792 25228 10804
rect 25183 10764 25228 10792
rect 25222 10752 25228 10764
rect 25280 10752 25286 10804
rect 25866 10792 25872 10804
rect 25827 10764 25872 10792
rect 25866 10752 25872 10764
rect 25924 10752 25930 10804
rect 26234 10792 26240 10804
rect 26195 10764 26240 10792
rect 26234 10752 26240 10764
rect 26292 10752 26298 10804
rect 26881 10795 26939 10801
rect 26881 10761 26893 10795
rect 26927 10792 26939 10795
rect 27062 10792 27068 10804
rect 26927 10764 27068 10792
rect 26927 10761 26939 10764
rect 26881 10755 26939 10761
rect 18138 10684 18144 10736
rect 18196 10724 18202 10736
rect 19978 10724 19984 10736
rect 18196 10696 19984 10724
rect 18196 10684 18202 10696
rect 8849 10659 8907 10665
rect 7432 10628 7477 10656
rect 7432 10616 7438 10628
rect 8849 10625 8861 10659
rect 8895 10625 8907 10659
rect 8849 10619 8907 10625
rect 8938 10616 8944 10668
rect 8996 10656 9002 10668
rect 8996 10628 9041 10656
rect 8996 10616 9002 10628
rect 12434 10616 12440 10668
rect 12492 10656 12498 10668
rect 12897 10659 12955 10665
rect 12897 10656 12909 10659
rect 12492 10628 12909 10656
rect 12492 10616 12498 10628
rect 12897 10625 12909 10628
rect 12943 10656 12955 10659
rect 12986 10656 12992 10668
rect 12943 10628 12992 10656
rect 12943 10625 12955 10628
rect 12897 10619 12955 10625
rect 12986 10616 12992 10628
rect 13044 10616 13050 10668
rect 13081 10659 13139 10665
rect 13081 10625 13093 10659
rect 13127 10656 13139 10659
rect 13262 10656 13268 10668
rect 13127 10628 13268 10656
rect 13127 10625 13139 10628
rect 13081 10619 13139 10625
rect 13262 10616 13268 10628
rect 13320 10616 13326 10668
rect 15194 10616 15200 10668
rect 15252 10656 15258 10668
rect 15473 10659 15531 10665
rect 15473 10656 15485 10659
rect 15252 10628 15485 10656
rect 15252 10616 15258 10628
rect 15473 10625 15485 10628
rect 15519 10625 15531 10659
rect 19702 10656 19708 10668
rect 19663 10628 19708 10656
rect 15473 10619 15531 10625
rect 19702 10616 19708 10628
rect 19760 10616 19766 10668
rect 19812 10665 19840 10696
rect 19978 10684 19984 10696
rect 20036 10684 20042 10736
rect 19797 10659 19855 10665
rect 19797 10625 19809 10659
rect 19843 10625 19855 10659
rect 19797 10619 19855 10625
rect 8754 10588 8760 10600
rect 8715 10560 8760 10588
rect 8754 10548 8760 10560
rect 8812 10548 8818 10600
rect 10686 10548 10692 10600
rect 10744 10588 10750 10600
rect 10781 10591 10839 10597
rect 10781 10588 10793 10591
rect 10744 10560 10793 10588
rect 10744 10548 10750 10560
rect 10781 10557 10793 10560
rect 10827 10557 10839 10591
rect 10781 10551 10839 10557
rect 12253 10591 12311 10597
rect 12253 10557 12265 10591
rect 12299 10588 12311 10591
rect 12805 10591 12863 10597
rect 12805 10588 12817 10591
rect 12299 10560 12817 10588
rect 12299 10557 12311 10560
rect 12253 10551 12311 10557
rect 12805 10557 12817 10560
rect 12851 10588 12863 10591
rect 13722 10588 13728 10600
rect 12851 10560 13728 10588
rect 12851 10557 12863 10560
rect 12805 10551 12863 10557
rect 13722 10548 13728 10560
rect 13780 10548 13786 10600
rect 18049 10591 18107 10597
rect 18049 10557 18061 10591
rect 18095 10588 18107 10591
rect 19610 10588 19616 10600
rect 18095 10560 18736 10588
rect 19571 10560 19616 10588
rect 18095 10557 18107 10560
rect 18049 10551 18107 10557
rect 6546 10480 6552 10532
rect 6604 10520 6610 10532
rect 6604 10492 6960 10520
rect 6604 10480 6610 10492
rect 6822 10452 6828 10464
rect 6783 10424 6828 10452
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 6932 10452 6960 10492
rect 7006 10480 7012 10532
rect 7064 10520 7070 10532
rect 7193 10523 7251 10529
rect 7193 10520 7205 10523
rect 7064 10492 7205 10520
rect 7064 10480 7070 10492
rect 7193 10489 7205 10492
rect 7239 10489 7251 10523
rect 7193 10483 7251 10489
rect 10597 10523 10655 10529
rect 10597 10489 10609 10523
rect 10643 10489 10655 10523
rect 10597 10483 10655 10489
rect 15013 10523 15071 10529
rect 15013 10489 15025 10523
rect 15059 10520 15071 10523
rect 15718 10523 15776 10529
rect 15718 10520 15730 10523
rect 15059 10492 15730 10520
rect 15059 10489 15071 10492
rect 15013 10483 15071 10489
rect 15718 10489 15730 10492
rect 15764 10520 15776 10523
rect 16298 10520 16304 10532
rect 15764 10492 16304 10520
rect 15764 10489 15776 10492
rect 15718 10483 15776 10489
rect 7374 10452 7380 10464
rect 6932 10424 7380 10452
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 7650 10412 7656 10464
rect 7708 10452 7714 10464
rect 8389 10455 8447 10461
rect 8389 10452 8401 10455
rect 7708 10424 8401 10452
rect 7708 10412 7714 10424
rect 8389 10421 8401 10424
rect 8435 10421 8447 10455
rect 10612 10452 10640 10483
rect 16298 10480 16304 10492
rect 16356 10480 16362 10532
rect 18708 10464 18736 10560
rect 19610 10548 19616 10560
rect 19668 10588 19674 10600
rect 20070 10588 20076 10600
rect 19668 10560 20076 10588
rect 19668 10548 19674 10560
rect 20070 10548 20076 10560
rect 20128 10548 20134 10600
rect 20806 10588 20812 10600
rect 20767 10560 20812 10588
rect 20806 10548 20812 10560
rect 20864 10548 20870 10600
rect 25685 10591 25743 10597
rect 25685 10557 25697 10591
rect 25731 10588 25743 10591
rect 26234 10588 26240 10600
rect 25731 10560 26240 10588
rect 25731 10557 25743 10560
rect 25685 10551 25743 10557
rect 26234 10548 26240 10560
rect 26292 10548 26298 10600
rect 26988 10597 27016 10764
rect 27062 10752 27068 10764
rect 27120 10752 27126 10804
rect 27154 10752 27160 10804
rect 27212 10792 27218 10804
rect 27890 10792 27896 10804
rect 27212 10764 27257 10792
rect 27851 10764 27896 10792
rect 27212 10752 27218 10764
rect 27890 10752 27896 10764
rect 27948 10752 27954 10804
rect 28353 10795 28411 10801
rect 28353 10761 28365 10795
rect 28399 10792 28411 10795
rect 28902 10792 28908 10804
rect 28399 10764 28908 10792
rect 28399 10761 28411 10764
rect 28353 10755 28411 10761
rect 28902 10752 28908 10764
rect 28960 10752 28966 10804
rect 29086 10792 29092 10804
rect 29047 10764 29092 10792
rect 29086 10752 29092 10764
rect 29144 10752 29150 10804
rect 29362 10752 29368 10804
rect 29420 10792 29426 10804
rect 29641 10795 29699 10801
rect 29641 10792 29653 10795
rect 29420 10764 29653 10792
rect 29420 10752 29426 10764
rect 29641 10761 29653 10764
rect 29687 10761 29699 10795
rect 32122 10792 32128 10804
rect 32083 10764 32128 10792
rect 29641 10755 29699 10761
rect 27246 10684 27252 10736
rect 27304 10724 27310 10736
rect 27617 10727 27675 10733
rect 27617 10724 27629 10727
rect 27304 10696 27629 10724
rect 27304 10684 27310 10696
rect 27617 10693 27629 10696
rect 27663 10693 27675 10727
rect 28718 10724 28724 10736
rect 28679 10696 28724 10724
rect 27617 10687 27675 10693
rect 28718 10684 28724 10696
rect 28776 10684 28782 10736
rect 29656 10656 29684 10755
rect 32122 10752 32128 10764
rect 32180 10752 32186 10804
rect 36814 10792 36820 10804
rect 36775 10764 36820 10792
rect 36814 10752 36820 10764
rect 36872 10752 36878 10804
rect 29825 10659 29883 10665
rect 29825 10656 29837 10659
rect 29656 10628 29837 10656
rect 29825 10625 29837 10628
rect 29871 10656 29883 10659
rect 29871 10628 29960 10656
rect 29871 10625 29883 10628
rect 29825 10619 29883 10625
rect 29932 10600 29960 10628
rect 26973 10591 27031 10597
rect 26973 10557 26985 10591
rect 27019 10557 27031 10591
rect 26973 10551 27031 10557
rect 29914 10548 29920 10600
rect 29972 10548 29978 10600
rect 32306 10588 32312 10600
rect 32267 10560 32312 10588
rect 32306 10548 32312 10560
rect 32364 10588 32370 10600
rect 32861 10591 32919 10597
rect 32861 10588 32873 10591
rect 32364 10560 32873 10588
rect 32364 10548 32370 10560
rect 32861 10557 32873 10560
rect 32907 10557 32919 10591
rect 35437 10591 35495 10597
rect 35437 10588 35449 10591
rect 32861 10551 32919 10557
rect 35268 10560 35449 10588
rect 30092 10523 30150 10529
rect 30092 10489 30104 10523
rect 30138 10520 30150 10523
rect 30282 10520 30288 10532
rect 30138 10492 30288 10520
rect 30138 10489 30150 10492
rect 30092 10483 30150 10489
rect 30282 10480 30288 10492
rect 30340 10480 30346 10532
rect 11330 10452 11336 10464
rect 10612 10424 11336 10452
rect 8389 10415 8447 10421
rect 11330 10412 11336 10424
rect 11388 10412 11394 10464
rect 12437 10455 12495 10461
rect 12437 10421 12449 10455
rect 12483 10452 12495 10455
rect 12526 10452 12532 10464
rect 12483 10424 12532 10452
rect 12483 10421 12495 10424
rect 12437 10415 12495 10421
rect 12526 10412 12532 10424
rect 12584 10412 12590 10464
rect 15194 10412 15200 10464
rect 15252 10452 15258 10464
rect 15289 10455 15347 10461
rect 15289 10452 15301 10455
rect 15252 10424 15301 10452
rect 15252 10412 15258 10424
rect 15289 10421 15301 10424
rect 15335 10421 15347 10455
rect 15289 10415 15347 10421
rect 18138 10412 18144 10464
rect 18196 10452 18202 10464
rect 18233 10455 18291 10461
rect 18233 10452 18245 10455
rect 18196 10424 18245 10452
rect 18196 10412 18202 10424
rect 18233 10421 18245 10424
rect 18279 10421 18291 10455
rect 18690 10452 18696 10464
rect 18651 10424 18696 10452
rect 18233 10415 18291 10421
rect 18690 10412 18696 10424
rect 18748 10412 18754 10464
rect 19242 10452 19248 10464
rect 19203 10424 19248 10452
rect 19242 10412 19248 10424
rect 19300 10412 19306 10464
rect 20717 10455 20775 10461
rect 20717 10421 20729 10455
rect 20763 10452 20775 10455
rect 20898 10452 20904 10464
rect 20763 10424 20904 10452
rect 20763 10421 20775 10424
rect 20717 10415 20775 10421
rect 20898 10412 20904 10424
rect 20956 10412 20962 10464
rect 21910 10412 21916 10464
rect 21968 10452 21974 10464
rect 22097 10455 22155 10461
rect 22097 10452 22109 10455
rect 21968 10424 22109 10452
rect 21968 10412 21974 10424
rect 22097 10421 22109 10424
rect 22143 10421 22155 10455
rect 31202 10452 31208 10464
rect 31163 10424 31208 10452
rect 22097 10415 22155 10421
rect 31202 10412 31208 10424
rect 31260 10412 31266 10464
rect 32490 10452 32496 10464
rect 32451 10424 32496 10452
rect 32490 10412 32496 10424
rect 32548 10412 32554 10464
rect 33318 10452 33324 10464
rect 33279 10424 33324 10452
rect 33318 10412 33324 10424
rect 33376 10412 33382 10464
rect 35158 10412 35164 10464
rect 35216 10452 35222 10464
rect 35268 10461 35296 10560
rect 35437 10557 35449 10560
rect 35483 10557 35495 10591
rect 35437 10551 35495 10557
rect 35526 10548 35532 10600
rect 35584 10588 35590 10600
rect 35693 10591 35751 10597
rect 35693 10588 35705 10591
rect 35584 10560 35705 10588
rect 35584 10548 35590 10560
rect 35693 10557 35705 10560
rect 35739 10557 35751 10591
rect 35693 10551 35751 10557
rect 35253 10455 35311 10461
rect 35253 10452 35265 10455
rect 35216 10424 35265 10452
rect 35216 10412 35222 10424
rect 35253 10421 35265 10424
rect 35299 10421 35311 10455
rect 35253 10415 35311 10421
rect 1104 10362 38824 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 38824 10362
rect 1104 10288 38824 10310
rect 6546 10248 6552 10260
rect 6507 10220 6552 10248
rect 6546 10208 6552 10220
rect 6604 10208 6610 10260
rect 6822 10208 6828 10260
rect 6880 10248 6886 10260
rect 7098 10248 7104 10260
rect 6880 10220 7104 10248
rect 6880 10208 6886 10220
rect 7098 10208 7104 10220
rect 7156 10248 7162 10260
rect 7650 10248 7656 10260
rect 7156 10220 7512 10248
rect 7611 10220 7656 10248
rect 7156 10208 7162 10220
rect 7484 10180 7512 10220
rect 7650 10208 7656 10220
rect 7708 10208 7714 10260
rect 8481 10251 8539 10257
rect 8481 10217 8493 10251
rect 8527 10248 8539 10251
rect 8754 10248 8760 10260
rect 8527 10220 8760 10248
rect 8527 10217 8539 10220
rect 8481 10211 8539 10217
rect 8754 10208 8760 10220
rect 8812 10208 8818 10260
rect 10686 10208 10692 10260
rect 10744 10248 10750 10260
rect 11057 10251 11115 10257
rect 11057 10248 11069 10251
rect 10744 10220 11069 10248
rect 10744 10208 10750 10220
rect 11057 10217 11069 10220
rect 11103 10217 11115 10251
rect 11057 10211 11115 10217
rect 12897 10251 12955 10257
rect 12897 10217 12909 10251
rect 12943 10248 12955 10251
rect 13262 10248 13268 10260
rect 12943 10220 13268 10248
rect 12943 10217 12955 10220
rect 12897 10211 12955 10217
rect 13262 10208 13268 10220
rect 13320 10208 13326 10260
rect 15194 10208 15200 10260
rect 15252 10248 15258 10260
rect 15473 10251 15531 10257
rect 15473 10248 15485 10251
rect 15252 10220 15485 10248
rect 15252 10208 15258 10220
rect 15473 10217 15485 10220
rect 15519 10217 15531 10251
rect 15473 10211 15531 10217
rect 15746 10208 15752 10260
rect 15804 10248 15810 10260
rect 15841 10251 15899 10257
rect 15841 10248 15853 10251
rect 15804 10220 15853 10248
rect 15804 10208 15810 10220
rect 15841 10217 15853 10220
rect 15887 10217 15899 10251
rect 15841 10211 15899 10217
rect 15930 10208 15936 10260
rect 15988 10248 15994 10260
rect 16393 10251 16451 10257
rect 16393 10248 16405 10251
rect 15988 10220 16405 10248
rect 15988 10208 15994 10220
rect 16393 10217 16405 10220
rect 16439 10248 16451 10251
rect 16574 10248 16580 10260
rect 16439 10220 16580 10248
rect 16439 10217 16451 10220
rect 16393 10211 16451 10217
rect 16574 10208 16580 10220
rect 16632 10208 16638 10260
rect 17957 10251 18015 10257
rect 17957 10217 17969 10251
rect 18003 10248 18015 10251
rect 18230 10248 18236 10260
rect 18003 10220 18236 10248
rect 18003 10217 18015 10220
rect 17957 10211 18015 10217
rect 18230 10208 18236 10220
rect 18288 10208 18294 10260
rect 29454 10248 29460 10260
rect 29415 10220 29460 10248
rect 29454 10208 29460 10220
rect 29512 10208 29518 10260
rect 29917 10251 29975 10257
rect 29917 10217 29929 10251
rect 29963 10248 29975 10251
rect 30282 10248 30288 10260
rect 29963 10220 30288 10248
rect 29963 10217 29975 10220
rect 29917 10211 29975 10217
rect 30282 10208 30288 10220
rect 30340 10208 30346 10260
rect 30374 10208 30380 10260
rect 30432 10248 30438 10260
rect 30469 10251 30527 10257
rect 30469 10248 30481 10251
rect 30432 10220 30481 10248
rect 30432 10208 30438 10220
rect 30469 10217 30481 10220
rect 30515 10248 30527 10251
rect 31662 10248 31668 10260
rect 30515 10220 31668 10248
rect 30515 10217 30527 10220
rect 30469 10211 30527 10217
rect 31662 10208 31668 10220
rect 31720 10208 31726 10260
rect 33226 10208 33232 10260
rect 33284 10248 33290 10260
rect 33689 10251 33747 10257
rect 33689 10248 33701 10251
rect 33284 10220 33701 10248
rect 33284 10208 33290 10220
rect 33689 10217 33701 10220
rect 33735 10248 33747 10251
rect 33778 10248 33784 10260
rect 33735 10220 33784 10248
rect 33735 10217 33747 10220
rect 33689 10211 33747 10217
rect 33778 10208 33784 10220
rect 33836 10208 33842 10260
rect 35526 10208 35532 10260
rect 35584 10248 35590 10260
rect 36541 10251 36599 10257
rect 36541 10248 36553 10251
rect 35584 10220 36553 10248
rect 35584 10208 35590 10220
rect 36541 10217 36553 10220
rect 36587 10217 36599 10251
rect 36541 10211 36599 10217
rect 7745 10183 7803 10189
rect 7745 10180 7757 10183
rect 7484 10152 7757 10180
rect 7745 10149 7757 10152
rect 7791 10149 7803 10183
rect 7745 10143 7803 10149
rect 11793 10183 11851 10189
rect 11793 10149 11805 10183
rect 11839 10180 11851 10183
rect 11882 10180 11888 10192
rect 11839 10152 11888 10180
rect 11839 10149 11851 10152
rect 11793 10143 11851 10149
rect 11882 10140 11888 10152
rect 11940 10140 11946 10192
rect 12986 10140 12992 10192
rect 13044 10180 13050 10192
rect 13173 10183 13231 10189
rect 13173 10180 13185 10183
rect 13044 10152 13185 10180
rect 13044 10140 13050 10152
rect 13173 10149 13185 10152
rect 13219 10149 13231 10183
rect 13173 10143 13231 10149
rect 20346 10140 20352 10192
rect 20404 10180 20410 10192
rect 21238 10183 21296 10189
rect 21238 10180 21250 10183
rect 20404 10152 21250 10180
rect 20404 10140 20410 10152
rect 21238 10149 21250 10152
rect 21284 10149 21296 10183
rect 21238 10143 21296 10149
rect 6822 10072 6828 10124
rect 6880 10112 6886 10124
rect 7650 10112 7656 10124
rect 6880 10084 7656 10112
rect 6880 10072 6886 10084
rect 7650 10072 7656 10084
rect 7708 10072 7714 10124
rect 9677 10115 9735 10121
rect 9677 10081 9689 10115
rect 9723 10112 9735 10115
rect 10410 10112 10416 10124
rect 9723 10084 10416 10112
rect 9723 10081 9735 10084
rect 9677 10075 9735 10081
rect 10410 10072 10416 10084
rect 10468 10072 10474 10124
rect 14093 10115 14151 10121
rect 14093 10081 14105 10115
rect 14139 10112 14151 10115
rect 14182 10112 14188 10124
rect 14139 10084 14188 10112
rect 14139 10081 14151 10084
rect 14093 10075 14151 10081
rect 14182 10072 14188 10084
rect 14240 10112 14246 10124
rect 19153 10115 19211 10121
rect 14240 10084 16068 10112
rect 14240 10072 14246 10084
rect 6917 10047 6975 10053
rect 6917 10013 6929 10047
rect 6963 10044 6975 10047
rect 7006 10044 7012 10056
rect 6963 10016 7012 10044
rect 6963 10013 6975 10016
rect 6917 10007 6975 10013
rect 7006 10004 7012 10016
rect 7064 10004 7070 10056
rect 7742 10004 7748 10056
rect 7800 10044 7806 10056
rect 7837 10047 7895 10053
rect 7837 10044 7849 10047
rect 7800 10016 7849 10044
rect 7800 10004 7806 10016
rect 7837 10013 7849 10016
rect 7883 10044 7895 10047
rect 8294 10044 8300 10056
rect 7883 10016 8300 10044
rect 7883 10013 7895 10016
rect 7837 10007 7895 10013
rect 8294 10004 8300 10016
rect 8352 10004 8358 10056
rect 10778 10044 10784 10056
rect 10691 10016 10784 10044
rect 10778 10004 10784 10016
rect 10836 10044 10842 10056
rect 11885 10047 11943 10053
rect 11885 10044 11897 10047
rect 10836 10016 11897 10044
rect 10836 10004 10842 10016
rect 11885 10013 11897 10016
rect 11931 10013 11943 10047
rect 11885 10007 11943 10013
rect 12069 10047 12127 10053
rect 12069 10013 12081 10047
rect 12115 10044 12127 10047
rect 12158 10044 12164 10056
rect 12115 10016 12164 10044
rect 12115 10013 12127 10016
rect 12069 10007 12127 10013
rect 12158 10004 12164 10016
rect 12216 10004 12222 10056
rect 7466 9936 7472 9988
rect 7524 9976 7530 9988
rect 8757 9979 8815 9985
rect 8757 9976 8769 9979
rect 7524 9948 8769 9976
rect 7524 9936 7530 9948
rect 8757 9945 8769 9948
rect 8803 9976 8815 9979
rect 8938 9976 8944 9988
rect 8803 9948 8944 9976
rect 8803 9945 8815 9948
rect 8757 9939 8815 9945
rect 8938 9936 8944 9948
rect 8996 9936 9002 9988
rect 14274 9976 14280 9988
rect 14235 9948 14280 9976
rect 14274 9936 14280 9948
rect 14332 9936 14338 9988
rect 16040 9985 16068 10084
rect 19153 10081 19165 10115
rect 19199 10112 19211 10115
rect 19242 10112 19248 10124
rect 19199 10084 19248 10112
rect 19199 10081 19211 10084
rect 19153 10075 19211 10081
rect 19242 10072 19248 10084
rect 19300 10072 19306 10124
rect 28902 10112 28908 10124
rect 28815 10084 28908 10112
rect 28902 10072 28908 10084
rect 28960 10112 28966 10124
rect 29472 10112 29500 10208
rect 28960 10084 29500 10112
rect 28960 10072 28966 10084
rect 29822 10072 29828 10124
rect 29880 10112 29886 10124
rect 30377 10115 30435 10121
rect 30377 10112 30389 10115
rect 29880 10084 30389 10112
rect 29880 10072 29886 10084
rect 30377 10081 30389 10084
rect 30423 10081 30435 10115
rect 30377 10075 30435 10081
rect 32490 10072 32496 10124
rect 32548 10112 32554 10124
rect 33042 10112 33048 10124
rect 32548 10084 33048 10112
rect 32548 10072 32554 10084
rect 33042 10072 33048 10084
rect 33100 10112 33106 10124
rect 33597 10115 33655 10121
rect 33597 10112 33609 10115
rect 33100 10084 33609 10112
rect 33100 10072 33106 10084
rect 33597 10081 33609 10084
rect 33643 10081 33655 10115
rect 33597 10075 33655 10081
rect 34606 10072 34612 10124
rect 34664 10112 34670 10124
rect 35158 10112 35164 10124
rect 34664 10084 35164 10112
rect 34664 10072 34670 10084
rect 35158 10072 35164 10084
rect 35216 10072 35222 10124
rect 35428 10115 35486 10121
rect 35428 10081 35440 10115
rect 35474 10112 35486 10115
rect 35802 10112 35808 10124
rect 35474 10084 35808 10112
rect 35474 10081 35486 10084
rect 35428 10075 35486 10081
rect 35802 10072 35808 10084
rect 35860 10072 35866 10124
rect 16482 10044 16488 10056
rect 16443 10016 16488 10044
rect 16482 10004 16488 10016
rect 16540 10004 16546 10056
rect 16577 10047 16635 10053
rect 16577 10013 16589 10047
rect 16623 10013 16635 10047
rect 18046 10044 18052 10056
rect 18007 10016 18052 10044
rect 16577 10007 16635 10013
rect 16025 9979 16083 9985
rect 16025 9945 16037 9979
rect 16071 9945 16083 9979
rect 16025 9939 16083 9945
rect 16114 9936 16120 9988
rect 16172 9976 16178 9988
rect 16592 9976 16620 10007
rect 18046 10004 18052 10016
rect 18104 10004 18110 10056
rect 18138 10004 18144 10056
rect 18196 10044 18202 10056
rect 20993 10047 21051 10053
rect 20993 10044 21005 10047
rect 18196 10016 18241 10044
rect 20916 10016 21005 10044
rect 18196 10004 18202 10016
rect 16172 9948 16620 9976
rect 16172 9936 16178 9948
rect 20916 9920 20944 10016
rect 20993 10013 21005 10016
rect 21039 10013 21051 10047
rect 20993 10007 21051 10013
rect 29089 9979 29147 9985
rect 29089 9945 29101 9979
rect 29135 9976 29147 9979
rect 29840 9976 29868 10072
rect 30558 10044 30564 10056
rect 30519 10016 30564 10044
rect 30558 10004 30564 10016
rect 30616 10044 30622 10056
rect 31021 10047 31079 10053
rect 31021 10044 31033 10047
rect 30616 10016 31033 10044
rect 30616 10004 30622 10016
rect 31021 10013 31033 10016
rect 31067 10044 31079 10047
rect 31202 10044 31208 10056
rect 31067 10016 31208 10044
rect 31067 10013 31079 10016
rect 31021 10007 31079 10013
rect 31202 10004 31208 10016
rect 31260 10004 31266 10056
rect 33318 10004 33324 10056
rect 33376 10044 33382 10056
rect 33781 10047 33839 10053
rect 33781 10044 33793 10047
rect 33376 10016 33793 10044
rect 33376 10004 33382 10016
rect 33781 10013 33793 10016
rect 33827 10044 33839 10047
rect 34790 10044 34796 10056
rect 33827 10016 34796 10044
rect 33827 10013 33839 10016
rect 33781 10007 33839 10013
rect 34790 10004 34796 10016
rect 34848 10044 34854 10056
rect 34885 10047 34943 10053
rect 34885 10044 34897 10047
rect 34848 10016 34897 10044
rect 34848 10004 34854 10016
rect 34885 10013 34897 10016
rect 34931 10013 34943 10047
rect 34885 10007 34943 10013
rect 33226 9976 33232 9988
rect 29135 9948 29868 9976
rect 33187 9948 33232 9976
rect 29135 9945 29147 9948
rect 29089 9939 29147 9945
rect 33226 9936 33232 9948
rect 33284 9936 33290 9988
rect 7285 9911 7343 9917
rect 7285 9877 7297 9911
rect 7331 9908 7343 9911
rect 7834 9908 7840 9920
rect 7331 9880 7840 9908
rect 7331 9877 7343 9880
rect 7285 9871 7343 9877
rect 7834 9868 7840 9880
rect 7892 9868 7898 9920
rect 9674 9868 9680 9920
rect 9732 9908 9738 9920
rect 9861 9911 9919 9917
rect 9861 9908 9873 9911
rect 9732 9880 9873 9908
rect 9732 9868 9738 9880
rect 9861 9877 9873 9880
rect 9907 9877 9919 9911
rect 9861 9871 9919 9877
rect 11425 9911 11483 9917
rect 11425 9877 11437 9911
rect 11471 9908 11483 9911
rect 12342 9908 12348 9920
rect 11471 9880 12348 9908
rect 11471 9877 11483 9880
rect 11425 9871 11483 9877
rect 12342 9868 12348 9880
rect 12400 9868 12406 9920
rect 12529 9911 12587 9917
rect 12529 9877 12541 9911
rect 12575 9908 12587 9911
rect 12894 9908 12900 9920
rect 12575 9880 12900 9908
rect 12575 9877 12587 9880
rect 12529 9871 12587 9877
rect 12894 9868 12900 9880
rect 12952 9868 12958 9920
rect 17589 9911 17647 9917
rect 17589 9877 17601 9911
rect 17635 9908 17647 9911
rect 17862 9908 17868 9920
rect 17635 9880 17868 9908
rect 17635 9877 17647 9880
rect 17589 9871 17647 9877
rect 17862 9868 17868 9880
rect 17920 9868 17926 9920
rect 18969 9911 19027 9917
rect 18969 9877 18981 9911
rect 19015 9908 19027 9911
rect 19242 9908 19248 9920
rect 19015 9880 19248 9908
rect 19015 9877 19027 9880
rect 18969 9871 19027 9877
rect 19242 9868 19248 9880
rect 19300 9908 19306 9920
rect 19337 9911 19395 9917
rect 19337 9908 19349 9911
rect 19300 9880 19349 9908
rect 19300 9868 19306 9880
rect 19337 9877 19349 9880
rect 19383 9877 19395 9911
rect 19794 9908 19800 9920
rect 19755 9880 19800 9908
rect 19337 9871 19395 9877
rect 19794 9868 19800 9880
rect 19852 9868 19858 9920
rect 20162 9908 20168 9920
rect 20123 9880 20168 9908
rect 20162 9868 20168 9880
rect 20220 9868 20226 9920
rect 20717 9911 20775 9917
rect 20717 9877 20729 9911
rect 20763 9908 20775 9911
rect 20898 9908 20904 9920
rect 20763 9880 20904 9908
rect 20763 9877 20775 9880
rect 20717 9871 20775 9877
rect 20898 9868 20904 9880
rect 20956 9868 20962 9920
rect 22002 9868 22008 9920
rect 22060 9908 22066 9920
rect 22373 9911 22431 9917
rect 22373 9908 22385 9911
rect 22060 9880 22385 9908
rect 22060 9868 22066 9880
rect 22373 9877 22385 9880
rect 22419 9877 22431 9911
rect 25406 9908 25412 9920
rect 25367 9880 25412 9908
rect 22373 9871 22431 9877
rect 25406 9868 25412 9880
rect 25464 9868 25470 9920
rect 30006 9908 30012 9920
rect 29967 9880 30012 9908
rect 30006 9868 30012 9880
rect 30064 9868 30070 9920
rect 32858 9908 32864 9920
rect 32819 9880 32864 9908
rect 32858 9868 32864 9880
rect 32916 9868 32922 9920
rect 1104 9818 38824 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 34966 9818
rect 35018 9766 35030 9818
rect 35082 9766 35094 9818
rect 35146 9766 35158 9818
rect 35210 9766 38824 9818
rect 1104 9744 38824 9766
rect 7098 9664 7104 9716
rect 7156 9704 7162 9716
rect 7285 9707 7343 9713
rect 7285 9704 7297 9707
rect 7156 9676 7297 9704
rect 7156 9664 7162 9676
rect 7285 9673 7297 9676
rect 7331 9673 7343 9707
rect 7285 9667 7343 9673
rect 7466 9664 7472 9716
rect 7524 9704 7530 9716
rect 7929 9707 7987 9713
rect 7929 9704 7941 9707
rect 7524 9676 7941 9704
rect 7524 9664 7530 9676
rect 7929 9673 7941 9676
rect 7975 9673 7987 9707
rect 10778 9704 10784 9716
rect 10739 9676 10784 9704
rect 7929 9667 7987 9673
rect 10778 9664 10784 9676
rect 10836 9664 10842 9716
rect 14182 9704 14188 9716
rect 14143 9676 14188 9704
rect 14182 9664 14188 9676
rect 14240 9664 14246 9716
rect 16114 9704 16120 9716
rect 15120 9676 16120 9704
rect 6641 9639 6699 9645
rect 6641 9605 6653 9639
rect 6687 9636 6699 9639
rect 6822 9636 6828 9648
rect 6687 9608 6828 9636
rect 6687 9605 6699 9608
rect 6641 9599 6699 9605
rect 6822 9596 6828 9608
rect 6880 9596 6886 9648
rect 8294 9596 8300 9648
rect 8352 9636 8358 9648
rect 8665 9639 8723 9645
rect 8665 9636 8677 9639
rect 8352 9608 8677 9636
rect 8352 9596 8358 9608
rect 8665 9605 8677 9608
rect 8711 9636 8723 9639
rect 9582 9636 9588 9648
rect 8711 9608 9588 9636
rect 8711 9605 8723 9608
rect 8665 9599 8723 9605
rect 9582 9596 9588 9608
rect 9640 9596 9646 9648
rect 13906 9636 13912 9648
rect 13096 9608 13912 9636
rect 13096 9580 13124 9608
rect 13906 9596 13912 9608
rect 13964 9596 13970 9648
rect 14645 9639 14703 9645
rect 14645 9605 14657 9639
rect 14691 9636 14703 9639
rect 15120 9636 15148 9676
rect 16114 9664 16120 9676
rect 16172 9664 16178 9716
rect 18230 9704 18236 9716
rect 18191 9676 18236 9704
rect 18230 9664 18236 9676
rect 18288 9664 18294 9716
rect 20070 9704 20076 9716
rect 20031 9676 20076 9704
rect 20070 9664 20076 9676
rect 20128 9664 20134 9716
rect 28902 9704 28908 9716
rect 28863 9676 28908 9704
rect 28902 9664 28908 9676
rect 28960 9664 28966 9716
rect 29822 9704 29828 9716
rect 29783 9676 29828 9704
rect 29822 9664 29828 9676
rect 29880 9664 29886 9716
rect 32490 9664 32496 9716
rect 32548 9704 32554 9716
rect 32585 9707 32643 9713
rect 32585 9704 32597 9707
rect 32548 9676 32597 9704
rect 32548 9664 32554 9676
rect 32585 9673 32597 9676
rect 32631 9673 32643 9707
rect 33778 9704 33784 9716
rect 33739 9676 33784 9704
rect 32585 9667 32643 9673
rect 33778 9664 33784 9676
rect 33836 9664 33842 9716
rect 17586 9636 17592 9648
rect 14691 9608 15148 9636
rect 17547 9608 17592 9636
rect 14691 9605 14703 9608
rect 14645 9599 14703 9605
rect 17586 9596 17592 9608
rect 17644 9596 17650 9648
rect 18782 9636 18788 9648
rect 18743 9608 18788 9636
rect 18782 9596 18788 9608
rect 18840 9596 18846 9648
rect 19981 9639 20039 9645
rect 19981 9605 19993 9639
rect 20027 9636 20039 9639
rect 20346 9636 20352 9648
rect 20027 9608 20352 9636
rect 20027 9605 20039 9608
rect 19981 9599 20039 9605
rect 20346 9596 20352 9608
rect 20404 9596 20410 9648
rect 11422 9568 11428 9580
rect 11383 9540 11428 9568
rect 11422 9528 11428 9540
rect 11480 9528 11486 9580
rect 12618 9528 12624 9580
rect 12676 9568 12682 9580
rect 12894 9568 12900 9580
rect 12676 9540 12900 9568
rect 12676 9528 12682 9540
rect 12894 9528 12900 9540
rect 12952 9528 12958 9580
rect 13078 9568 13084 9580
rect 12991 9540 13084 9568
rect 13078 9528 13084 9540
rect 13136 9528 13142 9580
rect 18800 9568 18828 9596
rect 19337 9571 19395 9577
rect 19337 9568 19349 9571
rect 18800 9540 19349 9568
rect 19337 9537 19349 9540
rect 19383 9537 19395 9571
rect 19337 9531 19395 9537
rect 19429 9571 19487 9577
rect 19429 9537 19441 9571
rect 19475 9537 19487 9571
rect 19429 9531 19487 9537
rect 7745 9503 7803 9509
rect 7745 9469 7757 9503
rect 7791 9500 7803 9503
rect 10689 9503 10747 9509
rect 7791 9472 8432 9500
rect 7791 9469 7803 9472
rect 7745 9463 7803 9469
rect 8404 9441 8432 9472
rect 10689 9469 10701 9503
rect 10735 9500 10747 9503
rect 11149 9503 11207 9509
rect 11149 9500 11161 9503
rect 10735 9472 11161 9500
rect 10735 9469 10747 9472
rect 10689 9463 10747 9469
rect 11149 9469 11161 9472
rect 11195 9500 11207 9503
rect 12250 9500 12256 9512
rect 11195 9472 12256 9500
rect 11195 9469 11207 9472
rect 11149 9463 11207 9469
rect 12250 9460 12256 9472
rect 12308 9460 12314 9512
rect 15473 9503 15531 9509
rect 15473 9500 15485 9503
rect 15304 9472 15485 9500
rect 8389 9435 8447 9441
rect 8389 9401 8401 9435
rect 8435 9432 8447 9435
rect 9398 9432 9404 9444
rect 8435 9404 9404 9432
rect 8435 9401 8447 9404
rect 8389 9395 8447 9401
rect 9398 9392 9404 9404
rect 9456 9392 9462 9444
rect 9769 9435 9827 9441
rect 9769 9401 9781 9435
rect 9815 9432 9827 9435
rect 10870 9432 10876 9444
rect 9815 9404 10876 9432
rect 9815 9401 9827 9404
rect 9769 9395 9827 9401
rect 10870 9392 10876 9404
rect 10928 9392 10934 9444
rect 12526 9432 12532 9444
rect 11256 9404 12532 9432
rect 11256 9376 11284 9404
rect 12526 9392 12532 9404
rect 12584 9432 12590 9444
rect 12805 9435 12863 9441
rect 12805 9432 12817 9435
rect 12584 9404 12817 9432
rect 12584 9392 12590 9404
rect 12805 9401 12817 9404
rect 12851 9432 12863 9435
rect 13449 9435 13507 9441
rect 13449 9432 13461 9435
rect 12851 9404 13461 9432
rect 12851 9401 12863 9404
rect 12805 9395 12863 9401
rect 13449 9401 13461 9404
rect 13495 9401 13507 9435
rect 13449 9395 13507 9401
rect 10321 9367 10379 9373
rect 10321 9333 10333 9367
rect 10367 9364 10379 9367
rect 10410 9364 10416 9376
rect 10367 9336 10416 9364
rect 10367 9333 10379 9336
rect 10321 9327 10379 9333
rect 10410 9324 10416 9336
rect 10468 9324 10474 9376
rect 11238 9324 11244 9376
rect 11296 9364 11302 9376
rect 11882 9364 11888 9376
rect 11296 9336 11341 9364
rect 11843 9336 11888 9364
rect 11296 9324 11302 9336
rect 11882 9324 11888 9336
rect 11940 9324 11946 9376
rect 12158 9364 12164 9376
rect 12119 9336 12164 9364
rect 12158 9324 12164 9336
rect 12216 9324 12222 9376
rect 12437 9367 12495 9373
rect 12437 9333 12449 9367
rect 12483 9364 12495 9367
rect 12710 9364 12716 9376
rect 12483 9336 12716 9364
rect 12483 9333 12495 9336
rect 12437 9327 12495 9333
rect 12710 9324 12716 9336
rect 12768 9324 12774 9376
rect 15010 9364 15016 9376
rect 14971 9336 15016 9364
rect 15010 9324 15016 9336
rect 15068 9324 15074 9376
rect 15194 9324 15200 9376
rect 15252 9364 15258 9376
rect 15304 9373 15332 9472
rect 15473 9469 15485 9472
rect 15519 9469 15531 9503
rect 19242 9500 19248 9512
rect 19203 9472 19248 9500
rect 15473 9463 15531 9469
rect 19242 9460 19248 9472
rect 19300 9460 19306 9512
rect 19444 9500 19472 9531
rect 19794 9528 19800 9580
rect 19852 9568 19858 9580
rect 20625 9571 20683 9577
rect 20625 9568 20637 9571
rect 19852 9540 20637 9568
rect 19852 9528 19858 9540
rect 20625 9537 20637 9540
rect 20671 9537 20683 9571
rect 20625 9531 20683 9537
rect 32490 9528 32496 9580
rect 32548 9568 32554 9580
rect 33413 9571 33471 9577
rect 33413 9568 33425 9571
rect 32548 9540 33425 9568
rect 32548 9528 32554 9540
rect 33413 9537 33425 9540
rect 33459 9568 33471 9571
rect 34149 9571 34207 9577
rect 34149 9568 34161 9571
rect 33459 9540 34161 9568
rect 33459 9537 33471 9540
rect 33413 9531 33471 9537
rect 34149 9537 34161 9540
rect 34195 9537 34207 9571
rect 34149 9531 34207 9537
rect 20898 9500 20904 9512
rect 19352 9472 19472 9500
rect 20859 9472 20904 9500
rect 15746 9441 15752 9444
rect 15740 9432 15752 9441
rect 15707 9404 15752 9432
rect 15740 9395 15752 9404
rect 15746 9392 15752 9395
rect 15804 9392 15810 9444
rect 18138 9392 18144 9444
rect 18196 9432 18202 9444
rect 19352 9432 19380 9472
rect 20898 9460 20904 9472
rect 20956 9460 20962 9512
rect 21168 9503 21226 9509
rect 21168 9500 21180 9503
rect 21008 9472 21180 9500
rect 18196 9404 19380 9432
rect 18196 9392 18202 9404
rect 20162 9392 20168 9444
rect 20220 9432 20226 9444
rect 20533 9435 20591 9441
rect 20533 9432 20545 9435
rect 20220 9404 20545 9432
rect 20220 9392 20226 9404
rect 20533 9401 20545 9404
rect 20579 9432 20591 9435
rect 21008 9432 21036 9472
rect 21168 9469 21180 9472
rect 21214 9500 21226 9503
rect 22002 9500 22008 9512
rect 21214 9472 22008 9500
rect 21214 9469 21226 9472
rect 21168 9463 21226 9469
rect 22002 9460 22008 9472
rect 22060 9460 22066 9512
rect 25317 9503 25375 9509
rect 25317 9469 25329 9503
rect 25363 9469 25375 9503
rect 25317 9463 25375 9469
rect 20579 9404 21036 9432
rect 20579 9401 20591 9404
rect 20533 9395 20591 9401
rect 15289 9367 15347 9373
rect 15289 9364 15301 9367
rect 15252 9336 15301 9364
rect 15252 9324 15258 9336
rect 15289 9333 15301 9336
rect 15335 9333 15347 9367
rect 15289 9327 15347 9333
rect 16298 9324 16304 9376
rect 16356 9364 16362 9376
rect 16853 9367 16911 9373
rect 16853 9364 16865 9367
rect 16356 9336 16865 9364
rect 16356 9324 16362 9336
rect 16853 9333 16865 9336
rect 16899 9333 16911 9367
rect 18874 9364 18880 9376
rect 18835 9336 18880 9364
rect 16853 9327 16911 9333
rect 18874 9324 18880 9336
rect 18932 9324 18938 9376
rect 20438 9364 20444 9376
rect 20399 9336 20444 9364
rect 20438 9324 20444 9336
rect 20496 9324 20502 9376
rect 22278 9364 22284 9376
rect 22239 9336 22284 9364
rect 22278 9324 22284 9336
rect 22336 9324 22342 9376
rect 25225 9367 25283 9373
rect 25225 9333 25237 9367
rect 25271 9364 25283 9367
rect 25332 9364 25360 9463
rect 25406 9460 25412 9512
rect 25464 9500 25470 9512
rect 25573 9503 25631 9509
rect 25573 9500 25585 9503
rect 25464 9472 25585 9500
rect 25464 9460 25470 9472
rect 25573 9469 25585 9472
rect 25619 9469 25631 9503
rect 25573 9463 25631 9469
rect 29914 9460 29920 9512
rect 29972 9500 29978 9512
rect 30285 9503 30343 9509
rect 30285 9500 30297 9503
rect 29972 9472 30297 9500
rect 29972 9460 29978 9472
rect 30285 9469 30297 9472
rect 30331 9500 30343 9503
rect 32306 9500 32312 9512
rect 30331 9472 30788 9500
rect 32219 9472 32312 9500
rect 30331 9469 30343 9472
rect 30285 9463 30343 9469
rect 29730 9392 29736 9444
rect 29788 9432 29794 9444
rect 30558 9441 30564 9444
rect 30530 9435 30564 9441
rect 30530 9432 30542 9435
rect 29788 9404 30542 9432
rect 29788 9392 29794 9404
rect 30530 9401 30542 9404
rect 30616 9432 30622 9444
rect 30616 9404 30678 9432
rect 30530 9395 30564 9401
rect 30558 9392 30564 9395
rect 30616 9392 30622 9404
rect 26510 9364 26516 9376
rect 25271 9336 26516 9364
rect 25271 9333 25283 9336
rect 25225 9327 25283 9333
rect 26510 9324 26516 9336
rect 26568 9324 26574 9376
rect 26694 9364 26700 9376
rect 26655 9336 26700 9364
rect 26694 9324 26700 9336
rect 26752 9324 26758 9376
rect 30193 9367 30251 9373
rect 30193 9333 30205 9367
rect 30239 9364 30251 9367
rect 30760 9364 30788 9472
rect 32306 9460 32312 9472
rect 32364 9500 32370 9512
rect 33137 9503 33195 9509
rect 33137 9500 33149 9503
rect 32364 9472 33149 9500
rect 32364 9460 32370 9472
rect 33137 9469 33149 9472
rect 33183 9500 33195 9503
rect 34514 9500 34520 9512
rect 33183 9472 34520 9500
rect 33183 9469 33195 9472
rect 33137 9463 33195 9469
rect 34514 9460 34520 9472
rect 34572 9460 34578 9512
rect 34882 9500 34888 9512
rect 34843 9472 34888 9500
rect 34882 9460 34888 9472
rect 34940 9460 34946 9512
rect 32858 9392 32864 9444
rect 32916 9432 32922 9444
rect 32916 9404 33272 9432
rect 32916 9392 32922 9404
rect 31018 9364 31024 9376
rect 30239 9336 31024 9364
rect 30239 9333 30251 9336
rect 30193 9327 30251 9333
rect 31018 9324 31024 9336
rect 31076 9324 31082 9376
rect 31110 9324 31116 9376
rect 31168 9364 31174 9376
rect 31665 9367 31723 9373
rect 31665 9364 31677 9367
rect 31168 9336 31677 9364
rect 31168 9324 31174 9336
rect 31665 9333 31677 9336
rect 31711 9333 31723 9367
rect 31665 9327 31723 9333
rect 32769 9367 32827 9373
rect 32769 9333 32781 9367
rect 32815 9364 32827 9367
rect 32950 9364 32956 9376
rect 32815 9336 32956 9364
rect 32815 9333 32827 9336
rect 32769 9327 32827 9333
rect 32950 9324 32956 9336
rect 33008 9324 33014 9376
rect 33244 9373 33272 9404
rect 34422 9392 34428 9444
rect 34480 9432 34486 9444
rect 34790 9432 34796 9444
rect 34480 9404 34796 9432
rect 34480 9392 34486 9404
rect 34790 9392 34796 9404
rect 34848 9432 34854 9444
rect 35130 9435 35188 9441
rect 35130 9432 35142 9435
rect 34848 9404 35142 9432
rect 34848 9392 34854 9404
rect 35130 9401 35142 9404
rect 35176 9401 35188 9435
rect 35130 9395 35188 9401
rect 33229 9367 33287 9373
rect 33229 9333 33241 9367
rect 33275 9364 33287 9367
rect 33318 9364 33324 9376
rect 33275 9336 33324 9364
rect 33275 9333 33287 9336
rect 33229 9327 33287 9333
rect 33318 9324 33324 9336
rect 33376 9324 33382 9376
rect 34606 9324 34612 9376
rect 34664 9364 34670 9376
rect 34701 9367 34759 9373
rect 34701 9364 34713 9367
rect 34664 9336 34713 9364
rect 34664 9324 34670 9336
rect 34701 9333 34713 9336
rect 34747 9364 34759 9367
rect 34882 9364 34888 9376
rect 34747 9336 34888 9364
rect 34747 9333 34759 9336
rect 34701 9327 34759 9333
rect 34882 9324 34888 9336
rect 34940 9324 34946 9376
rect 36262 9364 36268 9376
rect 36223 9336 36268 9364
rect 36262 9324 36268 9336
rect 36320 9324 36326 9376
rect 36814 9364 36820 9376
rect 36775 9336 36820 9364
rect 36814 9324 36820 9336
rect 36872 9324 36878 9376
rect 37090 9324 37096 9376
rect 37148 9364 37154 9376
rect 37369 9367 37427 9373
rect 37369 9364 37381 9367
rect 37148 9336 37381 9364
rect 37148 9324 37154 9336
rect 37369 9333 37381 9336
rect 37415 9333 37427 9367
rect 37369 9327 37427 9333
rect 1104 9274 38824 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 38824 9274
rect 1104 9200 38824 9222
rect 10873 9163 10931 9169
rect 10873 9129 10885 9163
rect 10919 9160 10931 9163
rect 11238 9160 11244 9172
rect 10919 9132 11244 9160
rect 10919 9129 10931 9132
rect 10873 9123 10931 9129
rect 11238 9120 11244 9132
rect 11296 9120 11302 9172
rect 12434 9120 12440 9172
rect 12492 9160 12498 9172
rect 13170 9160 13176 9172
rect 12492 9132 13176 9160
rect 12492 9120 12498 9132
rect 13170 9120 13176 9132
rect 13228 9160 13234 9172
rect 13633 9163 13691 9169
rect 13633 9160 13645 9163
rect 13228 9132 13645 9160
rect 13228 9120 13234 9132
rect 13633 9129 13645 9132
rect 13679 9129 13691 9163
rect 14182 9160 14188 9172
rect 14143 9132 14188 9160
rect 13633 9123 13691 9129
rect 14182 9120 14188 9132
rect 14240 9120 14246 9172
rect 15010 9120 15016 9172
rect 15068 9160 15074 9172
rect 15933 9163 15991 9169
rect 15933 9160 15945 9163
rect 15068 9132 15945 9160
rect 15068 9120 15074 9132
rect 15933 9129 15945 9132
rect 15979 9160 15991 9163
rect 16482 9160 16488 9172
rect 15979 9132 16488 9160
rect 15979 9129 15991 9132
rect 15933 9123 15991 9129
rect 16482 9120 16488 9132
rect 16540 9120 16546 9172
rect 16574 9120 16580 9172
rect 16632 9160 16638 9172
rect 16945 9163 17003 9169
rect 16945 9160 16957 9163
rect 16632 9132 16957 9160
rect 16632 9120 16638 9132
rect 16945 9129 16957 9132
rect 16991 9129 17003 9163
rect 16945 9123 17003 9129
rect 17954 9120 17960 9172
rect 18012 9160 18018 9172
rect 18322 9160 18328 9172
rect 18012 9132 18328 9160
rect 18012 9120 18018 9132
rect 18322 9120 18328 9132
rect 18380 9160 18386 9172
rect 18693 9163 18751 9169
rect 18693 9160 18705 9163
rect 18380 9132 18705 9160
rect 18380 9120 18386 9132
rect 18693 9129 18705 9132
rect 18739 9129 18751 9163
rect 19334 9160 19340 9172
rect 19295 9132 19340 9160
rect 18693 9123 18751 9129
rect 11609 9095 11667 9101
rect 11609 9061 11621 9095
rect 11655 9092 11667 9095
rect 11968 9095 12026 9101
rect 11968 9092 11980 9095
rect 11655 9064 11980 9092
rect 11655 9061 11667 9064
rect 11609 9055 11667 9061
rect 11968 9061 11980 9064
rect 12014 9092 12026 9095
rect 13078 9092 13084 9104
rect 12014 9064 13084 9092
rect 12014 9061 12026 9064
rect 11968 9055 12026 9061
rect 13078 9052 13084 9064
rect 13136 9052 13142 9104
rect 16298 9092 16304 9104
rect 16259 9064 16304 9092
rect 16298 9052 16304 9064
rect 16356 9052 16362 9104
rect 18708 9092 18736 9123
rect 19334 9120 19340 9132
rect 19392 9120 19398 9172
rect 20162 9120 20168 9172
rect 20220 9160 20226 9172
rect 20257 9163 20315 9169
rect 20257 9160 20269 9163
rect 20220 9132 20269 9160
rect 20220 9120 20226 9132
rect 20257 9129 20269 9132
rect 20303 9129 20315 9163
rect 20257 9123 20315 9129
rect 25317 9163 25375 9169
rect 25317 9129 25329 9163
rect 25363 9160 25375 9163
rect 25406 9160 25412 9172
rect 25363 9132 25412 9160
rect 25363 9129 25375 9132
rect 25317 9123 25375 9129
rect 25406 9120 25412 9132
rect 25464 9120 25470 9172
rect 29730 9160 29736 9172
rect 29691 9132 29736 9160
rect 29730 9120 29736 9132
rect 29788 9120 29794 9172
rect 30101 9163 30159 9169
rect 30101 9129 30113 9163
rect 30147 9160 30159 9163
rect 30282 9160 30288 9172
rect 30147 9132 30288 9160
rect 30147 9129 30159 9132
rect 30101 9123 30159 9129
rect 30282 9120 30288 9132
rect 30340 9120 30346 9172
rect 30469 9163 30527 9169
rect 30469 9129 30481 9163
rect 30515 9160 30527 9163
rect 32306 9160 32312 9172
rect 30515 9132 32312 9160
rect 30515 9129 30527 9132
rect 30469 9123 30527 9129
rect 32306 9120 32312 9132
rect 32364 9120 32370 9172
rect 32674 9120 32680 9172
rect 32732 9160 32738 9172
rect 33047 9163 33105 9169
rect 33047 9160 33059 9163
rect 32732 9132 33059 9160
rect 32732 9120 32738 9132
rect 33047 9129 33059 9132
rect 33093 9160 33105 9163
rect 33134 9160 33140 9172
rect 33093 9132 33140 9160
rect 33093 9129 33105 9132
rect 33047 9123 33105 9129
rect 33134 9120 33140 9132
rect 33192 9120 33198 9172
rect 33778 9120 33784 9172
rect 33836 9160 33842 9172
rect 34425 9163 34483 9169
rect 34425 9160 34437 9163
rect 33836 9132 34437 9160
rect 33836 9120 33842 9132
rect 34425 9129 34437 9132
rect 34471 9129 34483 9163
rect 35986 9160 35992 9172
rect 35947 9132 35992 9160
rect 34425 9123 34483 9129
rect 35986 9120 35992 9132
rect 36044 9120 36050 9172
rect 19426 9092 19432 9104
rect 18708 9064 19432 9092
rect 19426 9052 19432 9064
rect 19484 9052 19490 9104
rect 19981 9095 20039 9101
rect 19981 9061 19993 9095
rect 20027 9092 20039 9095
rect 20438 9092 20444 9104
rect 20027 9064 20444 9092
rect 20027 9061 20039 9064
rect 19981 9055 20039 9061
rect 20438 9052 20444 9064
rect 20496 9092 20502 9104
rect 21168 9095 21226 9101
rect 21168 9092 21180 9095
rect 20496 9064 21180 9092
rect 20496 9052 20502 9064
rect 21168 9061 21180 9064
rect 21214 9092 21226 9095
rect 21358 9092 21364 9104
rect 21214 9064 21364 9092
rect 21214 9061 21226 9064
rect 21168 9055 21226 9061
rect 21358 9052 21364 9064
rect 21416 9092 21422 9104
rect 22278 9092 22284 9104
rect 21416 9064 22284 9092
rect 21416 9052 21422 9064
rect 22278 9052 22284 9064
rect 22336 9052 22342 9104
rect 25225 9095 25283 9101
rect 25225 9061 25237 9095
rect 25271 9092 25283 9095
rect 26694 9092 26700 9104
rect 25271 9064 26700 9092
rect 25271 9061 25283 9064
rect 25225 9055 25283 9061
rect 26694 9052 26700 9064
rect 26752 9101 26758 9104
rect 26752 9095 26816 9101
rect 26752 9061 26770 9095
rect 26804 9061 26816 9095
rect 26752 9055 26816 9061
rect 26752 9052 26758 9055
rect 30006 9052 30012 9104
rect 30064 9092 30070 9104
rect 30929 9095 30987 9101
rect 30929 9092 30941 9095
rect 30064 9064 30941 9092
rect 30064 9052 30070 9064
rect 30929 9061 30941 9064
rect 30975 9061 30987 9095
rect 30929 9055 30987 9061
rect 6914 8984 6920 9036
rect 6972 9024 6978 9036
rect 7190 9033 7196 9036
rect 7184 9024 7196 9033
rect 6972 8996 7017 9024
rect 7151 8996 7196 9024
rect 6972 8984 6978 8996
rect 7184 8987 7196 8996
rect 7190 8984 7196 8987
rect 7248 8984 7254 9036
rect 11698 9024 11704 9036
rect 11659 8996 11704 9024
rect 11698 8984 11704 8996
rect 11756 8984 11762 9036
rect 17954 8984 17960 9036
rect 18012 9024 18018 9036
rect 18601 9027 18659 9033
rect 18601 9024 18613 9027
rect 18012 8996 18613 9024
rect 18012 8984 18018 8996
rect 18601 8993 18613 8996
rect 18647 9024 18659 9027
rect 18874 9024 18880 9036
rect 18647 8996 18880 9024
rect 18647 8993 18659 8996
rect 18601 8987 18659 8993
rect 18874 8984 18880 8996
rect 18932 8984 18938 9036
rect 30834 9024 30840 9036
rect 30795 8996 30840 9024
rect 30834 8984 30840 8996
rect 30892 8984 30898 9036
rect 32398 9024 32404 9036
rect 32359 8996 32404 9024
rect 32398 8984 32404 8996
rect 32456 9024 32462 9036
rect 32585 9027 32643 9033
rect 32585 9024 32597 9027
rect 32456 8996 32597 9024
rect 32456 8984 32462 8996
rect 32585 8993 32597 8996
rect 32631 8993 32643 9027
rect 32585 8987 32643 8993
rect 35897 9027 35955 9033
rect 35897 8993 35909 9027
rect 35943 9024 35955 9027
rect 37090 9024 37096 9036
rect 35943 8996 37096 9024
rect 35943 8993 35955 8996
rect 35897 8987 35955 8993
rect 37090 8984 37096 8996
rect 37148 8984 37154 9036
rect 9953 8959 10011 8965
rect 9953 8925 9965 8959
rect 9999 8956 10011 8959
rect 10134 8956 10140 8968
rect 9999 8928 10140 8956
rect 9999 8925 10011 8928
rect 9953 8919 10011 8925
rect 10134 8916 10140 8928
rect 10192 8916 10198 8968
rect 15565 8959 15623 8965
rect 15565 8925 15577 8959
rect 15611 8956 15623 8959
rect 15746 8956 15752 8968
rect 15611 8928 15752 8956
rect 15611 8925 15623 8928
rect 15565 8919 15623 8925
rect 15746 8916 15752 8928
rect 15804 8956 15810 8968
rect 16393 8959 16451 8965
rect 16393 8956 16405 8959
rect 15804 8928 16405 8956
rect 15804 8916 15810 8928
rect 16393 8925 16405 8928
rect 16439 8956 16451 8959
rect 16482 8956 16488 8968
rect 16439 8928 16488 8956
rect 16439 8925 16451 8928
rect 16393 8919 16451 8925
rect 16482 8916 16488 8928
rect 16540 8916 16546 8968
rect 16577 8959 16635 8965
rect 16577 8925 16589 8959
rect 16623 8956 16635 8959
rect 16666 8956 16672 8968
rect 16623 8928 16672 8956
rect 16623 8925 16635 8928
rect 16577 8919 16635 8925
rect 16666 8916 16672 8928
rect 16724 8916 16730 8968
rect 18782 8916 18788 8968
rect 18840 8956 18846 8968
rect 20717 8959 20775 8965
rect 18840 8928 18885 8956
rect 18840 8916 18846 8928
rect 20717 8925 20729 8959
rect 20763 8956 20775 8959
rect 20898 8956 20904 8968
rect 20763 8928 20904 8956
rect 20763 8925 20775 8928
rect 20717 8919 20775 8925
rect 20898 8916 20904 8928
rect 20956 8916 20962 8968
rect 25409 8959 25467 8965
rect 25409 8956 25421 8959
rect 24780 8928 25421 8956
rect 17862 8848 17868 8900
rect 17920 8888 17926 8900
rect 18233 8891 18291 8897
rect 18233 8888 18245 8891
rect 17920 8860 18245 8888
rect 17920 8848 17926 8860
rect 18233 8857 18245 8860
rect 18279 8857 18291 8891
rect 18233 8851 18291 8857
rect 24780 8832 24808 8928
rect 25409 8925 25421 8928
rect 25455 8925 25467 8959
rect 26510 8956 26516 8968
rect 26471 8928 26516 8956
rect 25409 8919 25467 8925
rect 26510 8916 26516 8928
rect 26568 8916 26574 8968
rect 31110 8956 31116 8968
rect 31071 8928 31116 8956
rect 31110 8916 31116 8928
rect 31168 8916 31174 8968
rect 33042 8956 33048 8968
rect 33003 8928 33048 8956
rect 33042 8916 33048 8928
rect 33100 8916 33106 8968
rect 33318 8956 33324 8968
rect 33279 8928 33324 8956
rect 33318 8916 33324 8928
rect 33376 8916 33382 8968
rect 34606 8916 34612 8968
rect 34664 8956 34670 8968
rect 35710 8956 35716 8968
rect 34664 8928 35716 8956
rect 34664 8916 34670 8928
rect 35710 8916 35716 8928
rect 35768 8916 35774 8968
rect 36173 8959 36231 8965
rect 36173 8925 36185 8959
rect 36219 8956 36231 8959
rect 36262 8956 36268 8968
rect 36219 8928 36268 8956
rect 36219 8925 36231 8928
rect 36173 8919 36231 8925
rect 36262 8916 36268 8928
rect 36320 8916 36326 8968
rect 8294 8820 8300 8832
rect 8255 8792 8300 8820
rect 8294 8780 8300 8792
rect 8352 8780 8358 8832
rect 11241 8823 11299 8829
rect 11241 8789 11253 8823
rect 11287 8820 11299 8823
rect 11422 8820 11428 8832
rect 11287 8792 11428 8820
rect 11287 8789 11299 8792
rect 11241 8783 11299 8789
rect 11422 8780 11428 8792
rect 11480 8780 11486 8832
rect 13081 8823 13139 8829
rect 13081 8789 13093 8823
rect 13127 8820 13139 8823
rect 13722 8820 13728 8832
rect 13127 8792 13728 8820
rect 13127 8789 13139 8792
rect 13081 8783 13139 8789
rect 13722 8780 13728 8792
rect 13780 8780 13786 8832
rect 17681 8823 17739 8829
rect 17681 8789 17693 8823
rect 17727 8820 17739 8823
rect 18138 8820 18144 8832
rect 17727 8792 18144 8820
rect 17727 8789 17739 8792
rect 17681 8783 17739 8789
rect 18138 8780 18144 8792
rect 18196 8780 18202 8832
rect 22278 8820 22284 8832
rect 22239 8792 22284 8820
rect 22278 8780 22284 8792
rect 22336 8780 22342 8832
rect 24302 8820 24308 8832
rect 24263 8792 24308 8820
rect 24302 8780 24308 8792
rect 24360 8780 24366 8832
rect 24762 8820 24768 8832
rect 24723 8792 24768 8820
rect 24762 8780 24768 8792
rect 24820 8780 24826 8832
rect 24857 8823 24915 8829
rect 24857 8789 24869 8823
rect 24903 8820 24915 8823
rect 25314 8820 25320 8832
rect 24903 8792 25320 8820
rect 24903 8789 24915 8792
rect 24857 8783 24915 8789
rect 25314 8780 25320 8792
rect 25372 8780 25378 8832
rect 26329 8823 26387 8829
rect 26329 8789 26341 8823
rect 26375 8820 26387 8823
rect 26878 8820 26884 8832
rect 26375 8792 26884 8820
rect 26375 8789 26387 8792
rect 26329 8783 26387 8789
rect 26878 8780 26884 8792
rect 26936 8820 26942 8832
rect 27893 8823 27951 8829
rect 27893 8820 27905 8823
rect 26936 8792 27905 8820
rect 26936 8780 26942 8792
rect 27893 8789 27905 8792
rect 27939 8789 27951 8823
rect 27893 8783 27951 8789
rect 34790 8780 34796 8832
rect 34848 8820 34854 8832
rect 35161 8823 35219 8829
rect 35161 8820 35173 8823
rect 34848 8792 35173 8820
rect 34848 8780 34854 8792
rect 35161 8789 35173 8792
rect 35207 8789 35219 8823
rect 35161 8783 35219 8789
rect 35434 8780 35440 8832
rect 35492 8820 35498 8832
rect 35529 8823 35587 8829
rect 35529 8820 35541 8823
rect 35492 8792 35541 8820
rect 35492 8780 35498 8792
rect 35529 8789 35541 8792
rect 35575 8820 35587 8823
rect 35710 8820 35716 8832
rect 35575 8792 35716 8820
rect 35575 8789 35587 8792
rect 35529 8783 35587 8789
rect 35710 8780 35716 8792
rect 35768 8780 35774 8832
rect 1104 8730 38824 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 34966 8730
rect 35018 8678 35030 8730
rect 35082 8678 35094 8730
rect 35146 8678 35158 8730
rect 35210 8678 38824 8730
rect 1104 8656 38824 8678
rect 6273 8619 6331 8625
rect 6273 8585 6285 8619
rect 6319 8616 6331 8619
rect 7190 8616 7196 8628
rect 6319 8588 7196 8616
rect 6319 8585 6331 8588
rect 6273 8579 6331 8585
rect 7190 8576 7196 8588
rect 7248 8576 7254 8628
rect 11238 8616 11244 8628
rect 11199 8588 11244 8616
rect 11238 8576 11244 8588
rect 11296 8616 11302 8628
rect 12158 8616 12164 8628
rect 11296 8588 12164 8616
rect 11296 8576 11302 8588
rect 12158 8576 12164 8588
rect 12216 8576 12222 8628
rect 12618 8576 12624 8628
rect 12676 8616 12682 8628
rect 14553 8619 14611 8625
rect 14553 8616 14565 8619
rect 12676 8588 14565 8616
rect 12676 8576 12682 8588
rect 14553 8585 14565 8588
rect 14599 8585 14611 8619
rect 16298 8616 16304 8628
rect 16259 8588 16304 8616
rect 14553 8579 14611 8585
rect 16298 8576 16304 8588
rect 16356 8576 16362 8628
rect 18322 8616 18328 8628
rect 18283 8588 18328 8616
rect 18322 8576 18328 8588
rect 18380 8576 18386 8628
rect 19334 8576 19340 8628
rect 19392 8616 19398 8628
rect 20441 8619 20499 8625
rect 20441 8616 20453 8619
rect 19392 8588 20453 8616
rect 19392 8576 19398 8588
rect 20441 8585 20453 8588
rect 20487 8585 20499 8619
rect 21358 8616 21364 8628
rect 21319 8588 21364 8616
rect 20441 8579 20499 8585
rect 21358 8576 21364 8588
rect 21416 8576 21422 8628
rect 25406 8576 25412 8628
rect 25464 8616 25470 8628
rect 25593 8619 25651 8625
rect 25593 8616 25605 8619
rect 25464 8588 25605 8616
rect 25464 8576 25470 8588
rect 25593 8585 25605 8588
rect 25639 8585 25651 8619
rect 25593 8579 25651 8585
rect 27614 8576 27620 8628
rect 27672 8616 27678 8628
rect 28077 8619 28135 8625
rect 28077 8616 28089 8619
rect 27672 8588 28089 8616
rect 27672 8576 27678 8588
rect 28077 8585 28089 8588
rect 28123 8585 28135 8619
rect 30006 8616 30012 8628
rect 29967 8588 30012 8616
rect 28077 8579 28135 8585
rect 30006 8576 30012 8588
rect 30064 8576 30070 8628
rect 30653 8619 30711 8625
rect 30653 8585 30665 8619
rect 30699 8616 30711 8619
rect 30834 8616 30840 8628
rect 30699 8588 30840 8616
rect 30699 8585 30711 8588
rect 30653 8579 30711 8585
rect 12250 8548 12256 8560
rect 12211 8520 12256 8548
rect 12250 8508 12256 8520
rect 12308 8508 12314 8560
rect 15657 8551 15715 8557
rect 15657 8517 15669 8551
rect 15703 8548 15715 8551
rect 16666 8548 16672 8560
rect 15703 8520 16672 8548
rect 15703 8517 15715 8520
rect 15657 8511 15715 8517
rect 16666 8508 16672 8520
rect 16724 8548 16730 8560
rect 16945 8551 17003 8557
rect 16945 8548 16957 8551
rect 16724 8520 16957 8548
rect 16724 8508 16730 8520
rect 16945 8517 16957 8520
rect 16991 8517 17003 8551
rect 16945 8511 17003 8517
rect 4706 8480 4712 8492
rect 4667 8452 4712 8480
rect 4706 8440 4712 8452
rect 4764 8440 4770 8492
rect 12713 8483 12771 8489
rect 12713 8449 12725 8483
rect 12759 8480 12771 8483
rect 12894 8480 12900 8492
rect 12759 8452 12900 8480
rect 12759 8449 12771 8452
rect 12713 8443 12771 8449
rect 12894 8440 12900 8452
rect 12952 8440 12958 8492
rect 13170 8480 13176 8492
rect 13131 8452 13176 8480
rect 13170 8440 13176 8452
rect 13228 8440 13234 8492
rect 13446 8480 13452 8492
rect 13407 8452 13452 8480
rect 13446 8440 13452 8452
rect 13504 8440 13510 8492
rect 30101 8483 30159 8489
rect 30101 8449 30113 8483
rect 30147 8480 30159 8483
rect 30668 8480 30696 8579
rect 30834 8576 30840 8588
rect 30892 8576 30898 8628
rect 32490 8616 32496 8628
rect 32451 8588 32496 8616
rect 32490 8576 32496 8588
rect 32548 8576 32554 8628
rect 33042 8576 33048 8628
rect 33100 8616 33106 8628
rect 33413 8619 33471 8625
rect 33413 8616 33425 8619
rect 33100 8588 33425 8616
rect 33100 8576 33106 8588
rect 33413 8585 33425 8588
rect 33459 8585 33471 8619
rect 33413 8579 33471 8585
rect 35802 8576 35808 8628
rect 35860 8616 35866 8628
rect 36449 8619 36507 8625
rect 36449 8616 36461 8619
rect 35860 8588 36461 8616
rect 35860 8576 35866 8588
rect 36449 8585 36461 8588
rect 36495 8616 36507 8619
rect 36814 8616 36820 8628
rect 36495 8588 36820 8616
rect 36495 8585 36507 8588
rect 36449 8579 36507 8585
rect 36814 8576 36820 8588
rect 36872 8576 36878 8628
rect 37090 8616 37096 8628
rect 37051 8588 37096 8616
rect 37090 8576 37096 8588
rect 37148 8576 37154 8628
rect 31018 8480 31024 8492
rect 30147 8452 30696 8480
rect 30931 8452 31024 8480
rect 30147 8449 30159 8452
rect 30101 8443 30159 8449
rect 31018 8440 31024 8452
rect 31076 8480 31082 8492
rect 31113 8483 31171 8489
rect 31113 8480 31125 8483
rect 31076 8452 31125 8480
rect 31076 8440 31082 8452
rect 31113 8449 31125 8452
rect 31159 8449 31171 8483
rect 31113 8443 31171 8449
rect 34333 8483 34391 8489
rect 34333 8449 34345 8483
rect 34379 8480 34391 8483
rect 34379 8452 35204 8480
rect 34379 8449 34391 8452
rect 34333 8443 34391 8449
rect 35176 8424 35204 8452
rect 3973 8415 4031 8421
rect 3973 8381 3985 8415
rect 4019 8412 4031 8415
rect 4525 8415 4583 8421
rect 4525 8412 4537 8415
rect 4019 8384 4537 8412
rect 4019 8381 4031 8384
rect 3973 8375 4031 8381
rect 4525 8381 4537 8384
rect 4571 8412 4583 8415
rect 5350 8412 5356 8424
rect 4571 8384 5356 8412
rect 4571 8381 4583 8384
rect 4525 8375 4583 8381
rect 5350 8372 5356 8384
rect 5408 8412 5414 8424
rect 6825 8415 6883 8421
rect 6825 8412 6837 8415
rect 5408 8384 5580 8412
rect 5408 8372 5414 8384
rect 3050 8304 3056 8356
rect 3108 8344 3114 8356
rect 3605 8347 3663 8353
rect 3605 8344 3617 8347
rect 3108 8316 3617 8344
rect 3108 8304 3114 8316
rect 3605 8313 3617 8316
rect 3651 8344 3663 8347
rect 4433 8347 4491 8353
rect 4433 8344 4445 8347
rect 3651 8316 4445 8344
rect 3651 8313 3663 8316
rect 3605 8307 3663 8313
rect 4433 8313 4445 8316
rect 4479 8344 4491 8347
rect 5442 8344 5448 8356
rect 4479 8316 5448 8344
rect 4479 8313 4491 8316
rect 4433 8307 4491 8313
rect 5442 8304 5448 8316
rect 5500 8304 5506 8356
rect 4062 8276 4068 8288
rect 4023 8248 4068 8276
rect 4062 8236 4068 8248
rect 4120 8236 4126 8288
rect 5552 8276 5580 8384
rect 6564 8384 6837 8412
rect 6564 8288 6592 8384
rect 6825 8381 6837 8384
rect 6871 8412 6883 8415
rect 6914 8412 6920 8424
rect 6871 8384 6920 8412
rect 6871 8381 6883 8384
rect 6825 8375 6883 8381
rect 6914 8372 6920 8384
rect 6972 8372 6978 8424
rect 9769 8415 9827 8421
rect 9769 8381 9781 8415
rect 9815 8412 9827 8415
rect 9861 8415 9919 8421
rect 9861 8412 9873 8415
rect 9815 8384 9873 8412
rect 9815 8381 9827 8384
rect 9769 8375 9827 8381
rect 9861 8381 9873 8384
rect 9907 8412 9919 8415
rect 10502 8412 10508 8424
rect 9907 8384 10508 8412
rect 9907 8381 9919 8384
rect 9861 8375 9919 8381
rect 10502 8372 10508 8384
rect 10560 8412 10566 8424
rect 11698 8412 11704 8424
rect 10560 8384 11704 8412
rect 10560 8372 10566 8384
rect 11698 8372 11704 8384
rect 11756 8412 11762 8424
rect 11793 8415 11851 8421
rect 11793 8412 11805 8415
rect 11756 8384 11805 8412
rect 11756 8372 11762 8384
rect 11793 8381 11805 8384
rect 11839 8381 11851 8415
rect 11793 8375 11851 8381
rect 12802 8372 12808 8424
rect 12860 8412 12866 8424
rect 13036 8415 13094 8421
rect 13036 8412 13048 8415
rect 12860 8384 13048 8412
rect 12860 8372 12866 8384
rect 13036 8381 13048 8384
rect 13082 8381 13094 8415
rect 13036 8375 13094 8381
rect 16761 8415 16819 8421
rect 16761 8381 16773 8415
rect 16807 8381 16819 8415
rect 16761 8375 16819 8381
rect 17865 8415 17923 8421
rect 17865 8381 17877 8415
rect 17911 8412 17923 8415
rect 17954 8412 17960 8424
rect 17911 8384 17960 8412
rect 17911 8381 17923 8384
rect 17865 8375 17923 8381
rect 7092 8347 7150 8353
rect 7092 8313 7104 8347
rect 7138 8344 7150 8347
rect 7282 8344 7288 8356
rect 7138 8316 7288 8344
rect 7138 8313 7150 8316
rect 7092 8307 7150 8313
rect 7282 8304 7288 8316
rect 7340 8304 7346 8356
rect 9950 8304 9956 8356
rect 10008 8344 10014 8356
rect 10128 8347 10186 8353
rect 10128 8344 10140 8347
rect 10008 8316 10140 8344
rect 10008 8304 10014 8316
rect 10128 8313 10140 8316
rect 10174 8344 10186 8347
rect 11422 8344 11428 8356
rect 10174 8316 11428 8344
rect 10174 8313 10186 8316
rect 10128 8307 10186 8313
rect 11422 8304 11428 8316
rect 11480 8304 11486 8356
rect 16025 8347 16083 8353
rect 16025 8313 16037 8347
rect 16071 8344 16083 8347
rect 16482 8344 16488 8356
rect 16071 8316 16488 8344
rect 16071 8313 16083 8316
rect 16025 8307 16083 8313
rect 16482 8304 16488 8316
rect 16540 8304 16546 8356
rect 16776 8344 16804 8375
rect 17954 8372 17960 8384
rect 18012 8372 18018 8424
rect 18046 8372 18052 8424
rect 18104 8412 18110 8424
rect 18969 8415 19027 8421
rect 18969 8412 18981 8415
rect 18104 8384 18981 8412
rect 18104 8372 18110 8384
rect 18969 8381 18981 8384
rect 19015 8412 19027 8415
rect 19061 8415 19119 8421
rect 19061 8412 19073 8415
rect 19015 8384 19073 8412
rect 19015 8381 19027 8384
rect 18969 8375 19027 8381
rect 19061 8381 19073 8384
rect 19107 8381 19119 8415
rect 19061 8375 19119 8381
rect 24213 8415 24271 8421
rect 24213 8381 24225 8415
rect 24259 8381 24271 8415
rect 24213 8375 24271 8381
rect 17405 8347 17463 8353
rect 17405 8344 17417 8347
rect 16776 8316 17417 8344
rect 17405 8313 17417 8316
rect 17451 8344 17463 8347
rect 18322 8344 18328 8356
rect 17451 8316 18328 8344
rect 17451 8313 17463 8316
rect 17405 8307 17463 8313
rect 18322 8304 18328 8316
rect 18380 8304 18386 8356
rect 19334 8353 19340 8356
rect 19328 8344 19340 8353
rect 19295 8316 19340 8344
rect 19328 8307 19340 8316
rect 19334 8304 19340 8307
rect 19392 8304 19398 8356
rect 20898 8304 20904 8356
rect 20956 8344 20962 8356
rect 21085 8347 21143 8353
rect 21085 8344 21097 8347
rect 20956 8316 21097 8344
rect 20956 8304 20962 8316
rect 21085 8313 21097 8316
rect 21131 8344 21143 8347
rect 21131 8316 22140 8344
rect 21131 8313 21143 8316
rect 21085 8307 21143 8313
rect 6362 8276 6368 8288
rect 5552 8248 6368 8276
rect 6362 8236 6368 8248
rect 6420 8236 6426 8288
rect 6546 8276 6552 8288
rect 6507 8248 6552 8276
rect 6546 8236 6552 8248
rect 6604 8236 6610 8288
rect 7926 8236 7932 8288
rect 7984 8276 7990 8288
rect 8205 8279 8263 8285
rect 8205 8276 8217 8279
rect 7984 8248 8217 8276
rect 7984 8236 7990 8248
rect 8205 8245 8217 8248
rect 8251 8245 8263 8279
rect 16500 8276 16528 8304
rect 22112 8288 22140 8316
rect 23474 8304 23480 8356
rect 23532 8344 23538 8356
rect 24121 8347 24179 8353
rect 24121 8344 24133 8347
rect 23532 8316 24133 8344
rect 23532 8304 23538 8316
rect 24121 8313 24133 8316
rect 24167 8344 24179 8347
rect 24228 8344 24256 8375
rect 24302 8372 24308 8424
rect 24360 8412 24366 8424
rect 24469 8415 24527 8421
rect 24469 8412 24481 8415
rect 24360 8384 24481 8412
rect 24360 8372 24366 8384
rect 24469 8381 24481 8384
rect 24515 8381 24527 8415
rect 26697 8415 26755 8421
rect 26697 8412 26709 8415
rect 24469 8375 24527 8381
rect 26528 8384 26709 8412
rect 24167 8316 26280 8344
rect 24167 8313 24179 8316
rect 24121 8307 24179 8313
rect 16666 8276 16672 8288
rect 16500 8248 16672 8276
rect 8205 8239 8263 8245
rect 16666 8236 16672 8248
rect 16724 8236 16730 8288
rect 22094 8236 22100 8288
rect 22152 8236 22158 8288
rect 26252 8285 26280 8316
rect 26528 8288 26556 8384
rect 26697 8381 26709 8384
rect 26743 8381 26755 8415
rect 26697 8375 26755 8381
rect 35069 8415 35127 8421
rect 35069 8381 35081 8415
rect 35115 8381 35127 8415
rect 35069 8375 35127 8381
rect 26878 8304 26884 8356
rect 26936 8353 26942 8356
rect 26936 8347 27000 8353
rect 26936 8313 26954 8347
rect 26988 8313 27000 8347
rect 31358 8347 31416 8353
rect 31358 8344 31370 8347
rect 26936 8307 27000 8313
rect 31128 8316 31370 8344
rect 26936 8304 26942 8307
rect 31128 8288 31156 8316
rect 31358 8313 31370 8316
rect 31404 8313 31416 8347
rect 33134 8344 33140 8356
rect 33047 8316 33140 8344
rect 31358 8307 31416 8313
rect 33134 8304 33140 8316
rect 33192 8344 33198 8356
rect 34330 8344 34336 8356
rect 33192 8316 34336 8344
rect 33192 8304 33198 8316
rect 34330 8304 34336 8316
rect 34388 8304 34394 8356
rect 34609 8347 34667 8353
rect 34609 8344 34621 8347
rect 34440 8316 34621 8344
rect 26237 8279 26295 8285
rect 26237 8245 26249 8279
rect 26283 8276 26295 8279
rect 26510 8276 26516 8288
rect 26283 8248 26516 8276
rect 26283 8245 26295 8248
rect 26237 8239 26295 8245
rect 26510 8236 26516 8248
rect 26568 8236 26574 8288
rect 31110 8236 31116 8288
rect 31168 8236 31174 8288
rect 33594 8276 33600 8288
rect 33555 8248 33600 8276
rect 33594 8236 33600 8248
rect 33652 8236 33658 8288
rect 33962 8236 33968 8288
rect 34020 8276 34026 8288
rect 34440 8276 34468 8316
rect 34609 8313 34621 8316
rect 34655 8344 34667 8347
rect 34790 8344 34796 8356
rect 34655 8316 34796 8344
rect 34655 8313 34667 8316
rect 34609 8307 34667 8313
rect 34790 8304 34796 8316
rect 34848 8344 34854 8356
rect 35084 8344 35112 8375
rect 35158 8372 35164 8424
rect 35216 8412 35222 8424
rect 35336 8415 35394 8421
rect 35336 8412 35348 8415
rect 35216 8384 35348 8412
rect 35216 8372 35222 8384
rect 35336 8381 35348 8384
rect 35382 8412 35394 8415
rect 36262 8412 36268 8424
rect 35382 8384 36268 8412
rect 35382 8381 35394 8384
rect 35336 8375 35394 8381
rect 36262 8372 36268 8384
rect 36320 8372 36326 8424
rect 34848 8316 35112 8344
rect 34848 8304 34854 8316
rect 34020 8248 34468 8276
rect 34020 8236 34026 8248
rect 1104 8186 38824 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 38824 8186
rect 1104 8112 38824 8134
rect 6362 8072 6368 8084
rect 6323 8044 6368 8072
rect 6362 8032 6368 8044
rect 6420 8032 6426 8084
rect 7926 8072 7932 8084
rect 7887 8044 7932 8072
rect 7926 8032 7932 8044
rect 7984 8032 7990 8084
rect 9950 8072 9956 8084
rect 9911 8044 9956 8072
rect 9950 8032 9956 8044
rect 10008 8032 10014 8084
rect 12802 8072 12808 8084
rect 12763 8044 12808 8072
rect 12802 8032 12808 8044
rect 12860 8032 12866 8084
rect 16666 8072 16672 8084
rect 16627 8044 16672 8072
rect 16666 8032 16672 8044
rect 16724 8032 16730 8084
rect 21082 8072 21088 8084
rect 21043 8044 21088 8072
rect 21082 8032 21088 8044
rect 21140 8032 21146 8084
rect 24302 8032 24308 8084
rect 24360 8072 24366 8084
rect 24670 8072 24676 8084
rect 24360 8044 24676 8072
rect 24360 8032 24366 8044
rect 24670 8032 24676 8044
rect 24728 8072 24734 8084
rect 24765 8075 24823 8081
rect 24765 8072 24777 8075
rect 24728 8044 24777 8072
rect 24728 8032 24734 8044
rect 24765 8041 24777 8044
rect 24811 8041 24823 8075
rect 25406 8072 25412 8084
rect 25367 8044 25412 8072
rect 24765 8035 24823 8041
rect 25406 8032 25412 8044
rect 25464 8032 25470 8084
rect 25777 8075 25835 8081
rect 25777 8041 25789 8075
rect 25823 8072 25835 8075
rect 26329 8075 26387 8081
rect 26329 8072 26341 8075
rect 25823 8044 26341 8072
rect 25823 8041 25835 8044
rect 25777 8035 25835 8041
rect 26329 8041 26341 8044
rect 26375 8072 26387 8075
rect 26694 8072 26700 8084
rect 26375 8044 26700 8072
rect 26375 8041 26387 8044
rect 26329 8035 26387 8041
rect 26694 8032 26700 8044
rect 26752 8032 26758 8084
rect 26878 8032 26884 8084
rect 26936 8072 26942 8084
rect 27065 8075 27123 8081
rect 27065 8072 27077 8075
rect 26936 8044 27077 8072
rect 26936 8032 26942 8044
rect 27065 8041 27077 8044
rect 27111 8041 27123 8075
rect 27065 8035 27123 8041
rect 30561 8075 30619 8081
rect 30561 8041 30573 8075
rect 30607 8072 30619 8075
rect 31110 8072 31116 8084
rect 30607 8044 31116 8072
rect 30607 8041 30619 8044
rect 30561 8035 30619 8041
rect 31110 8032 31116 8044
rect 31168 8032 31174 8084
rect 34333 8075 34391 8081
rect 34333 8041 34345 8075
rect 34379 8072 34391 8075
rect 34422 8072 34428 8084
rect 34379 8044 34428 8072
rect 34379 8041 34391 8044
rect 34333 8035 34391 8041
rect 34422 8032 34428 8044
rect 34480 8032 34486 8084
rect 34977 8075 35035 8081
rect 34977 8041 34989 8075
rect 35023 8072 35035 8075
rect 35158 8072 35164 8084
rect 35023 8044 35164 8072
rect 35023 8041 35035 8044
rect 34977 8035 35035 8041
rect 35158 8032 35164 8044
rect 35216 8032 35222 8084
rect 35345 8075 35403 8081
rect 35345 8041 35357 8075
rect 35391 8072 35403 8075
rect 35897 8075 35955 8081
rect 35897 8072 35909 8075
rect 35391 8044 35909 8072
rect 35391 8041 35403 8044
rect 35345 8035 35403 8041
rect 35897 8041 35909 8044
rect 35943 8041 35955 8075
rect 35897 8035 35955 8041
rect 12710 7964 12716 8016
rect 12768 8004 12774 8016
rect 13446 8004 13452 8016
rect 12768 7976 13452 8004
rect 12768 7964 12774 7976
rect 13446 7964 13452 7976
rect 13504 7964 13510 8016
rect 15470 7964 15476 8016
rect 15528 8013 15534 8016
rect 15528 8007 15592 8013
rect 15528 7973 15546 8007
rect 15580 7973 15592 8007
rect 17402 8004 17408 8016
rect 17363 7976 17408 8004
rect 15528 7967 15592 7973
rect 15528 7964 15534 7967
rect 17402 7964 17408 7976
rect 17460 7964 17466 8016
rect 19153 8007 19211 8013
rect 19153 7973 19165 8007
rect 19199 8004 19211 8007
rect 19334 8004 19340 8016
rect 19199 7976 19340 8004
rect 19199 7973 19211 7976
rect 19153 7967 19211 7973
rect 19334 7964 19340 7976
rect 19392 8004 19398 8016
rect 19705 8007 19763 8013
rect 19705 8004 19717 8007
rect 19392 7976 19717 8004
rect 19392 7964 19398 7976
rect 19705 7973 19717 7976
rect 19751 8004 19763 8007
rect 20438 8004 20444 8016
rect 19751 7976 20444 8004
rect 19751 7973 19763 7976
rect 19705 7967 19763 7973
rect 20438 7964 20444 7976
rect 20496 7964 20502 8016
rect 23293 8007 23351 8013
rect 23293 7973 23305 8007
rect 23339 8004 23351 8007
rect 23566 8004 23572 8016
rect 23339 7976 23572 8004
rect 23339 7973 23351 7976
rect 23293 7967 23351 7973
rect 23566 7964 23572 7976
rect 23624 8013 23630 8016
rect 23624 8007 23688 8013
rect 23624 7973 23642 8007
rect 23676 7973 23688 8007
rect 26970 8004 26976 8016
rect 26883 7976 26976 8004
rect 23624 7967 23688 7973
rect 23624 7964 23630 7967
rect 26970 7964 26976 7976
rect 27028 8004 27034 8016
rect 27522 8004 27528 8016
rect 27028 7976 27528 8004
rect 27028 7964 27034 7976
rect 27522 7964 27528 7976
rect 27580 7964 27586 8016
rect 34514 7964 34520 8016
rect 34572 8004 34578 8016
rect 35360 8004 35388 8035
rect 35986 8032 35992 8084
rect 36044 8072 36050 8084
rect 36449 8075 36507 8081
rect 36449 8072 36461 8075
rect 36044 8044 36461 8072
rect 36044 8032 36050 8044
rect 36449 8041 36461 8044
rect 36495 8041 36507 8075
rect 36449 8035 36507 8041
rect 34572 7976 35388 8004
rect 34572 7964 34578 7976
rect 5258 7945 5264 7948
rect 5252 7936 5264 7945
rect 5171 7908 5264 7936
rect 5252 7899 5264 7908
rect 5316 7936 5322 7948
rect 7837 7939 7895 7945
rect 7837 7936 7849 7939
rect 5316 7908 7849 7936
rect 5258 7896 5264 7899
rect 5316 7896 5322 7908
rect 7837 7905 7849 7908
rect 7883 7936 7895 7939
rect 8202 7936 8208 7948
rect 7883 7908 8208 7936
rect 7883 7905 7895 7908
rect 7837 7899 7895 7905
rect 8202 7896 8208 7908
rect 8260 7896 8266 7948
rect 10413 7939 10471 7945
rect 10413 7905 10425 7939
rect 10459 7936 10471 7939
rect 10772 7939 10830 7945
rect 10772 7936 10784 7939
rect 10459 7908 10784 7936
rect 10459 7905 10471 7908
rect 10413 7899 10471 7905
rect 10772 7905 10784 7908
rect 10818 7936 10830 7939
rect 10818 7908 11928 7936
rect 10818 7905 10830 7908
rect 10772 7899 10830 7905
rect 4982 7868 4988 7880
rect 4943 7840 4988 7868
rect 4982 7828 4988 7840
rect 5040 7828 5046 7880
rect 8021 7871 8079 7877
rect 8021 7837 8033 7871
rect 8067 7837 8079 7871
rect 10502 7868 10508 7880
rect 10463 7840 10508 7868
rect 8021 7831 8079 7837
rect 7374 7760 7380 7812
rect 7432 7800 7438 7812
rect 8036 7800 8064 7831
rect 10502 7828 10508 7840
rect 10560 7828 10566 7880
rect 11900 7868 11928 7908
rect 12158 7896 12164 7948
rect 12216 7936 12222 7948
rect 13357 7939 13415 7945
rect 13357 7936 13369 7939
rect 12216 7908 13369 7936
rect 12216 7896 12222 7908
rect 13357 7905 13369 7908
rect 13403 7905 13415 7939
rect 18230 7936 18236 7948
rect 18191 7908 18236 7936
rect 13357 7899 13415 7905
rect 18230 7896 18236 7908
rect 18288 7896 18294 7948
rect 19518 7936 19524 7948
rect 19479 7908 19524 7936
rect 19518 7896 19524 7908
rect 19576 7896 19582 7948
rect 19889 7939 19947 7945
rect 19889 7905 19901 7939
rect 19935 7936 19947 7939
rect 20901 7939 20959 7945
rect 20901 7936 20913 7939
rect 19935 7908 20913 7936
rect 19935 7905 19947 7908
rect 19889 7899 19947 7905
rect 20901 7905 20913 7908
rect 20947 7936 20959 7939
rect 21450 7936 21456 7948
rect 20947 7908 21456 7936
rect 20947 7905 20959 7908
rect 20901 7899 20959 7905
rect 21450 7896 21456 7908
rect 21508 7896 21514 7948
rect 23385 7939 23443 7945
rect 23385 7905 23397 7939
rect 23431 7936 23443 7939
rect 23474 7936 23480 7948
rect 23431 7908 23480 7936
rect 23431 7905 23443 7908
rect 23385 7899 23443 7905
rect 23474 7896 23480 7908
rect 23532 7896 23538 7948
rect 28534 7945 28540 7948
rect 28528 7936 28540 7945
rect 28495 7908 28540 7936
rect 28528 7899 28540 7908
rect 28534 7896 28540 7899
rect 28592 7896 28598 7948
rect 33220 7939 33278 7945
rect 33220 7905 33232 7939
rect 33266 7936 33278 7939
rect 33502 7936 33508 7948
rect 33266 7908 33508 7936
rect 33266 7905 33278 7908
rect 33220 7899 33278 7905
rect 33502 7896 33508 7908
rect 33560 7896 33566 7948
rect 35250 7896 35256 7948
rect 35308 7936 35314 7948
rect 35805 7939 35863 7945
rect 35805 7936 35817 7939
rect 35308 7908 35817 7936
rect 35308 7896 35314 7908
rect 35805 7905 35817 7908
rect 35851 7905 35863 7939
rect 35805 7899 35863 7905
rect 13633 7871 13691 7877
rect 13633 7868 13645 7871
rect 11900 7840 13645 7868
rect 13633 7837 13645 7840
rect 13679 7868 13691 7871
rect 13722 7868 13728 7880
rect 13679 7840 13728 7868
rect 13679 7837 13691 7840
rect 13633 7831 13691 7837
rect 13722 7828 13728 7840
rect 13780 7828 13786 7880
rect 15194 7828 15200 7880
rect 15252 7868 15258 7880
rect 15289 7871 15347 7877
rect 15289 7868 15301 7871
rect 15252 7840 15301 7868
rect 15252 7828 15258 7840
rect 15289 7837 15301 7840
rect 15335 7837 15347 7871
rect 15289 7831 15347 7837
rect 17034 7828 17040 7880
rect 17092 7868 17098 7880
rect 17773 7871 17831 7877
rect 17773 7868 17785 7871
rect 17092 7840 17785 7868
rect 17092 7828 17098 7840
rect 17773 7837 17785 7840
rect 17819 7868 17831 7871
rect 18325 7871 18383 7877
rect 18325 7868 18337 7871
rect 17819 7840 18337 7868
rect 17819 7837 17831 7840
rect 17773 7831 17831 7837
rect 18325 7837 18337 7840
rect 18371 7837 18383 7871
rect 18506 7868 18512 7880
rect 18419 7840 18512 7868
rect 18325 7831 18383 7837
rect 18506 7828 18512 7840
rect 18564 7868 18570 7880
rect 19242 7868 19248 7880
rect 18564 7840 19248 7868
rect 18564 7828 18570 7840
rect 19242 7828 19248 7840
rect 19300 7828 19306 7880
rect 27154 7868 27160 7880
rect 27115 7840 27160 7868
rect 27154 7828 27160 7840
rect 27212 7828 27218 7880
rect 28074 7828 28080 7880
rect 28132 7868 28138 7880
rect 28261 7871 28319 7877
rect 28261 7868 28273 7871
rect 28132 7840 28273 7868
rect 28132 7828 28138 7840
rect 28261 7837 28273 7840
rect 28307 7837 28319 7871
rect 32674 7868 32680 7880
rect 32635 7840 32680 7868
rect 28261 7831 28319 7837
rect 32674 7828 32680 7840
rect 32732 7828 32738 7880
rect 32953 7871 33011 7877
rect 32953 7837 32965 7871
rect 32999 7837 33011 7871
rect 32953 7831 33011 7837
rect 35989 7871 36047 7877
rect 35989 7837 36001 7871
rect 36035 7837 36047 7871
rect 35989 7831 36047 7837
rect 8481 7803 8539 7809
rect 8481 7800 8493 7803
rect 7432 7772 8493 7800
rect 7432 7760 7438 7772
rect 8481 7769 8493 7772
rect 8527 7769 8539 7803
rect 8481 7763 8539 7769
rect 12894 7760 12900 7812
rect 12952 7800 12958 7812
rect 14001 7803 14059 7809
rect 14001 7800 14013 7803
rect 12952 7772 14013 7800
rect 12952 7760 12958 7772
rect 14001 7769 14013 7772
rect 14047 7800 14059 7803
rect 14369 7803 14427 7809
rect 14369 7800 14381 7803
rect 14047 7772 14381 7800
rect 14047 7769 14059 7772
rect 14001 7763 14059 7769
rect 14369 7769 14381 7772
rect 14415 7769 14427 7803
rect 14369 7763 14427 7769
rect 3050 7732 3056 7744
rect 3011 7704 3056 7732
rect 3050 7692 3056 7704
rect 3108 7692 3114 7744
rect 4341 7735 4399 7741
rect 4341 7701 4353 7735
rect 4387 7732 4399 7735
rect 4706 7732 4712 7744
rect 4387 7704 4712 7732
rect 4387 7701 4399 7704
rect 4341 7695 4399 7701
rect 4706 7692 4712 7704
rect 4764 7732 4770 7744
rect 5166 7732 5172 7744
rect 4764 7704 5172 7732
rect 4764 7692 4770 7704
rect 5166 7692 5172 7704
rect 5224 7692 5230 7744
rect 6546 7692 6552 7744
rect 6604 7732 6610 7744
rect 6917 7735 6975 7741
rect 6917 7732 6929 7735
rect 6604 7704 6929 7732
rect 6604 7692 6610 7704
rect 6917 7701 6929 7704
rect 6963 7701 6975 7735
rect 7282 7732 7288 7744
rect 7243 7704 7288 7732
rect 6917 7695 6975 7701
rect 7282 7692 7288 7704
rect 7340 7692 7346 7744
rect 7466 7732 7472 7744
rect 7427 7704 7472 7732
rect 7466 7692 7472 7704
rect 7524 7692 7530 7744
rect 11885 7735 11943 7741
rect 11885 7701 11897 7735
rect 11931 7732 11943 7735
rect 12342 7732 12348 7744
rect 11931 7704 12348 7732
rect 11931 7701 11943 7704
rect 11885 7695 11943 7701
rect 12342 7692 12348 7704
rect 12400 7692 12406 7744
rect 12986 7732 12992 7744
rect 12947 7704 12992 7732
rect 12986 7692 12992 7704
rect 13044 7692 13050 7744
rect 17770 7692 17776 7744
rect 17828 7732 17834 7744
rect 17865 7735 17923 7741
rect 17865 7732 17877 7735
rect 17828 7704 17877 7732
rect 17828 7692 17834 7704
rect 17865 7701 17877 7704
rect 17911 7701 17923 7735
rect 26602 7732 26608 7744
rect 26563 7704 26608 7732
rect 17865 7695 17923 7701
rect 26602 7692 26608 7704
rect 26660 7692 26666 7744
rect 29638 7732 29644 7744
rect 29599 7704 29644 7732
rect 29638 7692 29644 7704
rect 29696 7692 29702 7744
rect 32122 7692 32128 7744
rect 32180 7732 32186 7744
rect 32968 7732 32996 7831
rect 34790 7760 34796 7812
rect 34848 7800 34854 7812
rect 35802 7800 35808 7812
rect 34848 7772 35808 7800
rect 34848 7760 34854 7772
rect 35802 7760 35808 7772
rect 35860 7800 35866 7812
rect 36004 7800 36032 7831
rect 35860 7772 36032 7800
rect 35860 7760 35866 7772
rect 33962 7732 33968 7744
rect 32180 7704 33968 7732
rect 32180 7692 32186 7704
rect 33962 7692 33968 7704
rect 34020 7692 34026 7744
rect 35434 7732 35440 7744
rect 35395 7704 35440 7732
rect 35434 7692 35440 7704
rect 35492 7692 35498 7744
rect 1104 7642 38824 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 34966 7642
rect 35018 7590 35030 7642
rect 35082 7590 35094 7642
rect 35146 7590 35158 7642
rect 35210 7590 38824 7642
rect 1104 7568 38824 7590
rect 5258 7488 5264 7540
rect 5316 7528 5322 7540
rect 5353 7531 5411 7537
rect 5353 7528 5365 7531
rect 5316 7500 5365 7528
rect 5316 7488 5322 7500
rect 5353 7497 5365 7500
rect 5399 7497 5411 7531
rect 5353 7491 5411 7497
rect 7926 7488 7932 7540
rect 7984 7528 7990 7540
rect 8757 7531 8815 7537
rect 8757 7528 8769 7531
rect 7984 7500 8769 7528
rect 7984 7488 7990 7500
rect 8757 7497 8769 7500
rect 8803 7497 8815 7531
rect 8757 7491 8815 7497
rect 9677 7531 9735 7537
rect 9677 7497 9689 7531
rect 9723 7528 9735 7531
rect 10042 7528 10048 7540
rect 9723 7500 10048 7528
rect 9723 7497 9735 7500
rect 9677 7491 9735 7497
rect 9784 7401 9812 7500
rect 10042 7488 10048 7500
rect 10100 7528 10106 7540
rect 10502 7528 10508 7540
rect 10100 7500 10508 7528
rect 10100 7488 10106 7500
rect 10502 7488 10508 7500
rect 10560 7488 10566 7540
rect 10870 7488 10876 7540
rect 10928 7528 10934 7540
rect 12158 7528 12164 7540
rect 10928 7500 12164 7528
rect 10928 7488 10934 7500
rect 12158 7488 12164 7500
rect 12216 7488 12222 7540
rect 12802 7528 12808 7540
rect 12763 7500 12808 7528
rect 12802 7488 12808 7500
rect 12860 7488 12866 7540
rect 17034 7528 17040 7540
rect 16995 7500 17040 7528
rect 17034 7488 17040 7500
rect 17092 7488 17098 7540
rect 17497 7531 17555 7537
rect 17497 7497 17509 7531
rect 17543 7528 17555 7531
rect 18230 7528 18236 7540
rect 17543 7500 18236 7528
rect 17543 7497 17555 7500
rect 17497 7491 17555 7497
rect 18230 7488 18236 7500
rect 18288 7488 18294 7540
rect 19518 7488 19524 7540
rect 19576 7528 19582 7540
rect 19981 7531 20039 7537
rect 19981 7528 19993 7531
rect 19576 7500 19993 7528
rect 19576 7488 19582 7500
rect 19981 7497 19993 7500
rect 20027 7528 20039 7531
rect 20070 7528 20076 7540
rect 20027 7500 20076 7528
rect 20027 7497 20039 7500
rect 19981 7491 20039 7497
rect 20070 7488 20076 7500
rect 20128 7488 20134 7540
rect 20438 7528 20444 7540
rect 20399 7500 20444 7528
rect 20438 7488 20444 7500
rect 20496 7488 20502 7540
rect 20714 7528 20720 7540
rect 20675 7500 20720 7528
rect 20714 7488 20720 7500
rect 20772 7488 20778 7540
rect 21450 7528 21456 7540
rect 21411 7500 21456 7528
rect 21450 7488 21456 7500
rect 21508 7488 21514 7540
rect 22094 7488 22100 7540
rect 22152 7528 22158 7540
rect 23109 7531 23167 7537
rect 23109 7528 23121 7531
rect 22152 7500 23121 7528
rect 22152 7488 22158 7500
rect 23109 7497 23121 7500
rect 23155 7528 23167 7531
rect 23474 7528 23480 7540
rect 23155 7500 23480 7528
rect 23155 7497 23167 7500
rect 23109 7491 23167 7497
rect 23474 7488 23480 7500
rect 23532 7488 23538 7540
rect 26237 7531 26295 7537
rect 26237 7497 26249 7531
rect 26283 7528 26295 7531
rect 26878 7528 26884 7540
rect 26283 7500 26884 7528
rect 26283 7497 26295 7500
rect 26237 7491 26295 7497
rect 26878 7488 26884 7500
rect 26936 7488 26942 7540
rect 33502 7528 33508 7540
rect 33463 7500 33508 7528
rect 33502 7488 33508 7500
rect 33560 7488 33566 7540
rect 37274 7528 37280 7540
rect 37235 7500 37280 7528
rect 37274 7488 37280 7500
rect 37332 7488 37338 7540
rect 11698 7460 11704 7472
rect 11659 7432 11704 7460
rect 11698 7420 11704 7432
rect 11756 7460 11762 7472
rect 11974 7460 11980 7472
rect 11756 7432 11980 7460
rect 11756 7420 11762 7432
rect 11974 7420 11980 7432
rect 12032 7420 12038 7472
rect 9769 7395 9827 7401
rect 9769 7361 9781 7395
rect 9815 7361 9827 7395
rect 12820 7392 12848 7488
rect 16761 7463 16819 7469
rect 16761 7429 16773 7463
rect 16807 7460 16819 7463
rect 17862 7460 17868 7472
rect 16807 7432 17868 7460
rect 16807 7429 16819 7432
rect 16761 7423 16819 7429
rect 13220 7395 13278 7401
rect 13220 7392 13232 7395
rect 12820 7364 13232 7392
rect 9769 7355 9827 7361
rect 13220 7361 13232 7364
rect 13266 7361 13278 7395
rect 13354 7392 13360 7404
rect 13315 7364 13360 7392
rect 13220 7355 13278 7361
rect 13354 7352 13360 7364
rect 13412 7352 13418 7404
rect 2961 7327 3019 7333
rect 2961 7324 2973 7327
rect 2792 7296 2973 7324
rect 2792 7200 2820 7296
rect 2961 7293 2973 7296
rect 3007 7293 3019 7327
rect 2961 7287 3019 7293
rect 3050 7284 3056 7336
rect 3108 7324 3114 7336
rect 3217 7327 3275 7333
rect 3217 7324 3229 7327
rect 3108 7296 3229 7324
rect 3108 7284 3114 7296
rect 3217 7293 3229 7296
rect 3263 7293 3275 7327
rect 3217 7287 3275 7293
rect 5534 7284 5540 7336
rect 5592 7324 5598 7336
rect 5629 7327 5687 7333
rect 5629 7324 5641 7327
rect 5592 7296 5641 7324
rect 5592 7284 5598 7296
rect 5629 7293 5641 7296
rect 5675 7293 5687 7327
rect 5629 7287 5687 7293
rect 6546 7284 6552 7336
rect 6604 7324 6610 7336
rect 6825 7327 6883 7333
rect 6825 7324 6837 7327
rect 6604 7296 6837 7324
rect 6604 7284 6610 7296
rect 6825 7293 6837 7296
rect 6871 7293 6883 7327
rect 10036 7327 10094 7333
rect 10036 7324 10048 7327
rect 6825 7287 6883 7293
rect 9968 7296 10048 7324
rect 3970 7216 3976 7268
rect 4028 7256 4034 7268
rect 4982 7256 4988 7268
rect 4028 7228 4988 7256
rect 4028 7216 4034 7228
rect 4982 7216 4988 7228
rect 5040 7216 5046 7268
rect 6273 7259 6331 7265
rect 6273 7225 6285 7259
rect 6319 7256 6331 7259
rect 7092 7259 7150 7265
rect 7092 7256 7104 7259
rect 6319 7228 7104 7256
rect 6319 7225 6331 7228
rect 6273 7219 6331 7225
rect 7092 7225 7104 7228
rect 7138 7256 7150 7259
rect 7926 7256 7932 7268
rect 7138 7228 7932 7256
rect 7138 7225 7150 7228
rect 7092 7219 7150 7225
rect 7926 7216 7932 7228
rect 7984 7216 7990 7268
rect 9309 7259 9367 7265
rect 9309 7225 9321 7259
rect 9355 7256 9367 7259
rect 9968 7256 9996 7296
rect 10036 7293 10048 7296
rect 10082 7324 10094 7327
rect 12342 7324 12348 7336
rect 10082 7296 12348 7324
rect 10082 7293 10094 7296
rect 10036 7287 10094 7293
rect 12342 7284 12348 7296
rect 12400 7284 12406 7336
rect 12894 7324 12900 7336
rect 12855 7296 12900 7324
rect 12894 7284 12900 7296
rect 12952 7284 12958 7336
rect 16868 7333 16896 7432
rect 17862 7420 17868 7432
rect 17920 7420 17926 7472
rect 17773 7395 17831 7401
rect 17773 7361 17785 7395
rect 17819 7392 17831 7395
rect 18046 7392 18052 7404
rect 17819 7364 18052 7392
rect 17819 7361 17831 7364
rect 17773 7355 17831 7361
rect 13633 7327 13691 7333
rect 13633 7324 13645 7327
rect 13004 7296 13645 7324
rect 9355 7228 9996 7256
rect 9355 7225 9367 7228
rect 9309 7219 9367 7225
rect 12618 7216 12624 7268
rect 12676 7256 12682 7268
rect 13004 7256 13032 7296
rect 13633 7293 13645 7296
rect 13679 7293 13691 7327
rect 13633 7287 13691 7293
rect 16853 7327 16911 7333
rect 16853 7293 16865 7327
rect 16899 7293 16911 7327
rect 16853 7287 16911 7293
rect 12676 7228 13032 7256
rect 12676 7216 12682 7228
rect 15194 7216 15200 7268
rect 15252 7256 15258 7268
rect 15289 7259 15347 7265
rect 15289 7256 15301 7259
rect 15252 7228 15301 7256
rect 15252 7216 15258 7228
rect 15289 7225 15301 7228
rect 15335 7256 15347 7259
rect 17788 7256 17816 7355
rect 18046 7352 18052 7364
rect 18104 7352 18110 7404
rect 23492 7392 23520 7488
rect 23661 7395 23719 7401
rect 23661 7392 23673 7395
rect 23492 7364 23673 7392
rect 23661 7361 23673 7364
rect 23707 7361 23719 7395
rect 23661 7355 23719 7361
rect 25869 7395 25927 7401
rect 25869 7361 25881 7395
rect 25915 7392 25927 7395
rect 32033 7395 32091 7401
rect 25915 7364 26832 7392
rect 25915 7361 25927 7364
rect 25869 7355 25927 7361
rect 19426 7284 19432 7336
rect 19484 7324 19490 7336
rect 20533 7327 20591 7333
rect 20533 7324 20545 7327
rect 19484 7296 20545 7324
rect 19484 7284 19490 7296
rect 20533 7293 20545 7296
rect 20579 7324 20591 7327
rect 21085 7327 21143 7333
rect 21085 7324 21097 7327
rect 20579 7296 21097 7324
rect 20579 7293 20591 7296
rect 20533 7287 20591 7293
rect 21085 7293 21097 7296
rect 21131 7293 21143 7327
rect 21085 7287 21143 7293
rect 22465 7327 22523 7333
rect 22465 7293 22477 7327
rect 22511 7293 22523 7327
rect 22465 7287 22523 7293
rect 26697 7327 26755 7333
rect 26697 7293 26709 7327
rect 26743 7293 26755 7327
rect 26804 7324 26832 7364
rect 32033 7361 32045 7395
rect 32079 7392 32091 7395
rect 32122 7392 32128 7404
rect 32079 7364 32128 7392
rect 32079 7361 32091 7364
rect 32033 7355 32091 7361
rect 32122 7352 32128 7364
rect 32180 7352 32186 7404
rect 34238 7352 34244 7404
rect 34296 7392 34302 7404
rect 35158 7392 35164 7404
rect 34296 7364 35164 7392
rect 34296 7352 34302 7364
rect 35158 7352 35164 7364
rect 35216 7392 35222 7404
rect 35437 7395 35495 7401
rect 35437 7392 35449 7395
rect 35216 7364 35449 7392
rect 35216 7352 35222 7364
rect 35437 7361 35449 7364
rect 35483 7361 35495 7395
rect 35437 7355 35495 7361
rect 35802 7352 35808 7404
rect 35860 7392 35866 7404
rect 35897 7395 35955 7401
rect 35897 7392 35909 7395
rect 35860 7364 35909 7392
rect 35860 7352 35866 7364
rect 35897 7361 35909 7364
rect 35943 7361 35955 7395
rect 35897 7355 35955 7361
rect 26970 7333 26976 7336
rect 26964 7324 26976 7333
rect 26804 7296 26976 7324
rect 26697 7287 26755 7293
rect 26964 7287 26976 7296
rect 15335 7228 17816 7256
rect 15335 7225 15347 7228
rect 15289 7219 15347 7225
rect 17862 7216 17868 7268
rect 17920 7256 17926 7268
rect 18316 7259 18374 7265
rect 18316 7256 18328 7259
rect 17920 7228 18328 7256
rect 17920 7216 17926 7228
rect 18316 7225 18328 7228
rect 18362 7256 18374 7259
rect 18506 7256 18512 7268
rect 18362 7228 18512 7256
rect 18362 7225 18374 7228
rect 18316 7219 18374 7225
rect 18506 7216 18512 7228
rect 18564 7216 18570 7268
rect 22480 7200 22508 7287
rect 23934 7265 23940 7268
rect 23928 7256 23940 7265
rect 23895 7228 23940 7256
rect 23928 7219 23940 7228
rect 23934 7216 23940 7219
rect 23992 7216 23998 7268
rect 26510 7216 26516 7268
rect 26568 7256 26574 7268
rect 26605 7259 26663 7265
rect 26605 7256 26617 7259
rect 26568 7228 26617 7256
rect 26568 7216 26574 7228
rect 26605 7225 26617 7228
rect 26651 7256 26663 7259
rect 26712 7256 26740 7287
rect 26970 7284 26976 7287
rect 27028 7284 27034 7336
rect 28074 7324 28080 7336
rect 27080 7296 28080 7324
rect 27080 7256 27108 7296
rect 28074 7284 28080 7296
rect 28132 7324 28138 7336
rect 28629 7327 28687 7333
rect 28629 7324 28641 7327
rect 28132 7296 28641 7324
rect 28132 7284 28138 7296
rect 28629 7293 28641 7296
rect 28675 7293 28687 7327
rect 28629 7287 28687 7293
rect 34701 7327 34759 7333
rect 34701 7293 34713 7327
rect 34747 7324 34759 7327
rect 35250 7324 35256 7336
rect 34747 7296 35256 7324
rect 34747 7293 34759 7296
rect 34701 7287 34759 7293
rect 35250 7284 35256 7296
rect 35308 7284 35314 7336
rect 36170 7324 36176 7336
rect 36131 7296 36176 7324
rect 36170 7284 36176 7296
rect 36228 7284 36234 7336
rect 28534 7256 28540 7268
rect 26651 7228 27108 7256
rect 28092 7228 28540 7256
rect 26651 7225 26663 7228
rect 26605 7219 26663 7225
rect 2498 7188 2504 7200
rect 2459 7160 2504 7188
rect 2498 7148 2504 7160
rect 2556 7148 2562 7200
rect 2774 7188 2780 7200
rect 2735 7160 2780 7188
rect 2774 7148 2780 7160
rect 2832 7148 2838 7200
rect 4154 7148 4160 7200
rect 4212 7188 4218 7200
rect 4341 7191 4399 7197
rect 4341 7188 4353 7191
rect 4212 7160 4353 7188
rect 4212 7148 4218 7160
rect 4341 7157 4353 7160
rect 4387 7157 4399 7191
rect 5810 7188 5816 7200
rect 5771 7160 5816 7188
rect 4341 7151 4399 7157
rect 5810 7148 5816 7160
rect 5868 7148 5874 7200
rect 6546 7188 6552 7200
rect 6507 7160 6552 7188
rect 6546 7148 6552 7160
rect 6604 7148 6610 7200
rect 8202 7188 8208 7200
rect 8163 7160 8208 7188
rect 8202 7148 8208 7160
rect 8260 7148 8266 7200
rect 11146 7188 11152 7200
rect 11107 7160 11152 7188
rect 11146 7148 11152 7160
rect 11204 7148 11210 7200
rect 14734 7188 14740 7200
rect 14695 7160 14740 7188
rect 14734 7148 14740 7160
rect 14792 7148 14798 7200
rect 15470 7148 15476 7200
rect 15528 7188 15534 7200
rect 15657 7191 15715 7197
rect 15657 7188 15669 7191
rect 15528 7160 15669 7188
rect 15528 7148 15534 7160
rect 15657 7157 15669 7160
rect 15703 7157 15715 7191
rect 19426 7188 19432 7200
rect 19387 7160 19432 7188
rect 15657 7151 15715 7157
rect 19426 7148 19432 7160
rect 19484 7148 19490 7200
rect 22373 7191 22431 7197
rect 22373 7157 22385 7191
rect 22419 7188 22431 7191
rect 22462 7188 22468 7200
rect 22419 7160 22468 7188
rect 22419 7157 22431 7160
rect 22373 7151 22431 7157
rect 22462 7148 22468 7160
rect 22520 7148 22526 7200
rect 22646 7188 22652 7200
rect 22607 7160 22652 7188
rect 22646 7148 22652 7160
rect 22704 7148 22710 7200
rect 23566 7148 23572 7200
rect 23624 7188 23630 7200
rect 25041 7191 25099 7197
rect 25041 7188 25053 7191
rect 23624 7160 25053 7188
rect 23624 7148 23630 7160
rect 25041 7157 25053 7160
rect 25087 7157 25099 7191
rect 25041 7151 25099 7157
rect 27982 7148 27988 7200
rect 28040 7188 28046 7200
rect 28092 7197 28120 7228
rect 28534 7216 28540 7228
rect 28592 7256 28598 7268
rect 28997 7259 29055 7265
rect 28997 7256 29009 7259
rect 28592 7228 29009 7256
rect 28592 7216 28598 7228
rect 28997 7225 29009 7228
rect 29043 7225 29055 7259
rect 28997 7219 29055 7225
rect 31665 7259 31723 7265
rect 31665 7225 31677 7259
rect 31711 7256 31723 7259
rect 32392 7259 32450 7265
rect 32392 7256 32404 7259
rect 31711 7228 32404 7256
rect 31711 7225 31723 7228
rect 31665 7219 31723 7225
rect 32392 7225 32404 7228
rect 32438 7256 32450 7259
rect 32490 7256 32496 7268
rect 32438 7228 32496 7256
rect 32438 7225 32450 7228
rect 32392 7219 32450 7225
rect 32490 7216 32496 7228
rect 32548 7216 32554 7268
rect 28077 7191 28135 7197
rect 28077 7188 28089 7191
rect 28040 7160 28089 7188
rect 28040 7148 28046 7160
rect 28077 7157 28089 7160
rect 28123 7157 28135 7191
rect 28077 7151 28135 7157
rect 28902 7148 28908 7200
rect 28960 7188 28966 7200
rect 29273 7191 29331 7197
rect 29273 7188 29285 7191
rect 28960 7160 29285 7188
rect 28960 7148 28966 7160
rect 29273 7157 29285 7160
rect 29319 7157 29331 7191
rect 29273 7151 29331 7157
rect 33962 7148 33968 7200
rect 34020 7188 34026 7200
rect 34057 7191 34115 7197
rect 34057 7188 34069 7191
rect 34020 7160 34069 7188
rect 34020 7148 34026 7160
rect 34057 7157 34069 7160
rect 34103 7157 34115 7191
rect 34057 7151 34115 7157
rect 34514 7148 34520 7200
rect 34572 7188 34578 7200
rect 35066 7188 35072 7200
rect 34572 7160 35072 7188
rect 34572 7148 34578 7160
rect 35066 7148 35072 7160
rect 35124 7188 35130 7200
rect 35253 7191 35311 7197
rect 35253 7188 35265 7191
rect 35124 7160 35265 7188
rect 35124 7148 35130 7160
rect 35253 7157 35265 7160
rect 35299 7188 35311 7191
rect 35899 7191 35957 7197
rect 35899 7188 35911 7191
rect 35299 7160 35911 7188
rect 35299 7157 35311 7160
rect 35253 7151 35311 7157
rect 35899 7157 35911 7160
rect 35945 7157 35957 7191
rect 35899 7151 35957 7157
rect 1104 7098 38824 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 38824 7098
rect 1104 7024 38824 7046
rect 2498 6944 2504 6996
rect 2556 6984 2562 6996
rect 2777 6987 2835 6993
rect 2777 6984 2789 6987
rect 2556 6956 2789 6984
rect 2556 6944 2562 6956
rect 2777 6953 2789 6956
rect 2823 6953 2835 6987
rect 5442 6984 5448 6996
rect 5403 6956 5448 6984
rect 2777 6947 2835 6953
rect 5442 6944 5448 6956
rect 5500 6944 5506 6996
rect 11422 6984 11428 6996
rect 11383 6956 11428 6984
rect 11422 6944 11428 6956
rect 11480 6944 11486 6996
rect 12437 6987 12495 6993
rect 12437 6953 12449 6987
rect 12483 6984 12495 6987
rect 12618 6984 12624 6996
rect 12483 6956 12624 6984
rect 12483 6953 12495 6956
rect 12437 6947 12495 6953
rect 12618 6944 12624 6956
rect 12676 6944 12682 6996
rect 12989 6987 13047 6993
rect 12989 6953 13001 6987
rect 13035 6984 13047 6987
rect 13170 6984 13176 6996
rect 13035 6956 13176 6984
rect 13035 6953 13047 6956
rect 12989 6947 13047 6953
rect 13170 6944 13176 6956
rect 13228 6984 13234 6996
rect 14734 6984 14740 6996
rect 13228 6956 14740 6984
rect 13228 6944 13234 6956
rect 14734 6944 14740 6956
rect 14792 6944 14798 6996
rect 15194 6944 15200 6996
rect 15252 6944 15258 6996
rect 25225 6987 25283 6993
rect 25225 6953 25237 6987
rect 25271 6984 25283 6987
rect 25498 6984 25504 6996
rect 25271 6956 25504 6984
rect 25271 6953 25283 6956
rect 25225 6947 25283 6953
rect 25498 6944 25504 6956
rect 25556 6984 25562 6996
rect 26602 6984 26608 6996
rect 25556 6956 26608 6984
rect 25556 6944 25562 6956
rect 26602 6944 26608 6956
rect 26660 6944 26666 6996
rect 26970 6944 26976 6996
rect 27028 6984 27034 6996
rect 27065 6987 27123 6993
rect 27065 6984 27077 6987
rect 27028 6956 27077 6984
rect 27028 6944 27034 6956
rect 27065 6953 27077 6956
rect 27111 6953 27123 6987
rect 27065 6947 27123 6953
rect 33042 6944 33048 6996
rect 33100 6984 33106 6996
rect 33229 6987 33287 6993
rect 33229 6984 33241 6987
rect 33100 6956 33241 6984
rect 33100 6944 33106 6956
rect 33229 6953 33241 6956
rect 33275 6984 33287 6987
rect 33594 6984 33600 6996
rect 33275 6956 33600 6984
rect 33275 6953 33287 6956
rect 33229 6947 33287 6953
rect 33594 6944 33600 6956
rect 33652 6944 33658 6996
rect 34790 6984 34796 6996
rect 34751 6956 34796 6984
rect 34790 6944 34796 6956
rect 34848 6944 34854 6996
rect 35434 6944 35440 6996
rect 35492 6984 35498 6996
rect 35713 6987 35771 6993
rect 35713 6984 35725 6987
rect 35492 6956 35725 6984
rect 35492 6944 35498 6956
rect 35713 6953 35725 6956
rect 35759 6953 35771 6987
rect 35713 6947 35771 6953
rect 4154 6916 4160 6928
rect 4080 6888 4160 6916
rect 2317 6851 2375 6857
rect 2317 6817 2329 6851
rect 2363 6848 2375 6851
rect 2590 6848 2596 6860
rect 2363 6820 2596 6848
rect 2363 6817 2375 6820
rect 2317 6811 2375 6817
rect 2590 6808 2596 6820
rect 2648 6848 2654 6860
rect 2869 6851 2927 6857
rect 2869 6848 2881 6851
rect 2648 6820 2881 6848
rect 2648 6808 2654 6820
rect 2869 6817 2881 6820
rect 2915 6848 2927 6851
rect 4080 6848 4108 6888
rect 4154 6876 4160 6888
rect 4212 6876 4218 6928
rect 11146 6916 11152 6928
rect 10980 6888 11152 6916
rect 2915 6820 4108 6848
rect 4332 6851 4390 6857
rect 2915 6817 2927 6820
rect 2869 6811 2927 6817
rect 4332 6817 4344 6851
rect 4378 6848 4390 6851
rect 4706 6848 4712 6860
rect 4378 6820 4712 6848
rect 4378 6817 4390 6820
rect 4332 6811 4390 6817
rect 4706 6808 4712 6820
rect 4764 6848 4770 6860
rect 5350 6848 5356 6860
rect 4764 6820 5356 6848
rect 4764 6808 4770 6820
rect 5350 6808 5356 6820
rect 5408 6808 5414 6860
rect 6638 6808 6644 6860
rect 6696 6848 6702 6860
rect 6805 6851 6863 6857
rect 6805 6848 6817 6851
rect 6696 6820 6817 6848
rect 6696 6808 6702 6820
rect 6805 6817 6817 6820
rect 6851 6848 6863 6851
rect 8294 6848 8300 6860
rect 6851 6820 8300 6848
rect 6851 6817 6863 6820
rect 6805 6811 6863 6817
rect 8294 6808 8300 6820
rect 8352 6808 8358 6860
rect 10042 6848 10048 6860
rect 10003 6820 10048 6848
rect 10042 6808 10048 6820
rect 10100 6808 10106 6860
rect 10312 6851 10370 6857
rect 10312 6817 10324 6851
rect 10358 6848 10370 6851
rect 10686 6848 10692 6860
rect 10358 6820 10692 6848
rect 10358 6817 10370 6820
rect 10312 6811 10370 6817
rect 10686 6808 10692 6820
rect 10744 6848 10750 6860
rect 10980 6848 11008 6888
rect 11146 6876 11152 6888
rect 11204 6876 11210 6928
rect 11974 6876 11980 6928
rect 12032 6916 12038 6928
rect 15212 6916 15240 6944
rect 18049 6919 18107 6925
rect 18049 6916 18061 6919
rect 12032 6888 15240 6916
rect 17880 6888 18061 6916
rect 12032 6876 12038 6888
rect 10744 6820 11008 6848
rect 10744 6808 10750 6820
rect 11790 6808 11796 6860
rect 11848 6848 11854 6860
rect 12897 6851 12955 6857
rect 12897 6848 12909 6851
rect 11848 6820 12909 6848
rect 11848 6808 11854 6820
rect 12897 6817 12909 6820
rect 12943 6848 12955 6851
rect 13354 6848 13360 6860
rect 12943 6820 13360 6848
rect 12943 6817 12955 6820
rect 12897 6811 12955 6817
rect 13354 6808 13360 6820
rect 13412 6848 13418 6860
rect 13541 6851 13599 6857
rect 13541 6848 13553 6851
rect 13412 6820 13553 6848
rect 13412 6808 13418 6820
rect 13541 6817 13553 6820
rect 13587 6817 13599 6851
rect 13541 6811 13599 6817
rect 13814 6808 13820 6860
rect 13872 6848 13878 6860
rect 13909 6851 13967 6857
rect 13909 6848 13921 6851
rect 13872 6820 13921 6848
rect 13872 6808 13878 6820
rect 13909 6817 13921 6820
rect 13955 6817 13967 6851
rect 13909 6811 13967 6817
rect 16669 6851 16727 6857
rect 16669 6817 16681 6851
rect 16715 6848 16727 6851
rect 17494 6848 17500 6860
rect 16715 6820 17500 6848
rect 16715 6817 16727 6820
rect 16669 6811 16727 6817
rect 17494 6808 17500 6820
rect 17552 6848 17558 6860
rect 17880 6848 17908 6888
rect 18049 6885 18061 6888
rect 18095 6885 18107 6919
rect 18049 6879 18107 6885
rect 35158 6876 35164 6928
rect 35216 6916 35222 6928
rect 35216 6888 35848 6916
rect 35216 6876 35222 6888
rect 17552 6820 17908 6848
rect 17552 6808 17558 6820
rect 17954 6808 17960 6860
rect 18012 6848 18018 6860
rect 19245 6851 19303 6857
rect 19245 6848 19257 6851
rect 18012 6820 19257 6848
rect 18012 6808 18018 6820
rect 19245 6817 19257 6820
rect 19291 6848 19303 6851
rect 19978 6848 19984 6860
rect 19291 6820 19984 6848
rect 19291 6817 19303 6820
rect 19245 6811 19303 6817
rect 19978 6808 19984 6820
rect 20036 6808 20042 6860
rect 22370 6857 22376 6860
rect 22364 6811 22376 6857
rect 22428 6848 22434 6860
rect 22428 6820 22464 6848
rect 22370 6808 22376 6811
rect 22428 6808 22434 6820
rect 25314 6808 25320 6860
rect 25372 6848 25378 6860
rect 26513 6851 26571 6857
rect 25372 6820 25417 6848
rect 25372 6808 25378 6820
rect 26513 6817 26525 6851
rect 26559 6848 26571 6851
rect 26970 6848 26976 6860
rect 26559 6820 26976 6848
rect 26559 6817 26571 6820
rect 26513 6811 26571 6817
rect 26970 6808 26976 6820
rect 27028 6808 27034 6860
rect 28528 6851 28586 6857
rect 28528 6817 28540 6851
rect 28574 6848 28586 6851
rect 28994 6848 29000 6860
rect 28574 6820 29000 6848
rect 28574 6817 28586 6820
rect 28528 6811 28586 6817
rect 28994 6808 29000 6820
rect 29052 6848 29058 6860
rect 29638 6848 29644 6860
rect 29052 6820 29644 6848
rect 29052 6808 29058 6820
rect 29638 6808 29644 6820
rect 29696 6808 29702 6860
rect 32950 6808 32956 6860
rect 33008 6848 33014 6860
rect 33321 6851 33379 6857
rect 33321 6848 33333 6851
rect 33008 6820 33333 6848
rect 33008 6808 33014 6820
rect 33321 6817 33333 6820
rect 33367 6848 33379 6851
rect 33594 6848 33600 6860
rect 33367 6820 33600 6848
rect 33367 6817 33379 6820
rect 33321 6811 33379 6817
rect 33594 6808 33600 6820
rect 33652 6808 33658 6860
rect 35618 6848 35624 6860
rect 35579 6820 35624 6848
rect 35618 6808 35624 6820
rect 35676 6808 35682 6860
rect 35820 6848 35848 6888
rect 36633 6851 36691 6857
rect 36633 6848 36645 6851
rect 35820 6820 36645 6848
rect 36633 6817 36645 6820
rect 36679 6817 36691 6851
rect 36633 6811 36691 6817
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6780 2007 6783
rect 3053 6783 3111 6789
rect 3053 6780 3065 6783
rect 1995 6752 3065 6780
rect 1995 6749 2007 6752
rect 1949 6743 2007 6749
rect 3053 6749 3065 6752
rect 3099 6780 3111 6783
rect 3099 6752 3556 6780
rect 3099 6749 3111 6752
rect 3053 6743 3111 6749
rect 3528 6656 3556 6752
rect 3970 6740 3976 6792
rect 4028 6780 4034 6792
rect 4065 6783 4123 6789
rect 4065 6780 4077 6783
rect 4028 6752 4077 6780
rect 4028 6740 4034 6752
rect 4065 6749 4077 6752
rect 4111 6749 4123 6783
rect 6546 6780 6552 6792
rect 6507 6752 6552 6780
rect 4065 6743 4123 6749
rect 6546 6740 6552 6752
rect 6604 6740 6610 6792
rect 12434 6740 12440 6792
rect 12492 6780 12498 6792
rect 12802 6780 12808 6792
rect 12492 6752 12808 6780
rect 12492 6740 12498 6752
rect 12802 6740 12808 6752
rect 12860 6780 12866 6792
rect 13081 6783 13139 6789
rect 13081 6780 13093 6783
rect 12860 6752 13093 6780
rect 12860 6740 12866 6752
rect 13081 6749 13093 6752
rect 13127 6749 13139 6783
rect 13081 6743 13139 6749
rect 13722 6740 13728 6792
rect 13780 6780 13786 6792
rect 14093 6783 14151 6789
rect 14093 6780 14105 6783
rect 13780 6752 14105 6780
rect 13780 6740 13786 6752
rect 14093 6749 14105 6752
rect 14139 6749 14151 6783
rect 15286 6780 15292 6792
rect 15247 6752 15292 6780
rect 14093 6743 14151 6749
rect 15286 6740 15292 6752
rect 15344 6740 15350 6792
rect 17221 6783 17279 6789
rect 17221 6749 17233 6783
rect 17267 6780 17279 6783
rect 17589 6783 17647 6789
rect 17589 6780 17601 6783
rect 17267 6752 17601 6780
rect 17267 6749 17279 6752
rect 17221 6743 17279 6749
rect 17589 6749 17601 6752
rect 17635 6780 17647 6783
rect 17862 6780 17868 6792
rect 17635 6752 17868 6780
rect 17635 6749 17647 6752
rect 17589 6743 17647 6749
rect 17862 6740 17868 6752
rect 17920 6740 17926 6792
rect 18141 6783 18199 6789
rect 18141 6749 18153 6783
rect 18187 6749 18199 6783
rect 18141 6743 18199 6749
rect 18325 6783 18383 6789
rect 18325 6749 18337 6783
rect 18371 6780 18383 6783
rect 18414 6780 18420 6792
rect 18371 6752 18420 6780
rect 18371 6749 18383 6752
rect 18325 6743 18383 6749
rect 5074 6672 5080 6724
rect 5132 6712 5138 6724
rect 6362 6712 6368 6724
rect 5132 6684 6368 6712
rect 5132 6672 5138 6684
rect 6362 6672 6368 6684
rect 6420 6672 6426 6724
rect 17770 6672 17776 6724
rect 17828 6712 17834 6724
rect 17954 6712 17960 6724
rect 17828 6684 17960 6712
rect 17828 6672 17834 6684
rect 17954 6672 17960 6684
rect 18012 6712 18018 6724
rect 18156 6712 18184 6743
rect 18414 6740 18420 6752
rect 18472 6780 18478 6792
rect 18693 6783 18751 6789
rect 18693 6780 18705 6783
rect 18472 6752 18705 6780
rect 18472 6740 18478 6752
rect 18693 6749 18705 6752
rect 18739 6780 18751 6783
rect 19426 6780 19432 6792
rect 18739 6752 19432 6780
rect 18739 6749 18751 6752
rect 18693 6743 18751 6749
rect 19426 6740 19432 6752
rect 19484 6740 19490 6792
rect 21910 6740 21916 6792
rect 21968 6780 21974 6792
rect 22094 6780 22100 6792
rect 21968 6752 22100 6780
rect 21968 6740 21974 6752
rect 22094 6740 22100 6752
rect 22152 6780 22158 6792
rect 25406 6780 25412 6792
rect 22152 6752 22197 6780
rect 25367 6752 25412 6780
rect 22152 6740 22158 6752
rect 25406 6740 25412 6752
rect 25464 6780 25470 6792
rect 25869 6783 25927 6789
rect 25869 6780 25881 6783
rect 25464 6752 25881 6780
rect 25464 6740 25470 6752
rect 25869 6749 25881 6752
rect 25915 6749 25927 6783
rect 25869 6743 25927 6749
rect 28074 6740 28080 6792
rect 28132 6780 28138 6792
rect 28261 6783 28319 6789
rect 28261 6780 28273 6783
rect 28132 6752 28273 6780
rect 28132 6740 28138 6752
rect 28261 6749 28273 6752
rect 28307 6749 28319 6783
rect 33502 6780 33508 6792
rect 33463 6752 33508 6780
rect 28261 6743 28319 6749
rect 33502 6740 33508 6752
rect 33560 6740 33566 6792
rect 35526 6740 35532 6792
rect 35584 6780 35590 6792
rect 35805 6783 35863 6789
rect 35805 6780 35817 6783
rect 35584 6752 35817 6780
rect 35584 6740 35590 6752
rect 35805 6749 35817 6752
rect 35851 6749 35863 6783
rect 35805 6743 35863 6749
rect 24762 6712 24768 6724
rect 18012 6684 18184 6712
rect 24412 6684 24768 6712
rect 18012 6672 18018 6684
rect 2406 6644 2412 6656
rect 2367 6616 2412 6644
rect 2406 6604 2412 6616
rect 2464 6604 2470 6656
rect 3510 6644 3516 6656
rect 3471 6616 3516 6644
rect 3510 6604 3516 6616
rect 3568 6604 3574 6656
rect 5534 6604 5540 6656
rect 5592 6644 5598 6656
rect 5997 6647 6055 6653
rect 5997 6644 6009 6647
rect 5592 6616 6009 6644
rect 5592 6604 5598 6616
rect 5997 6613 6009 6616
rect 6043 6613 6055 6647
rect 5997 6607 6055 6613
rect 7282 6604 7288 6656
rect 7340 6644 7346 6656
rect 7929 6647 7987 6653
rect 7929 6644 7941 6647
rect 7340 6616 7941 6644
rect 7340 6604 7346 6616
rect 7929 6613 7941 6616
rect 7975 6613 7987 6647
rect 7929 6607 7987 6613
rect 8386 6604 8392 6656
rect 8444 6644 8450 6656
rect 8481 6647 8539 6653
rect 8481 6644 8493 6647
rect 8444 6616 8493 6644
rect 8444 6604 8450 6616
rect 8481 6613 8493 6616
rect 8527 6613 8539 6647
rect 12066 6644 12072 6656
rect 12027 6616 12072 6644
rect 8481 6607 8539 6613
rect 12066 6604 12072 6616
rect 12124 6604 12130 6656
rect 12526 6644 12532 6656
rect 12487 6616 12532 6644
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 16942 6604 16948 6656
rect 17000 6644 17006 6656
rect 17681 6647 17739 6653
rect 17681 6644 17693 6647
rect 17000 6616 17693 6644
rect 17000 6604 17006 6616
rect 17681 6613 17693 6616
rect 17727 6613 17739 6647
rect 19426 6644 19432 6656
rect 19387 6616 19432 6644
rect 17681 6607 17739 6613
rect 19426 6604 19432 6616
rect 19484 6604 19490 6656
rect 22002 6644 22008 6656
rect 21963 6616 22008 6644
rect 22002 6604 22008 6616
rect 22060 6604 22066 6656
rect 23474 6644 23480 6656
rect 23435 6616 23480 6644
rect 23474 6604 23480 6616
rect 23532 6644 23538 6656
rect 23934 6644 23940 6656
rect 23532 6616 23940 6644
rect 23532 6604 23538 6616
rect 23934 6604 23940 6616
rect 23992 6644 23998 6656
rect 24029 6647 24087 6653
rect 24029 6644 24041 6647
rect 23992 6616 24041 6644
rect 23992 6604 23998 6616
rect 24029 6613 24041 6616
rect 24075 6613 24087 6647
rect 24029 6607 24087 6613
rect 24118 6604 24124 6656
rect 24176 6644 24182 6656
rect 24412 6653 24440 6684
rect 24762 6672 24768 6684
rect 24820 6712 24826 6724
rect 26237 6715 26295 6721
rect 26237 6712 26249 6715
rect 24820 6684 26249 6712
rect 24820 6672 24826 6684
rect 26237 6681 26249 6684
rect 26283 6712 26295 6715
rect 27154 6712 27160 6724
rect 26283 6684 27160 6712
rect 26283 6681 26295 6684
rect 26237 6675 26295 6681
rect 27154 6672 27160 6684
rect 27212 6712 27218 6724
rect 27525 6715 27583 6721
rect 27525 6712 27537 6715
rect 27212 6684 27537 6712
rect 27212 6672 27218 6684
rect 27525 6681 27537 6684
rect 27571 6712 27583 6715
rect 27890 6712 27896 6724
rect 27571 6684 27896 6712
rect 27571 6681 27583 6684
rect 27525 6675 27583 6681
rect 27890 6672 27896 6684
rect 27948 6672 27954 6724
rect 32769 6715 32827 6721
rect 32769 6681 32781 6715
rect 32815 6712 32827 6715
rect 33520 6712 33548 6740
rect 32815 6684 33548 6712
rect 32815 6681 32827 6684
rect 32769 6675 32827 6681
rect 24397 6647 24455 6653
rect 24397 6644 24409 6647
rect 24176 6616 24409 6644
rect 24176 6604 24182 6616
rect 24397 6613 24409 6616
rect 24443 6613 24455 6647
rect 24854 6644 24860 6656
rect 24815 6616 24860 6644
rect 24397 6607 24455 6613
rect 24854 6604 24860 6616
rect 24912 6604 24918 6656
rect 26602 6604 26608 6656
rect 26660 6644 26666 6656
rect 26697 6647 26755 6653
rect 26697 6644 26709 6647
rect 26660 6616 26709 6644
rect 26660 6604 26666 6616
rect 26697 6613 26709 6616
rect 26743 6613 26755 6647
rect 29638 6644 29644 6656
rect 29599 6616 29644 6644
rect 26697 6607 26755 6613
rect 29638 6604 29644 6616
rect 29696 6604 29702 6656
rect 32858 6644 32864 6656
rect 32819 6616 32864 6644
rect 32858 6604 32864 6616
rect 32916 6604 32922 6656
rect 35161 6647 35219 6653
rect 35161 6613 35173 6647
rect 35207 6644 35219 6647
rect 35253 6647 35311 6653
rect 35253 6644 35265 6647
rect 35207 6616 35265 6644
rect 35207 6613 35219 6616
rect 35161 6607 35219 6613
rect 35253 6613 35265 6616
rect 35299 6644 35311 6647
rect 35802 6644 35808 6656
rect 35299 6616 35808 6644
rect 35299 6613 35311 6616
rect 35253 6607 35311 6613
rect 35802 6604 35808 6616
rect 35860 6604 35866 6656
rect 35894 6604 35900 6656
rect 35952 6644 35958 6656
rect 36170 6644 36176 6656
rect 35952 6616 36176 6644
rect 35952 6604 35958 6616
rect 36170 6604 36176 6616
rect 36228 6644 36234 6656
rect 36265 6647 36323 6653
rect 36265 6644 36277 6647
rect 36228 6616 36277 6644
rect 36228 6604 36234 6616
rect 36265 6613 36277 6616
rect 36311 6613 36323 6647
rect 36265 6607 36323 6613
rect 1104 6554 38824 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 34966 6554
rect 35018 6502 35030 6554
rect 35082 6502 35094 6554
rect 35146 6502 35158 6554
rect 35210 6502 38824 6554
rect 1104 6480 38824 6502
rect 2222 6440 2228 6452
rect 2183 6412 2228 6440
rect 2222 6400 2228 6412
rect 2280 6400 2286 6452
rect 2498 6400 2504 6452
rect 2556 6440 2562 6452
rect 3234 6440 3240 6452
rect 2556 6412 3240 6440
rect 2556 6400 2562 6412
rect 3234 6400 3240 6412
rect 3292 6440 3298 6452
rect 3697 6443 3755 6449
rect 3697 6440 3709 6443
rect 3292 6412 3709 6440
rect 3292 6400 3298 6412
rect 3697 6409 3709 6412
rect 3743 6409 3755 6443
rect 3697 6403 3755 6409
rect 3970 6400 3976 6452
rect 4028 6440 4034 6452
rect 4249 6443 4307 6449
rect 4249 6440 4261 6443
rect 4028 6412 4261 6440
rect 4028 6400 4034 6412
rect 4249 6409 4261 6412
rect 4295 6409 4307 6443
rect 4706 6440 4712 6452
rect 4667 6412 4712 6440
rect 4249 6403 4307 6409
rect 4264 6372 4292 6403
rect 4706 6400 4712 6412
rect 4764 6400 4770 6452
rect 7929 6443 7987 6449
rect 7929 6409 7941 6443
rect 7975 6440 7987 6443
rect 8202 6440 8208 6452
rect 7975 6412 8208 6440
rect 7975 6409 7987 6412
rect 7929 6403 7987 6409
rect 8202 6400 8208 6412
rect 8260 6400 8266 6452
rect 10042 6440 10048 6452
rect 10003 6412 10048 6440
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 11790 6440 11796 6452
rect 11751 6412 11796 6440
rect 11790 6400 11796 6412
rect 11848 6400 11854 6452
rect 13446 6440 13452 6452
rect 13407 6412 13452 6440
rect 13446 6400 13452 6412
rect 13504 6400 13510 6452
rect 13909 6443 13967 6449
rect 13909 6409 13921 6443
rect 13955 6440 13967 6443
rect 15102 6440 15108 6452
rect 13955 6412 15108 6440
rect 13955 6409 13967 6412
rect 13909 6403 13967 6409
rect 6546 6372 6552 6384
rect 4264 6344 6552 6372
rect 6546 6332 6552 6344
rect 6604 6332 6610 6384
rect 9309 6375 9367 6381
rect 9309 6341 9321 6375
rect 9355 6372 9367 6375
rect 9355 6344 10732 6372
rect 9355 6341 9367 6344
rect 9309 6335 9367 6341
rect 10704 6316 10732 6344
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6304 1915 6307
rect 1903 6276 2452 6304
rect 1903 6273 1915 6276
rect 1857 6267 1915 6273
rect 2222 6196 2228 6248
rect 2280 6236 2286 6248
rect 2317 6239 2375 6245
rect 2317 6236 2329 6239
rect 2280 6208 2329 6236
rect 2280 6196 2286 6208
rect 2317 6205 2329 6208
rect 2363 6205 2375 6239
rect 2424 6236 2452 6276
rect 6362 6264 6368 6316
rect 6420 6304 6426 6316
rect 7377 6307 7435 6313
rect 7377 6304 7389 6307
rect 6420 6276 7389 6304
rect 6420 6264 6426 6276
rect 7377 6273 7389 6276
rect 7423 6304 7435 6307
rect 8294 6304 8300 6316
rect 7423 6276 8300 6304
rect 7423 6273 7435 6276
rect 7377 6267 7435 6273
rect 8294 6264 8300 6276
rect 8352 6264 8358 6316
rect 10594 6304 10600 6316
rect 10555 6276 10600 6304
rect 10594 6264 10600 6276
rect 10652 6264 10658 6316
rect 10686 6264 10692 6316
rect 10744 6304 10750 6316
rect 10744 6276 10789 6304
rect 10744 6264 10750 6276
rect 11698 6264 11704 6316
rect 11756 6304 11762 6316
rect 14016 6313 14044 6412
rect 15102 6400 15108 6412
rect 15160 6400 15166 6452
rect 17494 6440 17500 6452
rect 17455 6412 17500 6440
rect 17494 6400 17500 6412
rect 17552 6400 17558 6452
rect 19978 6440 19984 6452
rect 19939 6412 19984 6440
rect 19978 6400 19984 6412
rect 20036 6400 20042 6452
rect 21910 6440 21916 6452
rect 21871 6412 21916 6440
rect 21910 6400 21916 6412
rect 21968 6400 21974 6452
rect 23477 6443 23535 6449
rect 23477 6409 23489 6443
rect 23523 6440 23535 6443
rect 23566 6440 23572 6452
rect 23523 6412 23572 6440
rect 23523 6409 23535 6412
rect 23477 6403 23535 6409
rect 23566 6400 23572 6412
rect 23624 6440 23630 6452
rect 24670 6440 24676 6452
rect 23624 6412 24164 6440
rect 24631 6412 24676 6440
rect 23624 6400 23630 6412
rect 22002 6332 22008 6384
rect 22060 6372 22066 6384
rect 24026 6372 24032 6384
rect 22060 6344 24032 6372
rect 22060 6332 22066 6344
rect 22572 6316 22600 6344
rect 24026 6332 24032 6344
rect 24084 6332 24090 6384
rect 12989 6307 13047 6313
rect 12989 6304 13001 6307
rect 11756 6276 13001 6304
rect 11756 6264 11762 6276
rect 12989 6273 13001 6276
rect 13035 6273 13047 6307
rect 12989 6267 13047 6273
rect 14001 6307 14059 6313
rect 14001 6273 14013 6307
rect 14047 6273 14059 6307
rect 14001 6267 14059 6273
rect 17310 6264 17316 6316
rect 17368 6304 17374 6316
rect 17865 6307 17923 6313
rect 17865 6304 17877 6307
rect 17368 6276 17877 6304
rect 17368 6264 17374 6276
rect 17865 6273 17877 6276
rect 17911 6304 17923 6307
rect 18046 6304 18052 6316
rect 17911 6276 18052 6304
rect 17911 6273 17923 6276
rect 17865 6267 17923 6273
rect 18046 6264 18052 6276
rect 18104 6264 18110 6316
rect 21177 6307 21235 6313
rect 21177 6273 21189 6307
rect 21223 6304 21235 6307
rect 21545 6307 21603 6313
rect 21545 6304 21557 6307
rect 21223 6276 21557 6304
rect 21223 6273 21235 6276
rect 21177 6267 21235 6273
rect 21545 6273 21557 6276
rect 21591 6304 21603 6307
rect 22370 6304 22376 6316
rect 21591 6276 22376 6304
rect 21591 6273 21603 6276
rect 21545 6267 21603 6273
rect 22370 6264 22376 6276
rect 22428 6304 22434 6316
rect 22465 6307 22523 6313
rect 22465 6304 22477 6307
rect 22428 6276 22477 6304
rect 22428 6264 22434 6276
rect 22465 6273 22477 6276
rect 22511 6273 22523 6307
rect 22465 6267 22523 6273
rect 22554 6264 22560 6316
rect 22612 6304 22618 6316
rect 24136 6313 24164 6412
rect 24670 6400 24676 6412
rect 24728 6400 24734 6452
rect 25133 6443 25191 6449
rect 25133 6409 25145 6443
rect 25179 6440 25191 6443
rect 25314 6440 25320 6452
rect 25179 6412 25320 6440
rect 25179 6409 25191 6412
rect 25133 6403 25191 6409
rect 25314 6400 25320 6412
rect 25372 6400 25378 6452
rect 25498 6440 25504 6452
rect 25459 6412 25504 6440
rect 25498 6400 25504 6412
rect 25556 6400 25562 6452
rect 28994 6440 29000 6452
rect 28955 6412 29000 6440
rect 28994 6400 29000 6412
rect 29052 6400 29058 6452
rect 32953 6443 33011 6449
rect 32953 6409 32965 6443
rect 32999 6440 33011 6443
rect 33042 6440 33048 6452
rect 32999 6412 33048 6440
rect 32999 6409 33011 6412
rect 32953 6403 33011 6409
rect 33042 6400 33048 6412
rect 33100 6400 33106 6452
rect 33321 6443 33379 6449
rect 33321 6409 33333 6443
rect 33367 6440 33379 6443
rect 33502 6440 33508 6452
rect 33367 6412 33508 6440
rect 33367 6409 33379 6412
rect 33321 6403 33379 6409
rect 33502 6400 33508 6412
rect 33560 6400 33566 6452
rect 33594 6400 33600 6452
rect 33652 6440 33658 6452
rect 35345 6443 35403 6449
rect 33652 6412 33697 6440
rect 33652 6400 33658 6412
rect 35345 6409 35357 6443
rect 35391 6440 35403 6443
rect 35618 6440 35624 6452
rect 35391 6412 35624 6440
rect 35391 6409 35403 6412
rect 35345 6403 35403 6409
rect 27525 6375 27583 6381
rect 27525 6372 27537 6375
rect 26436 6344 27537 6372
rect 24121 6307 24179 6313
rect 22612 6276 22657 6304
rect 22612 6264 22618 6276
rect 24121 6273 24133 6307
rect 24167 6273 24179 6307
rect 24121 6267 24179 6273
rect 24210 6264 24216 6316
rect 24268 6304 24274 6316
rect 26436 6313 26464 6344
rect 27525 6341 27537 6344
rect 27571 6341 27583 6375
rect 27525 6335 27583 6341
rect 27890 6332 27896 6384
rect 27948 6372 27954 6384
rect 27948 6344 28120 6372
rect 27948 6332 27954 6344
rect 25869 6307 25927 6313
rect 24268 6276 24313 6304
rect 24268 6264 24274 6276
rect 25869 6273 25881 6307
rect 25915 6304 25927 6307
rect 26421 6307 26479 6313
rect 26421 6304 26433 6307
rect 25915 6276 26433 6304
rect 25915 6273 25927 6276
rect 25869 6267 25927 6273
rect 26421 6273 26433 6276
rect 26467 6273 26479 6307
rect 26421 6267 26479 6273
rect 26513 6307 26571 6313
rect 26513 6273 26525 6307
rect 26559 6273 26571 6307
rect 26513 6267 26571 6273
rect 27433 6307 27491 6313
rect 27433 6273 27445 6307
rect 27479 6304 27491 6307
rect 27982 6304 27988 6316
rect 27479 6276 27988 6304
rect 27479 6273 27491 6276
rect 27433 6267 27491 6273
rect 2590 6245 2596 6248
rect 2584 6236 2596 6245
rect 2424 6208 2596 6236
rect 2317 6199 2375 6205
rect 2584 6199 2596 6208
rect 2590 6196 2596 6199
rect 2648 6196 2654 6248
rect 3970 6196 3976 6248
rect 4028 6236 4034 6248
rect 5261 6239 5319 6245
rect 5261 6236 5273 6239
rect 4028 6208 5273 6236
rect 4028 6196 4034 6208
rect 5261 6205 5273 6208
rect 5307 6236 5319 6239
rect 5813 6239 5871 6245
rect 5813 6236 5825 6239
rect 5307 6208 5825 6236
rect 5307 6205 5319 6208
rect 5261 6199 5319 6205
rect 5813 6205 5825 6208
rect 5859 6205 5871 6239
rect 5813 6199 5871 6205
rect 7193 6239 7251 6245
rect 7193 6205 7205 6239
rect 7239 6236 7251 6239
rect 7466 6236 7472 6248
rect 7239 6208 7472 6236
rect 7239 6205 7251 6208
rect 7193 6199 7251 6205
rect 7466 6196 7472 6208
rect 7524 6196 7530 6248
rect 8386 6236 8392 6248
rect 8347 6208 8392 6236
rect 8386 6196 8392 6208
rect 8444 6196 8450 6248
rect 9677 6239 9735 6245
rect 9677 6205 9689 6239
rect 9723 6236 9735 6239
rect 10505 6239 10563 6245
rect 10505 6236 10517 6239
rect 9723 6208 10517 6236
rect 9723 6205 9735 6208
rect 9677 6199 9735 6205
rect 10505 6205 10517 6208
rect 10551 6236 10563 6239
rect 10778 6236 10784 6248
rect 10551 6208 10784 6236
rect 10551 6205 10563 6208
rect 10505 6199 10563 6205
rect 10778 6196 10784 6208
rect 10836 6196 10842 6248
rect 12253 6239 12311 6245
rect 12253 6205 12265 6239
rect 12299 6236 12311 6239
rect 13170 6236 13176 6248
rect 12299 6208 13176 6236
rect 12299 6205 12311 6208
rect 12253 6199 12311 6205
rect 13170 6196 13176 6208
rect 13228 6196 13234 6248
rect 18064 6236 18092 6264
rect 19150 6236 19156 6248
rect 18064 6208 19156 6236
rect 19150 6196 19156 6208
rect 19208 6196 19214 6248
rect 24029 6239 24087 6245
rect 24029 6205 24041 6239
rect 24075 6236 24087 6239
rect 24670 6236 24676 6248
rect 24075 6208 24676 6236
rect 24075 6205 24087 6208
rect 24029 6199 24087 6205
rect 24670 6196 24676 6208
rect 24728 6196 24734 6248
rect 25406 6196 25412 6248
rect 25464 6236 25470 6248
rect 26528 6236 26556 6267
rect 27982 6264 27988 6276
rect 28040 6264 28046 6316
rect 28092 6313 28120 6344
rect 35452 6313 35480 6412
rect 35618 6400 35624 6412
rect 35676 6400 35682 6452
rect 35526 6332 35532 6384
rect 35584 6372 35590 6384
rect 35897 6375 35955 6381
rect 35897 6372 35909 6375
rect 35584 6344 35909 6372
rect 35584 6332 35590 6344
rect 35897 6341 35909 6344
rect 35943 6341 35955 6375
rect 35897 6335 35955 6341
rect 28077 6307 28135 6313
rect 28077 6273 28089 6307
rect 28123 6273 28135 6307
rect 28077 6267 28135 6273
rect 35437 6307 35495 6313
rect 35437 6273 35449 6307
rect 35483 6273 35495 6307
rect 35437 6267 35495 6273
rect 25464 6208 26556 6236
rect 25464 6196 25470 6208
rect 27614 6196 27620 6248
rect 27672 6236 27678 6248
rect 27893 6239 27951 6245
rect 27893 6236 27905 6239
rect 27672 6208 27905 6236
rect 27672 6196 27678 6208
rect 27893 6205 27905 6208
rect 27939 6236 27951 6239
rect 28994 6236 29000 6248
rect 27939 6208 29000 6236
rect 27939 6205 27951 6208
rect 27893 6199 27951 6205
rect 28994 6196 29000 6208
rect 29052 6196 29058 6248
rect 29270 6236 29276 6248
rect 29231 6208 29276 6236
rect 29270 6196 29276 6208
rect 29328 6236 29334 6248
rect 29825 6239 29883 6245
rect 29825 6236 29837 6239
rect 29328 6208 29837 6236
rect 29328 6196 29334 6208
rect 29825 6205 29837 6208
rect 29871 6205 29883 6239
rect 29825 6199 29883 6205
rect 6273 6171 6331 6177
rect 6273 6137 6285 6171
rect 6319 6168 6331 6171
rect 6638 6168 6644 6180
rect 6319 6140 6644 6168
rect 6319 6137 6331 6140
rect 6273 6131 6331 6137
rect 6638 6128 6644 6140
rect 6696 6128 6702 6180
rect 12066 6128 12072 6180
rect 12124 6168 12130 6180
rect 12897 6171 12955 6177
rect 12897 6168 12909 6171
rect 12124 6140 12909 6168
rect 12124 6128 12130 6140
rect 12897 6137 12909 6140
rect 12943 6168 12955 6171
rect 13906 6168 13912 6180
rect 12943 6140 13912 6168
rect 12943 6137 12955 6140
rect 12897 6131 12955 6137
rect 13906 6128 13912 6140
rect 13964 6128 13970 6180
rect 14268 6171 14326 6177
rect 14268 6137 14280 6171
rect 14314 6168 14326 6171
rect 14366 6168 14372 6180
rect 14314 6140 14372 6168
rect 14314 6137 14326 6140
rect 14268 6131 14326 6137
rect 14366 6128 14372 6140
rect 14424 6128 14430 6180
rect 16853 6171 16911 6177
rect 16853 6137 16865 6171
rect 16899 6168 16911 6171
rect 18294 6171 18352 6177
rect 18294 6168 18306 6171
rect 16899 6140 18306 6168
rect 16899 6137 16911 6140
rect 16853 6131 16911 6137
rect 18294 6137 18306 6140
rect 18340 6168 18352 6171
rect 18414 6168 18420 6180
rect 18340 6140 18420 6168
rect 18340 6137 18352 6140
rect 18294 6131 18352 6137
rect 18414 6128 18420 6140
rect 18472 6128 18478 6180
rect 22373 6171 22431 6177
rect 22373 6137 22385 6171
rect 22419 6168 22431 6171
rect 23017 6171 23075 6177
rect 23017 6168 23029 6171
rect 22419 6140 23029 6168
rect 22419 6137 22431 6140
rect 22373 6131 22431 6137
rect 23017 6137 23029 6140
rect 23063 6168 23075 6171
rect 23474 6168 23480 6180
rect 23063 6140 23480 6168
rect 23063 6137 23075 6140
rect 23017 6131 23075 6137
rect 23474 6128 23480 6140
rect 23532 6128 23538 6180
rect 29730 6128 29736 6180
rect 29788 6168 29794 6180
rect 30561 6171 30619 6177
rect 30561 6168 30573 6171
rect 29788 6140 30573 6168
rect 29788 6128 29794 6140
rect 30561 6137 30573 6140
rect 30607 6137 30619 6171
rect 30561 6131 30619 6137
rect 5074 6100 5080 6112
rect 5035 6072 5080 6100
rect 5074 6060 5080 6072
rect 5132 6060 5138 6112
rect 5442 6100 5448 6112
rect 5403 6072 5448 6100
rect 5442 6060 5448 6072
rect 5500 6060 5506 6112
rect 6822 6100 6828 6112
rect 6783 6072 6828 6100
rect 6822 6060 6828 6072
rect 6880 6060 6886 6112
rect 7282 6060 7288 6112
rect 7340 6100 7346 6112
rect 8205 6103 8263 6109
rect 8205 6100 8217 6103
rect 7340 6072 8217 6100
rect 7340 6060 7346 6072
rect 8205 6069 8217 6072
rect 8251 6069 8263 6103
rect 8570 6100 8576 6112
rect 8531 6072 8576 6100
rect 8205 6063 8263 6069
rect 8570 6060 8576 6072
rect 8628 6060 8634 6112
rect 9766 6060 9772 6112
rect 9824 6100 9830 6112
rect 10137 6103 10195 6109
rect 10137 6100 10149 6103
rect 9824 6072 10149 6100
rect 9824 6060 9830 6072
rect 10137 6069 10149 6072
rect 10183 6069 10195 6103
rect 10137 6063 10195 6069
rect 10962 6060 10968 6112
rect 11020 6100 11026 6112
rect 11425 6103 11483 6109
rect 11425 6100 11437 6103
rect 11020 6072 11437 6100
rect 11020 6060 11026 6072
rect 11425 6069 11437 6072
rect 11471 6100 11483 6103
rect 12158 6100 12164 6112
rect 11471 6072 12164 6100
rect 11471 6069 11483 6072
rect 11425 6063 11483 6069
rect 12158 6060 12164 6072
rect 12216 6060 12222 6112
rect 12434 6100 12440 6112
rect 12395 6072 12440 6100
rect 12434 6060 12440 6072
rect 12492 6060 12498 6112
rect 12526 6060 12532 6112
rect 12584 6100 12590 6112
rect 12805 6103 12863 6109
rect 12805 6100 12817 6103
rect 12584 6072 12817 6100
rect 12584 6060 12590 6072
rect 12805 6069 12817 6072
rect 12851 6069 12863 6103
rect 12805 6063 12863 6069
rect 13998 6060 14004 6112
rect 14056 6100 14062 6112
rect 15381 6103 15439 6109
rect 15381 6100 15393 6103
rect 14056 6072 15393 6100
rect 14056 6060 14062 6072
rect 15381 6069 15393 6072
rect 15427 6100 15439 6103
rect 15470 6100 15476 6112
rect 15427 6072 15476 6100
rect 15427 6069 15439 6072
rect 15381 6063 15439 6069
rect 15470 6060 15476 6072
rect 15528 6060 15534 6112
rect 16206 6060 16212 6112
rect 16264 6100 16270 6112
rect 16945 6103 17003 6109
rect 16945 6100 16957 6103
rect 16264 6072 16957 6100
rect 16264 6060 16270 6072
rect 16945 6069 16957 6072
rect 16991 6069 17003 6103
rect 16945 6063 17003 6069
rect 19334 6060 19340 6112
rect 19392 6100 19398 6112
rect 19429 6103 19487 6109
rect 19429 6100 19441 6103
rect 19392 6072 19441 6100
rect 19392 6060 19398 6072
rect 19429 6069 19441 6072
rect 19475 6069 19487 6103
rect 22002 6100 22008 6112
rect 21963 6072 22008 6100
rect 19429 6063 19487 6069
rect 22002 6060 22008 6072
rect 22060 6060 22066 6112
rect 23658 6100 23664 6112
rect 23619 6072 23664 6100
rect 23658 6060 23664 6072
rect 23716 6060 23722 6112
rect 25958 6100 25964 6112
rect 25919 6072 25964 6100
rect 25958 6060 25964 6072
rect 26016 6060 26022 6112
rect 26234 6060 26240 6112
rect 26292 6100 26298 6112
rect 26329 6103 26387 6109
rect 26329 6100 26341 6103
rect 26292 6072 26341 6100
rect 26292 6060 26298 6072
rect 26329 6069 26341 6072
rect 26375 6069 26387 6103
rect 26970 6100 26976 6112
rect 26931 6072 26976 6100
rect 26329 6063 26387 6069
rect 26970 6060 26976 6072
rect 27028 6060 27034 6112
rect 28074 6060 28080 6112
rect 28132 6100 28138 6112
rect 28537 6103 28595 6109
rect 28537 6100 28549 6103
rect 28132 6072 28549 6100
rect 28132 6060 28138 6072
rect 28537 6069 28549 6072
rect 28583 6069 28595 6103
rect 29454 6100 29460 6112
rect 29415 6072 29460 6100
rect 28537 6063 28595 6069
rect 29454 6060 29460 6072
rect 29512 6060 29518 6112
rect 30282 6100 30288 6112
rect 30243 6072 30288 6100
rect 30282 6060 30288 6072
rect 30340 6060 30346 6112
rect 1104 6010 38824 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 38824 6010
rect 1104 5936 38824 5958
rect 3970 5856 3976 5908
rect 4028 5896 4034 5908
rect 4065 5899 4123 5905
rect 4065 5896 4077 5899
rect 4028 5868 4077 5896
rect 4028 5856 4034 5868
rect 4065 5865 4077 5868
rect 4111 5865 4123 5899
rect 4065 5859 4123 5865
rect 4154 5856 4160 5908
rect 4212 5896 4218 5908
rect 4525 5899 4583 5905
rect 4525 5896 4537 5899
rect 4212 5868 4537 5896
rect 4212 5856 4218 5868
rect 4525 5865 4537 5868
rect 4571 5896 4583 5899
rect 4614 5896 4620 5908
rect 4571 5868 4620 5896
rect 4571 5865 4583 5868
rect 4525 5859 4583 5865
rect 4614 5856 4620 5868
rect 4672 5856 4678 5908
rect 5994 5896 6000 5908
rect 5955 5868 6000 5896
rect 5994 5856 6000 5868
rect 6052 5856 6058 5908
rect 6549 5899 6607 5905
rect 6549 5865 6561 5899
rect 6595 5896 6607 5899
rect 7282 5896 7288 5908
rect 6595 5868 7288 5896
rect 6595 5865 6607 5868
rect 6549 5859 6607 5865
rect 7282 5856 7288 5868
rect 7340 5856 7346 5908
rect 7558 5896 7564 5908
rect 7519 5868 7564 5896
rect 7558 5856 7564 5868
rect 7616 5856 7622 5908
rect 8294 5896 8300 5908
rect 8255 5868 8300 5896
rect 8294 5856 8300 5868
rect 8352 5856 8358 5908
rect 10594 5896 10600 5908
rect 10555 5868 10600 5896
rect 10594 5856 10600 5868
rect 10652 5856 10658 5908
rect 11698 5896 11704 5908
rect 11659 5868 11704 5896
rect 11698 5856 11704 5868
rect 11756 5856 11762 5908
rect 12802 5896 12808 5908
rect 12763 5868 12808 5896
rect 12802 5856 12808 5868
rect 12860 5856 12866 5908
rect 13170 5896 13176 5908
rect 13131 5868 13176 5896
rect 13170 5856 13176 5868
rect 13228 5896 13234 5908
rect 13814 5896 13820 5908
rect 13228 5868 13820 5896
rect 13228 5856 13234 5868
rect 13814 5856 13820 5868
rect 13872 5856 13878 5908
rect 14366 5896 14372 5908
rect 14327 5868 14372 5896
rect 14366 5856 14372 5868
rect 14424 5856 14430 5908
rect 16485 5899 16543 5905
rect 16485 5865 16497 5899
rect 16531 5896 16543 5899
rect 16942 5896 16948 5908
rect 16531 5868 16948 5896
rect 16531 5865 16543 5868
rect 16485 5859 16543 5865
rect 16942 5856 16948 5868
rect 17000 5856 17006 5908
rect 17681 5899 17739 5905
rect 17681 5865 17693 5899
rect 17727 5896 17739 5899
rect 17954 5896 17960 5908
rect 17727 5868 17960 5896
rect 17727 5865 17739 5868
rect 17681 5859 17739 5865
rect 17954 5856 17960 5868
rect 18012 5856 18018 5908
rect 22281 5899 22339 5905
rect 22281 5865 22293 5899
rect 22327 5896 22339 5899
rect 22370 5896 22376 5908
rect 22327 5868 22376 5896
rect 22327 5865 22339 5868
rect 22281 5859 22339 5865
rect 22370 5856 22376 5868
rect 22428 5856 22434 5908
rect 23293 5899 23351 5905
rect 23293 5865 23305 5899
rect 23339 5896 23351 5899
rect 23658 5896 23664 5908
rect 23339 5868 23664 5896
rect 23339 5865 23351 5868
rect 23293 5859 23351 5865
rect 23658 5856 23664 5868
rect 23716 5896 23722 5908
rect 23753 5899 23811 5905
rect 23753 5896 23765 5899
rect 23716 5868 23765 5896
rect 23716 5856 23722 5868
rect 23753 5865 23765 5868
rect 23799 5865 23811 5899
rect 23753 5859 23811 5865
rect 23842 5856 23848 5908
rect 23900 5896 23906 5908
rect 25501 5899 25559 5905
rect 23900 5868 23945 5896
rect 23900 5856 23906 5868
rect 25501 5865 25513 5899
rect 25547 5865 25559 5899
rect 26510 5896 26516 5908
rect 26471 5868 26516 5896
rect 25501 5859 25559 5865
rect 1664 5831 1722 5837
rect 1664 5797 1676 5831
rect 1710 5828 1722 5831
rect 2498 5828 2504 5840
rect 1710 5800 2504 5828
rect 1710 5797 1722 5800
rect 1664 5791 1722 5797
rect 2498 5788 2504 5800
rect 2556 5788 2562 5840
rect 4430 5828 4436 5840
rect 4391 5800 4436 5828
rect 4430 5788 4436 5800
rect 4488 5828 4494 5840
rect 5534 5828 5540 5840
rect 4488 5800 5540 5828
rect 4488 5788 4494 5800
rect 5534 5788 5540 5800
rect 5592 5788 5598 5840
rect 6457 5831 6515 5837
rect 6457 5797 6469 5831
rect 6503 5828 6515 5831
rect 7466 5828 7472 5840
rect 6503 5800 7472 5828
rect 6503 5797 6515 5800
rect 6457 5791 6515 5797
rect 7466 5788 7472 5800
rect 7524 5788 7530 5840
rect 10321 5831 10379 5837
rect 10321 5797 10333 5831
rect 10367 5828 10379 5831
rect 10686 5828 10692 5840
rect 10367 5800 10692 5828
rect 10367 5797 10379 5800
rect 10321 5791 10379 5797
rect 10686 5788 10692 5800
rect 10744 5788 10750 5840
rect 11514 5788 11520 5840
rect 11572 5828 11578 5840
rect 12253 5831 12311 5837
rect 12253 5828 12265 5831
rect 11572 5800 12265 5828
rect 11572 5788 11578 5800
rect 12253 5797 12265 5800
rect 12299 5828 12311 5831
rect 12434 5828 12440 5840
rect 12299 5800 12440 5828
rect 12299 5797 12311 5800
rect 12253 5791 12311 5797
rect 12434 5788 12440 5800
rect 12492 5788 12498 5840
rect 16850 5828 16856 5840
rect 16811 5800 16856 5828
rect 16850 5788 16856 5800
rect 16908 5788 16914 5840
rect 17313 5831 17371 5837
rect 17313 5797 17325 5831
rect 17359 5828 17371 5831
rect 18233 5831 18291 5837
rect 18233 5828 18245 5831
rect 17359 5800 18245 5828
rect 17359 5797 17371 5800
rect 17313 5791 17371 5797
rect 18233 5797 18245 5800
rect 18279 5797 18291 5831
rect 25516 5828 25544 5859
rect 26510 5856 26516 5868
rect 26568 5856 26574 5908
rect 27614 5896 27620 5908
rect 27575 5868 27620 5896
rect 27614 5856 27620 5868
rect 27672 5856 27678 5908
rect 27890 5896 27896 5908
rect 27851 5868 27896 5896
rect 27890 5856 27896 5868
rect 27948 5856 27954 5908
rect 30282 5856 30288 5908
rect 30340 5896 30346 5908
rect 30377 5899 30435 5905
rect 30377 5896 30389 5899
rect 30340 5868 30389 5896
rect 30340 5856 30346 5868
rect 30377 5865 30389 5868
rect 30423 5865 30435 5899
rect 30742 5896 30748 5908
rect 30703 5868 30748 5896
rect 30377 5859 30435 5865
rect 30742 5856 30748 5868
rect 30800 5856 30806 5908
rect 35345 5899 35403 5905
rect 35345 5865 35357 5899
rect 35391 5896 35403 5899
rect 35434 5896 35440 5908
rect 35391 5868 35440 5896
rect 35391 5865 35403 5868
rect 35345 5859 35403 5865
rect 35434 5856 35440 5868
rect 35492 5856 35498 5908
rect 28344 5831 28402 5837
rect 25516 5800 27200 5828
rect 18233 5791 18291 5797
rect 1397 5763 1455 5769
rect 1397 5729 1409 5763
rect 1443 5760 1455 5763
rect 1486 5760 1492 5772
rect 1443 5732 1492 5760
rect 1443 5729 1455 5732
rect 1397 5723 1455 5729
rect 1486 5720 1492 5732
rect 1544 5760 1550 5772
rect 2222 5760 2228 5772
rect 1544 5732 2228 5760
rect 1544 5720 1550 5732
rect 2222 5720 2228 5732
rect 2280 5720 2286 5772
rect 6914 5720 6920 5772
rect 6972 5760 6978 5772
rect 7190 5760 7196 5772
rect 6972 5732 7196 5760
rect 6972 5720 6978 5732
rect 7190 5720 7196 5732
rect 7248 5720 7254 5772
rect 8110 5760 8116 5772
rect 8071 5732 8116 5760
rect 8110 5720 8116 5732
rect 8168 5720 8174 5772
rect 9674 5760 9680 5772
rect 9635 5732 9680 5760
rect 9674 5720 9680 5732
rect 9732 5720 9738 5772
rect 10781 5763 10839 5769
rect 10781 5729 10793 5763
rect 10827 5760 10839 5763
rect 11790 5760 11796 5772
rect 10827 5732 11796 5760
rect 10827 5729 10839 5732
rect 10781 5723 10839 5729
rect 11790 5720 11796 5732
rect 11848 5760 11854 5772
rect 12161 5763 12219 5769
rect 12161 5760 12173 5763
rect 11848 5732 12173 5760
rect 11848 5720 11854 5732
rect 12161 5729 12173 5732
rect 12207 5729 12219 5763
rect 13722 5760 13728 5772
rect 13683 5732 13728 5760
rect 12161 5723 12219 5729
rect 13722 5720 13728 5732
rect 13780 5720 13786 5772
rect 15657 5763 15715 5769
rect 15657 5729 15669 5763
rect 15703 5760 15715 5763
rect 15930 5760 15936 5772
rect 15703 5732 15936 5760
rect 15703 5729 15715 5732
rect 15657 5723 15715 5729
rect 15930 5720 15936 5732
rect 15988 5720 15994 5772
rect 17328 5760 17356 5791
rect 17236 5732 17356 5760
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5692 4767 5695
rect 4755 5664 5120 5692
rect 4755 5661 4767 5664
rect 4709 5655 4767 5661
rect 3050 5584 3056 5636
rect 3108 5624 3114 5636
rect 3510 5624 3516 5636
rect 3108 5596 3516 5624
rect 3108 5584 3114 5596
rect 3510 5584 3516 5596
rect 3568 5624 3574 5636
rect 3697 5627 3755 5633
rect 3697 5624 3709 5627
rect 3568 5596 3709 5624
rect 3568 5584 3574 5596
rect 3697 5593 3709 5596
rect 3743 5593 3755 5627
rect 3697 5587 3755 5593
rect 5092 5568 5120 5664
rect 6638 5652 6644 5704
rect 6696 5692 6702 5704
rect 7009 5695 7067 5701
rect 7009 5692 7021 5695
rect 6696 5664 7021 5692
rect 6696 5652 6702 5664
rect 7009 5661 7021 5664
rect 7055 5661 7067 5695
rect 7009 5655 7067 5661
rect 7101 5695 7159 5701
rect 7101 5661 7113 5695
rect 7147 5692 7159 5695
rect 7374 5692 7380 5704
rect 7147 5664 7380 5692
rect 7147 5661 7159 5664
rect 7101 5655 7159 5661
rect 5994 5584 6000 5636
rect 6052 5624 6058 5636
rect 7116 5624 7144 5655
rect 7374 5652 7380 5664
rect 7432 5692 7438 5704
rect 8202 5692 8208 5704
rect 7432 5664 8208 5692
rect 7432 5652 7438 5664
rect 8202 5652 8208 5664
rect 8260 5652 8266 5704
rect 12342 5692 12348 5704
rect 12303 5664 12348 5692
rect 12342 5652 12348 5664
rect 12400 5652 12406 5704
rect 13170 5652 13176 5704
rect 13228 5692 13234 5704
rect 13817 5695 13875 5701
rect 13817 5692 13829 5695
rect 13228 5664 13829 5692
rect 13228 5652 13234 5664
rect 13817 5661 13829 5664
rect 13863 5661 13875 5695
rect 13998 5692 14004 5704
rect 13959 5664 14004 5692
rect 13817 5655 13875 5661
rect 9858 5624 9864 5636
rect 6052 5596 7144 5624
rect 9819 5596 9864 5624
rect 6052 5584 6058 5596
rect 9858 5584 9864 5596
rect 9916 5584 9922 5636
rect 13832 5624 13860 5655
rect 13998 5652 14004 5664
rect 14056 5652 14062 5704
rect 15746 5692 15752 5704
rect 15707 5664 15752 5692
rect 15746 5652 15752 5664
rect 15804 5652 15810 5704
rect 15841 5695 15899 5701
rect 15841 5661 15853 5695
rect 15887 5661 15899 5695
rect 15841 5655 15899 5661
rect 14737 5627 14795 5633
rect 14737 5624 14749 5627
rect 13832 5596 14749 5624
rect 14737 5593 14749 5596
rect 14783 5593 14795 5627
rect 14737 5587 14795 5593
rect 15470 5584 15476 5636
rect 15528 5624 15534 5636
rect 15856 5624 15884 5655
rect 15528 5596 15884 5624
rect 15528 5584 15534 5596
rect 16482 5584 16488 5636
rect 16540 5624 16546 5636
rect 17236 5624 17264 5732
rect 18046 5720 18052 5772
rect 18104 5760 18110 5772
rect 18141 5763 18199 5769
rect 18141 5760 18153 5763
rect 18104 5732 18153 5760
rect 18104 5720 18110 5732
rect 18141 5729 18153 5732
rect 18187 5729 18199 5763
rect 18874 5760 18880 5772
rect 18835 5732 18880 5760
rect 18141 5723 18199 5729
rect 18874 5720 18880 5732
rect 18932 5720 18938 5772
rect 20714 5720 20720 5772
rect 20772 5760 20778 5772
rect 21157 5763 21215 5769
rect 21157 5760 21169 5763
rect 20772 5732 21169 5760
rect 20772 5720 20778 5732
rect 21157 5729 21169 5732
rect 21203 5729 21215 5763
rect 21157 5723 21215 5729
rect 25317 5763 25375 5769
rect 25317 5729 25329 5763
rect 25363 5760 25375 5763
rect 26326 5760 26332 5772
rect 25363 5732 26332 5760
rect 25363 5729 25375 5732
rect 25317 5723 25375 5729
rect 26326 5720 26332 5732
rect 26384 5720 26390 5772
rect 26694 5720 26700 5772
rect 26752 5760 26758 5772
rect 26881 5763 26939 5769
rect 26881 5760 26893 5763
rect 26752 5732 26893 5760
rect 26752 5720 26758 5732
rect 26881 5729 26893 5732
rect 26927 5729 26939 5763
rect 26881 5723 26939 5729
rect 27172 5704 27200 5800
rect 28344 5797 28356 5831
rect 28390 5828 28402 5831
rect 28718 5828 28724 5840
rect 28390 5800 28724 5828
rect 28390 5797 28402 5800
rect 28344 5791 28402 5797
rect 28718 5788 28724 5800
rect 28776 5828 28782 5840
rect 29638 5828 29644 5840
rect 28776 5800 29644 5828
rect 28776 5788 28782 5800
rect 29638 5788 29644 5800
rect 29696 5788 29702 5840
rect 30561 5763 30619 5769
rect 30561 5729 30573 5763
rect 30607 5760 30619 5763
rect 30834 5760 30840 5772
rect 30607 5732 30840 5760
rect 30607 5729 30619 5732
rect 30561 5723 30619 5729
rect 30834 5720 30840 5732
rect 30892 5720 30898 5772
rect 18325 5695 18383 5701
rect 18325 5661 18337 5695
rect 18371 5661 18383 5695
rect 18325 5655 18383 5661
rect 19429 5695 19487 5701
rect 19429 5661 19441 5695
rect 19475 5692 19487 5695
rect 20530 5692 20536 5704
rect 19475 5664 20536 5692
rect 19475 5661 19487 5664
rect 19429 5655 19487 5661
rect 16540 5596 17264 5624
rect 16540 5584 16546 5596
rect 17954 5584 17960 5636
rect 18012 5624 18018 5636
rect 18340 5624 18368 5655
rect 20530 5652 20536 5664
rect 20588 5652 20594 5704
rect 20898 5692 20904 5704
rect 20859 5664 20904 5692
rect 20898 5652 20904 5664
rect 20956 5652 20962 5704
rect 24029 5695 24087 5701
rect 24029 5661 24041 5695
rect 24075 5692 24087 5695
rect 24210 5692 24216 5704
rect 24075 5664 24216 5692
rect 24075 5661 24087 5664
rect 24029 5655 24087 5661
rect 24210 5652 24216 5664
rect 24268 5692 24274 5704
rect 25133 5695 25191 5701
rect 25133 5692 25145 5695
rect 24268 5664 25145 5692
rect 24268 5652 24274 5664
rect 25133 5661 25145 5664
rect 25179 5692 25191 5695
rect 25406 5692 25412 5704
rect 25179 5664 25412 5692
rect 25179 5661 25191 5664
rect 25133 5655 25191 5661
rect 25406 5652 25412 5664
rect 25464 5652 25470 5704
rect 26970 5692 26976 5704
rect 26931 5664 26976 5692
rect 26970 5652 26976 5664
rect 27028 5652 27034 5704
rect 27154 5652 27160 5704
rect 27212 5692 27218 5704
rect 28074 5692 28080 5704
rect 27212 5664 27305 5692
rect 28035 5664 28080 5692
rect 27212 5652 27218 5664
rect 28074 5652 28080 5664
rect 28132 5652 28138 5704
rect 32030 5652 32036 5704
rect 32088 5692 32094 5704
rect 32125 5695 32183 5701
rect 32125 5692 32137 5695
rect 32088 5664 32137 5692
rect 32088 5652 32094 5664
rect 32125 5661 32137 5664
rect 32171 5661 32183 5695
rect 32125 5655 32183 5661
rect 18012 5596 18368 5624
rect 18012 5584 18018 5596
rect 22462 5584 22468 5636
rect 22520 5624 22526 5636
rect 23385 5627 23443 5633
rect 23385 5624 23397 5627
rect 22520 5596 23397 5624
rect 22520 5584 22526 5596
rect 23385 5593 23397 5596
rect 23431 5593 23443 5627
rect 23385 5587 23443 5593
rect 2774 5556 2780 5568
rect 2735 5528 2780 5556
rect 2774 5516 2780 5528
rect 2832 5516 2838 5568
rect 3326 5556 3332 5568
rect 3287 5528 3332 5556
rect 3326 5516 3332 5528
rect 3384 5516 3390 5568
rect 5074 5556 5080 5568
rect 5035 5528 5080 5556
rect 5074 5516 5080 5528
rect 5132 5556 5138 5568
rect 5445 5559 5503 5565
rect 5445 5556 5457 5559
rect 5132 5528 5457 5556
rect 5132 5516 5138 5528
rect 5445 5525 5457 5528
rect 5491 5525 5503 5559
rect 5445 5519 5503 5525
rect 7466 5516 7472 5568
rect 7524 5556 7530 5568
rect 7929 5559 7987 5565
rect 7929 5556 7941 5559
rect 7524 5528 7941 5556
rect 7524 5516 7530 5528
rect 7929 5525 7941 5528
rect 7975 5525 7987 5559
rect 7929 5519 7987 5525
rect 11606 5516 11612 5568
rect 11664 5556 11670 5568
rect 11793 5559 11851 5565
rect 11793 5556 11805 5559
rect 11664 5528 11805 5556
rect 11664 5516 11670 5528
rect 11793 5525 11805 5528
rect 11839 5525 11851 5559
rect 13354 5556 13360 5568
rect 13315 5528 13360 5556
rect 11793 5519 11851 5525
rect 13354 5516 13360 5528
rect 13412 5516 13418 5568
rect 15286 5556 15292 5568
rect 15247 5528 15292 5556
rect 15286 5516 15292 5528
rect 15344 5516 15350 5568
rect 17773 5559 17831 5565
rect 17773 5525 17785 5559
rect 17819 5556 17831 5559
rect 17862 5556 17868 5568
rect 17819 5528 17868 5556
rect 17819 5525 17831 5528
rect 17773 5519 17831 5525
rect 17862 5516 17868 5528
rect 17920 5516 17926 5568
rect 19886 5556 19892 5568
rect 19847 5528 19892 5556
rect 19886 5516 19892 5528
rect 19944 5516 19950 5568
rect 22830 5556 22836 5568
rect 22791 5528 22836 5556
rect 22830 5516 22836 5528
rect 22888 5516 22894 5568
rect 24118 5516 24124 5568
rect 24176 5556 24182 5568
rect 24397 5559 24455 5565
rect 24397 5556 24409 5559
rect 24176 5528 24409 5556
rect 24176 5516 24182 5528
rect 24397 5525 24409 5528
rect 24443 5525 24455 5559
rect 24854 5556 24860 5568
rect 24815 5528 24860 5556
rect 24397 5519 24455 5525
rect 24854 5516 24860 5528
rect 24912 5516 24918 5568
rect 26053 5559 26111 5565
rect 26053 5525 26065 5559
rect 26099 5556 26111 5559
rect 26234 5556 26240 5568
rect 26099 5528 26240 5556
rect 26099 5525 26111 5528
rect 26053 5519 26111 5525
rect 26234 5516 26240 5528
rect 26292 5516 26298 5568
rect 28994 5516 29000 5568
rect 29052 5556 29058 5568
rect 29457 5559 29515 5565
rect 29457 5556 29469 5559
rect 29052 5528 29469 5556
rect 29052 5516 29058 5528
rect 29457 5525 29469 5528
rect 29503 5525 29515 5559
rect 30098 5556 30104 5568
rect 30059 5528 30104 5556
rect 29457 5519 29515 5525
rect 30098 5516 30104 5528
rect 30156 5516 30162 5568
rect 31202 5556 31208 5568
rect 31163 5528 31208 5556
rect 31202 5516 31208 5528
rect 31260 5516 31266 5568
rect 31754 5516 31760 5568
rect 31812 5556 31818 5568
rect 31812 5528 31857 5556
rect 31812 5516 31818 5528
rect 1104 5466 38824 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 34966 5466
rect 35018 5414 35030 5466
rect 35082 5414 35094 5466
rect 35146 5414 35158 5466
rect 35210 5414 38824 5466
rect 1104 5392 38824 5414
rect 1486 5312 1492 5364
rect 1544 5352 1550 5364
rect 1581 5355 1639 5361
rect 1581 5352 1593 5355
rect 1544 5324 1593 5352
rect 1544 5312 1550 5324
rect 1581 5321 1593 5324
rect 1627 5352 1639 5355
rect 1949 5355 2007 5361
rect 1949 5352 1961 5355
rect 1627 5324 1961 5352
rect 1627 5321 1639 5324
rect 1581 5315 1639 5321
rect 1949 5321 1961 5324
rect 1995 5321 2007 5355
rect 3234 5352 3240 5364
rect 3195 5324 3240 5352
rect 1949 5315 2007 5321
rect 3234 5312 3240 5324
rect 3292 5312 3298 5364
rect 4614 5352 4620 5364
rect 4575 5324 4620 5352
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 5534 5312 5540 5364
rect 5592 5352 5598 5364
rect 5721 5355 5779 5361
rect 5721 5352 5733 5355
rect 5592 5324 5733 5352
rect 5592 5312 5598 5324
rect 5721 5321 5733 5324
rect 5767 5321 5779 5355
rect 5721 5315 5779 5321
rect 6273 5355 6331 5361
rect 6273 5321 6285 5355
rect 6319 5352 6331 5355
rect 6730 5352 6736 5364
rect 6319 5324 6736 5352
rect 6319 5321 6331 5324
rect 6273 5315 6331 5321
rect 6730 5312 6736 5324
rect 6788 5312 6794 5364
rect 9674 5312 9680 5364
rect 9732 5352 9738 5364
rect 10045 5355 10103 5361
rect 10045 5352 10057 5355
rect 9732 5324 10057 5352
rect 9732 5312 9738 5324
rect 10045 5321 10057 5324
rect 10091 5321 10103 5355
rect 11790 5352 11796 5364
rect 11751 5324 11796 5352
rect 10045 5315 10103 5321
rect 11790 5312 11796 5324
rect 11848 5312 11854 5364
rect 12713 5355 12771 5361
rect 12713 5321 12725 5355
rect 12759 5352 12771 5355
rect 13722 5352 13728 5364
rect 12759 5324 13728 5352
rect 12759 5321 12771 5324
rect 12713 5315 12771 5321
rect 13722 5312 13728 5324
rect 13780 5312 13786 5364
rect 13906 5312 13912 5364
rect 13964 5352 13970 5364
rect 14550 5352 14556 5364
rect 13964 5324 14556 5352
rect 13964 5312 13970 5324
rect 14550 5312 14556 5324
rect 14608 5352 14614 5364
rect 15013 5355 15071 5361
rect 15013 5352 15025 5355
rect 14608 5324 15025 5352
rect 14608 5312 14614 5324
rect 15013 5321 15025 5324
rect 15059 5321 15071 5355
rect 15013 5315 15071 5321
rect 15657 5355 15715 5361
rect 15657 5321 15669 5355
rect 15703 5352 15715 5355
rect 15746 5352 15752 5364
rect 15703 5324 15752 5352
rect 15703 5321 15715 5324
rect 15657 5315 15715 5321
rect 15746 5312 15752 5324
rect 15804 5312 15810 5364
rect 15930 5352 15936 5364
rect 15891 5324 15936 5352
rect 15930 5312 15936 5324
rect 15988 5312 15994 5364
rect 17497 5355 17555 5361
rect 17497 5321 17509 5355
rect 17543 5352 17555 5355
rect 17770 5352 17776 5364
rect 17543 5324 17776 5352
rect 17543 5321 17555 5324
rect 17497 5315 17555 5321
rect 17770 5312 17776 5324
rect 17828 5312 17834 5364
rect 18138 5312 18144 5364
rect 18196 5352 18202 5364
rect 18417 5355 18475 5361
rect 18417 5352 18429 5355
rect 18196 5324 18429 5352
rect 18196 5312 18202 5324
rect 18417 5321 18429 5324
rect 18463 5321 18475 5355
rect 19150 5352 19156 5364
rect 19111 5324 19156 5352
rect 18417 5315 18475 5321
rect 19150 5312 19156 5324
rect 19208 5312 19214 5364
rect 20714 5352 20720 5364
rect 20675 5324 20720 5352
rect 20714 5312 20720 5324
rect 20772 5352 20778 5364
rect 21637 5355 21695 5361
rect 21637 5352 21649 5355
rect 20772 5324 21649 5352
rect 20772 5312 20778 5324
rect 21637 5321 21649 5324
rect 21683 5321 21695 5355
rect 21637 5315 21695 5321
rect 23477 5355 23535 5361
rect 23477 5321 23489 5355
rect 23523 5352 23535 5355
rect 23842 5352 23848 5364
rect 23523 5324 23848 5352
rect 23523 5321 23535 5324
rect 23477 5315 23535 5321
rect 23842 5312 23848 5324
rect 23900 5312 23906 5364
rect 25038 5352 25044 5364
rect 24999 5324 25044 5352
rect 25038 5312 25044 5324
rect 25096 5312 25102 5364
rect 26234 5312 26240 5364
rect 26292 5352 26298 5364
rect 27341 5355 27399 5361
rect 27341 5352 27353 5355
rect 26292 5324 27353 5352
rect 26292 5312 26298 5324
rect 27341 5321 27353 5324
rect 27387 5321 27399 5355
rect 28718 5352 28724 5364
rect 27341 5315 27399 5321
rect 27816 5324 28724 5352
rect 6638 5284 6644 5296
rect 6599 5256 6644 5284
rect 6638 5244 6644 5256
rect 6696 5244 6702 5296
rect 15102 5244 15108 5296
rect 15160 5284 15166 5296
rect 15948 5284 15976 5312
rect 15160 5256 15976 5284
rect 15160 5244 15166 5256
rect 2685 5219 2743 5225
rect 2685 5185 2697 5219
rect 2731 5216 2743 5219
rect 3050 5216 3056 5228
rect 2731 5188 3056 5216
rect 2731 5185 2743 5188
rect 2685 5179 2743 5185
rect 3050 5176 3056 5188
rect 3108 5176 3114 5228
rect 5442 5216 5448 5228
rect 4816 5188 5448 5216
rect 2590 5108 2596 5160
rect 2648 5148 2654 5160
rect 2774 5148 2780 5160
rect 2648 5120 2780 5148
rect 2648 5108 2654 5120
rect 2774 5108 2780 5120
rect 2832 5148 2838 5160
rect 4816 5157 4844 5188
rect 5442 5176 5448 5188
rect 5500 5176 5506 5228
rect 7282 5216 7288 5228
rect 7243 5188 7288 5216
rect 7282 5176 7288 5188
rect 7340 5176 7346 5228
rect 7466 5216 7472 5228
rect 7427 5188 7472 5216
rect 7466 5176 7472 5188
rect 7524 5176 7530 5228
rect 12253 5219 12311 5225
rect 12253 5185 12265 5219
rect 12299 5216 12311 5219
rect 13354 5216 13360 5228
rect 12299 5188 13360 5216
rect 12299 5185 12311 5188
rect 12253 5179 12311 5185
rect 13354 5176 13360 5188
rect 13412 5216 13418 5228
rect 13633 5219 13691 5225
rect 13633 5216 13645 5219
rect 13412 5188 13645 5216
rect 13412 5176 13418 5188
rect 13633 5185 13645 5188
rect 13679 5185 13691 5219
rect 13633 5179 13691 5185
rect 13814 5176 13820 5228
rect 13872 5216 13878 5228
rect 13909 5219 13967 5225
rect 13909 5216 13921 5219
rect 13872 5188 13921 5216
rect 13872 5176 13878 5188
rect 13909 5185 13921 5188
rect 13955 5185 13967 5219
rect 13909 5179 13967 5185
rect 16850 5176 16856 5228
rect 16908 5216 16914 5228
rect 16945 5219 17003 5225
rect 16945 5216 16957 5219
rect 16908 5188 16957 5216
rect 16908 5176 16914 5188
rect 16945 5185 16957 5188
rect 16991 5185 17003 5219
rect 16945 5179 17003 5185
rect 18966 5176 18972 5228
rect 19024 5216 19030 5228
rect 19168 5216 19196 5312
rect 22002 5284 22008 5296
rect 21963 5256 22008 5284
rect 22002 5244 22008 5256
rect 22060 5244 22066 5296
rect 23661 5287 23719 5293
rect 23661 5253 23673 5287
rect 23707 5284 23719 5287
rect 24762 5284 24768 5296
rect 23707 5256 24768 5284
rect 23707 5253 23719 5256
rect 23661 5247 23719 5253
rect 24762 5244 24768 5256
rect 24820 5244 24826 5296
rect 25225 5287 25283 5293
rect 25225 5253 25237 5287
rect 25271 5284 25283 5287
rect 26421 5287 26479 5293
rect 26421 5284 26433 5287
rect 25271 5256 26433 5284
rect 25271 5253 25283 5256
rect 25225 5247 25283 5253
rect 26421 5253 26433 5256
rect 26467 5284 26479 5287
rect 26970 5284 26976 5296
rect 26467 5256 26976 5284
rect 26467 5253 26479 5256
rect 26421 5247 26479 5253
rect 26970 5244 26976 5256
rect 27028 5244 27034 5296
rect 27249 5287 27307 5293
rect 27249 5253 27261 5287
rect 27295 5284 27307 5287
rect 27816 5284 27844 5324
rect 28718 5312 28724 5324
rect 28776 5312 28782 5364
rect 31202 5312 31208 5364
rect 31260 5352 31266 5364
rect 31665 5355 31723 5361
rect 31665 5352 31677 5355
rect 31260 5324 31677 5352
rect 31260 5312 31266 5324
rect 31665 5321 31677 5324
rect 31711 5321 31723 5355
rect 31665 5315 31723 5321
rect 27295 5256 27844 5284
rect 27295 5253 27307 5256
rect 27249 5247 27307 5253
rect 19337 5219 19395 5225
rect 19337 5216 19349 5219
rect 19024 5188 19349 5216
rect 19024 5176 19030 5188
rect 19337 5185 19349 5188
rect 19383 5185 19395 5219
rect 22554 5216 22560 5228
rect 22515 5188 22560 5216
rect 19337 5179 19395 5185
rect 3513 5151 3571 5157
rect 3513 5148 3525 5151
rect 2832 5120 3525 5148
rect 2832 5108 2838 5120
rect 3513 5117 3525 5120
rect 3559 5117 3571 5151
rect 3513 5111 3571 5117
rect 3697 5151 3755 5157
rect 3697 5117 3709 5151
rect 3743 5117 3755 5151
rect 3697 5111 3755 5117
rect 4801 5151 4859 5157
rect 4801 5117 4813 5151
rect 4847 5117 4859 5151
rect 4801 5111 4859 5117
rect 7193 5151 7251 5157
rect 7193 5117 7205 5151
rect 7239 5148 7251 5151
rect 7558 5148 7564 5160
rect 7239 5120 7564 5148
rect 7239 5117 7251 5120
rect 7193 5111 7251 5117
rect 2501 5083 2559 5089
rect 2501 5049 2513 5083
rect 2547 5080 2559 5083
rect 3326 5080 3332 5092
rect 2547 5052 3332 5080
rect 2547 5049 2559 5052
rect 2501 5043 2559 5049
rect 3326 5040 3332 5052
rect 3384 5040 3390 5092
rect 3712 5080 3740 5111
rect 7558 5108 7564 5120
rect 7616 5108 7622 5160
rect 8389 5151 8447 5157
rect 8389 5117 8401 5151
rect 8435 5148 8447 5151
rect 9493 5151 9551 5157
rect 9493 5148 9505 5151
rect 8435 5120 9076 5148
rect 8435 5117 8447 5120
rect 8389 5111 8447 5117
rect 4338 5080 4344 5092
rect 3712 5052 4344 5080
rect 4338 5040 4344 5052
rect 4396 5040 4402 5092
rect 9048 5024 9076 5120
rect 9324 5120 9505 5148
rect 9324 5024 9352 5120
rect 9493 5117 9505 5120
rect 9539 5117 9551 5151
rect 10594 5148 10600 5160
rect 10555 5120 10600 5148
rect 9493 5111 9551 5117
rect 10594 5108 10600 5120
rect 10652 5148 10658 5160
rect 11149 5151 11207 5157
rect 11149 5148 11161 5151
rect 10652 5120 11161 5148
rect 10652 5108 10658 5120
rect 11149 5117 11161 5120
rect 11195 5117 11207 5151
rect 11149 5111 11207 5117
rect 12894 5108 12900 5160
rect 12952 5148 12958 5160
rect 13173 5151 13231 5157
rect 13173 5148 13185 5151
rect 12952 5120 13185 5148
rect 12952 5108 12958 5120
rect 13173 5117 13185 5120
rect 13219 5148 13231 5151
rect 13446 5148 13452 5160
rect 13219 5120 13452 5148
rect 13219 5117 13231 5120
rect 13173 5111 13231 5117
rect 13446 5108 13452 5120
rect 13504 5108 13510 5160
rect 18233 5151 18291 5157
rect 18233 5117 18245 5151
rect 18279 5148 18291 5151
rect 19352 5148 19380 5179
rect 22554 5176 22560 5188
rect 22612 5176 22618 5228
rect 24118 5216 24124 5228
rect 24079 5188 24124 5216
rect 24118 5176 24124 5188
rect 24176 5176 24182 5228
rect 24210 5176 24216 5228
rect 24268 5216 24274 5228
rect 24268 5188 24313 5216
rect 24268 5176 24274 5188
rect 25590 5176 25596 5228
rect 25648 5216 25654 5228
rect 27816 5225 27844 5256
rect 31573 5287 31631 5293
rect 31573 5253 31585 5287
rect 31619 5284 31631 5287
rect 31619 5256 32352 5284
rect 31619 5253 31631 5256
rect 31573 5247 31631 5253
rect 32324 5228 32352 5256
rect 25777 5219 25835 5225
rect 25777 5216 25789 5219
rect 25648 5188 25789 5216
rect 25648 5176 25654 5188
rect 25777 5185 25789 5188
rect 25823 5185 25835 5219
rect 25777 5179 25835 5185
rect 27801 5219 27859 5225
rect 27801 5185 27813 5219
rect 27847 5185 27859 5219
rect 27801 5179 27859 5185
rect 27890 5176 27896 5228
rect 27948 5216 27954 5228
rect 27948 5188 27993 5216
rect 27948 5176 27954 5188
rect 31754 5176 31760 5228
rect 31812 5216 31818 5228
rect 32122 5216 32128 5228
rect 31812 5188 32128 5216
rect 31812 5176 31818 5188
rect 32122 5176 32128 5188
rect 32180 5176 32186 5228
rect 32306 5216 32312 5228
rect 32267 5188 32312 5216
rect 32306 5176 32312 5188
rect 32364 5176 32370 5228
rect 20898 5148 20904 5160
rect 18279 5120 18920 5148
rect 19352 5120 20904 5148
rect 18279 5117 18291 5120
rect 18233 5111 18291 5117
rect 10505 5083 10563 5089
rect 10505 5049 10517 5083
rect 10551 5080 10563 5083
rect 10870 5080 10876 5092
rect 10551 5052 10876 5080
rect 10551 5049 10563 5052
rect 10505 5043 10563 5049
rect 10870 5040 10876 5052
rect 10928 5040 10934 5092
rect 16761 5083 16819 5089
rect 16761 5049 16773 5083
rect 16807 5080 16819 5083
rect 16942 5080 16948 5092
rect 16807 5052 16948 5080
rect 16807 5049 16819 5052
rect 16761 5043 16819 5049
rect 16942 5040 16948 5052
rect 17000 5040 17006 5092
rect 18892 5024 18920 5120
rect 20898 5108 20904 5120
rect 20956 5148 20962 5160
rect 21269 5151 21327 5157
rect 21269 5148 21281 5151
rect 20956 5120 21281 5148
rect 20956 5108 20962 5120
rect 21269 5117 21281 5120
rect 21315 5117 21327 5151
rect 21269 5111 21327 5117
rect 22373 5151 22431 5157
rect 22373 5117 22385 5151
rect 22419 5148 22431 5151
rect 22830 5148 22836 5160
rect 22419 5120 22836 5148
rect 22419 5117 22431 5120
rect 22373 5111 22431 5117
rect 22830 5108 22836 5120
rect 22888 5148 22894 5160
rect 23382 5148 23388 5160
rect 22888 5120 23388 5148
rect 22888 5108 22894 5120
rect 23382 5108 23388 5120
rect 23440 5108 23446 5160
rect 25038 5108 25044 5160
rect 25096 5148 25102 5160
rect 25685 5151 25743 5157
rect 25685 5148 25697 5151
rect 25096 5120 25697 5148
rect 25096 5108 25102 5120
rect 25685 5117 25697 5120
rect 25731 5117 25743 5151
rect 26878 5148 26884 5160
rect 26791 5120 26884 5148
rect 25685 5111 25743 5117
rect 26878 5108 26884 5120
rect 26936 5148 26942 5160
rect 27709 5151 27767 5157
rect 27709 5148 27721 5151
rect 26936 5120 27721 5148
rect 26936 5108 26942 5120
rect 27709 5117 27721 5120
rect 27755 5148 27767 5151
rect 28994 5148 29000 5160
rect 27755 5120 29000 5148
rect 27755 5117 27767 5120
rect 27709 5111 27767 5117
rect 28994 5108 29000 5120
rect 29052 5108 29058 5160
rect 29270 5148 29276 5160
rect 29231 5120 29276 5148
rect 29270 5108 29276 5120
rect 29328 5148 29334 5160
rect 29825 5151 29883 5157
rect 29825 5148 29837 5151
rect 29328 5120 29837 5148
rect 29328 5108 29334 5120
rect 29825 5117 29837 5120
rect 29871 5117 29883 5151
rect 30377 5151 30435 5157
rect 30377 5148 30389 5151
rect 29825 5111 29883 5117
rect 30208 5120 30389 5148
rect 19604 5083 19662 5089
rect 19604 5049 19616 5083
rect 19650 5080 19662 5083
rect 19886 5080 19892 5092
rect 19650 5052 19892 5080
rect 19650 5049 19662 5052
rect 19604 5043 19662 5049
rect 19886 5040 19892 5052
rect 19944 5080 19950 5092
rect 20622 5080 20628 5092
rect 19944 5052 20628 5080
rect 19944 5040 19950 5052
rect 20622 5040 20628 5052
rect 20680 5040 20686 5092
rect 24765 5083 24823 5089
rect 24765 5049 24777 5083
rect 24811 5080 24823 5083
rect 25593 5083 25651 5089
rect 25593 5080 25605 5083
rect 24811 5052 25605 5080
rect 24811 5049 24823 5052
rect 24765 5043 24823 5049
rect 25593 5049 25605 5052
rect 25639 5080 25651 5083
rect 25774 5080 25780 5092
rect 25639 5052 25780 5080
rect 25639 5049 25651 5052
rect 25593 5043 25651 5049
rect 25774 5040 25780 5052
rect 25832 5040 25838 5092
rect 30208 5024 30236 5120
rect 30377 5117 30389 5120
rect 30423 5117 30435 5151
rect 32030 5148 32036 5160
rect 31991 5120 32036 5148
rect 30377 5111 30435 5117
rect 32030 5108 32036 5120
rect 32088 5108 32094 5160
rect 2133 5015 2191 5021
rect 2133 4981 2145 5015
rect 2179 5012 2191 5015
rect 2406 5012 2412 5024
rect 2179 4984 2412 5012
rect 2179 4981 2191 4984
rect 2133 4975 2191 4981
rect 2406 4972 2412 4984
rect 2464 4972 2470 5024
rect 2590 5012 2596 5024
rect 2551 4984 2596 5012
rect 2590 4972 2596 4984
rect 2648 4972 2654 5024
rect 2682 4972 2688 5024
rect 2740 5012 2746 5024
rect 3881 5015 3939 5021
rect 3881 5012 3893 5015
rect 2740 4984 3893 5012
rect 2740 4972 2746 4984
rect 3881 4981 3893 4984
rect 3927 4981 3939 5015
rect 3881 4975 3939 4981
rect 4614 4972 4620 5024
rect 4672 5012 4678 5024
rect 4985 5015 5043 5021
rect 4985 5012 4997 5015
rect 4672 4984 4997 5012
rect 4672 4972 4678 4984
rect 4985 4981 4997 4984
rect 5031 4981 5043 5015
rect 4985 4975 5043 4981
rect 6825 5015 6883 5021
rect 6825 4981 6837 5015
rect 6871 5012 6883 5015
rect 7926 5012 7932 5024
rect 6871 4984 7932 5012
rect 6871 4981 6883 4984
rect 6825 4975 6883 4981
rect 7926 4972 7932 4984
rect 7984 4972 7990 5024
rect 8110 5012 8116 5024
rect 8071 4984 8116 5012
rect 8110 4972 8116 4984
rect 8168 4972 8174 5024
rect 8386 4972 8392 5024
rect 8444 5012 8450 5024
rect 8573 5015 8631 5021
rect 8573 5012 8585 5015
rect 8444 4984 8585 5012
rect 8444 4972 8450 4984
rect 8573 4981 8585 4984
rect 8619 4981 8631 5015
rect 9030 5012 9036 5024
rect 8991 4984 9036 5012
rect 8573 4975 8631 4981
rect 9030 4972 9036 4984
rect 9088 4972 9094 5024
rect 9306 5012 9312 5024
rect 9267 4984 9312 5012
rect 9306 4972 9312 4984
rect 9364 4972 9370 5024
rect 9490 4972 9496 5024
rect 9548 5012 9554 5024
rect 9677 5015 9735 5021
rect 9677 5012 9689 5015
rect 9548 4984 9689 5012
rect 9548 4972 9554 4984
rect 9677 4981 9689 4984
rect 9723 4981 9735 5015
rect 10778 5012 10784 5024
rect 10739 4984 10784 5012
rect 9677 4975 9735 4981
rect 10778 4972 10784 4984
rect 10836 4972 10842 5024
rect 12710 4972 12716 5024
rect 12768 5012 12774 5024
rect 13081 5015 13139 5021
rect 13081 5012 13093 5015
rect 12768 4984 13093 5012
rect 12768 4972 12774 4984
rect 13081 4981 13093 4984
rect 13127 5012 13139 5015
rect 13635 5015 13693 5021
rect 13635 5012 13647 5015
rect 13127 4984 13647 5012
rect 13127 4981 13139 4984
rect 13081 4975 13139 4981
rect 13635 4981 13647 4984
rect 13681 5012 13693 5015
rect 14274 5012 14280 5024
rect 13681 4984 14280 5012
rect 13681 4981 13693 4984
rect 13635 4975 13693 4981
rect 14274 4972 14280 4984
rect 14332 4972 14338 5024
rect 16390 5012 16396 5024
rect 16351 4984 16396 5012
rect 16390 4972 16396 4984
rect 16448 4972 16454 5024
rect 16574 4972 16580 5024
rect 16632 5012 16638 5024
rect 16853 5015 16911 5021
rect 16853 5012 16865 5015
rect 16632 4984 16865 5012
rect 16632 4972 16638 4984
rect 16853 4981 16865 4984
rect 16899 4981 16911 5015
rect 17770 5012 17776 5024
rect 17731 4984 17776 5012
rect 16853 4975 16911 4981
rect 17770 4972 17776 4984
rect 17828 4972 17834 5024
rect 18874 5012 18880 5024
rect 18835 4984 18880 5012
rect 18874 4972 18880 4984
rect 18932 4972 18938 5024
rect 22465 5015 22523 5021
rect 22465 4981 22477 5015
rect 22511 5012 22523 5015
rect 23106 5012 23112 5024
rect 22511 4984 23112 5012
rect 22511 4981 22523 4984
rect 22465 4975 22523 4981
rect 23106 4972 23112 4984
rect 23164 4972 23170 5024
rect 24026 5012 24032 5024
rect 23987 4984 24032 5012
rect 24026 4972 24032 4984
rect 24084 4972 24090 5024
rect 28074 4972 28080 5024
rect 28132 5012 28138 5024
rect 28445 5015 28503 5021
rect 28445 5012 28457 5015
rect 28132 4984 28457 5012
rect 28132 4972 28138 4984
rect 28445 4981 28457 4984
rect 28491 5012 28503 5015
rect 29270 5012 29276 5024
rect 28491 4984 29276 5012
rect 28491 4981 28503 4984
rect 28445 4975 28503 4981
rect 29270 4972 29276 4984
rect 29328 4972 29334 5024
rect 29454 5012 29460 5024
rect 29415 4984 29460 5012
rect 29454 4972 29460 4984
rect 29512 4972 29518 5024
rect 30190 5012 30196 5024
rect 30151 4984 30196 5012
rect 30190 4972 30196 4984
rect 30248 4972 30254 5024
rect 30558 5012 30564 5024
rect 30519 4984 30564 5012
rect 30558 4972 30564 4984
rect 30616 4972 30622 5024
rect 30834 4972 30840 5024
rect 30892 5012 30898 5024
rect 30929 5015 30987 5021
rect 30929 5012 30941 5015
rect 30892 4984 30941 5012
rect 30892 4972 30898 4984
rect 30929 4981 30941 4984
rect 30975 4981 30987 5015
rect 30929 4975 30987 4981
rect 31662 4972 31668 5024
rect 31720 5012 31726 5024
rect 32766 5012 32772 5024
rect 31720 4984 32772 5012
rect 31720 4972 31726 4984
rect 32766 4972 32772 4984
rect 32824 4972 32830 5024
rect 33229 5015 33287 5021
rect 33229 4981 33241 5015
rect 33275 5012 33287 5015
rect 34514 5012 34520 5024
rect 33275 4984 34520 5012
rect 33275 4981 33287 4984
rect 33229 4975 33287 4981
rect 34514 4972 34520 4984
rect 34572 4972 34578 5024
rect 1104 4922 38824 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 38824 4922
rect 1104 4848 38824 4870
rect 3326 4808 3332 4820
rect 3287 4780 3332 4808
rect 3326 4768 3332 4780
rect 3384 4768 3390 4820
rect 5810 4768 5816 4820
rect 5868 4808 5874 4820
rect 6365 4811 6423 4817
rect 6365 4808 6377 4811
rect 5868 4780 6377 4808
rect 5868 4768 5874 4780
rect 6365 4777 6377 4780
rect 6411 4808 6423 4811
rect 6730 4808 6736 4820
rect 6411 4780 6736 4808
rect 6411 4777 6423 4780
rect 6365 4771 6423 4777
rect 6730 4768 6736 4780
rect 6788 4768 6794 4820
rect 7282 4768 7288 4820
rect 7340 4808 7346 4820
rect 7469 4811 7527 4817
rect 7469 4808 7481 4811
rect 7340 4780 7481 4808
rect 7340 4768 7346 4780
rect 7469 4777 7481 4780
rect 7515 4777 7527 4811
rect 8018 4808 8024 4820
rect 7979 4780 8024 4808
rect 7469 4771 7527 4777
rect 8018 4768 8024 4780
rect 8076 4768 8082 4820
rect 9490 4808 9496 4820
rect 9451 4780 9496 4808
rect 9490 4768 9496 4780
rect 9548 4768 9554 4820
rect 10137 4811 10195 4817
rect 10137 4777 10149 4811
rect 10183 4808 10195 4811
rect 10226 4808 10232 4820
rect 10183 4780 10232 4808
rect 10183 4777 10195 4780
rect 10137 4771 10195 4777
rect 10226 4768 10232 4780
rect 10284 4808 10290 4820
rect 10778 4808 10784 4820
rect 10284 4780 10784 4808
rect 10284 4768 10290 4780
rect 10778 4768 10784 4780
rect 10836 4768 10842 4820
rect 11514 4808 11520 4820
rect 11475 4780 11520 4808
rect 11514 4768 11520 4780
rect 11572 4768 11578 4820
rect 13998 4808 14004 4820
rect 13959 4780 14004 4808
rect 13998 4768 14004 4780
rect 14056 4768 14062 4820
rect 14737 4811 14795 4817
rect 14737 4777 14749 4811
rect 14783 4808 14795 4811
rect 15286 4808 15292 4820
rect 14783 4780 15292 4808
rect 14783 4777 14795 4780
rect 14737 4771 14795 4777
rect 15286 4768 15292 4780
rect 15344 4808 15350 4820
rect 15749 4811 15807 4817
rect 15749 4808 15761 4811
rect 15344 4780 15761 4808
rect 15344 4768 15350 4780
rect 15749 4777 15761 4780
rect 15795 4777 15807 4811
rect 15749 4771 15807 4777
rect 16853 4811 16911 4817
rect 16853 4777 16865 4811
rect 16899 4808 16911 4811
rect 16942 4808 16948 4820
rect 16899 4780 16948 4808
rect 16899 4777 16911 4780
rect 16853 4771 16911 4777
rect 16942 4768 16948 4780
rect 17000 4768 17006 4820
rect 17218 4808 17224 4820
rect 17179 4780 17224 4808
rect 17218 4768 17224 4780
rect 17276 4768 17282 4820
rect 19334 4768 19340 4820
rect 19392 4808 19398 4820
rect 19797 4811 19855 4817
rect 19797 4808 19809 4811
rect 19392 4780 19809 4808
rect 19392 4768 19398 4780
rect 19797 4777 19809 4780
rect 19843 4777 19855 4811
rect 19797 4771 19855 4777
rect 20349 4811 20407 4817
rect 20349 4777 20361 4811
rect 20395 4808 20407 4811
rect 20438 4808 20444 4820
rect 20395 4780 20444 4808
rect 20395 4777 20407 4780
rect 20349 4771 20407 4777
rect 1664 4743 1722 4749
rect 1664 4709 1676 4743
rect 1710 4740 1722 4743
rect 3344 4740 3372 4768
rect 1710 4712 3372 4740
rect 4709 4743 4767 4749
rect 1710 4709 1722 4712
rect 1664 4703 1722 4709
rect 4709 4709 4721 4743
rect 4755 4740 4767 4743
rect 4798 4740 4804 4752
rect 4755 4712 4804 4740
rect 4755 4709 4767 4712
rect 4709 4703 4767 4709
rect 4798 4700 4804 4712
rect 4856 4700 4862 4752
rect 7926 4740 7932 4752
rect 7839 4712 7932 4740
rect 7926 4700 7932 4712
rect 7984 4740 7990 4752
rect 7984 4712 8524 4740
rect 7984 4700 7990 4712
rect 8496 4684 8524 4712
rect 11698 4700 11704 4752
rect 11756 4740 11762 4752
rect 12066 4740 12072 4752
rect 11756 4712 12072 4740
rect 11756 4700 11762 4712
rect 12066 4700 12072 4712
rect 12124 4740 12130 4752
rect 12222 4743 12280 4749
rect 12222 4740 12234 4743
rect 12124 4712 12234 4740
rect 12124 4700 12130 4712
rect 12222 4709 12234 4712
rect 12268 4709 12280 4743
rect 12222 4703 12280 4709
rect 16485 4743 16543 4749
rect 16485 4709 16497 4743
rect 16531 4740 16543 4743
rect 16574 4740 16580 4752
rect 16531 4712 16580 4740
rect 16531 4709 16543 4712
rect 16485 4703 16543 4709
rect 16574 4700 16580 4712
rect 16632 4740 16638 4752
rect 17770 4740 17776 4752
rect 16632 4712 17776 4740
rect 16632 4700 16638 4712
rect 17770 4700 17776 4712
rect 17828 4700 17834 4752
rect 19426 4700 19432 4752
rect 19484 4740 19490 4752
rect 19521 4743 19579 4749
rect 19521 4740 19533 4743
rect 19484 4712 19533 4740
rect 19484 4700 19490 4712
rect 19521 4709 19533 4712
rect 19567 4709 19579 4743
rect 19521 4703 19579 4709
rect 19610 4700 19616 4752
rect 19668 4740 19674 4752
rect 20364 4740 20392 4771
rect 20438 4768 20444 4780
rect 20496 4768 20502 4820
rect 21818 4808 21824 4820
rect 21779 4780 21824 4808
rect 21818 4768 21824 4780
rect 21876 4768 21882 4820
rect 24210 4768 24216 4820
rect 24268 4808 24274 4820
rect 25317 4811 25375 4817
rect 25317 4808 25329 4811
rect 24268 4780 25329 4808
rect 24268 4768 24274 4780
rect 25317 4777 25329 4780
rect 25363 4808 25375 4811
rect 25685 4811 25743 4817
rect 25685 4808 25697 4811
rect 25363 4780 25697 4808
rect 25363 4777 25375 4780
rect 25317 4771 25375 4777
rect 25685 4777 25697 4780
rect 25731 4777 25743 4811
rect 27154 4808 27160 4820
rect 27115 4780 27160 4808
rect 25685 4771 25743 4777
rect 27154 4768 27160 4780
rect 27212 4768 27218 4820
rect 30282 4768 30288 4820
rect 30340 4808 30346 4820
rect 30653 4811 30711 4817
rect 30653 4808 30665 4811
rect 30340 4780 30665 4808
rect 30340 4768 30346 4780
rect 30653 4777 30665 4780
rect 30699 4777 30711 4811
rect 32122 4808 32128 4820
rect 32083 4780 32128 4808
rect 30653 4771 30711 4777
rect 32122 4768 32128 4780
rect 32180 4768 32186 4820
rect 32766 4768 32772 4820
rect 32824 4808 32830 4820
rect 33597 4811 33655 4817
rect 33597 4808 33609 4811
rect 32824 4780 33609 4808
rect 32824 4768 32830 4780
rect 33597 4777 33609 4780
rect 33643 4808 33655 4811
rect 34238 4808 34244 4820
rect 33643 4780 34244 4808
rect 33643 4777 33655 4780
rect 33597 4771 33655 4777
rect 34238 4768 34244 4780
rect 34296 4768 34302 4820
rect 34606 4768 34612 4820
rect 34664 4808 34670 4820
rect 35345 4811 35403 4817
rect 35345 4808 35357 4811
rect 34664 4780 35357 4808
rect 34664 4768 34670 4780
rect 35345 4777 35357 4780
rect 35391 4777 35403 4811
rect 35345 4771 35403 4777
rect 19668 4712 20392 4740
rect 19668 4700 19674 4712
rect 23290 4700 23296 4752
rect 23348 4740 23354 4752
rect 23658 4749 23664 4752
rect 23652 4740 23664 4749
rect 23348 4712 23664 4740
rect 23348 4700 23354 4712
rect 23652 4703 23664 4712
rect 23658 4700 23664 4703
rect 23716 4700 23722 4752
rect 31757 4743 31815 4749
rect 31757 4709 31769 4743
rect 31803 4740 31815 4743
rect 32030 4740 32036 4752
rect 31803 4712 32036 4740
rect 31803 4709 31815 4712
rect 31757 4703 31815 4709
rect 32030 4700 32036 4712
rect 32088 4700 32094 4752
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4672 1455 4675
rect 1486 4672 1492 4684
rect 1443 4644 1492 4672
rect 1443 4641 1455 4644
rect 1397 4635 1455 4641
rect 1486 4632 1492 4644
rect 1544 4632 1550 4684
rect 4617 4675 4675 4681
rect 4617 4641 4629 4675
rect 4663 4672 4675 4675
rect 5166 4672 5172 4684
rect 4663 4644 5172 4672
rect 4663 4641 4675 4644
rect 4617 4635 4675 4641
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 5813 4675 5871 4681
rect 5813 4641 5825 4675
rect 5859 4672 5871 4675
rect 6178 4672 6184 4684
rect 5859 4644 6184 4672
rect 5859 4641 5871 4644
rect 5813 4635 5871 4641
rect 6178 4632 6184 4644
rect 6236 4632 6242 4684
rect 6822 4672 6828 4684
rect 6783 4644 6828 4672
rect 6822 4632 6828 4644
rect 6880 4632 6886 4684
rect 6917 4675 6975 4681
rect 6917 4641 6929 4675
rect 6963 4672 6975 4675
rect 7006 4672 7012 4684
rect 6963 4644 7012 4672
rect 6963 4641 6975 4644
rect 6917 4635 6975 4641
rect 7006 4632 7012 4644
rect 7064 4632 7070 4684
rect 8389 4675 8447 4681
rect 8389 4641 8401 4675
rect 8435 4641 8447 4675
rect 8389 4635 8447 4641
rect 4801 4607 4859 4613
rect 4801 4604 4813 4607
rect 3804 4576 4813 4604
rect 2774 4468 2780 4480
rect 2735 4440 2780 4468
rect 2774 4428 2780 4440
rect 2832 4428 2838 4480
rect 3050 4428 3056 4480
rect 3108 4468 3114 4480
rect 3804 4477 3832 4576
rect 4801 4573 4813 4576
rect 4847 4573 4859 4607
rect 8404 4604 8432 4635
rect 8478 4632 8484 4684
rect 8536 4672 8542 4684
rect 10045 4675 10103 4681
rect 8536 4644 8581 4672
rect 8536 4632 8542 4644
rect 10045 4641 10057 4675
rect 10091 4672 10103 4675
rect 10594 4672 10600 4684
rect 10091 4644 10600 4672
rect 10091 4641 10103 4644
rect 10045 4635 10103 4641
rect 10594 4632 10600 4644
rect 10652 4632 10658 4684
rect 11974 4672 11980 4684
rect 11935 4644 11980 4672
rect 11974 4632 11980 4644
rect 12032 4632 12038 4684
rect 15654 4672 15660 4684
rect 15615 4644 15660 4672
rect 15654 4632 15660 4644
rect 15712 4632 15718 4684
rect 16850 4632 16856 4684
rect 16908 4672 16914 4684
rect 17586 4681 17592 4684
rect 17569 4675 17592 4681
rect 17569 4672 17581 4675
rect 16908 4644 17581 4672
rect 16908 4632 16914 4644
rect 17569 4641 17581 4644
rect 17644 4672 17650 4684
rect 22186 4672 22192 4684
rect 17644 4644 17717 4672
rect 22147 4644 22192 4672
rect 17569 4635 17592 4641
rect 17586 4632 17592 4635
rect 17644 4632 17650 4644
rect 22186 4632 22192 4644
rect 22244 4632 22250 4684
rect 27798 4672 27804 4684
rect 27759 4644 27804 4672
rect 27798 4632 27804 4644
rect 27856 4632 27862 4684
rect 27893 4675 27951 4681
rect 27893 4641 27905 4675
rect 27939 4672 27951 4675
rect 28350 4672 28356 4684
rect 27939 4644 28356 4672
rect 27939 4641 27951 4644
rect 27893 4635 27951 4641
rect 28350 4632 28356 4644
rect 28408 4632 28414 4684
rect 29362 4632 29368 4684
rect 29420 4672 29426 4684
rect 29529 4675 29587 4681
rect 29529 4672 29541 4675
rect 29420 4644 29541 4672
rect 29420 4632 29426 4644
rect 29529 4641 29541 4644
rect 29575 4641 29587 4675
rect 32490 4672 32496 4684
rect 32451 4644 32496 4672
rect 29529 4635 29587 4641
rect 32490 4632 32496 4644
rect 32548 4632 32554 4684
rect 32585 4675 32643 4681
rect 32585 4641 32597 4675
rect 32631 4672 32643 4675
rect 33042 4672 33048 4684
rect 32631 4644 33048 4672
rect 32631 4641 32643 4644
rect 32585 4635 32643 4641
rect 8665 4607 8723 4613
rect 8404 4576 8524 4604
rect 4801 4567 4859 4573
rect 8496 4548 8524 4576
rect 8665 4573 8677 4607
rect 8711 4604 8723 4607
rect 9490 4604 9496 4616
rect 8711 4576 9496 4604
rect 8711 4573 8723 4576
rect 8665 4567 8723 4573
rect 9490 4564 9496 4576
rect 9548 4564 9554 4616
rect 9950 4564 9956 4616
rect 10008 4604 10014 4616
rect 10229 4607 10287 4613
rect 10229 4604 10241 4607
rect 10008 4576 10241 4604
rect 10008 4564 10014 4576
rect 10229 4573 10241 4576
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 14090 4564 14096 4616
rect 14148 4604 14154 4616
rect 14369 4607 14427 4613
rect 14369 4604 14381 4607
rect 14148 4576 14381 4604
rect 14148 4564 14154 4576
rect 14369 4573 14381 4576
rect 14415 4604 14427 4607
rect 15838 4604 15844 4616
rect 14415 4576 15844 4604
rect 14415 4573 14427 4576
rect 14369 4567 14427 4573
rect 15838 4564 15844 4576
rect 15896 4564 15902 4616
rect 17310 4604 17316 4616
rect 17271 4576 17316 4604
rect 17310 4564 17316 4576
rect 17368 4564 17374 4616
rect 22278 4604 22284 4616
rect 22239 4576 22284 4604
rect 22278 4564 22284 4576
rect 22336 4564 22342 4616
rect 22373 4607 22431 4613
rect 22373 4573 22385 4607
rect 22419 4604 22431 4607
rect 22554 4604 22560 4616
rect 22419 4576 22560 4604
rect 22419 4573 22431 4576
rect 22373 4567 22431 4573
rect 5994 4536 6000 4548
rect 5955 4508 6000 4536
rect 5994 4496 6000 4508
rect 6052 4496 6058 4548
rect 8478 4496 8484 4548
rect 8536 4496 8542 4548
rect 15194 4496 15200 4548
rect 15252 4536 15258 4548
rect 15289 4539 15347 4545
rect 15289 4536 15301 4539
rect 15252 4508 15301 4536
rect 15252 4496 15258 4508
rect 15289 4505 15301 4508
rect 15335 4505 15347 4539
rect 22388 4536 22416 4567
rect 22554 4564 22560 4576
rect 22612 4564 22618 4616
rect 23198 4564 23204 4616
rect 23256 4604 23262 4616
rect 23385 4607 23443 4613
rect 23385 4604 23397 4607
rect 23256 4576 23397 4604
rect 23256 4564 23262 4576
rect 23385 4573 23397 4576
rect 23431 4573 23443 4607
rect 23385 4567 23443 4573
rect 27982 4564 27988 4616
rect 28040 4604 28046 4616
rect 29270 4604 29276 4616
rect 28040 4576 28085 4604
rect 29231 4576 29276 4604
rect 28040 4564 28046 4576
rect 29270 4564 29276 4576
rect 29328 4564 29334 4616
rect 15289 4499 15347 4505
rect 21652 4508 22416 4536
rect 22925 4539 22983 4545
rect 3789 4471 3847 4477
rect 3789 4468 3801 4471
rect 3108 4440 3801 4468
rect 3108 4428 3114 4440
rect 3789 4437 3801 4440
rect 3835 4437 3847 4471
rect 3789 4431 3847 4437
rect 4249 4471 4307 4477
rect 4249 4437 4261 4471
rect 4295 4468 4307 4471
rect 5261 4471 5319 4477
rect 5261 4468 5273 4471
rect 4295 4440 5273 4468
rect 4295 4437 4307 4440
rect 4249 4431 4307 4437
rect 5261 4437 5273 4440
rect 5307 4468 5319 4471
rect 5534 4468 5540 4480
rect 5307 4440 5540 4468
rect 5307 4437 5319 4440
rect 5261 4431 5319 4437
rect 5534 4428 5540 4440
rect 5592 4428 5598 4480
rect 5626 4428 5632 4480
rect 5684 4468 5690 4480
rect 7098 4468 7104 4480
rect 5684 4440 5729 4468
rect 7059 4440 7104 4468
rect 5684 4428 5690 4440
rect 7098 4428 7104 4440
rect 7156 4428 7162 4480
rect 7558 4428 7564 4480
rect 7616 4468 7622 4480
rect 9122 4468 9128 4480
rect 7616 4440 9128 4468
rect 7616 4428 7622 4440
rect 9122 4428 9128 4440
rect 9180 4428 9186 4480
rect 9677 4471 9735 4477
rect 9677 4437 9689 4471
rect 9723 4468 9735 4471
rect 10318 4468 10324 4480
rect 9723 4440 10324 4468
rect 9723 4437 9735 4440
rect 9677 4431 9735 4437
rect 10318 4428 10324 4440
rect 10376 4428 10382 4480
rect 11885 4471 11943 4477
rect 11885 4437 11897 4471
rect 11931 4468 11943 4471
rect 12342 4468 12348 4480
rect 11931 4440 12348 4468
rect 11931 4437 11943 4440
rect 11885 4431 11943 4437
rect 12342 4428 12348 4440
rect 12400 4468 12406 4480
rect 13357 4471 13415 4477
rect 13357 4468 13369 4471
rect 12400 4440 13369 4468
rect 12400 4428 12406 4440
rect 13357 4437 13369 4440
rect 13403 4468 13415 4471
rect 13630 4468 13636 4480
rect 13403 4440 13636 4468
rect 13403 4437 13415 4440
rect 13357 4431 13415 4437
rect 13630 4428 13636 4440
rect 13688 4428 13694 4480
rect 13814 4428 13820 4480
rect 13872 4468 13878 4480
rect 15013 4471 15071 4477
rect 15013 4468 15025 4471
rect 13872 4440 15025 4468
rect 13872 4428 13878 4440
rect 15013 4437 15025 4440
rect 15059 4468 15071 4471
rect 15470 4468 15476 4480
rect 15059 4440 15476 4468
rect 15059 4437 15071 4440
rect 15013 4431 15071 4437
rect 15470 4428 15476 4440
rect 15528 4428 15534 4480
rect 18693 4471 18751 4477
rect 18693 4437 18705 4471
rect 18739 4468 18751 4471
rect 19150 4468 19156 4480
rect 18739 4440 19156 4468
rect 18739 4437 18751 4440
rect 18693 4431 18751 4437
rect 19150 4428 19156 4440
rect 19208 4428 19214 4480
rect 21266 4468 21272 4480
rect 21227 4440 21272 4468
rect 21266 4428 21272 4440
rect 21324 4468 21330 4480
rect 21652 4477 21680 4508
rect 22925 4505 22937 4539
rect 22971 4536 22983 4539
rect 23106 4536 23112 4548
rect 22971 4508 23112 4536
rect 22971 4505 22983 4508
rect 22925 4499 22983 4505
rect 23106 4496 23112 4508
rect 23164 4536 23170 4548
rect 23164 4508 23428 4536
rect 23164 4496 23170 4508
rect 21637 4471 21695 4477
rect 21637 4468 21649 4471
rect 21324 4440 21649 4468
rect 21324 4428 21330 4440
rect 21637 4437 21649 4440
rect 21683 4437 21695 4471
rect 23198 4468 23204 4480
rect 23159 4440 23204 4468
rect 21637 4431 21695 4437
rect 23198 4428 23204 4440
rect 23256 4428 23262 4480
rect 23400 4468 23428 4508
rect 25590 4496 25596 4548
rect 25648 4536 25654 4548
rect 26145 4539 26203 4545
rect 26145 4536 26157 4539
rect 25648 4508 26157 4536
rect 25648 4496 25654 4508
rect 26145 4505 26157 4508
rect 26191 4505 26203 4539
rect 26145 4499 26203 4505
rect 27614 4496 27620 4548
rect 27672 4536 27678 4548
rect 28813 4539 28871 4545
rect 28813 4536 28825 4539
rect 27672 4508 28825 4536
rect 27672 4496 27678 4508
rect 28813 4505 28825 4508
rect 28859 4505 28871 4539
rect 28813 4499 28871 4505
rect 24762 4468 24768 4480
rect 23400 4440 24768 4468
rect 24762 4428 24768 4440
rect 24820 4428 24826 4480
rect 26694 4468 26700 4480
rect 26655 4440 26700 4468
rect 26694 4428 26700 4440
rect 26752 4428 26758 4480
rect 27433 4471 27491 4477
rect 27433 4437 27445 4471
rect 27479 4468 27491 4471
rect 27522 4468 27528 4480
rect 27479 4440 27528 4468
rect 27479 4437 27491 4440
rect 27433 4431 27491 4437
rect 27522 4428 27528 4440
rect 27580 4428 27586 4480
rect 28442 4468 28448 4480
rect 28403 4440 28448 4468
rect 28442 4428 28448 4440
rect 28500 4428 28506 4480
rect 30374 4428 30380 4480
rect 30432 4468 30438 4480
rect 31205 4471 31263 4477
rect 31205 4468 31217 4471
rect 30432 4440 31217 4468
rect 30432 4428 30438 4440
rect 31205 4437 31217 4440
rect 31251 4468 31263 4471
rect 32600 4468 32628 4635
rect 33042 4632 33048 4644
rect 33100 4632 33106 4684
rect 34238 4681 34244 4684
rect 33229 4675 33287 4681
rect 33229 4641 33241 4675
rect 33275 4672 33287 4675
rect 34232 4672 34244 4681
rect 33275 4644 34244 4672
rect 33275 4641 33287 4644
rect 33229 4635 33287 4641
rect 34232 4635 34244 4644
rect 32769 4607 32827 4613
rect 32769 4573 32781 4607
rect 32815 4604 32827 4607
rect 33244 4604 33272 4635
rect 34238 4632 34244 4635
rect 34296 4632 34302 4684
rect 33962 4604 33968 4616
rect 32815 4576 33272 4604
rect 33923 4576 33968 4604
rect 32815 4573 32827 4576
rect 32769 4567 32827 4573
rect 33962 4564 33968 4576
rect 34020 4564 34026 4616
rect 31251 4440 32628 4468
rect 31251 4437 31263 4440
rect 31205 4431 31263 4437
rect 1104 4378 38824 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 34966 4378
rect 35018 4326 35030 4378
rect 35082 4326 35094 4378
rect 35146 4326 35158 4378
rect 35210 4326 38824 4378
rect 1104 4304 38824 4326
rect 2777 4267 2835 4273
rect 2777 4233 2789 4267
rect 2823 4264 2835 4267
rect 3326 4264 3332 4276
rect 2823 4236 3332 4264
rect 2823 4233 2835 4236
rect 2777 4227 2835 4233
rect 3326 4224 3332 4236
rect 3384 4224 3390 4276
rect 6178 4264 6184 4276
rect 6139 4236 6184 4264
rect 6178 4224 6184 4236
rect 6236 4224 6242 4276
rect 11974 4264 11980 4276
rect 11935 4236 11980 4264
rect 11974 4224 11980 4236
rect 12032 4224 12038 4276
rect 15746 4224 15752 4276
rect 15804 4264 15810 4276
rect 16209 4267 16267 4273
rect 16209 4264 16221 4267
rect 15804 4236 16221 4264
rect 15804 4224 15810 4236
rect 16209 4233 16221 4236
rect 16255 4233 16267 4267
rect 16209 4227 16267 4233
rect 4614 4196 4620 4208
rect 4080 4168 4620 4196
rect 2866 4088 2872 4140
rect 2924 4128 2930 4140
rect 4080 4128 4108 4168
rect 4614 4156 4620 4168
rect 4672 4156 4678 4208
rect 6730 4156 6736 4208
rect 6788 4156 6794 4208
rect 7558 4156 7564 4208
rect 7616 4156 7622 4208
rect 5534 4128 5540 4140
rect 2924 4100 4108 4128
rect 5495 4100 5540 4128
rect 2924 4088 2930 4100
rect 5534 4088 5540 4100
rect 5592 4088 5598 4140
rect 5629 4131 5687 4137
rect 5629 4097 5641 4131
rect 5675 4097 5687 4131
rect 6748 4128 6776 4156
rect 7469 4131 7527 4137
rect 6748 4100 7236 4128
rect 5629 4091 5687 4097
rect 1397 4063 1455 4069
rect 1397 4029 1409 4063
rect 1443 4060 1455 4063
rect 1486 4060 1492 4072
rect 1443 4032 1492 4060
rect 1443 4029 1455 4032
rect 1397 4023 1455 4029
rect 1486 4020 1492 4032
rect 1544 4020 1550 4072
rect 1664 4063 1722 4069
rect 1664 4029 1676 4063
rect 1710 4060 1722 4063
rect 2590 4060 2596 4072
rect 1710 4032 2596 4060
rect 1710 4029 1722 4032
rect 1664 4023 1722 4029
rect 2590 4020 2596 4032
rect 2648 4060 2654 4072
rect 3329 4063 3387 4069
rect 3329 4060 3341 4063
rect 2648 4032 3341 4060
rect 2648 4020 2654 4032
rect 3329 4029 3341 4032
rect 3375 4029 3387 4063
rect 3329 4023 3387 4029
rect 3881 4063 3939 4069
rect 3881 4029 3893 4063
rect 3927 4060 3939 4063
rect 3927 4032 4568 4060
rect 3927 4029 3939 4032
rect 3881 4023 3939 4029
rect 3786 3924 3792 3936
rect 3747 3896 3792 3924
rect 3786 3884 3792 3896
rect 3844 3884 3850 3936
rect 4062 3924 4068 3936
rect 4023 3896 4068 3924
rect 4062 3884 4068 3896
rect 4120 3884 4126 3936
rect 4540 3933 4568 4032
rect 4706 4020 4712 4072
rect 4764 4060 4770 4072
rect 5074 4060 5080 4072
rect 4764 4032 5080 4060
rect 4764 4020 4770 4032
rect 5074 4020 5080 4032
rect 5132 4060 5138 4072
rect 5644 4060 5672 4091
rect 5132 4032 5672 4060
rect 6641 4063 6699 4069
rect 5132 4020 5138 4032
rect 6641 4029 6653 4063
rect 6687 4060 6699 4063
rect 7098 4060 7104 4072
rect 6687 4032 7104 4060
rect 6687 4029 6699 4032
rect 6641 4023 6699 4029
rect 7098 4020 7104 4032
rect 7156 4020 7162 4072
rect 7208 4069 7236 4100
rect 7469 4097 7481 4131
rect 7515 4128 7527 4131
rect 7576 4128 7604 4156
rect 7515 4100 7604 4128
rect 7515 4097 7527 4100
rect 7469 4091 7527 4097
rect 7193 4063 7251 4069
rect 7193 4029 7205 4063
rect 7239 4029 7251 4063
rect 7193 4023 7251 4029
rect 8481 4063 8539 4069
rect 8481 4029 8493 4063
rect 8527 4060 8539 4063
rect 8573 4063 8631 4069
rect 8573 4060 8585 4063
rect 8527 4032 8585 4060
rect 8527 4029 8539 4032
rect 8481 4023 8539 4029
rect 8573 4029 8585 4032
rect 8619 4060 8631 4063
rect 9582 4060 9588 4072
rect 8619 4032 9588 4060
rect 8619 4029 8631 4032
rect 8573 4023 8631 4029
rect 9582 4020 9588 4032
rect 9640 4020 9646 4072
rect 11057 4063 11115 4069
rect 11057 4029 11069 4063
rect 11103 4060 11115 4063
rect 12434 4060 12440 4072
rect 11103 4032 11744 4060
rect 12395 4032 12440 4060
rect 11103 4029 11115 4032
rect 11057 4023 11115 4029
rect 5350 3992 5356 4004
rect 5092 3964 5356 3992
rect 4525 3927 4583 3933
rect 4525 3893 4537 3927
rect 4571 3924 4583 3927
rect 4614 3924 4620 3936
rect 4571 3896 4620 3924
rect 4571 3893 4583 3896
rect 4525 3887 4583 3893
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 4798 3924 4804 3936
rect 4759 3896 4804 3924
rect 4798 3884 4804 3896
rect 4856 3884 4862 3936
rect 5092 3933 5120 3964
rect 5350 3952 5356 3964
rect 5408 3952 5414 4004
rect 6914 3952 6920 4004
rect 6972 3992 6978 4004
rect 7285 3995 7343 4001
rect 7285 3992 7297 3995
rect 6972 3964 7297 3992
rect 6972 3952 6978 3964
rect 7285 3961 7297 3964
rect 7331 3961 7343 3995
rect 7285 3955 7343 3961
rect 8113 3995 8171 4001
rect 8113 3961 8125 3995
rect 8159 3992 8171 3995
rect 8294 3992 8300 4004
rect 8159 3964 8300 3992
rect 8159 3961 8171 3964
rect 8113 3955 8171 3961
rect 8294 3952 8300 3964
rect 8352 3992 8358 4004
rect 8818 3995 8876 4001
rect 8818 3992 8830 3995
rect 8352 3964 8830 3992
rect 8352 3952 8358 3964
rect 8818 3961 8830 3964
rect 8864 3961 8876 3995
rect 10873 3995 10931 4001
rect 10873 3992 10885 3995
rect 8818 3955 8876 3961
rect 9968 3964 10885 3992
rect 9968 3936 9996 3964
rect 10873 3961 10885 3964
rect 10919 3961 10931 3995
rect 10873 3955 10931 3961
rect 11716 3936 11744 4032
rect 12434 4020 12440 4032
rect 12492 4060 12498 4072
rect 14090 4069 14096 4072
rect 12989 4063 13047 4069
rect 12989 4060 13001 4063
rect 12492 4032 13001 4060
rect 12492 4020 12498 4032
rect 12989 4029 13001 4032
rect 13035 4029 13047 4063
rect 12989 4023 13047 4029
rect 13817 4063 13875 4069
rect 13817 4029 13829 4063
rect 13863 4029 13875 4063
rect 14084 4060 14096 4069
rect 14051 4032 14096 4060
rect 13817 4023 13875 4029
rect 14084 4023 14096 4032
rect 11974 3952 11980 4004
rect 12032 3992 12038 4004
rect 13633 3995 13691 4001
rect 13633 3992 13645 3995
rect 12032 3964 13645 3992
rect 12032 3952 12038 3964
rect 13633 3961 13645 3964
rect 13679 3992 13691 3995
rect 13832 3992 13860 4023
rect 14090 4020 14096 4023
rect 14148 4020 14154 4072
rect 16224 4060 16252 4227
rect 17310 4224 17316 4276
rect 17368 4264 17374 4276
rect 17405 4267 17463 4273
rect 17405 4264 17417 4267
rect 17368 4236 17417 4264
rect 17368 4224 17374 4236
rect 17405 4233 17417 4236
rect 17451 4233 17463 4267
rect 17405 4227 17463 4233
rect 17586 4224 17592 4276
rect 17644 4264 17650 4276
rect 17773 4267 17831 4273
rect 17773 4264 17785 4267
rect 17644 4236 17785 4264
rect 17644 4224 17650 4236
rect 17773 4233 17785 4236
rect 17819 4233 17831 4267
rect 18598 4264 18604 4276
rect 18559 4236 18604 4264
rect 17773 4227 17831 4233
rect 18598 4224 18604 4236
rect 18656 4224 18662 4276
rect 19978 4224 19984 4276
rect 20036 4264 20042 4276
rect 20162 4264 20168 4276
rect 20036 4236 20168 4264
rect 20036 4224 20042 4236
rect 20162 4224 20168 4236
rect 20220 4224 20226 4276
rect 22186 4224 22192 4276
rect 22244 4264 22250 4276
rect 22373 4267 22431 4273
rect 22373 4264 22385 4267
rect 22244 4236 22385 4264
rect 22244 4224 22250 4236
rect 22373 4233 22385 4236
rect 22419 4233 22431 4267
rect 22373 4227 22431 4233
rect 23198 4224 23204 4276
rect 23256 4264 23262 4276
rect 23385 4267 23443 4273
rect 23385 4264 23397 4267
rect 23256 4236 23397 4264
rect 23256 4224 23262 4236
rect 23385 4233 23397 4236
rect 23431 4233 23443 4267
rect 23385 4227 23443 4233
rect 26145 4267 26203 4273
rect 26145 4233 26157 4267
rect 26191 4264 26203 4267
rect 26694 4264 26700 4276
rect 26191 4236 26700 4264
rect 26191 4233 26203 4236
rect 26145 4227 26203 4233
rect 26694 4224 26700 4236
rect 26752 4224 26758 4276
rect 27525 4267 27583 4273
rect 27525 4233 27537 4267
rect 27571 4264 27583 4267
rect 27798 4264 27804 4276
rect 27571 4236 27804 4264
rect 27571 4233 27583 4236
rect 27525 4227 27583 4233
rect 27798 4224 27804 4236
rect 27856 4264 27862 4276
rect 27893 4267 27951 4273
rect 27893 4264 27905 4267
rect 27856 4236 27905 4264
rect 27856 4224 27862 4236
rect 27893 4233 27905 4236
rect 27939 4233 27951 4267
rect 27893 4227 27951 4233
rect 17218 4196 17224 4208
rect 17052 4168 17224 4196
rect 17052 4137 17080 4168
rect 17218 4156 17224 4168
rect 17276 4156 17282 4208
rect 22278 4196 22284 4208
rect 22112 4168 22284 4196
rect 17037 4131 17095 4137
rect 17037 4097 17049 4131
rect 17083 4097 17095 4131
rect 17037 4091 17095 4097
rect 17402 4088 17408 4140
rect 17460 4128 17466 4140
rect 18325 4131 18383 4137
rect 18325 4128 18337 4131
rect 17460 4100 18337 4128
rect 17460 4088 17466 4100
rect 18325 4097 18337 4100
rect 18371 4128 18383 4131
rect 18371 4100 19196 4128
rect 18371 4097 18383 4100
rect 18325 4091 18383 4097
rect 16761 4063 16819 4069
rect 16761 4060 16773 4063
rect 16224 4032 16773 4060
rect 16761 4029 16773 4032
rect 16807 4029 16819 4063
rect 16761 4023 16819 4029
rect 18417 4063 18475 4069
rect 18417 4029 18429 4063
rect 18463 4060 18475 4063
rect 19168 4060 19196 4100
rect 19426 4088 19432 4140
rect 19484 4128 19490 4140
rect 19981 4131 20039 4137
rect 19981 4128 19993 4131
rect 19484 4100 19993 4128
rect 19484 4088 19490 4100
rect 19981 4097 19993 4100
rect 20027 4128 20039 4131
rect 20622 4128 20628 4140
rect 20027 4100 20628 4128
rect 20027 4097 20039 4100
rect 19981 4091 20039 4097
rect 20622 4088 20628 4100
rect 20680 4088 20686 4140
rect 22005 4131 22063 4137
rect 22005 4097 22017 4131
rect 22051 4128 22063 4131
rect 22112 4128 22140 4168
rect 22278 4156 22284 4168
rect 22336 4196 22342 4208
rect 25590 4196 25596 4208
rect 22336 4168 23428 4196
rect 25551 4168 25596 4196
rect 22336 4156 22342 4168
rect 22051 4100 22140 4128
rect 23400 4128 23428 4168
rect 25590 4156 25596 4168
rect 25648 4196 25654 4208
rect 25648 4168 26740 4196
rect 25648 4156 25654 4168
rect 23566 4128 23572 4140
rect 23400 4100 23572 4128
rect 22051 4097 22063 4100
rect 22005 4091 22063 4097
rect 23566 4088 23572 4100
rect 23624 4088 23630 4140
rect 26712 4137 26740 4168
rect 26970 4156 26976 4208
rect 27028 4196 27034 4208
rect 28442 4196 28448 4208
rect 27028 4168 28448 4196
rect 27028 4156 27034 4168
rect 26697 4131 26755 4137
rect 26697 4097 26709 4131
rect 26743 4097 26755 4131
rect 26697 4091 26755 4097
rect 19521 4063 19579 4069
rect 19521 4060 19533 4063
rect 18463 4032 19104 4060
rect 19168 4032 19533 4060
rect 18463 4029 18475 4032
rect 18417 4023 18475 4029
rect 13679 3964 13860 3992
rect 16853 3995 16911 4001
rect 13679 3961 13691 3964
rect 13633 3955 13691 3961
rect 16853 3961 16865 3995
rect 16899 3992 16911 3995
rect 16942 3992 16948 4004
rect 16899 3964 16948 3992
rect 16899 3961 16911 3964
rect 16853 3955 16911 3961
rect 16942 3952 16948 3964
rect 17000 3952 17006 4004
rect 19076 3936 19104 4032
rect 19521 4029 19533 4032
rect 19567 4060 19579 4063
rect 19610 4060 19616 4072
rect 19567 4032 19616 4060
rect 19567 4029 19579 4032
rect 19521 4023 19579 4029
rect 19610 4020 19616 4032
rect 19668 4020 19674 4072
rect 20162 4020 20168 4072
rect 20220 4060 20226 4072
rect 20257 4063 20315 4069
rect 20257 4060 20269 4063
rect 20220 4032 20269 4060
rect 20220 4020 20226 4032
rect 20257 4029 20269 4032
rect 20303 4029 20315 4063
rect 20257 4023 20315 4029
rect 22465 4063 22523 4069
rect 22465 4029 22477 4063
rect 22511 4060 22523 4063
rect 22511 4032 23152 4060
rect 22511 4029 22523 4032
rect 22465 4023 22523 4029
rect 23124 3936 23152 4032
rect 23198 4020 23204 4072
rect 23256 4060 23262 4072
rect 23661 4063 23719 4069
rect 23661 4060 23673 4063
rect 23256 4032 23673 4060
rect 23256 4020 23262 4032
rect 23661 4029 23673 4032
rect 23707 4029 23719 4063
rect 23661 4023 23719 4029
rect 23928 4063 23986 4069
rect 23928 4029 23940 4063
rect 23974 4060 23986 4063
rect 24762 4060 24768 4072
rect 23974 4032 24768 4060
rect 23974 4029 23986 4032
rect 23928 4023 23986 4029
rect 24762 4020 24768 4032
rect 24820 4020 24826 4072
rect 26513 4063 26571 4069
rect 26513 4029 26525 4063
rect 26559 4060 26571 4063
rect 26602 4060 26608 4072
rect 26559 4032 26608 4060
rect 26559 4029 26571 4032
rect 26513 4023 26571 4029
rect 26602 4020 26608 4032
rect 26660 4020 26666 4072
rect 27724 4069 27752 4168
rect 28442 4156 28448 4168
rect 28500 4156 28506 4208
rect 29089 4131 29147 4137
rect 29089 4097 29101 4131
rect 29135 4128 29147 4131
rect 29270 4128 29276 4140
rect 29135 4100 29276 4128
rect 29135 4097 29147 4100
rect 29089 4091 29147 4097
rect 29270 4088 29276 4100
rect 29328 4128 29334 4140
rect 29638 4128 29644 4140
rect 29328 4100 29644 4128
rect 29328 4088 29334 4100
rect 29638 4088 29644 4100
rect 29696 4088 29702 4140
rect 30101 4131 30159 4137
rect 30101 4097 30113 4131
rect 30147 4128 30159 4131
rect 30282 4128 30288 4140
rect 30147 4100 30288 4128
rect 30147 4097 30159 4100
rect 30101 4091 30159 4097
rect 30282 4088 30288 4100
rect 30340 4088 30346 4140
rect 31202 4088 31208 4140
rect 31260 4128 31266 4140
rect 31481 4131 31539 4137
rect 31481 4128 31493 4131
rect 31260 4100 31493 4128
rect 31260 4088 31266 4100
rect 31481 4097 31493 4100
rect 31527 4097 31539 4131
rect 31481 4091 31539 4097
rect 33042 4088 33048 4140
rect 33100 4128 33106 4140
rect 33413 4131 33471 4137
rect 33413 4128 33425 4131
rect 33100 4100 33425 4128
rect 33100 4088 33106 4100
rect 33413 4097 33425 4100
rect 33459 4097 33471 4131
rect 33413 4091 33471 4097
rect 27709 4063 27767 4069
rect 27709 4029 27721 4063
rect 27755 4029 27767 4063
rect 27709 4023 27767 4029
rect 28258 4020 28264 4072
rect 28316 4060 28322 4072
rect 29825 4063 29883 4069
rect 29825 4060 29837 4063
rect 28316 4032 29837 4060
rect 28316 4020 28322 4032
rect 29825 4029 29837 4032
rect 29871 4060 29883 4063
rect 30374 4060 30380 4072
rect 29871 4032 30380 4060
rect 29871 4029 29883 4032
rect 29825 4023 29883 4029
rect 30374 4020 30380 4032
rect 30432 4020 30438 4072
rect 31021 4063 31079 4069
rect 31021 4029 31033 4063
rect 31067 4060 31079 4063
rect 31110 4060 31116 4072
rect 31067 4032 31116 4060
rect 31067 4029 31079 4032
rect 31021 4023 31079 4029
rect 31110 4020 31116 4032
rect 31168 4060 31174 4072
rect 31662 4060 31668 4072
rect 31168 4032 31668 4060
rect 31168 4020 31174 4032
rect 31662 4020 31668 4032
rect 31720 4020 31726 4072
rect 31757 4063 31815 4069
rect 31757 4029 31769 4063
rect 31803 4060 31815 4063
rect 32490 4060 32496 4072
rect 31803 4032 32496 4060
rect 31803 4029 31815 4032
rect 31757 4023 31815 4029
rect 32490 4020 32496 4032
rect 32548 4020 32554 4072
rect 26053 3995 26111 4001
rect 26053 3961 26065 3995
rect 26099 3992 26111 3995
rect 28721 3995 28779 4001
rect 26099 3964 26648 3992
rect 26099 3961 26111 3964
rect 26053 3955 26111 3961
rect 5077 3927 5135 3933
rect 5077 3893 5089 3927
rect 5123 3893 5135 3927
rect 5077 3887 5135 3893
rect 5445 3927 5503 3933
rect 5445 3893 5457 3927
rect 5491 3924 5503 3927
rect 5534 3924 5540 3936
rect 5491 3896 5540 3924
rect 5491 3893 5503 3896
rect 5445 3887 5503 3893
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 6822 3924 6828 3936
rect 6783 3896 6828 3924
rect 6822 3884 6828 3896
rect 6880 3884 6886 3936
rect 9950 3924 9956 3936
rect 9911 3896 9956 3924
rect 9950 3884 9956 3896
rect 10008 3884 10014 3936
rect 10594 3924 10600 3936
rect 10555 3896 10600 3924
rect 10594 3884 10600 3896
rect 10652 3884 10658 3936
rect 11238 3924 11244 3936
rect 11199 3896 11244 3924
rect 11238 3884 11244 3896
rect 11296 3884 11302 3936
rect 11698 3924 11704 3936
rect 11659 3896 11704 3924
rect 11698 3884 11704 3896
rect 11756 3884 11762 3936
rect 12621 3927 12679 3933
rect 12621 3893 12633 3927
rect 12667 3924 12679 3927
rect 12710 3924 12716 3936
rect 12667 3896 12716 3924
rect 12667 3893 12679 3896
rect 12621 3887 12679 3893
rect 12710 3884 12716 3896
rect 12768 3884 12774 3936
rect 14366 3884 14372 3936
rect 14424 3924 14430 3936
rect 14918 3924 14924 3936
rect 14424 3896 14924 3924
rect 14424 3884 14430 3896
rect 14918 3884 14924 3896
rect 14976 3924 14982 3936
rect 15197 3927 15255 3933
rect 15197 3924 15209 3927
rect 14976 3896 15209 3924
rect 14976 3884 14982 3896
rect 15197 3893 15209 3896
rect 15243 3893 15255 3927
rect 15197 3887 15255 3893
rect 15654 3884 15660 3936
rect 15712 3924 15718 3936
rect 15749 3927 15807 3933
rect 15749 3924 15761 3927
rect 15712 3896 15761 3924
rect 15712 3884 15718 3896
rect 15749 3893 15761 3896
rect 15795 3893 15807 3927
rect 15749 3887 15807 3893
rect 16393 3927 16451 3933
rect 16393 3893 16405 3927
rect 16439 3924 16451 3927
rect 16482 3924 16488 3936
rect 16439 3896 16488 3924
rect 16439 3893 16451 3896
rect 16393 3887 16451 3893
rect 16482 3884 16488 3896
rect 16540 3884 16546 3936
rect 19058 3924 19064 3936
rect 19019 3896 19064 3924
rect 19058 3884 19064 3896
rect 19116 3884 19122 3936
rect 19426 3924 19432 3936
rect 19339 3896 19432 3924
rect 19426 3884 19432 3896
rect 19484 3924 19490 3936
rect 19978 3924 19984 3936
rect 19484 3896 19984 3924
rect 19484 3884 19490 3896
rect 19978 3884 19984 3896
rect 20036 3924 20042 3936
rect 21358 3924 21364 3936
rect 20036 3896 20081 3924
rect 21319 3896 21364 3924
rect 20036 3884 20042 3896
rect 21358 3884 21364 3896
rect 21416 3884 21422 3936
rect 22646 3924 22652 3936
rect 22607 3896 22652 3924
rect 22646 3884 22652 3896
rect 22704 3884 22710 3936
rect 23106 3924 23112 3936
rect 23067 3896 23112 3924
rect 23106 3884 23112 3896
rect 23164 3884 23170 3936
rect 25038 3924 25044 3936
rect 24999 3896 25044 3924
rect 25038 3884 25044 3896
rect 25096 3884 25102 3936
rect 26620 3933 26648 3964
rect 28721 3961 28733 3995
rect 28767 3992 28779 3995
rect 28767 3964 29960 3992
rect 28767 3961 28779 3964
rect 28721 3955 28779 3961
rect 29932 3936 29960 3964
rect 26605 3927 26663 3933
rect 26605 3893 26617 3927
rect 26651 3924 26663 3927
rect 26694 3924 26700 3936
rect 26651 3896 26700 3924
rect 26651 3893 26663 3896
rect 26605 3887 26663 3893
rect 26694 3884 26700 3896
rect 26752 3884 26758 3936
rect 28350 3924 28356 3936
rect 28311 3896 28356 3924
rect 28350 3884 28356 3896
rect 28408 3884 28414 3936
rect 29457 3927 29515 3933
rect 29457 3893 29469 3927
rect 29503 3924 29515 3927
rect 29730 3924 29736 3936
rect 29503 3896 29736 3924
rect 29503 3893 29515 3896
rect 29457 3887 29515 3893
rect 29730 3884 29736 3896
rect 29788 3884 29794 3936
rect 29914 3884 29920 3936
rect 29972 3924 29978 3936
rect 30466 3924 30472 3936
rect 29972 3896 30017 3924
rect 30427 3896 30472 3924
rect 29972 3884 29978 3896
rect 30466 3884 30472 3896
rect 30524 3884 30530 3936
rect 30929 3927 30987 3933
rect 30929 3893 30941 3927
rect 30975 3924 30987 3927
rect 31018 3924 31024 3936
rect 30975 3896 31024 3924
rect 30975 3893 30987 3896
rect 30929 3887 30987 3893
rect 31018 3884 31024 3896
rect 31076 3924 31082 3936
rect 31483 3927 31541 3933
rect 31483 3924 31495 3927
rect 31076 3896 31495 3924
rect 31076 3884 31082 3896
rect 31483 3893 31495 3896
rect 31529 3893 31541 3927
rect 31483 3887 31541 3893
rect 32030 3884 32036 3936
rect 32088 3924 32094 3936
rect 32861 3927 32919 3933
rect 32861 3924 32873 3927
rect 32088 3896 32873 3924
rect 32088 3884 32094 3896
rect 32861 3893 32873 3896
rect 32907 3893 32919 3927
rect 32861 3887 32919 3893
rect 33594 3884 33600 3936
rect 33652 3924 33658 3936
rect 33962 3924 33968 3936
rect 33652 3896 33968 3924
rect 33652 3884 33658 3896
rect 33962 3884 33968 3896
rect 34020 3884 34026 3936
rect 34238 3884 34244 3936
rect 34296 3924 34302 3936
rect 34425 3927 34483 3933
rect 34425 3924 34437 3927
rect 34296 3896 34437 3924
rect 34296 3884 34302 3896
rect 34425 3893 34437 3896
rect 34471 3924 34483 3927
rect 34606 3924 34612 3936
rect 34471 3896 34612 3924
rect 34471 3893 34483 3896
rect 34425 3887 34483 3893
rect 34606 3884 34612 3896
rect 34664 3884 34670 3936
rect 1104 3834 38824 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 38824 3834
rect 1104 3760 38824 3782
rect 2406 3680 2412 3732
rect 2464 3720 2470 3732
rect 3789 3723 3847 3729
rect 3789 3720 3801 3723
rect 2464 3692 3801 3720
rect 2464 3680 2470 3692
rect 3789 3689 3801 3692
rect 3835 3720 3847 3723
rect 4525 3723 4583 3729
rect 4525 3720 4537 3723
rect 3835 3692 4537 3720
rect 3835 3689 3847 3692
rect 3789 3683 3847 3689
rect 4525 3689 4537 3692
rect 4571 3689 4583 3723
rect 4525 3683 4583 3689
rect 8478 3680 8484 3732
rect 8536 3720 8542 3732
rect 9033 3723 9091 3729
rect 9033 3720 9045 3723
rect 8536 3692 9045 3720
rect 8536 3680 8542 3692
rect 9033 3689 9045 3692
rect 9079 3689 9091 3723
rect 9490 3720 9496 3732
rect 9451 3692 9496 3720
rect 9033 3683 9091 3689
rect 9490 3680 9496 3692
rect 9548 3680 9554 3732
rect 9674 3720 9680 3732
rect 9635 3692 9680 3720
rect 9674 3680 9680 3692
rect 9732 3680 9738 3732
rect 10226 3720 10232 3732
rect 10187 3692 10232 3720
rect 10226 3680 10232 3692
rect 10284 3680 10290 3732
rect 12066 3720 12072 3732
rect 12027 3692 12072 3720
rect 12066 3680 12072 3692
rect 12124 3720 12130 3732
rect 12621 3723 12679 3729
rect 12621 3720 12633 3723
rect 12124 3692 12633 3720
rect 12124 3680 12130 3692
rect 12621 3689 12633 3692
rect 12667 3689 12679 3723
rect 13170 3720 13176 3732
rect 13131 3692 13176 3720
rect 12621 3683 12679 3689
rect 13170 3680 13176 3692
rect 13228 3680 13234 3732
rect 13541 3723 13599 3729
rect 13541 3689 13553 3723
rect 13587 3720 13599 3723
rect 13722 3720 13728 3732
rect 13587 3692 13728 3720
rect 13587 3689 13599 3692
rect 13541 3683 13599 3689
rect 13722 3680 13728 3692
rect 13780 3680 13786 3732
rect 14550 3720 14556 3732
rect 14511 3692 14556 3720
rect 14550 3680 14556 3692
rect 14608 3680 14614 3732
rect 14918 3720 14924 3732
rect 14879 3692 14924 3720
rect 14918 3680 14924 3692
rect 14976 3680 14982 3732
rect 15565 3723 15623 3729
rect 15565 3689 15577 3723
rect 15611 3720 15623 3723
rect 15838 3720 15844 3732
rect 15611 3692 15844 3720
rect 15611 3689 15623 3692
rect 15565 3683 15623 3689
rect 15838 3680 15844 3692
rect 15896 3680 15902 3732
rect 16206 3720 16212 3732
rect 16167 3692 16212 3720
rect 16206 3680 16212 3692
rect 16264 3680 16270 3732
rect 16301 3723 16359 3729
rect 16301 3689 16313 3723
rect 16347 3720 16359 3723
rect 16390 3720 16396 3732
rect 16347 3692 16396 3720
rect 16347 3689 16359 3692
rect 16301 3683 16359 3689
rect 16390 3680 16396 3692
rect 16448 3720 16454 3732
rect 17221 3723 17279 3729
rect 17221 3720 17233 3723
rect 16448 3692 17233 3720
rect 16448 3680 16454 3692
rect 17221 3689 17233 3692
rect 17267 3689 17279 3723
rect 17221 3683 17279 3689
rect 17770 3680 17776 3732
rect 17828 3720 17834 3732
rect 19245 3723 19303 3729
rect 19245 3720 19257 3723
rect 17828 3692 19257 3720
rect 17828 3680 17834 3692
rect 19245 3689 19257 3692
rect 19291 3720 19303 3723
rect 19797 3723 19855 3729
rect 19797 3720 19809 3723
rect 19291 3692 19809 3720
rect 19291 3689 19303 3692
rect 19245 3683 19303 3689
rect 19797 3689 19809 3692
rect 19843 3720 19855 3723
rect 20162 3720 20168 3732
rect 19843 3692 20168 3720
rect 19843 3689 19855 3692
rect 19797 3683 19855 3689
rect 20162 3680 20168 3692
rect 20220 3680 20226 3732
rect 20622 3720 20628 3732
rect 20583 3692 20628 3720
rect 20622 3680 20628 3692
rect 20680 3720 20686 3732
rect 21269 3723 21327 3729
rect 21269 3720 21281 3723
rect 20680 3692 21281 3720
rect 20680 3680 20686 3692
rect 21269 3689 21281 3692
rect 21315 3689 21327 3723
rect 21269 3683 21327 3689
rect 23201 3723 23259 3729
rect 23201 3689 23213 3723
rect 23247 3720 23259 3723
rect 23290 3720 23296 3732
rect 23247 3692 23296 3720
rect 23247 3689 23259 3692
rect 23201 3683 23259 3689
rect 23290 3680 23296 3692
rect 23348 3680 23354 3732
rect 26237 3723 26295 3729
rect 26237 3689 26249 3723
rect 26283 3720 26295 3723
rect 26602 3720 26608 3732
rect 26283 3692 26608 3720
rect 26283 3689 26295 3692
rect 26237 3683 26295 3689
rect 26602 3680 26608 3692
rect 26660 3680 26666 3732
rect 27985 3723 28043 3729
rect 27985 3689 27997 3723
rect 28031 3720 28043 3723
rect 28258 3720 28264 3732
rect 28031 3692 28264 3720
rect 28031 3689 28043 3692
rect 27985 3683 28043 3689
rect 28258 3680 28264 3692
rect 28316 3680 28322 3732
rect 28353 3723 28411 3729
rect 28353 3689 28365 3723
rect 28399 3720 28411 3723
rect 28626 3720 28632 3732
rect 28399 3692 28632 3720
rect 28399 3689 28411 3692
rect 28353 3683 28411 3689
rect 28626 3680 28632 3692
rect 28684 3720 28690 3732
rect 28902 3720 28908 3732
rect 28684 3692 28908 3720
rect 28684 3680 28690 3692
rect 28902 3680 28908 3692
rect 28960 3680 28966 3732
rect 29362 3720 29368 3732
rect 29323 3692 29368 3720
rect 29362 3680 29368 3692
rect 29420 3680 29426 3732
rect 30558 3680 30564 3732
rect 30616 3720 30622 3732
rect 31481 3723 31539 3729
rect 31481 3720 31493 3723
rect 30616 3692 31493 3720
rect 30616 3680 30622 3692
rect 31481 3689 31493 3692
rect 31527 3720 31539 3723
rect 31570 3720 31576 3732
rect 31527 3692 31576 3720
rect 31527 3689 31539 3692
rect 31481 3683 31539 3689
rect 31570 3680 31576 3692
rect 31628 3680 31634 3732
rect 31941 3723 31999 3729
rect 31941 3689 31953 3723
rect 31987 3720 31999 3723
rect 32030 3720 32036 3732
rect 31987 3692 32036 3720
rect 31987 3689 31999 3692
rect 31941 3683 31999 3689
rect 32030 3680 32036 3692
rect 32088 3680 32094 3732
rect 32306 3720 32312 3732
rect 32267 3692 32312 3720
rect 32306 3680 32312 3692
rect 32364 3680 32370 3732
rect 32490 3680 32496 3732
rect 32548 3720 32554 3732
rect 32677 3723 32735 3729
rect 32677 3720 32689 3723
rect 32548 3692 32689 3720
rect 32548 3680 32554 3692
rect 32677 3689 32689 3692
rect 32723 3689 32735 3723
rect 34606 3720 34612 3732
rect 34567 3692 34612 3720
rect 32677 3683 32735 3689
rect 34606 3680 34612 3692
rect 34664 3680 34670 3732
rect 1756 3655 1814 3661
rect 1756 3621 1768 3655
rect 1802 3652 1814 3655
rect 2774 3652 2780 3664
rect 1802 3624 2780 3652
rect 1802 3621 1814 3624
rect 1756 3615 1814 3621
rect 2774 3612 2780 3624
rect 2832 3612 2838 3664
rect 8202 3612 8208 3664
rect 8260 3652 8266 3664
rect 9508 3652 9536 3680
rect 8260 3624 9536 3652
rect 8260 3612 8266 3624
rect 9950 3612 9956 3664
rect 10008 3652 10014 3664
rect 10505 3655 10563 3661
rect 10505 3652 10517 3655
rect 10008 3624 10517 3652
rect 10008 3612 10014 3624
rect 10505 3621 10517 3624
rect 10551 3621 10563 3655
rect 11974 3652 11980 3664
rect 10505 3615 10563 3621
rect 10704 3624 11980 3652
rect 1486 3584 1492 3596
rect 1447 3556 1492 3584
rect 1486 3544 1492 3556
rect 1544 3544 1550 3596
rect 4430 3584 4436 3596
rect 4391 3556 4436 3584
rect 4430 3544 4436 3556
rect 4488 3584 4494 3596
rect 5445 3587 5503 3593
rect 5445 3584 5457 3587
rect 4488 3556 5457 3584
rect 4488 3544 4494 3556
rect 5445 3553 5457 3556
rect 5491 3553 5503 3587
rect 5445 3547 5503 3553
rect 5626 3544 5632 3596
rect 5684 3584 5690 3596
rect 5905 3587 5963 3593
rect 5905 3584 5917 3587
rect 5684 3556 5917 3584
rect 5684 3544 5690 3556
rect 5905 3553 5917 3556
rect 5951 3584 5963 3587
rect 6264 3587 6322 3593
rect 6264 3584 6276 3587
rect 5951 3556 6276 3584
rect 5951 3553 5963 3556
rect 5905 3547 5963 3553
rect 6264 3553 6276 3556
rect 6310 3584 6322 3587
rect 6822 3584 6828 3596
rect 6310 3556 6828 3584
rect 6310 3553 6322 3556
rect 6264 3547 6322 3553
rect 6822 3544 6828 3556
rect 6880 3544 6886 3596
rect 8481 3587 8539 3593
rect 8481 3553 8493 3587
rect 8527 3584 8539 3587
rect 8938 3584 8944 3596
rect 8527 3556 8944 3584
rect 8527 3553 8539 3556
rect 8481 3547 8539 3553
rect 8938 3544 8944 3556
rect 8996 3544 9002 3596
rect 9490 3544 9496 3596
rect 9548 3584 9554 3596
rect 10704 3593 10732 3624
rect 11974 3612 11980 3624
rect 12032 3612 12038 3664
rect 12710 3612 12716 3664
rect 12768 3652 12774 3664
rect 14277 3655 14335 3661
rect 14277 3652 14289 3655
rect 12768 3624 14289 3652
rect 12768 3612 12774 3624
rect 14277 3621 14289 3624
rect 14323 3652 14335 3655
rect 14458 3652 14464 3664
rect 14323 3624 14464 3652
rect 14323 3621 14335 3624
rect 14277 3615 14335 3621
rect 14458 3612 14464 3624
rect 14516 3652 14522 3664
rect 15102 3652 15108 3664
rect 14516 3624 15108 3652
rect 14516 3612 14522 3624
rect 15102 3612 15108 3624
rect 15160 3612 15166 3664
rect 16945 3655 17003 3661
rect 16945 3652 16957 3655
rect 16868 3624 16957 3652
rect 10689 3587 10747 3593
rect 10689 3584 10701 3587
rect 9548 3556 10701 3584
rect 9548 3544 9554 3556
rect 10689 3553 10701 3556
rect 10735 3553 10747 3587
rect 10689 3547 10747 3553
rect 10778 3544 10784 3596
rect 10836 3584 10842 3596
rect 10945 3587 11003 3593
rect 10945 3584 10957 3587
rect 10836 3556 10957 3584
rect 10836 3544 10842 3556
rect 10945 3553 10957 3556
rect 10991 3553 11003 3587
rect 10945 3547 11003 3553
rect 4706 3516 4712 3528
rect 4667 3488 4712 3516
rect 4706 3476 4712 3488
rect 4764 3476 4770 3528
rect 5994 3516 6000 3528
rect 5955 3488 6000 3516
rect 5994 3476 6000 3488
rect 6052 3476 6058 3528
rect 13633 3519 13691 3525
rect 13633 3516 13645 3519
rect 13004 3488 13645 3516
rect 3970 3408 3976 3460
rect 4028 3448 4034 3460
rect 4065 3451 4123 3457
rect 4065 3448 4077 3451
rect 4028 3420 4077 3448
rect 4028 3408 4034 3420
rect 4065 3417 4077 3420
rect 4111 3417 4123 3451
rect 4065 3411 4123 3417
rect 2869 3383 2927 3389
rect 2869 3349 2881 3383
rect 2915 3380 2927 3383
rect 2958 3380 2964 3392
rect 2915 3352 2964 3380
rect 2915 3349 2927 3352
rect 2869 3343 2927 3349
rect 2958 3340 2964 3352
rect 3016 3380 3022 3392
rect 3421 3383 3479 3389
rect 3421 3380 3433 3383
rect 3016 3352 3433 3380
rect 3016 3340 3022 3352
rect 3421 3349 3433 3352
rect 3467 3349 3479 3383
rect 5166 3380 5172 3392
rect 5079 3352 5172 3380
rect 3421 3343 3479 3349
rect 5166 3340 5172 3352
rect 5224 3380 5230 3392
rect 5442 3380 5448 3392
rect 5224 3352 5448 3380
rect 5224 3340 5230 3352
rect 5442 3340 5448 3352
rect 5500 3340 5506 3392
rect 7190 3340 7196 3392
rect 7248 3380 7254 3392
rect 7377 3383 7435 3389
rect 7377 3380 7389 3383
rect 7248 3352 7389 3380
rect 7248 3340 7254 3352
rect 7377 3349 7389 3352
rect 7423 3380 7435 3383
rect 8021 3383 8079 3389
rect 8021 3380 8033 3383
rect 7423 3352 8033 3380
rect 7423 3349 7435 3352
rect 7377 3343 7435 3349
rect 8021 3349 8033 3352
rect 8067 3380 8079 3383
rect 8297 3383 8355 3389
rect 8297 3380 8309 3383
rect 8067 3352 8309 3380
rect 8067 3349 8079 3352
rect 8021 3343 8079 3349
rect 8297 3349 8309 3352
rect 8343 3349 8355 3383
rect 8662 3380 8668 3392
rect 8623 3352 8668 3380
rect 8297 3343 8355 3349
rect 8662 3340 8668 3352
rect 8720 3340 8726 3392
rect 10962 3340 10968 3392
rect 11020 3380 11026 3392
rect 13004 3389 13032 3488
rect 13633 3485 13645 3488
rect 13679 3485 13691 3519
rect 13633 3479 13691 3485
rect 13817 3519 13875 3525
rect 13817 3485 13829 3519
rect 13863 3516 13875 3519
rect 14366 3516 14372 3528
rect 13863 3488 14372 3516
rect 13863 3485 13875 3488
rect 13817 3479 13875 3485
rect 14366 3476 14372 3488
rect 14424 3476 14430 3528
rect 16485 3519 16543 3525
rect 16485 3485 16497 3519
rect 16531 3485 16543 3519
rect 16485 3479 16543 3485
rect 16500 3448 16528 3479
rect 16868 3448 16896 3624
rect 16945 3621 16957 3624
rect 16991 3652 17003 3655
rect 17310 3652 17316 3664
rect 16991 3624 17316 3652
rect 16991 3621 17003 3624
rect 16945 3615 17003 3621
rect 17310 3612 17316 3624
rect 17368 3612 17374 3664
rect 23474 3612 23480 3664
rect 23532 3661 23538 3664
rect 23532 3655 23596 3661
rect 23532 3621 23550 3655
rect 23584 3652 23596 3655
rect 25038 3652 25044 3664
rect 23584 3624 25044 3652
rect 23584 3621 23596 3624
rect 23532 3615 23596 3621
rect 23532 3612 23538 3615
rect 25038 3612 25044 3624
rect 25096 3652 25102 3664
rect 25225 3655 25283 3661
rect 25225 3652 25237 3655
rect 25096 3624 25237 3652
rect 25096 3612 25102 3624
rect 25225 3621 25237 3624
rect 25271 3621 25283 3655
rect 25225 3615 25283 3621
rect 29816 3655 29874 3661
rect 29816 3621 29828 3655
rect 29862 3652 29874 3655
rect 30282 3652 30288 3664
rect 29862 3624 30288 3652
rect 29862 3621 29874 3624
rect 29816 3615 29874 3621
rect 30282 3612 30288 3624
rect 30340 3612 30346 3664
rect 30466 3612 30472 3664
rect 30524 3652 30530 3664
rect 32508 3652 32536 3680
rect 33134 3652 33140 3664
rect 30524 3624 32536 3652
rect 33095 3624 33140 3652
rect 30524 3612 30530 3624
rect 33134 3612 33140 3624
rect 33192 3612 33198 3664
rect 17402 3584 17408 3596
rect 17363 3556 17408 3584
rect 17402 3544 17408 3556
rect 17460 3544 17466 3596
rect 17678 3544 17684 3596
rect 17736 3593 17742 3596
rect 17736 3587 17786 3593
rect 17736 3553 17740 3587
rect 17774 3553 17786 3587
rect 21358 3584 21364 3596
rect 21319 3556 21364 3584
rect 17736 3547 17786 3553
rect 17736 3544 17742 3547
rect 21358 3544 21364 3556
rect 21416 3544 21422 3596
rect 23198 3544 23204 3596
rect 23256 3584 23262 3596
rect 23293 3587 23351 3593
rect 23293 3584 23305 3587
rect 23256 3556 23305 3584
rect 23256 3544 23262 3556
rect 23293 3553 23305 3556
rect 23339 3553 23351 3587
rect 26510 3584 26516 3596
rect 26471 3556 26516 3584
rect 23293 3547 23351 3553
rect 26510 3544 26516 3556
rect 26568 3544 26574 3596
rect 26697 3587 26755 3593
rect 26697 3553 26709 3587
rect 26743 3584 26755 3587
rect 26878 3584 26884 3596
rect 26743 3556 26884 3584
rect 26743 3553 26755 3556
rect 26697 3547 26755 3553
rect 26878 3544 26884 3556
rect 26936 3584 26942 3596
rect 27157 3587 27215 3593
rect 27157 3584 27169 3587
rect 26936 3556 27169 3584
rect 26936 3544 26942 3556
rect 27157 3553 27169 3556
rect 27203 3553 27215 3587
rect 27157 3547 27215 3553
rect 27893 3587 27951 3593
rect 27893 3553 27905 3587
rect 27939 3584 27951 3587
rect 29549 3587 29607 3593
rect 27939 3556 28672 3584
rect 27939 3553 27951 3556
rect 27893 3547 27951 3553
rect 17862 3516 17868 3528
rect 17823 3488 17868 3516
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 18138 3516 18144 3528
rect 18099 3488 18144 3516
rect 18138 3476 18144 3488
rect 18196 3476 18202 3528
rect 21450 3476 21456 3528
rect 21508 3516 21514 3528
rect 22373 3519 22431 3525
rect 22373 3516 22385 3519
rect 21508 3488 22385 3516
rect 21508 3476 21514 3488
rect 22373 3485 22385 3488
rect 22419 3516 22431 3519
rect 22554 3516 22560 3528
rect 22419 3488 22560 3516
rect 22419 3485 22431 3488
rect 22373 3479 22431 3485
rect 22554 3476 22560 3488
rect 22612 3476 22618 3528
rect 27522 3476 27528 3528
rect 27580 3516 27586 3528
rect 28442 3516 28448 3528
rect 27580 3488 28448 3516
rect 27580 3476 27586 3488
rect 28442 3476 28448 3488
rect 28500 3476 28506 3528
rect 28644 3525 28672 3556
rect 29549 3553 29561 3587
rect 29595 3584 29607 3587
rect 29638 3584 29644 3596
rect 29595 3556 29644 3584
rect 29595 3553 29607 3556
rect 29549 3547 29607 3553
rect 29638 3544 29644 3556
rect 29696 3544 29702 3596
rect 31938 3544 31944 3596
rect 31996 3584 32002 3596
rect 32125 3587 32183 3593
rect 32125 3584 32137 3587
rect 31996 3556 32137 3584
rect 31996 3544 32002 3556
rect 32125 3553 32137 3556
rect 32171 3553 32183 3587
rect 32125 3547 32183 3553
rect 33496 3587 33554 3593
rect 33496 3553 33508 3587
rect 33542 3584 33554 3587
rect 34054 3584 34060 3596
rect 33542 3556 34060 3584
rect 33542 3553 33554 3556
rect 33496 3547 33554 3553
rect 34054 3544 34060 3556
rect 34112 3584 34118 3596
rect 35161 3587 35219 3593
rect 35161 3584 35173 3587
rect 34112 3556 35173 3584
rect 34112 3544 34118 3556
rect 35161 3553 35173 3556
rect 35207 3584 35219 3587
rect 35434 3584 35440 3596
rect 35207 3556 35440 3584
rect 35207 3553 35219 3556
rect 35161 3547 35219 3553
rect 35434 3544 35440 3556
rect 35492 3544 35498 3596
rect 28629 3519 28687 3525
rect 28629 3485 28641 3519
rect 28675 3516 28687 3519
rect 28718 3516 28724 3528
rect 28675 3488 28724 3516
rect 28675 3485 28687 3488
rect 28629 3479 28687 3485
rect 28718 3476 28724 3488
rect 28776 3516 28782 3528
rect 29362 3516 29368 3528
rect 28776 3488 29368 3516
rect 28776 3476 28782 3488
rect 29362 3476 29368 3488
rect 29420 3476 29426 3528
rect 33229 3519 33287 3525
rect 33229 3485 33241 3519
rect 33275 3485 33287 3519
rect 33229 3479 33287 3485
rect 16500 3420 16896 3448
rect 19978 3408 19984 3460
rect 20036 3448 20042 3460
rect 20257 3451 20315 3457
rect 20257 3448 20269 3451
rect 20036 3420 20269 3448
rect 20036 3408 20042 3420
rect 20257 3417 20269 3420
rect 20303 3448 20315 3451
rect 22005 3451 22063 3457
rect 22005 3448 22017 3451
rect 20303 3420 22017 3448
rect 20303 3417 20315 3420
rect 20257 3411 20315 3417
rect 22005 3417 22017 3420
rect 22051 3448 22063 3451
rect 22462 3448 22468 3460
rect 22051 3420 22468 3448
rect 22051 3417 22063 3420
rect 22005 3411 22063 3417
rect 22462 3408 22468 3420
rect 22520 3408 22526 3460
rect 26326 3408 26332 3460
rect 26384 3448 26390 3460
rect 26881 3451 26939 3457
rect 26881 3448 26893 3451
rect 26384 3420 26893 3448
rect 26384 3408 26390 3420
rect 26881 3417 26893 3420
rect 26927 3448 26939 3451
rect 27430 3448 27436 3460
rect 26927 3420 27436 3448
rect 26927 3417 26939 3420
rect 26881 3411 26939 3417
rect 27430 3408 27436 3420
rect 27488 3408 27494 3460
rect 12989 3383 13047 3389
rect 12989 3380 13001 3383
rect 11020 3352 13001 3380
rect 11020 3340 11026 3352
rect 12989 3349 13001 3352
rect 13035 3349 13047 3383
rect 15838 3380 15844 3392
rect 15799 3352 15844 3380
rect 12989 3343 13047 3349
rect 15838 3340 15844 3352
rect 15896 3340 15902 3392
rect 20898 3380 20904 3392
rect 20859 3352 20904 3380
rect 20898 3340 20904 3352
rect 20956 3340 20962 3392
rect 22646 3380 22652 3392
rect 22607 3352 22652 3380
rect 22646 3340 22652 3352
rect 22704 3340 22710 3392
rect 23566 3340 23572 3392
rect 23624 3380 23630 3392
rect 24673 3383 24731 3389
rect 24673 3380 24685 3383
rect 23624 3352 24685 3380
rect 23624 3340 23630 3352
rect 24673 3349 24685 3352
rect 24719 3380 24731 3383
rect 25593 3383 25651 3389
rect 25593 3380 25605 3383
rect 24719 3352 25605 3380
rect 24719 3349 24731 3352
rect 24673 3343 24731 3349
rect 25593 3349 25605 3352
rect 25639 3349 25651 3383
rect 25593 3343 25651 3349
rect 30190 3340 30196 3392
rect 30248 3380 30254 3392
rect 30926 3380 30932 3392
rect 30248 3352 30932 3380
rect 30248 3340 30254 3352
rect 30926 3340 30932 3352
rect 30984 3340 30990 3392
rect 33244 3380 33272 3479
rect 33594 3380 33600 3392
rect 33244 3352 33600 3380
rect 33594 3340 33600 3352
rect 33652 3340 33658 3392
rect 35342 3340 35348 3392
rect 35400 3380 35406 3392
rect 35529 3383 35587 3389
rect 35529 3380 35541 3383
rect 35400 3352 35541 3380
rect 35400 3340 35406 3352
rect 35529 3349 35541 3352
rect 35575 3349 35587 3383
rect 35529 3343 35587 3349
rect 1104 3290 38824 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 34966 3290
rect 35018 3238 35030 3290
rect 35082 3238 35094 3290
rect 35146 3238 35158 3290
rect 35210 3238 38824 3290
rect 1104 3216 38824 3238
rect 1486 3136 1492 3188
rect 1544 3176 1550 3188
rect 1581 3179 1639 3185
rect 1581 3176 1593 3179
rect 1544 3148 1593 3176
rect 1544 3136 1550 3148
rect 1581 3145 1593 3148
rect 1627 3145 1639 3179
rect 5626 3176 5632 3188
rect 1581 3139 1639 3145
rect 4172 3148 5488 3176
rect 5587 3148 5632 3176
rect 1596 3040 1624 3139
rect 4172 3120 4200 3148
rect 4154 3068 4160 3120
rect 4212 3068 4218 3120
rect 5460 3108 5488 3148
rect 5626 3136 5632 3148
rect 5684 3136 5690 3188
rect 8294 3176 8300 3188
rect 8255 3148 8300 3176
rect 8294 3136 8300 3148
rect 8352 3136 8358 3188
rect 10778 3176 10784 3188
rect 10739 3148 10784 3176
rect 10778 3136 10784 3148
rect 10836 3136 10842 3188
rect 11425 3179 11483 3185
rect 11425 3145 11437 3179
rect 11471 3176 11483 3179
rect 11974 3176 11980 3188
rect 11471 3148 11980 3176
rect 11471 3145 11483 3148
rect 11425 3139 11483 3145
rect 11974 3136 11980 3148
rect 12032 3136 12038 3188
rect 12618 3176 12624 3188
rect 12579 3148 12624 3176
rect 12618 3136 12624 3148
rect 12676 3136 12682 3188
rect 13449 3179 13507 3185
rect 13449 3145 13461 3179
rect 13495 3176 13507 3179
rect 13722 3176 13728 3188
rect 13495 3148 13728 3176
rect 13495 3145 13507 3148
rect 13449 3139 13507 3145
rect 13722 3136 13728 3148
rect 13780 3136 13786 3188
rect 15746 3176 15752 3188
rect 15707 3148 15752 3176
rect 15746 3136 15752 3148
rect 15804 3136 15810 3188
rect 16206 3136 16212 3188
rect 16264 3176 16270 3188
rect 16301 3179 16359 3185
rect 16301 3176 16313 3179
rect 16264 3148 16313 3176
rect 16264 3136 16270 3148
rect 16301 3145 16313 3148
rect 16347 3145 16359 3179
rect 16666 3176 16672 3188
rect 16627 3148 16672 3176
rect 16301 3139 16359 3145
rect 16666 3136 16672 3148
rect 16724 3136 16730 3188
rect 17034 3176 17040 3188
rect 16995 3148 17040 3176
rect 17034 3136 17040 3148
rect 17092 3136 17098 3188
rect 17497 3179 17555 3185
rect 17497 3145 17509 3179
rect 17543 3176 17555 3179
rect 17678 3176 17684 3188
rect 17543 3148 17684 3176
rect 17543 3145 17555 3148
rect 17497 3139 17555 3145
rect 17678 3136 17684 3148
rect 17736 3136 17742 3188
rect 17865 3179 17923 3185
rect 17865 3145 17877 3179
rect 17911 3176 17923 3179
rect 18138 3176 18144 3188
rect 17911 3148 18144 3176
rect 17911 3145 17923 3148
rect 17865 3139 17923 3145
rect 5994 3108 6000 3120
rect 5460 3080 6000 3108
rect 5994 3068 6000 3080
rect 6052 3108 6058 3120
rect 6181 3111 6239 3117
rect 6181 3108 6193 3111
rect 6052 3080 6193 3108
rect 6052 3068 6058 3080
rect 6181 3077 6193 3080
rect 6227 3108 6239 3111
rect 6549 3111 6607 3117
rect 6549 3108 6561 3111
rect 6227 3080 6561 3108
rect 6227 3077 6239 3080
rect 6181 3071 6239 3077
rect 6549 3077 6561 3080
rect 6595 3077 6607 3111
rect 11992 3108 12020 3136
rect 12526 3108 12532 3120
rect 11992 3080 12532 3108
rect 6549 3071 6607 3077
rect 1762 3040 1768 3052
rect 1596 3012 1768 3040
rect 1762 3000 1768 3012
rect 1820 3000 1826 3052
rect 3786 3000 3792 3052
rect 3844 3040 3850 3052
rect 3844 3012 4384 3040
rect 3844 3000 3850 3012
rect 4154 2972 4160 2984
rect 4115 2944 4160 2972
rect 4154 2932 4160 2944
rect 4212 2972 4218 2984
rect 4249 2975 4307 2981
rect 4249 2972 4261 2975
rect 4212 2944 4261 2972
rect 4212 2932 4218 2944
rect 4249 2941 4261 2944
rect 4295 2941 4307 2975
rect 4356 2972 4384 3012
rect 4516 2975 4574 2981
rect 4516 2972 4528 2975
rect 4356 2944 4528 2972
rect 4249 2935 4307 2941
rect 4516 2941 4528 2944
rect 4562 2972 4574 2975
rect 5442 2972 5448 2984
rect 4562 2944 5448 2972
rect 4562 2941 4574 2944
rect 4516 2935 4574 2941
rect 5442 2932 5448 2944
rect 5500 2932 5506 2984
rect 6564 2972 6592 3071
rect 12526 3068 12532 3080
rect 12584 3068 12590 3120
rect 15764 3108 15792 3136
rect 17880 3108 17908 3139
rect 18138 3136 18144 3148
rect 18196 3136 18202 3188
rect 18414 3176 18420 3188
rect 18375 3148 18420 3176
rect 18414 3136 18420 3148
rect 18472 3136 18478 3188
rect 18966 3136 18972 3188
rect 19024 3176 19030 3188
rect 19153 3179 19211 3185
rect 19153 3176 19165 3179
rect 19024 3148 19165 3176
rect 19024 3136 19030 3148
rect 19153 3145 19165 3148
rect 19199 3145 19211 3179
rect 19153 3139 19211 3145
rect 15764 3080 17908 3108
rect 14274 3049 14280 3052
rect 13817 3043 13875 3049
rect 13817 3009 13829 3043
rect 13863 3040 13875 3043
rect 14232 3043 14280 3049
rect 14232 3040 14244 3043
rect 13863 3012 14244 3040
rect 13863 3009 13875 3012
rect 13817 3003 13875 3009
rect 14232 3009 14244 3012
rect 14278 3009 14280 3043
rect 14232 3003 14280 3009
rect 14274 3000 14280 3003
rect 14332 3000 14338 3052
rect 14369 3043 14427 3049
rect 14369 3009 14381 3043
rect 14415 3040 14427 3043
rect 14458 3040 14464 3052
rect 14415 3012 14464 3040
rect 14415 3009 14427 3012
rect 14369 3003 14427 3009
rect 14458 3000 14464 3012
rect 14516 3000 14522 3052
rect 14550 3000 14556 3052
rect 14608 3040 14614 3052
rect 14645 3043 14703 3049
rect 14645 3040 14657 3043
rect 14608 3012 14657 3040
rect 14608 3000 14614 3012
rect 14645 3009 14657 3012
rect 14691 3009 14703 3043
rect 18874 3040 18880 3052
rect 14645 3003 14703 3009
rect 18248 3012 18880 3040
rect 7190 2981 7196 2984
rect 6917 2975 6975 2981
rect 6917 2972 6929 2975
rect 6564 2944 6929 2972
rect 6917 2941 6929 2944
rect 6963 2941 6975 2975
rect 7184 2972 7196 2981
rect 7151 2944 7196 2972
rect 6917 2935 6975 2941
rect 7184 2935 7196 2944
rect 2032 2907 2090 2913
rect 2032 2873 2044 2907
rect 2078 2904 2090 2907
rect 2958 2904 2964 2916
rect 2078 2876 2964 2904
rect 2078 2873 2090 2876
rect 2032 2867 2090 2873
rect 2958 2864 2964 2876
rect 3016 2864 3022 2916
rect 4798 2904 4804 2916
rect 3160 2876 4804 2904
rect 1670 2796 1676 2848
rect 1728 2836 1734 2848
rect 2682 2836 2688 2848
rect 1728 2808 2688 2836
rect 1728 2796 1734 2808
rect 2682 2796 2688 2808
rect 2740 2796 2746 2848
rect 3160 2845 3188 2876
rect 4798 2864 4804 2876
rect 4856 2864 4862 2916
rect 6932 2904 6960 2935
rect 7190 2932 7196 2935
rect 7248 2932 7254 2984
rect 8938 2972 8944 2984
rect 8899 2944 8944 2972
rect 8938 2932 8944 2944
rect 8996 2932 9002 2984
rect 9309 2975 9367 2981
rect 9309 2941 9321 2975
rect 9355 2972 9367 2975
rect 9401 2975 9459 2981
rect 9401 2972 9413 2975
rect 9355 2944 9413 2972
rect 9355 2941 9367 2944
rect 9309 2935 9367 2941
rect 9401 2941 9413 2944
rect 9447 2972 9459 2975
rect 9490 2972 9496 2984
rect 9447 2944 9496 2972
rect 9447 2941 9459 2944
rect 9401 2935 9459 2941
rect 9324 2904 9352 2935
rect 9490 2932 9496 2944
rect 9548 2932 9554 2984
rect 9668 2975 9726 2981
rect 9668 2941 9680 2975
rect 9714 2972 9726 2975
rect 9950 2972 9956 2984
rect 9714 2944 9956 2972
rect 9714 2941 9726 2944
rect 9668 2935 9726 2941
rect 9950 2932 9956 2944
rect 10008 2932 10014 2984
rect 12437 2975 12495 2981
rect 12437 2941 12449 2975
rect 12483 2972 12495 2975
rect 13909 2975 13967 2981
rect 12483 2944 13124 2972
rect 12483 2941 12495 2944
rect 12437 2935 12495 2941
rect 6932 2876 9352 2904
rect 10318 2864 10324 2916
rect 10376 2904 10382 2916
rect 11701 2907 11759 2913
rect 11701 2904 11713 2907
rect 10376 2876 11713 2904
rect 10376 2864 10382 2876
rect 11701 2873 11713 2876
rect 11747 2873 11759 2907
rect 11701 2867 11759 2873
rect 13096 2848 13124 2944
rect 13909 2941 13921 2975
rect 13955 2972 13967 2975
rect 13998 2972 14004 2984
rect 13955 2944 14004 2972
rect 13955 2941 13967 2944
rect 13909 2935 13967 2941
rect 13998 2932 14004 2944
rect 14056 2932 14062 2984
rect 16666 2932 16672 2984
rect 16724 2972 16730 2984
rect 18248 2981 18276 3012
rect 18874 3000 18880 3012
rect 18932 3000 18938 3052
rect 19168 3040 19196 3139
rect 20714 3136 20720 3188
rect 20772 3176 20778 3188
rect 21545 3179 21603 3185
rect 21545 3176 21557 3179
rect 20772 3148 21557 3176
rect 20772 3136 20778 3148
rect 21545 3145 21557 3148
rect 21591 3176 21603 3179
rect 21637 3179 21695 3185
rect 21637 3176 21649 3179
rect 21591 3148 21649 3176
rect 21591 3145 21603 3148
rect 21545 3139 21603 3145
rect 21637 3145 21649 3148
rect 21683 3145 21695 3179
rect 21637 3139 21695 3145
rect 24578 3136 24584 3188
rect 24636 3176 24642 3188
rect 25041 3179 25099 3185
rect 25041 3176 25053 3179
rect 24636 3148 25053 3176
rect 24636 3136 24642 3148
rect 25041 3145 25053 3148
rect 25087 3145 25099 3179
rect 25041 3139 25099 3145
rect 21358 3108 21364 3120
rect 21319 3080 21364 3108
rect 21358 3068 21364 3080
rect 21416 3068 21422 3120
rect 25056 3108 25084 3139
rect 26050 3136 26056 3188
rect 26108 3176 26114 3188
rect 26510 3176 26516 3188
rect 26108 3148 26516 3176
rect 26108 3136 26114 3148
rect 26510 3136 26516 3148
rect 26568 3136 26574 3188
rect 27614 3136 27620 3188
rect 27672 3176 27678 3188
rect 27982 3176 27988 3188
rect 27672 3148 27988 3176
rect 27672 3136 27678 3148
rect 27982 3136 27988 3148
rect 28040 3176 28046 3188
rect 28902 3176 28908 3188
rect 28040 3148 28908 3176
rect 28040 3136 28046 3148
rect 28902 3136 28908 3148
rect 28960 3136 28966 3188
rect 31018 3176 31024 3188
rect 30979 3148 31024 3176
rect 31018 3136 31024 3148
rect 31076 3136 31082 3188
rect 31938 3136 31944 3188
rect 31996 3176 32002 3188
rect 33873 3179 33931 3185
rect 33873 3176 33885 3179
rect 31996 3148 33885 3176
rect 31996 3136 32002 3148
rect 33873 3145 33885 3148
rect 33919 3145 33931 3179
rect 34238 3176 34244 3188
rect 34199 3148 34244 3176
rect 33873 3139 33931 3145
rect 34238 3136 34244 3148
rect 34296 3136 34302 3188
rect 34514 3136 34520 3188
rect 34572 3176 34578 3188
rect 34609 3179 34667 3185
rect 34609 3176 34621 3179
rect 34572 3148 34621 3176
rect 34572 3136 34578 3148
rect 34609 3145 34621 3148
rect 34655 3145 34667 3179
rect 34609 3139 34667 3145
rect 26234 3108 26240 3120
rect 25056 3080 26240 3108
rect 26234 3068 26240 3080
rect 26292 3068 26298 3120
rect 28626 3108 28632 3120
rect 28587 3080 28632 3108
rect 28626 3068 28632 3080
rect 28684 3068 28690 3120
rect 19337 3043 19395 3049
rect 19337 3040 19349 3043
rect 19168 3012 19349 3040
rect 19337 3009 19349 3012
rect 19383 3009 19395 3043
rect 19337 3003 19395 3009
rect 16853 2975 16911 2981
rect 16853 2972 16865 2975
rect 16724 2944 16865 2972
rect 16724 2932 16730 2944
rect 16853 2941 16865 2944
rect 16899 2941 16911 2975
rect 16853 2935 16911 2941
rect 18233 2975 18291 2981
rect 18233 2941 18245 2975
rect 18279 2941 18291 2975
rect 18233 2935 18291 2941
rect 19352 2904 19380 3003
rect 20898 3000 20904 3052
rect 20956 3040 20962 3052
rect 22462 3040 22468 3052
rect 20956 3012 22324 3040
rect 22423 3012 22468 3040
rect 20956 3000 20962 3012
rect 19604 2975 19662 2981
rect 19604 2941 19616 2975
rect 19650 2972 19662 2975
rect 19978 2972 19984 2984
rect 19650 2944 19984 2972
rect 19650 2941 19662 2944
rect 19604 2935 19662 2941
rect 19978 2932 19984 2944
rect 20036 2932 20042 2984
rect 22296 2981 22324 3012
rect 22462 3000 22468 3012
rect 22520 3000 22526 3052
rect 29730 3000 29736 3052
rect 29788 3040 29794 3052
rect 30009 3043 30067 3049
rect 30009 3040 30021 3043
rect 29788 3012 30021 3040
rect 29788 3000 29794 3012
rect 30009 3009 30021 3012
rect 30055 3009 30067 3043
rect 30009 3003 30067 3009
rect 30098 3000 30104 3052
rect 30156 3040 30162 3052
rect 31036 3040 31064 3136
rect 31436 3043 31494 3049
rect 31436 3040 31448 3043
rect 30156 3012 30201 3040
rect 31036 3012 31448 3040
rect 30156 3000 30162 3012
rect 21545 2975 21603 2981
rect 21545 2941 21557 2975
rect 21591 2972 21603 2975
rect 22189 2975 22247 2981
rect 22189 2972 22201 2975
rect 21591 2944 22201 2972
rect 21591 2941 21603 2944
rect 21545 2935 21603 2941
rect 22189 2941 22201 2944
rect 22235 2941 22247 2975
rect 22189 2935 22247 2941
rect 22281 2975 22339 2981
rect 22281 2941 22293 2975
rect 22327 2972 22339 2975
rect 22646 2972 22652 2984
rect 22327 2944 22652 2972
rect 22327 2941 22339 2944
rect 22281 2935 22339 2941
rect 22646 2932 22652 2944
rect 22704 2932 22710 2984
rect 23109 2975 23167 2981
rect 23109 2941 23121 2975
rect 23155 2972 23167 2975
rect 23198 2972 23204 2984
rect 23155 2944 23204 2972
rect 23155 2941 23167 2944
rect 23109 2935 23167 2941
rect 20622 2904 20628 2916
rect 19352 2876 20628 2904
rect 20622 2864 20628 2876
rect 20680 2864 20686 2916
rect 22094 2864 22100 2916
rect 22152 2904 22158 2916
rect 23124 2904 23152 2935
rect 23198 2932 23204 2944
rect 23256 2972 23262 2984
rect 23477 2975 23535 2981
rect 23477 2972 23489 2975
rect 23256 2944 23489 2972
rect 23256 2932 23262 2944
rect 23477 2941 23489 2944
rect 23523 2972 23535 2975
rect 23661 2975 23719 2981
rect 23661 2972 23673 2975
rect 23523 2944 23673 2972
rect 23523 2941 23535 2944
rect 23477 2935 23535 2941
rect 23661 2941 23673 2944
rect 23707 2972 23719 2975
rect 23750 2972 23756 2984
rect 23707 2944 23756 2972
rect 23707 2941 23719 2944
rect 23661 2935 23719 2941
rect 23750 2932 23756 2944
rect 23808 2972 23814 2984
rect 26145 2975 26203 2981
rect 26145 2972 26157 2975
rect 23808 2944 26157 2972
rect 23808 2932 23814 2944
rect 26145 2941 26157 2944
rect 26191 2972 26203 2975
rect 26602 2972 26608 2984
rect 26660 2981 26666 2984
rect 26878 2981 26884 2984
rect 26191 2944 26608 2972
rect 26191 2941 26203 2944
rect 26145 2935 26203 2941
rect 26602 2932 26608 2944
rect 26660 2972 26670 2981
rect 26872 2972 26884 2981
rect 26660 2944 26705 2972
rect 26804 2944 26884 2972
rect 26660 2935 26670 2944
rect 26660 2932 26666 2935
rect 22152 2876 23152 2904
rect 22152 2864 22158 2876
rect 23566 2864 23572 2916
rect 23624 2904 23630 2916
rect 23906 2907 23964 2913
rect 23906 2904 23918 2907
rect 23624 2876 23918 2904
rect 23624 2864 23630 2876
rect 23906 2873 23918 2876
rect 23952 2873 23964 2907
rect 23906 2867 23964 2873
rect 25682 2864 25688 2916
rect 25740 2904 25746 2916
rect 25777 2907 25835 2913
rect 25777 2904 25789 2907
rect 25740 2876 25789 2904
rect 25740 2864 25746 2876
rect 25777 2873 25789 2876
rect 25823 2904 25835 2907
rect 26804 2904 26832 2944
rect 26872 2935 26884 2944
rect 26878 2932 26884 2935
rect 26936 2932 26942 2984
rect 31110 2972 31116 2984
rect 31071 2944 31116 2972
rect 31110 2932 31116 2944
rect 31168 2932 31174 2984
rect 25823 2876 26832 2904
rect 29089 2907 29147 2913
rect 25823 2873 25835 2876
rect 25777 2867 25835 2873
rect 29089 2873 29101 2907
rect 29135 2904 29147 2907
rect 29638 2904 29644 2916
rect 29135 2876 29644 2904
rect 29135 2873 29147 2876
rect 29089 2867 29147 2873
rect 3145 2839 3203 2845
rect 3145 2805 3157 2839
rect 3191 2805 3203 2839
rect 3694 2836 3700 2848
rect 3655 2808 3700 2836
rect 3145 2799 3203 2805
rect 3694 2796 3700 2808
rect 3752 2796 3758 2848
rect 12253 2839 12311 2845
rect 12253 2805 12265 2839
rect 12299 2836 12311 2839
rect 12434 2836 12440 2848
rect 12299 2808 12440 2836
rect 12299 2805 12311 2808
rect 12253 2799 12311 2805
rect 12434 2796 12440 2808
rect 12492 2796 12498 2848
rect 13078 2836 13084 2848
rect 13039 2808 13084 2836
rect 13078 2796 13084 2808
rect 13136 2796 13142 2848
rect 20717 2839 20775 2845
rect 20717 2805 20729 2839
rect 20763 2836 20775 2839
rect 20806 2836 20812 2848
rect 20763 2808 20812 2836
rect 20763 2805 20775 2808
rect 20717 2799 20775 2805
rect 20806 2796 20812 2808
rect 20864 2796 20870 2848
rect 21818 2836 21824 2848
rect 21779 2808 21824 2836
rect 21818 2796 21824 2808
rect 21876 2796 21882 2848
rect 26602 2796 26608 2848
rect 26660 2836 26666 2848
rect 29104 2836 29132 2867
rect 29638 2864 29644 2876
rect 29696 2864 29702 2916
rect 29917 2907 29975 2913
rect 29917 2873 29929 2907
rect 29963 2904 29975 2907
rect 30561 2907 30619 2913
rect 30561 2904 30573 2907
rect 29963 2876 30573 2904
rect 29963 2873 29975 2876
rect 29917 2867 29975 2873
rect 30561 2873 30573 2876
rect 30607 2904 30619 2907
rect 30650 2904 30656 2916
rect 30607 2876 30656 2904
rect 30607 2873 30619 2876
rect 30561 2867 30619 2873
rect 30650 2864 30656 2876
rect 30708 2864 30714 2916
rect 29546 2836 29552 2848
rect 26660 2808 29132 2836
rect 29507 2808 29552 2836
rect 26660 2796 26666 2808
rect 29546 2796 29552 2808
rect 29604 2796 29610 2848
rect 31220 2836 31248 3012
rect 31436 3009 31448 3012
rect 31482 3009 31494 3043
rect 31570 3040 31576 3052
rect 31531 3012 31576 3040
rect 31436 3003 31494 3009
rect 31570 3000 31576 3012
rect 31628 3000 31634 3052
rect 31849 3043 31907 3049
rect 31849 3009 31861 3043
rect 31895 3040 31907 3043
rect 32030 3040 32036 3052
rect 31895 3012 32036 3040
rect 31895 3009 31907 3012
rect 31849 3003 31907 3009
rect 32030 3000 32036 3012
rect 32088 3000 32094 3052
rect 32950 3040 32956 3052
rect 32911 3012 32956 3040
rect 32950 3000 32956 3012
rect 33008 3000 33014 3052
rect 34624 2972 34652 3139
rect 35342 3040 35348 3052
rect 35303 3012 35348 3040
rect 35342 3000 35348 3012
rect 35400 3000 35406 3052
rect 35434 3000 35440 3052
rect 35492 3040 35498 3052
rect 35897 3043 35955 3049
rect 35897 3040 35909 3043
rect 35492 3012 35909 3040
rect 35492 3000 35498 3012
rect 35897 3009 35909 3012
rect 35943 3009 35955 3043
rect 35897 3003 35955 3009
rect 35253 2975 35311 2981
rect 35253 2972 35265 2975
rect 34624 2944 35265 2972
rect 35253 2941 35265 2944
rect 35299 2941 35311 2975
rect 35253 2935 35311 2941
rect 37274 2904 37280 2916
rect 32508 2876 37280 2904
rect 32508 2836 32536 2876
rect 37274 2864 37280 2876
rect 37332 2904 37338 2916
rect 38286 2904 38292 2916
rect 37332 2876 38292 2904
rect 37332 2864 37338 2876
rect 38286 2864 38292 2876
rect 38344 2864 38350 2916
rect 33594 2836 33600 2848
rect 31220 2808 32536 2836
rect 33555 2808 33600 2836
rect 33594 2796 33600 2808
rect 33652 2796 33658 2848
rect 34882 2836 34888 2848
rect 34843 2808 34888 2836
rect 34882 2796 34888 2808
rect 34940 2796 34946 2848
rect 1104 2746 38824 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 38824 2746
rect 1104 2672 38824 2694
rect 1762 2632 1768 2644
rect 1723 2604 1768 2632
rect 1762 2592 1768 2604
rect 1820 2632 1826 2644
rect 2133 2635 2191 2641
rect 2133 2632 2145 2635
rect 1820 2604 2145 2632
rect 1820 2592 1826 2604
rect 2133 2601 2145 2604
rect 2179 2601 2191 2635
rect 2406 2632 2412 2644
rect 2367 2604 2412 2632
rect 2133 2595 2191 2601
rect 2148 2360 2176 2595
rect 2406 2592 2412 2604
rect 2464 2592 2470 2644
rect 2774 2592 2780 2644
rect 2832 2632 2838 2644
rect 2869 2635 2927 2641
rect 2869 2632 2881 2635
rect 2832 2604 2881 2632
rect 2832 2592 2838 2604
rect 2869 2601 2881 2604
rect 2915 2632 2927 2635
rect 3421 2635 3479 2641
rect 3421 2632 3433 2635
rect 2915 2604 3433 2632
rect 2915 2601 2927 2604
rect 2869 2595 2927 2601
rect 3421 2601 3433 2604
rect 3467 2632 3479 2635
rect 3694 2632 3700 2644
rect 3467 2604 3700 2632
rect 3467 2601 3479 2604
rect 3421 2595 3479 2601
rect 3694 2592 3700 2604
rect 3752 2592 3758 2644
rect 5442 2632 5448 2644
rect 5403 2604 5448 2632
rect 5442 2592 5448 2604
rect 5500 2592 5506 2644
rect 6917 2635 6975 2641
rect 6917 2601 6929 2635
rect 6963 2632 6975 2635
rect 7006 2632 7012 2644
rect 6963 2604 7012 2632
rect 6963 2601 6975 2604
rect 6917 2595 6975 2601
rect 7006 2592 7012 2604
rect 7064 2592 7070 2644
rect 7190 2592 7196 2644
rect 7248 2632 7254 2644
rect 7285 2635 7343 2641
rect 7285 2632 7297 2635
rect 7248 2604 7297 2632
rect 7248 2592 7254 2604
rect 7285 2601 7297 2604
rect 7331 2601 7343 2635
rect 8294 2632 8300 2644
rect 8255 2604 8300 2632
rect 7285 2595 7343 2601
rect 8294 2592 8300 2604
rect 8352 2632 8358 2644
rect 8849 2635 8907 2641
rect 8352 2604 8708 2632
rect 8352 2592 8358 2604
rect 2958 2564 2964 2576
rect 2792 2536 2964 2564
rect 2792 2505 2820 2536
rect 2958 2524 2964 2536
rect 3016 2564 3022 2576
rect 8680 2573 8708 2604
rect 8849 2601 8861 2635
rect 8895 2632 8907 2635
rect 9306 2632 9312 2644
rect 8895 2604 9312 2632
rect 8895 2601 8907 2604
rect 8849 2595 8907 2601
rect 9306 2592 9312 2604
rect 9364 2592 9370 2644
rect 10318 2632 10324 2644
rect 10279 2604 10324 2632
rect 10318 2592 10324 2604
rect 10376 2592 10382 2644
rect 10778 2592 10784 2644
rect 10836 2632 10842 2644
rect 10873 2635 10931 2641
rect 10873 2632 10885 2635
rect 10836 2604 10885 2632
rect 10836 2592 10842 2604
rect 10873 2601 10885 2604
rect 10919 2632 10931 2635
rect 11241 2635 11299 2641
rect 11241 2632 11253 2635
rect 10919 2604 11253 2632
rect 10919 2601 10931 2604
rect 10873 2595 10931 2601
rect 11241 2601 11253 2604
rect 11287 2601 11299 2635
rect 11241 2595 11299 2601
rect 14090 2592 14096 2644
rect 14148 2632 14154 2644
rect 14277 2635 14335 2641
rect 14277 2632 14289 2635
rect 14148 2604 14289 2632
rect 14148 2592 14154 2604
rect 14277 2601 14289 2604
rect 14323 2601 14335 2635
rect 16850 2632 16856 2644
rect 16811 2604 16856 2632
rect 14277 2595 14335 2601
rect 16850 2592 16856 2604
rect 16908 2592 16914 2644
rect 17497 2635 17555 2641
rect 17497 2601 17509 2635
rect 17543 2632 17555 2635
rect 17862 2632 17868 2644
rect 17543 2604 17868 2632
rect 17543 2601 17555 2604
rect 17497 2595 17555 2601
rect 17862 2592 17868 2604
rect 17920 2592 17926 2644
rect 18141 2635 18199 2641
rect 18141 2601 18153 2635
rect 18187 2632 18199 2635
rect 18966 2632 18972 2644
rect 18187 2604 18972 2632
rect 18187 2601 18199 2604
rect 18141 2595 18199 2601
rect 5997 2567 6055 2573
rect 5997 2564 6009 2567
rect 3016 2536 6009 2564
rect 3016 2524 3022 2536
rect 5997 2533 6009 2536
rect 6043 2533 6055 2567
rect 5997 2527 6055 2533
rect 8665 2567 8723 2573
rect 8665 2533 8677 2567
rect 8711 2533 8723 2567
rect 8665 2527 8723 2533
rect 9585 2567 9643 2573
rect 9585 2533 9597 2567
rect 9631 2564 9643 2567
rect 10134 2564 10140 2576
rect 9631 2536 10140 2564
rect 9631 2533 9643 2536
rect 9585 2527 9643 2533
rect 10134 2524 10140 2536
rect 10192 2564 10198 2576
rect 10229 2567 10287 2573
rect 10229 2564 10241 2567
rect 10192 2536 10241 2564
rect 10192 2524 10198 2536
rect 10229 2533 10241 2536
rect 10275 2533 10287 2567
rect 10229 2527 10287 2533
rect 12434 2524 12440 2576
rect 12492 2564 12498 2576
rect 13142 2567 13200 2573
rect 13142 2564 13154 2567
rect 12492 2536 13154 2564
rect 12492 2524 12498 2536
rect 13142 2533 13154 2536
rect 13188 2564 13200 2567
rect 13722 2564 13728 2576
rect 13188 2536 13728 2564
rect 13188 2533 13200 2536
rect 13142 2527 13200 2533
rect 13722 2524 13728 2536
rect 13780 2524 13786 2576
rect 15488 2536 15884 2564
rect 2777 2499 2835 2505
rect 2777 2465 2789 2499
rect 2823 2465 2835 2499
rect 2777 2459 2835 2465
rect 4332 2499 4390 2505
rect 4332 2465 4344 2499
rect 4378 2496 4390 2499
rect 4798 2496 4804 2508
rect 4378 2468 4804 2496
rect 4378 2465 4390 2468
rect 4332 2459 4390 2465
rect 4798 2456 4804 2468
rect 4856 2496 4862 2508
rect 6365 2499 6423 2505
rect 6365 2496 6377 2499
rect 4856 2468 6377 2496
rect 4856 2456 4862 2468
rect 6365 2465 6377 2468
rect 6411 2465 6423 2499
rect 6365 2459 6423 2465
rect 6914 2456 6920 2508
rect 6972 2496 6978 2508
rect 7377 2499 7435 2505
rect 7377 2496 7389 2499
rect 6972 2468 7389 2496
rect 6972 2456 6978 2468
rect 7377 2465 7389 2468
rect 7423 2496 7435 2499
rect 7929 2499 7987 2505
rect 7929 2496 7941 2499
rect 7423 2468 7941 2496
rect 7423 2465 7435 2468
rect 7377 2459 7435 2465
rect 7929 2465 7941 2468
rect 7975 2465 7987 2499
rect 7929 2459 7987 2465
rect 8481 2499 8539 2505
rect 8481 2465 8493 2499
rect 8527 2465 8539 2499
rect 8481 2459 8539 2465
rect 11425 2499 11483 2505
rect 11425 2465 11437 2499
rect 11471 2496 11483 2499
rect 12066 2496 12072 2508
rect 11471 2468 12072 2496
rect 11471 2465 11483 2468
rect 11425 2459 11483 2465
rect 3050 2428 3056 2440
rect 3011 2400 3056 2428
rect 3050 2388 3056 2400
rect 3108 2388 3114 2440
rect 4062 2428 4068 2440
rect 3975 2400 4068 2428
rect 4062 2388 4068 2400
rect 4120 2388 4126 2440
rect 7561 2431 7619 2437
rect 7561 2397 7573 2431
rect 7607 2428 7619 2431
rect 8202 2428 8208 2440
rect 7607 2400 8208 2428
rect 7607 2397 7619 2400
rect 7561 2391 7619 2397
rect 8202 2388 8208 2400
rect 8260 2388 8266 2440
rect 8496 2428 8524 2459
rect 12066 2456 12072 2468
rect 12124 2456 12130 2508
rect 13630 2456 13636 2508
rect 13688 2496 13694 2508
rect 15488 2505 15516 2536
rect 15289 2499 15347 2505
rect 13688 2468 14964 2496
rect 13688 2456 13694 2468
rect 9214 2428 9220 2440
rect 8496 2400 9220 2428
rect 9214 2388 9220 2400
rect 9272 2388 9278 2440
rect 10505 2431 10563 2437
rect 10505 2397 10517 2431
rect 10551 2428 10563 2431
rect 10778 2428 10784 2440
rect 10551 2400 10784 2428
rect 10551 2397 10563 2400
rect 10505 2391 10563 2397
rect 10778 2388 10784 2400
rect 10836 2388 10842 2440
rect 12437 2431 12495 2437
rect 12437 2397 12449 2431
rect 12483 2428 12495 2431
rect 12526 2428 12532 2440
rect 12483 2400 12532 2428
rect 12483 2397 12495 2400
rect 12437 2391 12495 2397
rect 12526 2388 12532 2400
rect 12584 2428 12590 2440
rect 14936 2437 14964 2468
rect 15289 2465 15301 2499
rect 15335 2496 15347 2499
rect 15473 2499 15531 2505
rect 15473 2496 15485 2499
rect 15335 2468 15485 2496
rect 15335 2465 15347 2468
rect 15289 2459 15347 2465
rect 15473 2465 15485 2468
rect 15519 2465 15531 2499
rect 15729 2499 15787 2505
rect 15729 2496 15741 2499
rect 15473 2459 15531 2465
rect 15580 2468 15741 2496
rect 12897 2431 12955 2437
rect 12897 2428 12909 2431
rect 12584 2400 12909 2428
rect 12584 2388 12590 2400
rect 12897 2397 12909 2400
rect 12943 2397 12955 2431
rect 12897 2391 12955 2397
rect 14921 2431 14979 2437
rect 14921 2397 14933 2431
rect 14967 2428 14979 2431
rect 15580 2428 15608 2468
rect 15729 2465 15741 2468
rect 15775 2465 15787 2499
rect 15856 2496 15884 2536
rect 18156 2496 18184 2595
rect 18616 2505 18644 2604
rect 18966 2592 18972 2604
rect 19024 2592 19030 2644
rect 19150 2592 19156 2644
rect 19208 2632 19214 2644
rect 19978 2632 19984 2644
rect 19208 2604 19380 2632
rect 19939 2604 19984 2632
rect 19208 2592 19214 2604
rect 18868 2567 18926 2573
rect 18868 2533 18880 2567
rect 18914 2564 18926 2567
rect 19242 2564 19248 2576
rect 18914 2536 19248 2564
rect 18914 2533 18926 2536
rect 18868 2527 18926 2533
rect 19242 2524 19248 2536
rect 19300 2524 19306 2576
rect 19352 2564 19380 2604
rect 19978 2592 19984 2604
rect 20036 2592 20042 2644
rect 20714 2592 20720 2644
rect 20772 2632 20778 2644
rect 20901 2635 20959 2641
rect 20901 2632 20913 2635
rect 20772 2604 20913 2632
rect 20772 2592 20778 2604
rect 20901 2601 20913 2604
rect 20947 2601 20959 2635
rect 22554 2632 22560 2644
rect 22515 2604 22560 2632
rect 20901 2595 20959 2601
rect 22554 2592 22560 2604
rect 22612 2632 22618 2644
rect 23109 2635 23167 2641
rect 23109 2632 23121 2635
rect 22612 2604 23121 2632
rect 22612 2592 22618 2604
rect 23109 2601 23121 2604
rect 23155 2601 23167 2635
rect 23750 2632 23756 2644
rect 23711 2604 23756 2632
rect 23109 2595 23167 2601
rect 23750 2592 23756 2604
rect 23808 2592 23814 2644
rect 25682 2632 25688 2644
rect 25643 2604 25688 2632
rect 25682 2592 25688 2604
rect 25740 2592 25746 2644
rect 26234 2592 26240 2644
rect 26292 2632 26298 2644
rect 26602 2632 26608 2644
rect 26292 2604 26337 2632
rect 26563 2604 26608 2632
rect 26292 2592 26298 2604
rect 26602 2592 26608 2604
rect 26660 2592 26666 2644
rect 28537 2635 28595 2641
rect 28537 2601 28549 2635
rect 28583 2632 28595 2635
rect 28626 2632 28632 2644
rect 28583 2604 28632 2632
rect 28583 2601 28595 2604
rect 28537 2595 28595 2601
rect 28626 2592 28632 2604
rect 28684 2592 28690 2644
rect 31389 2635 31447 2641
rect 31389 2601 31401 2635
rect 31435 2601 31447 2635
rect 31389 2595 31447 2601
rect 20625 2567 20683 2573
rect 20625 2564 20637 2567
rect 19352 2536 20637 2564
rect 20625 2533 20637 2536
rect 20671 2564 20683 2567
rect 21422 2567 21480 2573
rect 21422 2564 21434 2567
rect 20671 2536 21434 2564
rect 20671 2533 20683 2536
rect 20625 2527 20683 2533
rect 21422 2533 21434 2536
rect 21468 2533 21480 2567
rect 21422 2527 21480 2533
rect 15856 2468 18184 2496
rect 18601 2499 18659 2505
rect 15729 2459 15787 2465
rect 18601 2465 18613 2499
rect 18647 2465 18659 2499
rect 18601 2459 18659 2465
rect 20714 2456 20720 2508
rect 20772 2496 20778 2508
rect 21177 2499 21235 2505
rect 21177 2496 21189 2499
rect 20772 2468 21189 2496
rect 20772 2456 20778 2468
rect 21177 2465 21189 2468
rect 21223 2496 21235 2499
rect 22002 2496 22008 2508
rect 21223 2468 22008 2496
rect 21223 2465 21235 2468
rect 21177 2459 21235 2465
rect 22002 2456 22008 2468
rect 22060 2456 22066 2508
rect 23768 2496 23796 2592
rect 24578 2573 24584 2576
rect 24572 2564 24584 2573
rect 24539 2536 24584 2564
rect 24572 2527 24584 2536
rect 24578 2524 24584 2527
rect 24636 2524 24642 2576
rect 24305 2499 24363 2505
rect 24305 2496 24317 2499
rect 23768 2468 24317 2496
rect 24305 2465 24317 2468
rect 24351 2465 24363 2499
rect 26620 2496 26648 2592
rect 27424 2567 27482 2573
rect 27424 2533 27436 2567
rect 27470 2564 27482 2567
rect 27522 2564 27528 2576
rect 27470 2536 27528 2564
rect 27470 2533 27482 2536
rect 27424 2527 27482 2533
rect 27522 2524 27528 2536
rect 27580 2524 27586 2576
rect 30190 2524 30196 2576
rect 30248 2573 30254 2576
rect 30248 2567 30312 2573
rect 30248 2533 30266 2567
rect 30300 2533 30312 2567
rect 31404 2564 31432 2595
rect 34054 2592 34060 2644
rect 34112 2632 34118 2644
rect 34149 2635 34207 2641
rect 34149 2632 34161 2635
rect 34112 2604 34161 2632
rect 34112 2592 34118 2604
rect 34149 2601 34161 2604
rect 34195 2601 34207 2635
rect 34790 2632 34796 2644
rect 34751 2604 34796 2632
rect 34149 2595 34207 2601
rect 34790 2592 34796 2604
rect 34848 2592 34854 2644
rect 35158 2632 35164 2644
rect 35119 2604 35164 2632
rect 35158 2592 35164 2604
rect 35216 2592 35222 2644
rect 35342 2592 35348 2644
rect 35400 2632 35406 2644
rect 35437 2635 35495 2641
rect 35437 2632 35449 2635
rect 35400 2604 35449 2632
rect 35400 2592 35406 2604
rect 35437 2601 35449 2604
rect 35483 2601 35495 2635
rect 36998 2632 37004 2644
rect 36959 2604 37004 2632
rect 35437 2595 35495 2601
rect 36998 2592 37004 2604
rect 37056 2592 37062 2644
rect 33036 2567 33094 2573
rect 33036 2564 33048 2567
rect 31404 2536 33048 2564
rect 30248 2527 30312 2533
rect 33036 2533 33048 2536
rect 33082 2564 33094 2567
rect 33082 2536 36124 2564
rect 33082 2533 33094 2536
rect 33036 2527 33094 2533
rect 30248 2524 30254 2527
rect 27157 2499 27215 2505
rect 27157 2496 27169 2499
rect 26620 2468 27169 2496
rect 24305 2459 24363 2465
rect 27157 2465 27169 2468
rect 27203 2465 27215 2499
rect 27157 2459 27215 2465
rect 29549 2499 29607 2505
rect 29549 2465 29561 2499
rect 29595 2496 29607 2499
rect 29638 2496 29644 2508
rect 29595 2468 29644 2496
rect 29595 2465 29607 2468
rect 29549 2459 29607 2465
rect 29638 2456 29644 2468
rect 29696 2496 29702 2508
rect 30009 2499 30067 2505
rect 30009 2496 30021 2499
rect 29696 2468 30021 2496
rect 29696 2456 29702 2468
rect 30009 2465 30021 2468
rect 30055 2496 30067 2499
rect 32401 2499 32459 2505
rect 32401 2496 32413 2499
rect 30055 2468 32413 2496
rect 30055 2465 30067 2468
rect 30009 2459 30067 2465
rect 32401 2465 32413 2468
rect 32447 2496 32459 2499
rect 32769 2499 32827 2505
rect 32769 2496 32781 2499
rect 32447 2468 32781 2496
rect 32447 2465 32459 2468
rect 32401 2459 32459 2465
rect 32769 2465 32781 2468
rect 32815 2496 32827 2499
rect 33594 2496 33600 2508
rect 32815 2468 33600 2496
rect 32815 2465 32827 2468
rect 32769 2459 32827 2465
rect 33594 2456 33600 2468
rect 33652 2456 33658 2508
rect 34790 2456 34796 2508
rect 34848 2496 34854 2508
rect 35805 2499 35863 2505
rect 35805 2496 35817 2499
rect 34848 2468 35817 2496
rect 34848 2456 34854 2468
rect 35805 2465 35817 2468
rect 35851 2465 35863 2499
rect 35805 2459 35863 2465
rect 14967 2400 15608 2428
rect 14967 2397 14979 2400
rect 14921 2391 14979 2397
rect 35158 2388 35164 2440
rect 35216 2428 35222 2440
rect 36096 2437 36124 2536
rect 35897 2431 35955 2437
rect 35897 2428 35909 2431
rect 35216 2400 35909 2428
rect 35216 2388 35222 2400
rect 35897 2397 35909 2400
rect 35943 2397 35955 2431
rect 35897 2391 35955 2397
rect 36081 2431 36139 2437
rect 36081 2397 36093 2431
rect 36127 2428 36139 2431
rect 36541 2431 36599 2437
rect 36541 2428 36553 2431
rect 36127 2400 36553 2428
rect 36127 2397 36139 2400
rect 36081 2391 36139 2397
rect 36541 2397 36553 2400
rect 36587 2428 36599 2431
rect 36817 2431 36875 2437
rect 36817 2428 36829 2431
rect 36587 2400 36829 2428
rect 36587 2397 36599 2400
rect 36541 2391 36599 2397
rect 36817 2397 36829 2400
rect 36863 2397 36875 2431
rect 36817 2391 36875 2397
rect 3789 2363 3847 2369
rect 3789 2360 3801 2363
rect 2148 2332 3801 2360
rect 3789 2329 3801 2332
rect 3835 2360 3847 2363
rect 4080 2360 4108 2388
rect 3835 2332 4108 2360
rect 9861 2363 9919 2369
rect 3835 2329 3847 2332
rect 3789 2323 3847 2329
rect 9861 2329 9873 2363
rect 9907 2360 9919 2363
rect 10962 2360 10968 2372
rect 9907 2332 10968 2360
rect 9907 2329 9919 2332
rect 9861 2323 9919 2329
rect 10962 2320 10968 2332
rect 11020 2320 11026 2372
rect 28902 2320 28908 2372
rect 28960 2360 28966 2372
rect 29181 2363 29239 2369
rect 29181 2360 29193 2363
rect 28960 2332 29193 2360
rect 28960 2320 28966 2332
rect 29181 2329 29193 2332
rect 29227 2360 29239 2363
rect 29227 2332 29592 2360
rect 29227 2329 29239 2332
rect 29181 2323 29239 2329
rect 11054 2252 11060 2304
rect 11112 2292 11118 2304
rect 11609 2295 11667 2301
rect 11609 2292 11621 2295
rect 11112 2264 11621 2292
rect 11112 2252 11118 2264
rect 11609 2261 11621 2264
rect 11655 2261 11667 2295
rect 29564 2292 29592 2332
rect 31941 2295 31999 2301
rect 31941 2292 31953 2295
rect 29564 2264 31953 2292
rect 11609 2255 11667 2261
rect 31941 2261 31953 2264
rect 31987 2261 31999 2295
rect 31941 2255 31999 2261
rect 1104 2202 38824 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 34966 2202
rect 35018 2150 35030 2202
rect 35082 2150 35094 2202
rect 35146 2150 35158 2202
rect 35210 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 35624 35819 35676 35828
rect 35624 35785 35633 35819
rect 35633 35785 35667 35819
rect 35667 35785 35676 35819
rect 35624 35776 35676 35785
rect 35440 35615 35492 35624
rect 35440 35581 35449 35615
rect 35449 35581 35483 35615
rect 35483 35581 35492 35615
rect 35440 35572 35492 35581
rect 30472 35547 30524 35556
rect 30472 35513 30506 35547
rect 30506 35513 30524 35547
rect 30472 35504 30524 35513
rect 30012 35479 30064 35488
rect 30012 35445 30021 35479
rect 30021 35445 30055 35479
rect 30055 35445 30064 35479
rect 30012 35436 30064 35445
rect 30840 35436 30892 35488
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 30288 35232 30340 35284
rect 30840 35275 30892 35284
rect 30840 35241 30849 35275
rect 30849 35241 30883 35275
rect 30883 35241 30892 35275
rect 30840 35232 30892 35241
rect 36176 35275 36228 35284
rect 36176 35241 36185 35275
rect 36185 35241 36219 35275
rect 36219 35241 36228 35275
rect 36176 35232 36228 35241
rect 30472 35096 30524 35148
rect 32036 35096 32088 35148
rect 34704 35096 34756 35148
rect 36176 35096 36228 35148
rect 29092 35028 29144 35080
rect 32772 35028 32824 35080
rect 34796 34960 34848 35012
rect 31668 34892 31720 34944
rect 33324 34935 33376 34944
rect 33324 34901 33333 34935
rect 33333 34901 33367 34935
rect 33367 34901 33376 34935
rect 33324 34892 33376 34901
rect 33692 34892 33744 34944
rect 34520 34892 34572 34944
rect 35532 34935 35584 34944
rect 35532 34901 35541 34935
rect 35541 34901 35575 34935
rect 35575 34901 35584 34935
rect 35532 34892 35584 34901
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 29092 34731 29144 34740
rect 29092 34697 29101 34731
rect 29101 34697 29135 34731
rect 29135 34697 29144 34731
rect 29092 34688 29144 34697
rect 30380 34688 30432 34740
rect 32772 34731 32824 34740
rect 32772 34697 32781 34731
rect 32781 34697 32815 34731
rect 32815 34697 32824 34731
rect 32772 34688 32824 34697
rect 33140 34688 33192 34740
rect 34152 34688 34204 34740
rect 34796 34688 34848 34740
rect 37556 34731 37608 34740
rect 37556 34697 37565 34731
rect 37565 34697 37599 34731
rect 37599 34697 37608 34731
rect 37556 34688 37608 34697
rect 32036 34663 32088 34672
rect 32036 34629 32045 34663
rect 32045 34629 32079 34663
rect 32079 34629 32088 34663
rect 32036 34620 32088 34629
rect 34428 34620 34480 34672
rect 36268 34663 36320 34672
rect 36268 34629 36277 34663
rect 36277 34629 36311 34663
rect 36311 34629 36320 34663
rect 36268 34620 36320 34629
rect 30012 34527 30064 34536
rect 29368 34348 29420 34400
rect 30012 34493 30021 34527
rect 30021 34493 30055 34527
rect 30055 34493 30064 34527
rect 30012 34484 30064 34493
rect 34152 34552 34204 34604
rect 34520 34552 34572 34604
rect 30288 34527 30340 34536
rect 30288 34493 30322 34527
rect 30322 34493 30340 34527
rect 30288 34484 30340 34493
rect 33324 34484 33376 34536
rect 35532 34484 35584 34536
rect 35900 34484 35952 34536
rect 36176 34484 36228 34536
rect 37924 34527 37976 34536
rect 37924 34493 37933 34527
rect 37933 34493 37967 34527
rect 37967 34493 37976 34527
rect 37924 34484 37976 34493
rect 33232 34391 33284 34400
rect 33232 34357 33241 34391
rect 33241 34357 33275 34391
rect 33275 34357 33284 34391
rect 33232 34348 33284 34357
rect 34612 34391 34664 34400
rect 34612 34357 34621 34391
rect 34621 34357 34655 34391
rect 34655 34357 34664 34391
rect 34612 34348 34664 34357
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 27712 34144 27764 34196
rect 29736 34144 29788 34196
rect 34152 34187 34204 34196
rect 34152 34153 34161 34187
rect 34161 34153 34195 34187
rect 34195 34153 34204 34187
rect 34152 34144 34204 34153
rect 35900 34144 35952 34196
rect 34520 34076 34572 34128
rect 36268 34076 36320 34128
rect 28724 34008 28776 34060
rect 30288 34008 30340 34060
rect 31576 34008 31628 34060
rect 28908 33940 28960 33992
rect 29368 33940 29420 33992
rect 32128 33983 32180 33992
rect 32128 33949 32137 33983
rect 32137 33949 32171 33983
rect 32171 33949 32180 33983
rect 32128 33940 32180 33949
rect 34612 33940 34664 33992
rect 27988 33847 28040 33856
rect 27988 33813 27997 33847
rect 27997 33813 28031 33847
rect 28031 33813 28040 33847
rect 27988 33804 28040 33813
rect 30932 33847 30984 33856
rect 30932 33813 30941 33847
rect 30941 33813 30975 33847
rect 30975 33813 30984 33847
rect 30932 33804 30984 33813
rect 32772 33804 32824 33856
rect 33508 33847 33560 33856
rect 33508 33813 33517 33847
rect 33517 33813 33551 33847
rect 33551 33813 33560 33847
rect 33508 33804 33560 33813
rect 34704 33804 34756 33856
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 34966 33702 35018 33754
rect 35030 33702 35082 33754
rect 35094 33702 35146 33754
rect 35158 33702 35210 33754
rect 27712 33643 27764 33652
rect 27712 33609 27721 33643
rect 27721 33609 27755 33643
rect 27755 33609 27764 33643
rect 27712 33600 27764 33609
rect 28724 33643 28776 33652
rect 28724 33609 28733 33643
rect 28733 33609 28767 33643
rect 28767 33609 28776 33643
rect 28724 33600 28776 33609
rect 32128 33600 32180 33652
rect 33876 33643 33928 33652
rect 33876 33609 33885 33643
rect 33885 33609 33919 33643
rect 33919 33609 33928 33643
rect 33876 33600 33928 33609
rect 36268 33643 36320 33652
rect 36268 33609 36277 33643
rect 36277 33609 36311 33643
rect 36311 33609 36320 33643
rect 36268 33600 36320 33609
rect 34244 33575 34296 33584
rect 34244 33541 34253 33575
rect 34253 33541 34287 33575
rect 34287 33541 34296 33575
rect 34612 33575 34664 33584
rect 34244 33532 34296 33541
rect 34612 33541 34621 33575
rect 34621 33541 34655 33575
rect 34655 33541 34664 33575
rect 34612 33532 34664 33541
rect 31760 33464 31812 33516
rect 32772 33507 32824 33516
rect 29736 33396 29788 33448
rect 30932 33396 30984 33448
rect 32772 33473 32781 33507
rect 32781 33473 32815 33507
rect 32815 33473 32824 33507
rect 32772 33464 32824 33473
rect 29368 33260 29420 33312
rect 31852 33328 31904 33380
rect 30472 33260 30524 33312
rect 31576 33303 31628 33312
rect 31576 33269 31585 33303
rect 31585 33269 31619 33303
rect 31619 33269 31628 33303
rect 31576 33260 31628 33269
rect 32128 33303 32180 33312
rect 32128 33269 32137 33303
rect 32137 33269 32171 33303
rect 32171 33269 32180 33303
rect 32128 33260 32180 33269
rect 34704 33328 34756 33380
rect 35808 33328 35860 33380
rect 34796 33260 34848 33312
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 28908 33056 28960 33108
rect 29736 33056 29788 33108
rect 31852 33099 31904 33108
rect 31852 33065 31861 33099
rect 31861 33065 31895 33099
rect 31895 33065 31904 33099
rect 31852 33056 31904 33065
rect 33232 33099 33284 33108
rect 33232 33065 33241 33099
rect 33241 33065 33275 33099
rect 33275 33065 33284 33099
rect 33232 33056 33284 33065
rect 34336 33056 34388 33108
rect 35808 33056 35860 33108
rect 29828 33031 29880 33040
rect 29828 32997 29862 33031
rect 29862 32997 29880 33031
rect 29828 32988 29880 32997
rect 34888 32988 34940 33040
rect 32036 32920 32088 32972
rect 36268 32920 36320 32972
rect 29368 32852 29420 32904
rect 32588 32895 32640 32904
rect 32588 32861 32597 32895
rect 32597 32861 32631 32895
rect 32631 32861 32640 32895
rect 32588 32852 32640 32861
rect 33140 32852 33192 32904
rect 34244 32852 34296 32904
rect 31760 32784 31812 32836
rect 30932 32759 30984 32768
rect 30932 32725 30941 32759
rect 30941 32725 30975 32759
rect 30975 32725 30984 32759
rect 30932 32716 30984 32725
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 34966 32614 35018 32666
rect 35030 32614 35082 32666
rect 35094 32614 35146 32666
rect 35158 32614 35210 32666
rect 29828 32512 29880 32564
rect 32036 32555 32088 32564
rect 32036 32521 32045 32555
rect 32045 32521 32079 32555
rect 32079 32521 32088 32555
rect 32036 32512 32088 32521
rect 32588 32512 32640 32564
rect 34244 32555 34296 32564
rect 34244 32521 34253 32555
rect 34253 32521 34287 32555
rect 34287 32521 34296 32555
rect 34244 32512 34296 32521
rect 34428 32512 34480 32564
rect 36268 32555 36320 32564
rect 32772 32444 32824 32496
rect 33416 32444 33468 32496
rect 33692 32419 33744 32428
rect 33692 32385 33701 32419
rect 33701 32385 33735 32419
rect 33735 32385 33744 32419
rect 33692 32376 33744 32385
rect 36268 32521 36277 32555
rect 36277 32521 36311 32555
rect 36311 32521 36320 32555
rect 36268 32512 36320 32521
rect 37556 32555 37608 32564
rect 37556 32521 37565 32555
rect 37565 32521 37599 32555
rect 37599 32521 37608 32555
rect 37556 32512 37608 32521
rect 29368 32308 29420 32360
rect 32128 32351 32180 32360
rect 32128 32317 32137 32351
rect 32137 32317 32171 32351
rect 32171 32317 32180 32351
rect 32128 32308 32180 32317
rect 33232 32308 33284 32360
rect 37372 32351 37424 32360
rect 37372 32317 37381 32351
rect 37381 32317 37415 32351
rect 37415 32317 37424 32351
rect 37372 32308 37424 32317
rect 30932 32240 30984 32292
rect 32588 32240 32640 32292
rect 35164 32283 35216 32292
rect 35164 32249 35198 32283
rect 35198 32249 35216 32283
rect 35164 32240 35216 32249
rect 29368 32172 29420 32224
rect 30104 32172 30156 32224
rect 32036 32172 32088 32224
rect 33232 32215 33284 32224
rect 33232 32181 33241 32215
rect 33241 32181 33275 32215
rect 33275 32181 33284 32215
rect 33232 32172 33284 32181
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 30380 31968 30432 32020
rect 33416 32011 33468 32020
rect 33416 31977 33425 32011
rect 33425 31977 33459 32011
rect 33459 31977 33468 32011
rect 33416 31968 33468 31977
rect 33784 31968 33836 32020
rect 35992 32011 36044 32020
rect 35992 31977 36001 32011
rect 36001 31977 36035 32011
rect 36035 31977 36044 32011
rect 35992 31968 36044 31977
rect 30288 31900 30340 31952
rect 28908 31875 28960 31884
rect 28908 31841 28917 31875
rect 28917 31841 28951 31875
rect 28951 31841 28960 31875
rect 28908 31832 28960 31841
rect 29828 31832 29880 31884
rect 30472 31807 30524 31816
rect 29368 31696 29420 31748
rect 29920 31696 29972 31748
rect 30472 31773 30481 31807
rect 30481 31773 30515 31807
rect 30515 31773 30524 31807
rect 30472 31764 30524 31773
rect 33140 31900 33192 31952
rect 34152 31900 34204 31952
rect 32956 31832 33008 31884
rect 33232 31832 33284 31884
rect 34520 31832 34572 31884
rect 35164 31832 35216 31884
rect 34152 31764 34204 31816
rect 34704 31807 34756 31816
rect 34704 31773 34713 31807
rect 34713 31773 34747 31807
rect 34747 31773 34756 31807
rect 34704 31764 34756 31773
rect 35348 31832 35400 31884
rect 32128 31628 32180 31680
rect 33048 31671 33100 31680
rect 33048 31637 33057 31671
rect 33057 31637 33091 31671
rect 33091 31637 33100 31671
rect 33048 31628 33100 31637
rect 34244 31671 34296 31680
rect 34244 31637 34253 31671
rect 34253 31637 34287 31671
rect 34287 31637 34296 31671
rect 34244 31628 34296 31637
rect 34428 31628 34480 31680
rect 34612 31628 34664 31680
rect 36820 31696 36872 31748
rect 36268 31628 36320 31680
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 34966 31526 35018 31578
rect 35030 31526 35082 31578
rect 35094 31526 35146 31578
rect 35158 31526 35210 31578
rect 29000 31467 29052 31476
rect 29000 31433 29009 31467
rect 29009 31433 29043 31467
rect 29043 31433 29052 31467
rect 29000 31424 29052 31433
rect 29828 31424 29880 31476
rect 29920 31467 29972 31476
rect 29920 31433 29929 31467
rect 29929 31433 29963 31467
rect 29963 31433 29972 31467
rect 32956 31467 33008 31476
rect 29920 31424 29972 31433
rect 32956 31433 32965 31467
rect 32965 31433 32999 31467
rect 32999 31433 33008 31467
rect 32956 31424 33008 31433
rect 34428 31424 34480 31476
rect 34612 31467 34664 31476
rect 34612 31433 34621 31467
rect 34621 31433 34655 31467
rect 34655 31433 34664 31467
rect 34612 31424 34664 31433
rect 36268 31467 36320 31476
rect 36268 31433 36277 31467
rect 36277 31433 36311 31467
rect 36311 31433 36320 31467
rect 36268 31424 36320 31433
rect 36820 31467 36872 31476
rect 36820 31433 36829 31467
rect 36829 31433 36863 31467
rect 36863 31433 36872 31467
rect 36820 31424 36872 31433
rect 30380 31288 30432 31340
rect 30564 31331 30616 31340
rect 30564 31297 30573 31331
rect 30573 31297 30607 31331
rect 30607 31297 30616 31331
rect 30564 31288 30616 31297
rect 32036 31331 32088 31340
rect 32036 31297 32045 31331
rect 32045 31297 32079 31331
rect 32079 31297 32088 31331
rect 32036 31288 32088 31297
rect 32128 31331 32180 31340
rect 32128 31297 32137 31331
rect 32137 31297 32171 31331
rect 32171 31297 32180 31331
rect 32128 31288 32180 31297
rect 31668 31152 31720 31204
rect 34704 31152 34756 31204
rect 35164 31195 35216 31204
rect 35164 31161 35198 31195
rect 35198 31161 35216 31195
rect 35164 31152 35216 31161
rect 31576 31127 31628 31136
rect 31576 31093 31585 31127
rect 31585 31093 31619 31127
rect 31619 31093 31628 31127
rect 31576 31084 31628 31093
rect 31944 31127 31996 31136
rect 31944 31093 31953 31127
rect 31953 31093 31987 31127
rect 31987 31093 31996 31127
rect 31944 31084 31996 31093
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 30380 30880 30432 30932
rect 31944 30880 31996 30932
rect 33048 30880 33100 30932
rect 33600 30880 33652 30932
rect 34244 30880 34296 30932
rect 35164 30880 35216 30932
rect 30104 30812 30156 30864
rect 34612 30812 34664 30864
rect 29368 30744 29420 30796
rect 34520 30744 34572 30796
rect 32680 30719 32732 30728
rect 32680 30685 32689 30719
rect 32689 30685 32723 30719
rect 32723 30685 32732 30719
rect 32680 30676 32732 30685
rect 31668 30608 31720 30660
rect 32128 30608 32180 30660
rect 33140 30676 33192 30728
rect 29552 30540 29604 30592
rect 30840 30540 30892 30592
rect 31760 30540 31812 30592
rect 34612 30540 34664 30592
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 34966 30438 35018 30490
rect 35030 30438 35082 30490
rect 35094 30438 35146 30490
rect 35158 30438 35210 30490
rect 32680 30379 32732 30388
rect 32680 30345 32689 30379
rect 32689 30345 32723 30379
rect 32723 30345 32732 30379
rect 32680 30336 32732 30345
rect 33048 30379 33100 30388
rect 33048 30345 33057 30379
rect 33057 30345 33091 30379
rect 33091 30345 33100 30379
rect 33048 30336 33100 30345
rect 34520 30379 34572 30388
rect 34520 30345 34529 30379
rect 34529 30345 34563 30379
rect 34563 30345 34572 30379
rect 34520 30336 34572 30345
rect 28816 30268 28868 30320
rect 31668 30311 31720 30320
rect 31668 30277 31677 30311
rect 31677 30277 31711 30311
rect 31711 30277 31720 30311
rect 31668 30268 31720 30277
rect 28724 30243 28776 30252
rect 28724 30209 28733 30243
rect 28733 30209 28767 30243
rect 28767 30209 28776 30243
rect 28724 30200 28776 30209
rect 29368 30243 29420 30252
rect 29368 30209 29377 30243
rect 29377 30209 29411 30243
rect 29411 30209 29420 30243
rect 29368 30200 29420 30209
rect 33876 30243 33928 30252
rect 33876 30209 33885 30243
rect 33885 30209 33919 30243
rect 33919 30209 33928 30243
rect 33876 30200 33928 30209
rect 34888 30243 34940 30252
rect 34888 30209 34897 30243
rect 34897 30209 34931 30243
rect 34931 30209 34940 30243
rect 34888 30200 34940 30209
rect 33600 30175 33652 30184
rect 33600 30141 33609 30175
rect 33609 30141 33643 30175
rect 33643 30141 33652 30175
rect 33600 30132 33652 30141
rect 29552 30064 29604 30116
rect 34520 30064 34572 30116
rect 27988 30039 28040 30048
rect 27988 30005 27997 30039
rect 27997 30005 28031 30039
rect 28031 30005 28040 30039
rect 27988 29996 28040 30005
rect 29092 29996 29144 30048
rect 33692 30039 33744 30048
rect 33692 30005 33701 30039
rect 33701 30005 33735 30039
rect 33735 30005 33744 30039
rect 33692 29996 33744 30005
rect 34612 29996 34664 30048
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 30104 29835 30156 29844
rect 30104 29801 30113 29835
rect 30113 29801 30147 29835
rect 30147 29801 30156 29835
rect 30104 29792 30156 29801
rect 33692 29792 33744 29844
rect 34888 29792 34940 29844
rect 35900 29792 35952 29844
rect 29092 29724 29144 29776
rect 30656 29767 30708 29776
rect 30656 29733 30665 29767
rect 30665 29733 30699 29767
rect 30699 29733 30708 29767
rect 30656 29724 30708 29733
rect 34152 29767 34204 29776
rect 34152 29733 34161 29767
rect 34161 29733 34195 29767
rect 34195 29733 34204 29767
rect 34152 29724 34204 29733
rect 28724 29656 28776 29708
rect 30840 29699 30892 29708
rect 30840 29665 30849 29699
rect 30849 29665 30883 29699
rect 30883 29665 30892 29699
rect 30840 29656 30892 29665
rect 32128 29699 32180 29708
rect 32128 29665 32137 29699
rect 32137 29665 32171 29699
rect 32171 29665 32180 29699
rect 32128 29656 32180 29665
rect 34612 29699 34664 29708
rect 34612 29665 34621 29699
rect 34621 29665 34655 29699
rect 34655 29665 34664 29699
rect 34612 29656 34664 29665
rect 34520 29588 34572 29640
rect 35808 29699 35860 29708
rect 35808 29665 35817 29699
rect 35817 29665 35851 29699
rect 35851 29665 35860 29699
rect 35808 29656 35860 29665
rect 35256 29588 35308 29640
rect 36268 29520 36320 29572
rect 27712 29495 27764 29504
rect 27712 29461 27721 29495
rect 27721 29461 27755 29495
rect 27755 29461 27764 29495
rect 27712 29452 27764 29461
rect 28448 29452 28500 29504
rect 30748 29452 30800 29504
rect 33876 29452 33928 29504
rect 36084 29452 36136 29504
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 34966 29350 35018 29402
rect 35030 29350 35082 29402
rect 35094 29350 35146 29402
rect 35158 29350 35210 29402
rect 27988 29248 28040 29300
rect 30656 29248 30708 29300
rect 32128 29291 32180 29300
rect 32128 29257 32137 29291
rect 32137 29257 32171 29291
rect 32171 29257 32180 29291
rect 32128 29248 32180 29257
rect 34612 29248 34664 29300
rect 34796 29248 34848 29300
rect 36268 29291 36320 29300
rect 36268 29257 36277 29291
rect 36277 29257 36311 29291
rect 36311 29257 36320 29291
rect 36268 29248 36320 29257
rect 28724 29223 28776 29232
rect 28724 29189 28733 29223
rect 28733 29189 28767 29223
rect 28767 29189 28776 29223
rect 28724 29180 28776 29189
rect 29092 29223 29144 29232
rect 29092 29189 29101 29223
rect 29101 29189 29135 29223
rect 29135 29189 29144 29223
rect 29092 29180 29144 29189
rect 29828 29180 29880 29232
rect 30840 29180 30892 29232
rect 33140 29180 33192 29232
rect 28448 29112 28500 29164
rect 30748 29112 30800 29164
rect 34336 29155 34388 29164
rect 27712 29044 27764 29096
rect 28908 29044 28960 29096
rect 30472 29087 30524 29096
rect 30472 29053 30481 29087
rect 30481 29053 30515 29087
rect 30515 29053 30524 29087
rect 30472 29044 30524 29053
rect 31668 29044 31720 29096
rect 34336 29121 34345 29155
rect 34345 29121 34379 29155
rect 34379 29121 34388 29155
rect 34336 29112 34388 29121
rect 28172 28976 28224 29028
rect 30380 29019 30432 29028
rect 30380 28985 30389 29019
rect 30389 28985 30423 29019
rect 30423 28985 30432 29019
rect 30380 28976 30432 28985
rect 31576 28976 31628 29028
rect 34980 28976 35032 29028
rect 35808 28976 35860 29028
rect 27620 28951 27672 28960
rect 27620 28917 27629 28951
rect 27629 28917 27663 28951
rect 27663 28917 27672 28951
rect 27620 28908 27672 28917
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 29092 28704 29144 28756
rect 30288 28704 30340 28756
rect 34428 28704 34480 28756
rect 34980 28747 35032 28756
rect 34980 28713 34989 28747
rect 34989 28713 35023 28747
rect 35023 28713 35032 28747
rect 34980 28704 35032 28713
rect 35624 28747 35676 28756
rect 35624 28713 35633 28747
rect 35633 28713 35667 28747
rect 35667 28713 35676 28747
rect 35624 28704 35676 28713
rect 36084 28704 36136 28756
rect 28448 28636 28500 28688
rect 27988 28611 28040 28620
rect 27988 28577 27997 28611
rect 27997 28577 28031 28611
rect 28031 28577 28040 28611
rect 27988 28568 28040 28577
rect 28724 28568 28776 28620
rect 30472 28611 30524 28620
rect 30472 28577 30481 28611
rect 30481 28577 30515 28611
rect 30515 28577 30524 28611
rect 30472 28568 30524 28577
rect 35440 28611 35492 28620
rect 35440 28577 35449 28611
rect 35449 28577 35483 28611
rect 35483 28577 35492 28611
rect 35440 28568 35492 28577
rect 36636 28568 36688 28620
rect 32220 28500 32272 28552
rect 28632 28364 28684 28416
rect 30656 28407 30708 28416
rect 30656 28373 30665 28407
rect 30665 28373 30699 28407
rect 30699 28373 30708 28407
rect 30656 28364 30708 28373
rect 35992 28407 36044 28416
rect 35992 28373 36001 28407
rect 36001 28373 36035 28407
rect 36035 28373 36044 28407
rect 35992 28364 36044 28373
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 34966 28262 35018 28314
rect 35030 28262 35082 28314
rect 35094 28262 35146 28314
rect 35158 28262 35210 28314
rect 27988 28203 28040 28212
rect 27988 28169 27997 28203
rect 27997 28169 28031 28203
rect 28031 28169 28040 28203
rect 27988 28160 28040 28169
rect 28448 28160 28500 28212
rect 29000 28160 29052 28212
rect 30472 28160 30524 28212
rect 32220 28203 32272 28212
rect 32220 28169 32229 28203
rect 32229 28169 32263 28203
rect 32263 28169 32272 28203
rect 32220 28160 32272 28169
rect 32312 28203 32364 28212
rect 32312 28169 32321 28203
rect 32321 28169 32355 28203
rect 32355 28169 32364 28203
rect 32312 28160 32364 28169
rect 35256 28160 35308 28212
rect 28172 28067 28224 28076
rect 28172 28033 28181 28067
rect 28181 28033 28215 28067
rect 28215 28033 28224 28067
rect 28172 28024 28224 28033
rect 29000 28024 29052 28076
rect 29828 28067 29880 28076
rect 29828 28033 29837 28067
rect 29837 28033 29871 28067
rect 29871 28033 29880 28067
rect 29828 28024 29880 28033
rect 32864 28067 32916 28076
rect 32864 28033 32873 28067
rect 32873 28033 32907 28067
rect 32907 28033 32916 28067
rect 32864 28024 32916 28033
rect 30656 27956 30708 28008
rect 32220 27956 32272 28008
rect 36636 27999 36688 28008
rect 31668 27888 31720 27940
rect 36636 27965 36645 27999
rect 36645 27965 36679 27999
rect 36679 27965 36688 27999
rect 36636 27956 36688 27965
rect 35440 27820 35492 27872
rect 35808 27820 35860 27872
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 29828 27616 29880 27668
rect 31668 27616 31720 27668
rect 34244 27548 34296 27600
rect 23112 27523 23164 27532
rect 23112 27489 23121 27523
rect 23121 27489 23155 27523
rect 23155 27489 23164 27523
rect 23112 27480 23164 27489
rect 24308 27480 24360 27532
rect 28908 27523 28960 27532
rect 28908 27489 28917 27523
rect 28917 27489 28951 27523
rect 28951 27489 28960 27523
rect 28908 27480 28960 27489
rect 31852 27480 31904 27532
rect 29000 27455 29052 27464
rect 29000 27421 29009 27455
rect 29009 27421 29043 27455
rect 29043 27421 29052 27455
rect 29000 27412 29052 27421
rect 30104 27455 30156 27464
rect 30104 27421 30113 27455
rect 30113 27421 30147 27455
rect 30147 27421 30156 27455
rect 30104 27412 30156 27421
rect 31300 27412 31352 27464
rect 32588 27455 32640 27464
rect 32588 27421 32597 27455
rect 32597 27421 32631 27455
rect 32631 27421 32640 27455
rect 32588 27412 32640 27421
rect 33876 27455 33928 27464
rect 29552 27387 29604 27396
rect 29552 27353 29561 27387
rect 29561 27353 29595 27387
rect 29595 27353 29604 27387
rect 29552 27344 29604 27353
rect 32036 27344 32088 27396
rect 33876 27421 33885 27455
rect 33885 27421 33919 27455
rect 33919 27421 33928 27455
rect 33876 27412 33928 27421
rect 35716 27412 35768 27464
rect 21916 27319 21968 27328
rect 21916 27285 21925 27319
rect 21925 27285 21959 27319
rect 21959 27285 21968 27319
rect 21916 27276 21968 27285
rect 23296 27319 23348 27328
rect 23296 27285 23305 27319
rect 23305 27285 23339 27319
rect 23339 27285 23348 27319
rect 23296 27276 23348 27285
rect 24768 27276 24820 27328
rect 28816 27276 28868 27328
rect 35256 27319 35308 27328
rect 35256 27285 35265 27319
rect 35265 27285 35299 27319
rect 35299 27285 35308 27319
rect 35256 27276 35308 27285
rect 35532 27276 35584 27328
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 34966 27174 35018 27226
rect 35030 27174 35082 27226
rect 35094 27174 35146 27226
rect 35158 27174 35210 27226
rect 28724 27072 28776 27124
rect 31300 27115 31352 27124
rect 21824 26936 21876 26988
rect 31300 27081 31309 27115
rect 31309 27081 31343 27115
rect 31343 27081 31352 27115
rect 31300 27072 31352 27081
rect 32864 27072 32916 27124
rect 35900 27072 35952 27124
rect 29184 26936 29236 26988
rect 21916 26868 21968 26920
rect 24676 26911 24728 26920
rect 24676 26877 24685 26911
rect 24685 26877 24719 26911
rect 24719 26877 24728 26911
rect 24676 26868 24728 26877
rect 29552 26911 29604 26920
rect 25320 26800 25372 26852
rect 27896 26843 27948 26852
rect 27896 26809 27905 26843
rect 27905 26809 27939 26843
rect 27939 26809 27948 26843
rect 27896 26800 27948 26809
rect 29552 26877 29586 26911
rect 29586 26877 29604 26911
rect 29552 26868 29604 26877
rect 32036 26911 32088 26920
rect 32036 26877 32070 26911
rect 32070 26877 32088 26911
rect 32036 26868 32088 26877
rect 32404 26800 32456 26852
rect 33876 26800 33928 26852
rect 35532 26868 35584 26920
rect 35624 26800 35676 26852
rect 22008 26732 22060 26784
rect 22284 26775 22336 26784
rect 22284 26741 22293 26775
rect 22293 26741 22327 26775
rect 22327 26741 22336 26775
rect 22284 26732 22336 26741
rect 22744 26732 22796 26784
rect 23112 26775 23164 26784
rect 23112 26741 23121 26775
rect 23121 26741 23155 26775
rect 23155 26741 23164 26775
rect 23112 26732 23164 26741
rect 26056 26775 26108 26784
rect 26056 26741 26065 26775
rect 26065 26741 26099 26775
rect 26099 26741 26108 26775
rect 26056 26732 26108 26741
rect 27528 26732 27580 26784
rect 28724 26775 28776 26784
rect 28724 26741 28733 26775
rect 28733 26741 28767 26775
rect 28767 26741 28776 26775
rect 28724 26732 28776 26741
rect 29184 26732 29236 26784
rect 30656 26775 30708 26784
rect 30656 26741 30665 26775
rect 30665 26741 30699 26775
rect 30699 26741 30708 26775
rect 30656 26732 30708 26741
rect 34244 26775 34296 26784
rect 34244 26741 34253 26775
rect 34253 26741 34287 26775
rect 34287 26741 34296 26775
rect 34244 26732 34296 26741
rect 34612 26775 34664 26784
rect 34612 26741 34621 26775
rect 34621 26741 34655 26775
rect 34655 26741 34664 26775
rect 34612 26732 34664 26741
rect 35808 26732 35860 26784
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 21916 26528 21968 26580
rect 27896 26571 27948 26580
rect 22284 26460 22336 26512
rect 27896 26537 27905 26571
rect 27905 26537 27939 26571
rect 27939 26537 27948 26571
rect 27896 26528 27948 26537
rect 29552 26528 29604 26580
rect 33876 26528 33928 26580
rect 35532 26528 35584 26580
rect 20904 26324 20956 26376
rect 24676 26392 24728 26444
rect 26516 26435 26568 26444
rect 26516 26401 26525 26435
rect 26525 26401 26559 26435
rect 26559 26401 26568 26435
rect 26516 26392 26568 26401
rect 26792 26435 26844 26444
rect 26792 26401 26826 26435
rect 26826 26401 26844 26435
rect 26792 26392 26844 26401
rect 29368 26460 29420 26512
rect 32036 26460 32088 26512
rect 32864 26460 32916 26512
rect 35256 26460 35308 26512
rect 28448 26392 28500 26444
rect 32404 26367 32456 26376
rect 32404 26333 32413 26367
rect 32413 26333 32447 26367
rect 32447 26333 32456 26367
rect 32404 26324 32456 26333
rect 34612 26324 34664 26376
rect 21180 26231 21232 26240
rect 21180 26197 21189 26231
rect 21189 26197 21223 26231
rect 21223 26197 21232 26231
rect 21180 26188 21232 26197
rect 24584 26188 24636 26240
rect 27436 26188 27488 26240
rect 28908 26256 28960 26308
rect 31852 26299 31904 26308
rect 31852 26265 31861 26299
rect 31861 26265 31895 26299
rect 31895 26265 31904 26299
rect 31852 26256 31904 26265
rect 33416 26256 33468 26308
rect 34244 26256 34296 26308
rect 34704 26231 34756 26240
rect 34704 26197 34713 26231
rect 34713 26197 34747 26231
rect 34747 26197 34756 26231
rect 34704 26188 34756 26197
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 34966 26086 35018 26138
rect 35030 26086 35082 26138
rect 35094 26086 35146 26138
rect 35158 26086 35210 26138
rect 20904 25984 20956 26036
rect 22284 26027 22336 26036
rect 22284 25993 22293 26027
rect 22293 25993 22327 26027
rect 22327 25993 22336 26027
rect 22284 25984 22336 25993
rect 25320 26027 25372 26036
rect 25320 25993 25329 26027
rect 25329 25993 25363 26027
rect 25363 25993 25372 26027
rect 25320 25984 25372 25993
rect 27896 25984 27948 26036
rect 29000 25984 29052 26036
rect 32036 25984 32088 26036
rect 34796 25916 34848 25968
rect 36084 25916 36136 25968
rect 33876 25891 33928 25900
rect 33876 25857 33885 25891
rect 33885 25857 33919 25891
rect 33919 25857 33928 25891
rect 33876 25848 33928 25857
rect 35256 25848 35308 25900
rect 24032 25780 24084 25832
rect 24676 25780 24728 25832
rect 26516 25780 26568 25832
rect 29276 25823 29328 25832
rect 29276 25789 29285 25823
rect 29285 25789 29319 25823
rect 29319 25789 29328 25823
rect 29276 25780 29328 25789
rect 30380 25823 30432 25832
rect 30380 25789 30389 25823
rect 30389 25789 30423 25823
rect 30423 25789 30432 25823
rect 30380 25780 30432 25789
rect 30656 25823 30708 25832
rect 21180 25755 21232 25764
rect 21180 25721 21214 25755
rect 21214 25721 21232 25755
rect 21180 25712 21232 25721
rect 21548 25712 21600 25764
rect 24584 25712 24636 25764
rect 26056 25712 26108 25764
rect 30288 25712 30340 25764
rect 30656 25789 30690 25823
rect 30690 25789 30708 25823
rect 30656 25780 30708 25789
rect 32404 25780 32456 25832
rect 34612 25823 34664 25832
rect 34612 25789 34621 25823
rect 34621 25789 34655 25823
rect 34655 25789 34664 25823
rect 34612 25780 34664 25789
rect 34704 25780 34756 25832
rect 27804 25687 27856 25696
rect 27804 25653 27813 25687
rect 27813 25653 27847 25687
rect 27847 25653 27856 25687
rect 27804 25644 27856 25653
rect 29184 25644 29236 25696
rect 30380 25644 30432 25696
rect 32128 25644 32180 25696
rect 33232 25687 33284 25696
rect 33232 25653 33241 25687
rect 33241 25653 33275 25687
rect 33275 25653 33284 25687
rect 33232 25644 33284 25653
rect 33692 25687 33744 25696
rect 33692 25653 33701 25687
rect 33701 25653 33735 25687
rect 33735 25653 33744 25687
rect 33692 25644 33744 25653
rect 35164 25644 35216 25696
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 24032 25483 24084 25492
rect 24032 25449 24041 25483
rect 24041 25449 24075 25483
rect 24075 25449 24084 25483
rect 24032 25440 24084 25449
rect 24676 25440 24728 25492
rect 25320 25440 25372 25492
rect 26056 25440 26108 25492
rect 27436 25440 27488 25492
rect 29276 25483 29328 25492
rect 29276 25449 29285 25483
rect 29285 25449 29319 25483
rect 29319 25449 29328 25483
rect 29276 25440 29328 25449
rect 29552 25483 29604 25492
rect 29552 25449 29561 25483
rect 29561 25449 29595 25483
rect 29595 25449 29604 25483
rect 29552 25440 29604 25449
rect 30104 25440 30156 25492
rect 32680 25483 32732 25492
rect 32680 25449 32689 25483
rect 32689 25449 32723 25483
rect 32723 25449 32732 25483
rect 32680 25440 32732 25449
rect 33692 25483 33744 25492
rect 33692 25449 33701 25483
rect 33701 25449 33735 25483
rect 33735 25449 33744 25483
rect 33692 25440 33744 25449
rect 24584 25415 24636 25424
rect 24584 25381 24593 25415
rect 24593 25381 24627 25415
rect 24627 25381 24636 25415
rect 24584 25372 24636 25381
rect 25504 25372 25556 25424
rect 29000 25372 29052 25424
rect 30472 25372 30524 25424
rect 32864 25372 32916 25424
rect 20904 25347 20956 25356
rect 20904 25313 20913 25347
rect 20913 25313 20947 25347
rect 20947 25313 20956 25347
rect 20904 25304 20956 25313
rect 21180 25347 21232 25356
rect 21180 25313 21214 25347
rect 21214 25313 21232 25347
rect 21180 25304 21232 25313
rect 26700 25304 26752 25356
rect 28264 25347 28316 25356
rect 28264 25313 28273 25347
rect 28273 25313 28307 25347
rect 28307 25313 28316 25347
rect 28264 25304 28316 25313
rect 33048 25347 33100 25356
rect 33048 25313 33057 25347
rect 33057 25313 33091 25347
rect 33091 25313 33100 25347
rect 33048 25304 33100 25313
rect 24124 25236 24176 25288
rect 25596 25236 25648 25288
rect 28356 25279 28408 25288
rect 28356 25245 28365 25279
rect 28365 25245 28399 25279
rect 28399 25245 28408 25279
rect 28356 25236 28408 25245
rect 28724 25236 28776 25288
rect 30288 25236 30340 25288
rect 32680 25236 32732 25288
rect 33324 25279 33376 25288
rect 33324 25245 33333 25279
rect 33333 25245 33367 25279
rect 33367 25245 33376 25279
rect 33324 25236 33376 25245
rect 34060 25236 34112 25288
rect 34612 25236 34664 25288
rect 34888 25279 34940 25288
rect 34888 25245 34897 25279
rect 34897 25245 34931 25279
rect 34931 25245 34940 25279
rect 35164 25279 35216 25288
rect 34888 25236 34940 25245
rect 35164 25245 35173 25279
rect 35173 25245 35207 25279
rect 35207 25245 35216 25279
rect 35164 25236 35216 25245
rect 35624 25236 35676 25288
rect 36268 25279 36320 25288
rect 36268 25245 36277 25279
rect 36277 25245 36311 25279
rect 36311 25245 36320 25279
rect 36268 25236 36320 25245
rect 31944 25211 31996 25220
rect 31944 25177 31953 25211
rect 31953 25177 31987 25211
rect 31987 25177 31996 25211
rect 31944 25168 31996 25177
rect 20628 25143 20680 25152
rect 20628 25109 20637 25143
rect 20637 25109 20671 25143
rect 20671 25109 20680 25143
rect 20628 25100 20680 25109
rect 21548 25100 21600 25152
rect 24768 25100 24820 25152
rect 26240 25100 26292 25152
rect 26792 25100 26844 25152
rect 27804 25100 27856 25152
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 34966 24998 35018 25050
rect 35030 24998 35082 25050
rect 35094 24998 35146 25050
rect 35158 24998 35210 25050
rect 20904 24896 20956 24948
rect 24676 24939 24728 24948
rect 24676 24905 24685 24939
rect 24685 24905 24719 24939
rect 24719 24905 24728 24939
rect 24676 24896 24728 24905
rect 26700 24896 26752 24948
rect 28356 24896 28408 24948
rect 30104 24896 30156 24948
rect 24584 24828 24636 24880
rect 30288 24828 30340 24880
rect 20536 24803 20588 24812
rect 20536 24769 20545 24803
rect 20545 24769 20579 24803
rect 20579 24769 20588 24803
rect 20536 24760 20588 24769
rect 25596 24803 25648 24812
rect 25596 24769 25605 24803
rect 25605 24769 25639 24803
rect 25639 24769 25648 24803
rect 25596 24760 25648 24769
rect 26424 24803 26476 24812
rect 26424 24769 26433 24803
rect 26433 24769 26467 24803
rect 26467 24769 26476 24803
rect 27160 24803 27212 24812
rect 26424 24760 26476 24769
rect 20720 24624 20772 24676
rect 24860 24692 24912 24744
rect 26884 24692 26936 24744
rect 27160 24769 27169 24803
rect 27169 24769 27203 24803
rect 27203 24769 27212 24803
rect 27160 24760 27212 24769
rect 34612 24896 34664 24948
rect 34796 24896 34848 24948
rect 33232 24828 33284 24880
rect 32312 24803 32364 24812
rect 32312 24769 32321 24803
rect 32321 24769 32355 24803
rect 32355 24769 32364 24803
rect 32588 24803 32640 24812
rect 32312 24760 32364 24769
rect 32588 24769 32597 24803
rect 32597 24769 32631 24803
rect 32631 24769 32640 24803
rect 32588 24760 32640 24769
rect 35900 24803 35952 24812
rect 26148 24624 26200 24676
rect 20260 24556 20312 24608
rect 21916 24599 21968 24608
rect 21916 24565 21925 24599
rect 21925 24565 21959 24599
rect 21959 24565 21968 24599
rect 21916 24556 21968 24565
rect 23480 24599 23532 24608
rect 23480 24565 23489 24599
rect 23489 24565 23523 24599
rect 23523 24565 23532 24599
rect 23480 24556 23532 24565
rect 23848 24599 23900 24608
rect 23848 24565 23857 24599
rect 23857 24565 23891 24599
rect 23891 24565 23900 24599
rect 23848 24556 23900 24565
rect 25044 24599 25096 24608
rect 25044 24565 25053 24599
rect 25053 24565 25087 24599
rect 25087 24565 25096 24599
rect 25044 24556 25096 24565
rect 25412 24599 25464 24608
rect 25412 24565 25421 24599
rect 25421 24565 25455 24599
rect 25455 24565 25464 24599
rect 25412 24556 25464 24565
rect 25504 24599 25556 24608
rect 25504 24565 25513 24599
rect 25513 24565 25547 24599
rect 25547 24565 25556 24599
rect 28264 24624 28316 24676
rect 30932 24624 30984 24676
rect 35900 24769 35909 24803
rect 35909 24769 35943 24803
rect 35943 24769 35952 24803
rect 35900 24760 35952 24769
rect 34980 24624 35032 24676
rect 35716 24624 35768 24676
rect 25504 24556 25556 24565
rect 26884 24556 26936 24608
rect 28724 24599 28776 24608
rect 28724 24565 28733 24599
rect 28733 24565 28767 24599
rect 28767 24565 28776 24599
rect 28724 24556 28776 24565
rect 30380 24599 30432 24608
rect 30380 24565 30389 24599
rect 30389 24565 30423 24599
rect 30423 24565 30432 24599
rect 30380 24556 30432 24565
rect 32680 24556 32732 24608
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 20536 24395 20588 24404
rect 20536 24361 20545 24395
rect 20545 24361 20579 24395
rect 20579 24361 20588 24395
rect 20536 24352 20588 24361
rect 22744 24395 22796 24404
rect 22744 24361 22753 24395
rect 22753 24361 22787 24395
rect 22787 24361 22796 24395
rect 22744 24352 22796 24361
rect 24308 24395 24360 24404
rect 24308 24361 24317 24395
rect 24317 24361 24351 24395
rect 24351 24361 24360 24395
rect 24308 24352 24360 24361
rect 25044 24352 25096 24404
rect 25412 24395 25464 24404
rect 25412 24361 25421 24395
rect 25421 24361 25455 24395
rect 25455 24361 25464 24395
rect 25412 24352 25464 24361
rect 26148 24352 26200 24404
rect 27160 24352 27212 24404
rect 28724 24352 28776 24404
rect 30380 24352 30432 24404
rect 32312 24352 32364 24404
rect 33048 24395 33100 24404
rect 33048 24361 33057 24395
rect 33057 24361 33091 24395
rect 33091 24361 33100 24395
rect 33048 24352 33100 24361
rect 33324 24352 33376 24404
rect 34980 24395 35032 24404
rect 34980 24361 34989 24395
rect 34989 24361 35023 24395
rect 35023 24361 35032 24395
rect 34980 24352 35032 24361
rect 35348 24395 35400 24404
rect 35348 24361 35357 24395
rect 35357 24361 35391 24395
rect 35391 24361 35400 24395
rect 35348 24352 35400 24361
rect 20260 24284 20312 24336
rect 21180 24284 21232 24336
rect 21916 24284 21968 24336
rect 22100 24284 22152 24336
rect 23112 24327 23164 24336
rect 23112 24293 23121 24327
rect 23121 24293 23155 24327
rect 23155 24293 23164 24327
rect 23112 24284 23164 24293
rect 24768 24327 24820 24336
rect 24768 24293 24777 24327
rect 24777 24293 24811 24327
rect 24811 24293 24820 24327
rect 24768 24284 24820 24293
rect 28264 24284 28316 24336
rect 28632 24284 28684 24336
rect 30472 24327 30524 24336
rect 30472 24293 30481 24327
rect 30481 24293 30515 24327
rect 30515 24293 30524 24327
rect 30472 24284 30524 24293
rect 21548 24259 21600 24268
rect 21548 24225 21557 24259
rect 21557 24225 21591 24259
rect 21591 24225 21600 24259
rect 21548 24216 21600 24225
rect 27528 24216 27580 24268
rect 28448 24259 28500 24268
rect 28448 24225 28457 24259
rect 28457 24225 28491 24259
rect 28491 24225 28500 24259
rect 28448 24216 28500 24225
rect 35716 24259 35768 24268
rect 35716 24225 35725 24259
rect 35725 24225 35759 24259
rect 35759 24225 35768 24259
rect 35716 24216 35768 24225
rect 21824 24191 21876 24200
rect 21824 24157 21833 24191
rect 21833 24157 21867 24191
rect 21867 24157 21876 24191
rect 21824 24148 21876 24157
rect 22836 24148 22888 24200
rect 25412 24148 25464 24200
rect 35808 24191 35860 24200
rect 35808 24157 35817 24191
rect 35817 24157 35851 24191
rect 35851 24157 35860 24191
rect 35808 24148 35860 24157
rect 36268 24148 36320 24200
rect 22836 24012 22888 24064
rect 24124 24055 24176 24064
rect 24124 24021 24133 24055
rect 24133 24021 24167 24055
rect 24167 24021 24176 24055
rect 24124 24012 24176 24021
rect 29828 24055 29880 24064
rect 29828 24021 29837 24055
rect 29837 24021 29871 24055
rect 29871 24021 29880 24055
rect 29828 24012 29880 24021
rect 32680 24055 32732 24064
rect 32680 24021 32689 24055
rect 32689 24021 32723 24055
rect 32723 24021 32732 24055
rect 32680 24012 32732 24021
rect 34060 24055 34112 24064
rect 34060 24021 34069 24055
rect 34069 24021 34103 24055
rect 34103 24021 34112 24055
rect 34060 24012 34112 24021
rect 34612 24012 34664 24064
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 34966 23910 35018 23962
rect 35030 23910 35082 23962
rect 35094 23910 35146 23962
rect 35158 23910 35210 23962
rect 20260 23851 20312 23860
rect 20260 23817 20269 23851
rect 20269 23817 20303 23851
rect 20303 23817 20312 23851
rect 20260 23808 20312 23817
rect 20720 23851 20772 23860
rect 20720 23817 20729 23851
rect 20729 23817 20763 23851
rect 20763 23817 20772 23851
rect 20720 23808 20772 23817
rect 21548 23808 21600 23860
rect 22836 23851 22888 23860
rect 22836 23817 22845 23851
rect 22845 23817 22879 23851
rect 22879 23817 22888 23851
rect 22836 23808 22888 23817
rect 23112 23851 23164 23860
rect 23112 23817 23121 23851
rect 23121 23817 23155 23851
rect 23155 23817 23164 23851
rect 23112 23808 23164 23817
rect 24768 23808 24820 23860
rect 26148 23851 26200 23860
rect 24400 23783 24452 23792
rect 24400 23749 24409 23783
rect 24409 23749 24443 23783
rect 24443 23749 24452 23783
rect 24400 23740 24452 23749
rect 21824 23715 21876 23724
rect 21824 23681 21833 23715
rect 21833 23681 21867 23715
rect 21867 23681 21876 23715
rect 21824 23672 21876 23681
rect 26148 23817 26157 23851
rect 26157 23817 26191 23851
rect 26191 23817 26200 23851
rect 26148 23808 26200 23817
rect 26608 23851 26660 23860
rect 26608 23817 26617 23851
rect 26617 23817 26651 23851
rect 26651 23817 26660 23851
rect 26608 23808 26660 23817
rect 27528 23808 27580 23860
rect 28448 23808 28500 23860
rect 28264 23715 28316 23724
rect 28264 23681 28273 23715
rect 28273 23681 28307 23715
rect 28307 23681 28316 23715
rect 28264 23672 28316 23681
rect 35808 23808 35860 23860
rect 36176 23740 36228 23792
rect 29828 23715 29880 23724
rect 29828 23681 29837 23715
rect 29837 23681 29871 23715
rect 29871 23681 29880 23715
rect 29828 23672 29880 23681
rect 35624 23672 35676 23724
rect 20720 23604 20772 23656
rect 22100 23604 22152 23656
rect 23848 23604 23900 23656
rect 26608 23604 26660 23656
rect 26976 23604 27028 23656
rect 27620 23604 27672 23656
rect 34244 23604 34296 23656
rect 35716 23604 35768 23656
rect 24860 23579 24912 23588
rect 24860 23545 24869 23579
rect 24869 23545 24903 23579
rect 24903 23545 24912 23579
rect 24860 23536 24912 23545
rect 34796 23536 34848 23588
rect 19984 23511 20036 23520
rect 19984 23477 19993 23511
rect 19993 23477 20027 23511
rect 20027 23477 20036 23511
rect 19984 23468 20036 23477
rect 20996 23511 21048 23520
rect 20996 23477 21005 23511
rect 21005 23477 21039 23511
rect 21039 23477 21048 23511
rect 20996 23468 21048 23477
rect 21180 23511 21232 23520
rect 21180 23477 21189 23511
rect 21189 23477 21223 23511
rect 21223 23477 21232 23511
rect 21180 23468 21232 23477
rect 25412 23511 25464 23520
rect 25412 23477 25421 23511
rect 25421 23477 25455 23511
rect 25455 23477 25464 23511
rect 25412 23468 25464 23477
rect 28172 23468 28224 23520
rect 34612 23468 34664 23520
rect 35532 23468 35584 23520
rect 36268 23511 36320 23520
rect 36268 23477 36277 23511
rect 36277 23477 36311 23511
rect 36311 23477 36320 23511
rect 36268 23468 36320 23477
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 19984 23264 20036 23316
rect 21824 23264 21876 23316
rect 22100 23264 22152 23316
rect 23388 23307 23440 23316
rect 23388 23273 23397 23307
rect 23397 23273 23431 23307
rect 23431 23273 23440 23307
rect 23388 23264 23440 23273
rect 23756 23307 23808 23316
rect 23756 23273 23765 23307
rect 23765 23273 23799 23307
rect 23799 23273 23808 23307
rect 23756 23264 23808 23273
rect 23848 23264 23900 23316
rect 24860 23264 24912 23316
rect 26976 23307 27028 23316
rect 26976 23273 26985 23307
rect 26985 23273 27019 23307
rect 27019 23273 27028 23307
rect 26976 23264 27028 23273
rect 28264 23264 28316 23316
rect 34244 23264 34296 23316
rect 35624 23264 35676 23316
rect 36728 23264 36780 23316
rect 28908 23196 28960 23248
rect 20628 23128 20680 23180
rect 20996 23128 21048 23180
rect 24952 23171 25004 23180
rect 24952 23137 24961 23171
rect 24961 23137 24995 23171
rect 24995 23137 25004 23171
rect 24952 23128 25004 23137
rect 27896 23171 27948 23180
rect 27896 23137 27905 23171
rect 27905 23137 27939 23171
rect 27939 23137 27948 23171
rect 27896 23128 27948 23137
rect 28356 23128 28408 23180
rect 29828 23128 29880 23180
rect 35808 23128 35860 23180
rect 20904 23103 20956 23112
rect 20904 23069 20913 23103
rect 20913 23069 20947 23103
rect 20947 23069 20956 23103
rect 20904 23060 20956 23069
rect 23848 23103 23900 23112
rect 23848 23069 23857 23103
rect 23857 23069 23891 23103
rect 23891 23069 23900 23103
rect 23848 23060 23900 23069
rect 24032 23103 24084 23112
rect 24032 23069 24041 23103
rect 24041 23069 24075 23103
rect 24075 23069 24084 23103
rect 24032 23060 24084 23069
rect 25044 23060 25096 23112
rect 28448 23060 28500 23112
rect 28172 22992 28224 23044
rect 28080 22967 28132 22976
rect 28080 22933 28089 22967
rect 28089 22933 28123 22967
rect 28123 22933 28132 22967
rect 28080 22924 28132 22933
rect 29368 22924 29420 22976
rect 30656 22924 30708 22976
rect 34796 22924 34848 22976
rect 35348 22924 35400 22976
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 34966 22822 35018 22874
rect 35030 22822 35082 22874
rect 35094 22822 35146 22874
rect 35158 22822 35210 22874
rect 20904 22763 20956 22772
rect 20904 22729 20913 22763
rect 20913 22729 20947 22763
rect 20947 22729 20956 22763
rect 20904 22720 20956 22729
rect 21548 22763 21600 22772
rect 21548 22729 21557 22763
rect 21557 22729 21591 22763
rect 21591 22729 21600 22763
rect 21548 22720 21600 22729
rect 23848 22720 23900 22772
rect 25412 22763 25464 22772
rect 24952 22652 25004 22704
rect 21824 22584 21876 22636
rect 24032 22584 24084 22636
rect 25412 22729 25421 22763
rect 25421 22729 25455 22763
rect 25455 22729 25464 22763
rect 25412 22720 25464 22729
rect 27896 22763 27948 22772
rect 27896 22729 27905 22763
rect 27905 22729 27939 22763
rect 27939 22729 27948 22763
rect 27896 22720 27948 22729
rect 28356 22763 28408 22772
rect 28356 22729 28365 22763
rect 28365 22729 28399 22763
rect 28399 22729 28408 22763
rect 28356 22720 28408 22729
rect 28448 22720 28500 22772
rect 28632 22763 28684 22772
rect 28632 22729 28641 22763
rect 28641 22729 28675 22763
rect 28675 22729 28684 22763
rect 28632 22720 28684 22729
rect 25872 22627 25924 22636
rect 23664 22516 23716 22568
rect 25872 22593 25881 22627
rect 25881 22593 25915 22627
rect 25915 22593 25924 22627
rect 25872 22584 25924 22593
rect 26240 22584 26292 22636
rect 27528 22584 27580 22636
rect 32956 22720 33008 22772
rect 36268 22720 36320 22772
rect 26976 22516 27028 22568
rect 29368 22516 29420 22568
rect 32128 22516 32180 22568
rect 35164 22516 35216 22568
rect 35348 22559 35400 22568
rect 35348 22525 35357 22559
rect 35357 22525 35391 22559
rect 35391 22525 35400 22559
rect 35348 22516 35400 22525
rect 35624 22559 35676 22568
rect 35624 22525 35658 22559
rect 35658 22525 35676 22559
rect 35624 22516 35676 22525
rect 27160 22448 27212 22500
rect 32956 22448 33008 22500
rect 20628 22423 20680 22432
rect 20628 22389 20637 22423
rect 20637 22389 20671 22423
rect 20671 22389 20680 22423
rect 20628 22380 20680 22389
rect 21364 22423 21416 22432
rect 21364 22389 21373 22423
rect 21373 22389 21407 22423
rect 21407 22389 21416 22423
rect 21364 22380 21416 22389
rect 21916 22423 21968 22432
rect 21916 22389 21925 22423
rect 21925 22389 21959 22423
rect 21959 22389 21968 22423
rect 21916 22380 21968 22389
rect 23112 22423 23164 22432
rect 23112 22389 23121 22423
rect 23121 22389 23155 22423
rect 23155 22389 23164 22423
rect 23112 22380 23164 22389
rect 23756 22380 23808 22432
rect 26884 22423 26936 22432
rect 26884 22389 26893 22423
rect 26893 22389 26927 22423
rect 26927 22389 26936 22423
rect 26884 22380 26936 22389
rect 30472 22380 30524 22432
rect 32128 22423 32180 22432
rect 32128 22389 32137 22423
rect 32137 22389 32171 22423
rect 32171 22389 32180 22423
rect 32128 22380 32180 22389
rect 33600 22423 33652 22432
rect 33600 22389 33609 22423
rect 33609 22389 33643 22423
rect 33643 22389 33652 22423
rect 33600 22380 33652 22389
rect 34244 22380 34296 22432
rect 35164 22423 35216 22432
rect 35164 22389 35173 22423
rect 35173 22389 35207 22423
rect 35207 22389 35216 22423
rect 35164 22380 35216 22389
rect 35808 22380 35860 22432
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 20628 22176 20680 22228
rect 23112 22176 23164 22228
rect 21824 22108 21876 22160
rect 20720 22040 20772 22092
rect 21916 22040 21968 22092
rect 24032 22176 24084 22228
rect 24952 22219 25004 22228
rect 24952 22185 24961 22219
rect 24961 22185 24995 22219
rect 24995 22185 25004 22219
rect 24952 22176 25004 22185
rect 27436 22176 27488 22228
rect 34336 22176 34388 22228
rect 34704 22176 34756 22228
rect 35532 22176 35584 22228
rect 35716 22176 35768 22228
rect 36728 22219 36780 22228
rect 36728 22185 36737 22219
rect 36737 22185 36771 22219
rect 36771 22185 36780 22219
rect 36728 22176 36780 22185
rect 23756 22151 23808 22160
rect 23756 22117 23765 22151
rect 23765 22117 23799 22151
rect 23799 22117 23808 22151
rect 23756 22108 23808 22117
rect 24768 22108 24820 22160
rect 23204 22040 23256 22092
rect 25320 22083 25372 22092
rect 20904 22015 20956 22024
rect 20904 21981 20913 22015
rect 20913 21981 20947 22015
rect 20947 21981 20956 22015
rect 20904 21972 20956 21981
rect 25320 22049 25329 22083
rect 25329 22049 25363 22083
rect 25363 22049 25372 22083
rect 25320 22040 25372 22049
rect 25780 22040 25832 22092
rect 27160 22040 27212 22092
rect 24216 21972 24268 22024
rect 26792 22015 26844 22024
rect 26792 21981 26801 22015
rect 26801 21981 26835 22015
rect 26835 21981 26844 22015
rect 26792 21972 26844 21981
rect 27252 22015 27304 22024
rect 27252 21981 27261 22015
rect 27261 21981 27295 22015
rect 27295 21981 27304 22015
rect 27252 21972 27304 21981
rect 29552 22040 29604 22092
rect 31760 22040 31812 22092
rect 34428 22040 34480 22092
rect 35808 22040 35860 22092
rect 36268 22040 36320 22092
rect 27712 21972 27764 22024
rect 28172 21972 28224 22024
rect 30012 21972 30064 22024
rect 30288 21972 30340 22024
rect 30656 21972 30708 22024
rect 32588 22015 32640 22024
rect 32588 21981 32597 22015
rect 32597 21981 32631 22015
rect 32631 21981 32640 22015
rect 32588 21972 32640 21981
rect 29276 21904 29328 21956
rect 30932 21904 30984 21956
rect 32312 21904 32364 21956
rect 34796 22015 34848 22024
rect 34796 21981 34805 22015
rect 34805 21981 34839 22015
rect 34839 21981 34848 22015
rect 34796 21972 34848 21981
rect 35900 21972 35952 22024
rect 24676 21836 24728 21888
rect 26516 21836 26568 21888
rect 29552 21879 29604 21888
rect 29552 21845 29561 21879
rect 29561 21845 29595 21879
rect 29595 21845 29604 21879
rect 29552 21836 29604 21845
rect 29736 21879 29788 21888
rect 29736 21845 29745 21879
rect 29745 21845 29779 21879
rect 29779 21845 29788 21879
rect 29736 21836 29788 21845
rect 32956 21836 33008 21888
rect 33140 21836 33192 21888
rect 34060 21904 34112 21956
rect 33876 21836 33928 21888
rect 34796 21836 34848 21888
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 34966 21734 35018 21786
rect 35030 21734 35082 21786
rect 35094 21734 35146 21786
rect 35158 21734 35210 21786
rect 20904 21675 20956 21684
rect 20904 21641 20913 21675
rect 20913 21641 20947 21675
rect 20947 21641 20956 21675
rect 20904 21632 20956 21641
rect 21916 21632 21968 21684
rect 23664 21675 23716 21684
rect 23664 21641 23673 21675
rect 23673 21641 23707 21675
rect 23707 21641 23716 21675
rect 23664 21632 23716 21641
rect 24768 21632 24820 21684
rect 25320 21632 25372 21684
rect 27620 21675 27672 21684
rect 27620 21641 27629 21675
rect 27629 21641 27663 21675
rect 27663 21641 27672 21675
rect 27620 21632 27672 21641
rect 28080 21632 28132 21684
rect 29552 21632 29604 21684
rect 31760 21675 31812 21684
rect 31760 21641 31769 21675
rect 31769 21641 31803 21675
rect 31803 21641 31812 21675
rect 34336 21675 34388 21684
rect 31760 21632 31812 21641
rect 34336 21641 34345 21675
rect 34345 21641 34379 21675
rect 34379 21641 34388 21675
rect 34336 21632 34388 21641
rect 36268 21675 36320 21684
rect 36268 21641 36277 21675
rect 36277 21641 36311 21675
rect 36311 21641 36320 21675
rect 36268 21632 36320 21641
rect 24216 21539 24268 21548
rect 24216 21505 24225 21539
rect 24225 21505 24259 21539
rect 24259 21505 24268 21539
rect 24216 21496 24268 21505
rect 29276 21539 29328 21548
rect 29276 21505 29285 21539
rect 29285 21505 29319 21539
rect 29319 21505 29328 21539
rect 29276 21496 29328 21505
rect 29552 21496 29604 21548
rect 30012 21539 30064 21548
rect 30012 21505 30021 21539
rect 30021 21505 30055 21539
rect 30055 21505 30064 21539
rect 30012 21496 30064 21505
rect 32128 21496 32180 21548
rect 26332 21428 26384 21480
rect 31944 21428 31996 21480
rect 33232 21428 33284 21480
rect 33600 21428 33652 21480
rect 34244 21428 34296 21480
rect 34888 21471 34940 21480
rect 34888 21437 34897 21471
rect 34897 21437 34931 21471
rect 34931 21437 34940 21471
rect 34888 21428 34940 21437
rect 35624 21428 35676 21480
rect 36176 21428 36228 21480
rect 21364 21360 21416 21412
rect 22284 21360 22336 21412
rect 23940 21360 23992 21412
rect 24768 21360 24820 21412
rect 26516 21403 26568 21412
rect 26516 21369 26550 21403
rect 26550 21369 26568 21403
rect 26516 21360 26568 21369
rect 27252 21360 27304 21412
rect 32128 21403 32180 21412
rect 32128 21369 32137 21403
rect 32137 21369 32171 21403
rect 32171 21369 32180 21403
rect 32128 21360 32180 21369
rect 35348 21360 35400 21412
rect 23664 21292 23716 21344
rect 24124 21335 24176 21344
rect 24124 21301 24133 21335
rect 24133 21301 24167 21335
rect 24167 21301 24176 21335
rect 24124 21292 24176 21301
rect 24676 21335 24728 21344
rect 24676 21301 24685 21335
rect 24685 21301 24719 21335
rect 24719 21301 24728 21335
rect 24676 21292 24728 21301
rect 25228 21335 25280 21344
rect 25228 21301 25237 21335
rect 25237 21301 25271 21335
rect 25271 21301 25280 21335
rect 25228 21292 25280 21301
rect 26056 21335 26108 21344
rect 26056 21301 26065 21335
rect 26065 21301 26099 21335
rect 26099 21301 26108 21335
rect 26056 21292 26108 21301
rect 29092 21335 29144 21344
rect 29092 21301 29101 21335
rect 29101 21301 29135 21335
rect 29135 21301 29144 21335
rect 29092 21292 29144 21301
rect 29828 21292 29880 21344
rect 30380 21292 30432 21344
rect 32312 21292 32364 21344
rect 37372 21335 37424 21344
rect 37372 21301 37381 21335
rect 37381 21301 37415 21335
rect 37415 21301 37424 21335
rect 37372 21292 37424 21301
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 20720 21131 20772 21140
rect 20720 21097 20729 21131
rect 20729 21097 20763 21131
rect 20763 21097 20772 21131
rect 20720 21088 20772 21097
rect 22284 21131 22336 21140
rect 22284 21097 22293 21131
rect 22293 21097 22327 21131
rect 22327 21097 22336 21131
rect 22284 21088 22336 21097
rect 23204 21131 23256 21140
rect 23204 21097 23213 21131
rect 23213 21097 23247 21131
rect 23247 21097 23256 21131
rect 23204 21088 23256 21097
rect 24768 21131 24820 21140
rect 24768 21097 24777 21131
rect 24777 21097 24811 21131
rect 24811 21097 24820 21131
rect 24768 21088 24820 21097
rect 26792 21088 26844 21140
rect 26884 21088 26936 21140
rect 27712 21088 27764 21140
rect 29000 21088 29052 21140
rect 30656 21131 30708 21140
rect 30656 21097 30665 21131
rect 30665 21097 30699 21131
rect 30699 21097 30708 21131
rect 30656 21088 30708 21097
rect 31944 21131 31996 21140
rect 31944 21097 31953 21131
rect 31953 21097 31987 21131
rect 31987 21097 31996 21131
rect 31944 21088 31996 21097
rect 21364 21020 21416 21072
rect 23480 21020 23532 21072
rect 23664 21063 23716 21072
rect 23664 21029 23698 21063
rect 23698 21029 23716 21063
rect 23664 21020 23716 21029
rect 26148 21020 26200 21072
rect 26332 21063 26384 21072
rect 26332 21029 26341 21063
rect 26341 21029 26375 21063
rect 26375 21029 26384 21063
rect 26332 21020 26384 21029
rect 20904 20995 20956 21004
rect 20904 20961 20913 20995
rect 20913 20961 20947 20995
rect 20947 20961 20956 20995
rect 20904 20952 20956 20961
rect 25228 20952 25280 21004
rect 26700 20952 26752 21004
rect 29828 21020 29880 21072
rect 32772 21088 32824 21140
rect 34244 21088 34296 21140
rect 34428 21088 34480 21140
rect 34612 21088 34664 21140
rect 34888 21131 34940 21140
rect 34888 21097 34897 21131
rect 34897 21097 34931 21131
rect 34931 21097 34940 21131
rect 34888 21088 34940 21097
rect 35348 21131 35400 21140
rect 35348 21097 35357 21131
rect 35357 21097 35391 21131
rect 35391 21097 35400 21131
rect 35348 21088 35400 21097
rect 35808 21131 35860 21140
rect 35808 21097 35817 21131
rect 35817 21097 35851 21131
rect 35851 21097 35860 21131
rect 35808 21088 35860 21097
rect 28448 20952 28500 21004
rect 28632 20995 28684 21004
rect 28632 20961 28666 20995
rect 28666 20961 28684 20995
rect 28632 20952 28684 20961
rect 30932 20952 30984 21004
rect 33140 20952 33192 21004
rect 23296 20884 23348 20936
rect 27160 20927 27212 20936
rect 27160 20893 27169 20927
rect 27169 20893 27203 20927
rect 27203 20893 27212 20927
rect 27160 20884 27212 20893
rect 30288 20884 30340 20936
rect 32312 20927 32364 20936
rect 32312 20893 32321 20927
rect 32321 20893 32355 20927
rect 32355 20893 32364 20927
rect 32312 20884 32364 20893
rect 32404 20884 32456 20936
rect 32956 20927 33008 20936
rect 32956 20893 32965 20927
rect 32965 20893 32999 20927
rect 32999 20893 33008 20927
rect 32956 20884 33008 20893
rect 33324 20884 33376 20936
rect 35716 20884 35768 20936
rect 36268 20884 36320 20936
rect 27252 20816 27304 20868
rect 37464 20816 37516 20868
rect 29644 20748 29696 20800
rect 30380 20748 30432 20800
rect 36084 20748 36136 20800
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 34966 20646 35018 20698
rect 35030 20646 35082 20698
rect 35094 20646 35146 20698
rect 35158 20646 35210 20698
rect 20904 20587 20956 20596
rect 20904 20553 20913 20587
rect 20913 20553 20947 20587
rect 20947 20553 20956 20587
rect 20904 20544 20956 20553
rect 21364 20587 21416 20596
rect 21364 20553 21373 20587
rect 21373 20553 21407 20587
rect 21407 20553 21416 20587
rect 21364 20544 21416 20553
rect 23388 20544 23440 20596
rect 25872 20544 25924 20596
rect 27160 20544 27212 20596
rect 32588 20587 32640 20596
rect 32588 20553 32597 20587
rect 32597 20553 32631 20587
rect 32631 20553 32640 20587
rect 32588 20544 32640 20553
rect 33140 20544 33192 20596
rect 34612 20587 34664 20596
rect 34612 20553 34621 20587
rect 34621 20553 34655 20587
rect 34655 20553 34664 20587
rect 34612 20544 34664 20553
rect 35900 20587 35952 20596
rect 35900 20553 35909 20587
rect 35909 20553 35943 20587
rect 35943 20553 35952 20587
rect 35900 20544 35952 20553
rect 36268 20587 36320 20596
rect 36268 20553 36277 20587
rect 36277 20553 36311 20587
rect 36311 20553 36320 20587
rect 36268 20544 36320 20553
rect 22468 20476 22520 20528
rect 29368 20519 29420 20528
rect 29368 20485 29377 20519
rect 29377 20485 29411 20519
rect 29411 20485 29420 20519
rect 29368 20476 29420 20485
rect 26148 20451 26200 20460
rect 23940 20383 23992 20392
rect 23940 20349 23974 20383
rect 23974 20349 23992 20383
rect 23296 20272 23348 20324
rect 23940 20340 23992 20349
rect 26148 20417 26157 20451
rect 26157 20417 26191 20451
rect 26191 20417 26200 20451
rect 26148 20408 26200 20417
rect 29736 20408 29788 20460
rect 32772 20476 32824 20528
rect 35716 20476 35768 20528
rect 30012 20451 30064 20460
rect 30012 20417 30021 20451
rect 30021 20417 30055 20451
rect 30055 20417 30064 20451
rect 30012 20408 30064 20417
rect 30472 20408 30524 20460
rect 31668 20408 31720 20460
rect 32588 20408 32640 20460
rect 33232 20451 33284 20460
rect 33232 20417 33241 20451
rect 33241 20417 33275 20451
rect 33275 20417 33284 20451
rect 33232 20408 33284 20417
rect 35348 20408 35400 20460
rect 26240 20340 26292 20392
rect 30288 20272 30340 20324
rect 33324 20272 33376 20324
rect 34612 20272 34664 20324
rect 25044 20247 25096 20256
rect 25044 20213 25053 20247
rect 25053 20213 25087 20247
rect 25087 20213 25096 20247
rect 25044 20204 25096 20213
rect 28448 20247 28500 20256
rect 28448 20213 28457 20247
rect 28457 20213 28491 20247
rect 28491 20213 28500 20247
rect 28448 20204 28500 20213
rect 28816 20204 28868 20256
rect 32956 20247 33008 20256
rect 32956 20213 32965 20247
rect 32965 20213 32999 20247
rect 32999 20213 33008 20247
rect 32956 20204 33008 20213
rect 33048 20247 33100 20256
rect 33048 20213 33057 20247
rect 33057 20213 33091 20247
rect 33091 20213 33100 20247
rect 33048 20204 33100 20213
rect 34428 20204 34480 20256
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 23756 20000 23808 20052
rect 23940 20000 23992 20052
rect 26240 20043 26292 20052
rect 26240 20009 26249 20043
rect 26249 20009 26283 20043
rect 26283 20009 26292 20043
rect 26240 20000 26292 20009
rect 26700 20043 26752 20052
rect 26700 20009 26709 20043
rect 26709 20009 26743 20043
rect 26743 20009 26752 20043
rect 26700 20000 26752 20009
rect 26884 20000 26936 20052
rect 28632 20000 28684 20052
rect 30012 20000 30064 20052
rect 33048 20043 33100 20052
rect 33048 20009 33057 20043
rect 33057 20009 33091 20043
rect 33091 20009 33100 20043
rect 33048 20000 33100 20009
rect 33232 20000 33284 20052
rect 35348 20000 35400 20052
rect 22744 19907 22796 19916
rect 22744 19873 22778 19907
rect 22778 19873 22796 19907
rect 22744 19864 22796 19873
rect 35532 19864 35584 19916
rect 22468 19839 22520 19848
rect 22468 19805 22477 19839
rect 22477 19805 22511 19839
rect 22511 19805 22520 19839
rect 22468 19796 22520 19805
rect 34612 19796 34664 19848
rect 30012 19660 30064 19712
rect 33048 19660 33100 19712
rect 34612 19703 34664 19712
rect 34612 19669 34621 19703
rect 34621 19669 34655 19703
rect 34655 19669 34664 19703
rect 34612 19660 34664 19669
rect 35348 19660 35400 19712
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 34966 19558 35018 19610
rect 35030 19558 35082 19610
rect 35094 19558 35146 19610
rect 35158 19558 35210 19610
rect 22744 19456 22796 19508
rect 33876 19499 33928 19508
rect 33876 19465 33885 19499
rect 33885 19465 33919 19499
rect 33919 19465 33928 19499
rect 33876 19456 33928 19465
rect 34428 19456 34480 19508
rect 22468 19388 22520 19440
rect 23296 19388 23348 19440
rect 34612 19320 34664 19372
rect 35164 19320 35216 19372
rect 35532 19363 35584 19372
rect 35532 19329 35541 19363
rect 35541 19329 35575 19363
rect 35575 19329 35584 19363
rect 35532 19320 35584 19329
rect 28816 19116 28868 19168
rect 30012 19227 30064 19236
rect 30012 19193 30046 19227
rect 30046 19193 30064 19227
rect 30012 19184 30064 19193
rect 34704 19184 34756 19236
rect 31024 19116 31076 19168
rect 32404 19116 32456 19168
rect 33508 19159 33560 19168
rect 33508 19125 33517 19159
rect 33517 19125 33551 19159
rect 33551 19125 33560 19159
rect 33508 19116 33560 19125
rect 34336 19116 34388 19168
rect 35348 19116 35400 19168
rect 37188 19295 37240 19304
rect 37188 19261 37197 19295
rect 37197 19261 37231 19295
rect 37231 19261 37240 19295
rect 37188 19252 37240 19261
rect 35992 19159 36044 19168
rect 35992 19125 36001 19159
rect 36001 19125 36035 19159
rect 36035 19125 36044 19159
rect 35992 19116 36044 19125
rect 36268 19159 36320 19168
rect 36268 19125 36277 19159
rect 36277 19125 36311 19159
rect 36311 19125 36320 19159
rect 36268 19116 36320 19125
rect 36820 19159 36872 19168
rect 36820 19125 36829 19159
rect 36829 19125 36863 19159
rect 36863 19125 36872 19159
rect 36820 19116 36872 19125
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 25872 18955 25924 18964
rect 25872 18921 25881 18955
rect 25881 18921 25915 18955
rect 25915 18921 25924 18955
rect 25872 18912 25924 18921
rect 34704 18912 34756 18964
rect 35164 18955 35216 18964
rect 35164 18921 35173 18955
rect 35173 18921 35207 18955
rect 35207 18921 35216 18955
rect 35164 18912 35216 18921
rect 28264 18844 28316 18896
rect 29920 18844 29972 18896
rect 28172 18776 28224 18828
rect 32772 18776 32824 18828
rect 32956 18819 33008 18828
rect 32956 18785 32990 18819
rect 32990 18785 33008 18819
rect 32956 18776 33008 18785
rect 34244 18776 34296 18828
rect 28816 18751 28868 18760
rect 28816 18717 28825 18751
rect 28825 18717 28859 18751
rect 28859 18717 28868 18751
rect 28816 18708 28868 18717
rect 34428 18708 34480 18760
rect 35716 18751 35768 18760
rect 35716 18717 35725 18751
rect 35725 18717 35759 18751
rect 35759 18717 35768 18751
rect 35716 18708 35768 18717
rect 36820 18640 36872 18692
rect 29000 18572 29052 18624
rect 30012 18572 30064 18624
rect 31024 18615 31076 18624
rect 31024 18581 31033 18615
rect 31033 18581 31067 18615
rect 31067 18581 31076 18615
rect 31024 18572 31076 18581
rect 34060 18615 34112 18624
rect 34060 18581 34069 18615
rect 34069 18581 34103 18615
rect 34103 18581 34112 18615
rect 34060 18572 34112 18581
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 34966 18470 35018 18522
rect 35030 18470 35082 18522
rect 35094 18470 35146 18522
rect 35158 18470 35210 18522
rect 24492 18232 24544 18284
rect 26148 18368 26200 18420
rect 35992 18368 36044 18420
rect 36820 18411 36872 18420
rect 36820 18377 36829 18411
rect 36829 18377 36863 18411
rect 36863 18377 36872 18411
rect 36820 18368 36872 18377
rect 29920 18275 29972 18284
rect 29920 18241 29929 18275
rect 29929 18241 29963 18275
rect 29963 18241 29972 18275
rect 29920 18232 29972 18241
rect 34612 18300 34664 18352
rect 18880 18207 18932 18216
rect 18880 18173 18889 18207
rect 18889 18173 18923 18207
rect 18923 18173 18932 18207
rect 18880 18164 18932 18173
rect 25872 18164 25924 18216
rect 28540 18207 28592 18216
rect 28540 18173 28549 18207
rect 28549 18173 28583 18207
rect 28583 18173 28592 18207
rect 29736 18207 29788 18216
rect 28540 18164 28592 18173
rect 29736 18173 29745 18207
rect 29745 18173 29779 18207
rect 29779 18173 29788 18207
rect 29736 18164 29788 18173
rect 32772 18164 32824 18216
rect 33692 18207 33744 18216
rect 18696 18139 18748 18148
rect 18696 18105 18705 18139
rect 18705 18105 18739 18139
rect 18739 18105 18748 18139
rect 18696 18096 18748 18105
rect 28080 18096 28132 18148
rect 28816 18139 28868 18148
rect 28816 18105 28825 18139
rect 28825 18105 28859 18139
rect 28859 18105 28868 18139
rect 28816 18096 28868 18105
rect 31024 18096 31076 18148
rect 31668 18096 31720 18148
rect 32956 18096 33008 18148
rect 33692 18173 33701 18207
rect 33701 18173 33735 18207
rect 33735 18173 33744 18207
rect 33692 18164 33744 18173
rect 34336 18096 34388 18148
rect 35072 18096 35124 18148
rect 20260 18071 20312 18080
rect 20260 18037 20269 18071
rect 20269 18037 20303 18071
rect 20303 18037 20312 18071
rect 20260 18028 20312 18037
rect 27160 18071 27212 18080
rect 27160 18037 27169 18071
rect 27169 18037 27203 18071
rect 27203 18037 27212 18071
rect 27160 18028 27212 18037
rect 28172 18071 28224 18080
rect 28172 18037 28181 18071
rect 28181 18037 28215 18071
rect 28215 18037 28224 18071
rect 28172 18028 28224 18037
rect 29276 18071 29328 18080
rect 29276 18037 29285 18071
rect 29285 18037 29319 18071
rect 29319 18037 29328 18071
rect 29276 18028 29328 18037
rect 30288 18071 30340 18080
rect 30288 18037 30297 18071
rect 30297 18037 30331 18071
rect 30331 18037 30340 18071
rect 30288 18028 30340 18037
rect 32312 18071 32364 18080
rect 32312 18037 32321 18071
rect 32321 18037 32355 18071
rect 32355 18037 32364 18071
rect 32312 18028 32364 18037
rect 33140 18028 33192 18080
rect 34244 18071 34296 18080
rect 34244 18037 34253 18071
rect 34253 18037 34287 18071
rect 34287 18037 34296 18071
rect 34244 18028 34296 18037
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 29552 17867 29604 17876
rect 29552 17833 29561 17867
rect 29561 17833 29595 17867
rect 29595 17833 29604 17867
rect 29552 17824 29604 17833
rect 30288 17824 30340 17876
rect 33140 17824 33192 17876
rect 33692 17824 33744 17876
rect 35072 17824 35124 17876
rect 35716 17824 35768 17876
rect 28540 17756 28592 17808
rect 11612 17731 11664 17740
rect 11612 17697 11646 17731
rect 11646 17697 11664 17731
rect 11612 17688 11664 17697
rect 22652 17688 22704 17740
rect 23112 17688 23164 17740
rect 30932 17731 30984 17740
rect 30932 17697 30941 17731
rect 30941 17697 30975 17731
rect 30975 17697 30984 17731
rect 30932 17688 30984 17697
rect 33600 17688 33652 17740
rect 34060 17688 34112 17740
rect 11336 17663 11388 17672
rect 11336 17629 11345 17663
rect 11345 17629 11379 17663
rect 11379 17629 11388 17663
rect 11336 17620 11388 17629
rect 21456 17663 21508 17672
rect 21456 17629 21465 17663
rect 21465 17629 21499 17663
rect 21499 17629 21508 17663
rect 21456 17620 21508 17629
rect 8024 17527 8076 17536
rect 8024 17493 8033 17527
rect 8033 17493 8067 17527
rect 8067 17493 8076 17527
rect 8024 17484 8076 17493
rect 10876 17527 10928 17536
rect 10876 17493 10885 17527
rect 10885 17493 10919 17527
rect 10919 17493 10928 17527
rect 10876 17484 10928 17493
rect 12808 17484 12860 17536
rect 13268 17527 13320 17536
rect 13268 17493 13277 17527
rect 13277 17493 13311 17527
rect 13311 17493 13320 17527
rect 13268 17484 13320 17493
rect 18880 17527 18932 17536
rect 18880 17493 18889 17527
rect 18889 17493 18923 17527
rect 18923 17493 18932 17527
rect 18880 17484 18932 17493
rect 23756 17484 23808 17536
rect 28080 17620 28132 17672
rect 33324 17663 33376 17672
rect 33324 17629 33333 17663
rect 33333 17629 33367 17663
rect 33367 17629 33376 17663
rect 33324 17620 33376 17629
rect 34336 17620 34388 17672
rect 34060 17552 34112 17604
rect 24308 17484 24360 17536
rect 25320 17527 25372 17536
rect 25320 17493 25329 17527
rect 25329 17493 25363 17527
rect 25363 17493 25372 17527
rect 25320 17484 25372 17493
rect 27988 17484 28040 17536
rect 28908 17484 28960 17536
rect 30380 17484 30432 17536
rect 31852 17527 31904 17536
rect 31852 17493 31861 17527
rect 31861 17493 31895 17527
rect 31895 17493 31904 17527
rect 31852 17484 31904 17493
rect 32864 17527 32916 17536
rect 32864 17493 32873 17527
rect 32873 17493 32907 17527
rect 32907 17493 32916 17527
rect 32864 17484 32916 17493
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 34966 17382 35018 17434
rect 35030 17382 35082 17434
rect 35094 17382 35146 17434
rect 35158 17382 35210 17434
rect 11336 17280 11388 17332
rect 11888 17280 11940 17332
rect 22652 17323 22704 17332
rect 22652 17289 22661 17323
rect 22661 17289 22695 17323
rect 22695 17289 22704 17323
rect 22652 17280 22704 17289
rect 23112 17323 23164 17332
rect 23112 17289 23121 17323
rect 23121 17289 23155 17323
rect 23155 17289 23164 17323
rect 23112 17280 23164 17289
rect 24584 17280 24636 17332
rect 30932 17280 30984 17332
rect 28172 17212 28224 17264
rect 10876 17144 10928 17196
rect 13268 17144 13320 17196
rect 28264 17187 28316 17196
rect 28264 17153 28273 17187
rect 28273 17153 28307 17187
rect 28307 17153 28316 17187
rect 28264 17144 28316 17153
rect 31852 17144 31904 17196
rect 32772 17144 32824 17196
rect 7104 16940 7156 16992
rect 8024 17076 8076 17128
rect 11520 17076 11572 17128
rect 11612 17076 11664 17128
rect 13544 17119 13596 17128
rect 13544 17085 13553 17119
rect 13553 17085 13587 17119
rect 13587 17085 13596 17119
rect 13544 17076 13596 17085
rect 21456 17076 21508 17128
rect 20260 17051 20312 17060
rect 20260 17017 20269 17051
rect 20269 17017 20303 17051
rect 20303 17017 20312 17051
rect 20260 17008 20312 17017
rect 22192 17008 22244 17060
rect 23756 17076 23808 17128
rect 27988 17119 28040 17128
rect 27988 17085 27997 17119
rect 27997 17085 28031 17119
rect 28031 17085 28040 17119
rect 27988 17076 28040 17085
rect 28172 17076 28224 17128
rect 29552 17119 29604 17128
rect 29552 17085 29586 17119
rect 29586 17085 29604 17119
rect 29552 17076 29604 17085
rect 31116 17076 31168 17128
rect 33324 17280 33376 17332
rect 33600 17323 33652 17332
rect 33600 17289 33609 17323
rect 33609 17289 33643 17323
rect 33643 17289 33652 17323
rect 33600 17280 33652 17289
rect 34428 17280 34480 17332
rect 37096 17323 37148 17332
rect 37096 17289 37105 17323
rect 37105 17289 37139 17323
rect 37139 17289 37148 17323
rect 37096 17280 37148 17289
rect 34336 17144 34388 17196
rect 34612 17144 34664 17196
rect 35624 17144 35676 17196
rect 33784 17076 33836 17128
rect 24492 17008 24544 17060
rect 8300 16940 8352 16992
rect 10692 16940 10744 16992
rect 11152 16983 11204 16992
rect 11152 16949 11161 16983
rect 11161 16949 11195 16983
rect 11195 16949 11204 16983
rect 11152 16940 11204 16949
rect 12440 16983 12492 16992
rect 12440 16949 12449 16983
rect 12449 16949 12483 16983
rect 12483 16949 12492 16983
rect 12440 16940 12492 16949
rect 12808 16983 12860 16992
rect 12808 16949 12817 16983
rect 12817 16949 12851 16983
rect 12851 16949 12860 16983
rect 12808 16940 12860 16949
rect 22100 16983 22152 16992
rect 22100 16949 22109 16983
rect 22109 16949 22143 16983
rect 22143 16949 22152 16983
rect 22100 16940 22152 16949
rect 28080 16940 28132 16992
rect 28356 16940 28408 16992
rect 30656 16983 30708 16992
rect 30656 16949 30665 16983
rect 30665 16949 30699 16983
rect 30699 16949 30708 16983
rect 30656 16940 30708 16949
rect 32128 16983 32180 16992
rect 32128 16949 32137 16983
rect 32137 16949 32171 16983
rect 32171 16949 32180 16983
rect 32128 16940 32180 16949
rect 34980 17076 35032 17128
rect 37096 17076 37148 17128
rect 35348 16983 35400 16992
rect 35348 16949 35357 16983
rect 35357 16949 35391 16983
rect 35391 16949 35400 16983
rect 35348 16940 35400 16949
rect 36452 16940 36504 16992
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 7472 16736 7524 16788
rect 8300 16779 8352 16788
rect 8300 16745 8309 16779
rect 8309 16745 8343 16779
rect 8343 16745 8352 16779
rect 8300 16736 8352 16745
rect 11612 16736 11664 16788
rect 22652 16736 22704 16788
rect 7748 16643 7800 16652
rect 7748 16609 7757 16643
rect 7757 16609 7791 16643
rect 7791 16609 7800 16643
rect 7748 16600 7800 16609
rect 8024 16668 8076 16720
rect 8208 16643 8260 16652
rect 8208 16609 8217 16643
rect 8217 16609 8251 16643
rect 8251 16609 8260 16643
rect 8208 16600 8260 16609
rect 11152 16668 11204 16720
rect 12532 16668 12584 16720
rect 22100 16668 22152 16720
rect 23480 16736 23532 16788
rect 29736 16779 29788 16788
rect 29736 16745 29745 16779
rect 29745 16745 29779 16779
rect 29779 16745 29788 16779
rect 29736 16736 29788 16745
rect 30380 16779 30432 16788
rect 30380 16745 30389 16779
rect 30389 16745 30423 16779
rect 30423 16745 30432 16779
rect 30380 16736 30432 16745
rect 31116 16779 31168 16788
rect 31116 16745 31125 16779
rect 31125 16745 31159 16779
rect 31159 16745 31168 16779
rect 31116 16736 31168 16745
rect 32128 16779 32180 16788
rect 32128 16745 32137 16779
rect 32137 16745 32171 16779
rect 32171 16745 32180 16779
rect 32128 16736 32180 16745
rect 33140 16779 33192 16788
rect 33140 16745 33149 16779
rect 33149 16745 33183 16779
rect 33183 16745 33192 16779
rect 33140 16736 33192 16745
rect 33784 16779 33836 16788
rect 33784 16745 33793 16779
rect 33793 16745 33827 16779
rect 33827 16745 33836 16779
rect 33784 16736 33836 16745
rect 33968 16736 34020 16788
rect 35348 16779 35400 16788
rect 35348 16745 35357 16779
rect 35357 16745 35391 16779
rect 35391 16745 35400 16779
rect 35348 16736 35400 16745
rect 35624 16779 35676 16788
rect 35624 16745 35633 16779
rect 35633 16745 35667 16779
rect 35667 16745 35676 16779
rect 35624 16736 35676 16745
rect 23664 16668 23716 16720
rect 23756 16668 23808 16720
rect 24308 16668 24360 16720
rect 31760 16668 31812 16720
rect 32220 16668 32272 16720
rect 34060 16711 34112 16720
rect 34060 16677 34069 16711
rect 34069 16677 34103 16711
rect 34103 16677 34112 16711
rect 34060 16668 34112 16677
rect 10140 16575 10192 16584
rect 10140 16541 10149 16575
rect 10149 16541 10183 16575
rect 10183 16541 10192 16575
rect 10140 16532 10192 16541
rect 9128 16464 9180 16516
rect 10876 16532 10928 16584
rect 11244 16600 11296 16652
rect 12808 16600 12860 16652
rect 24860 16600 24912 16652
rect 25320 16600 25372 16652
rect 26516 16643 26568 16652
rect 26516 16609 26525 16643
rect 26525 16609 26559 16643
rect 26559 16609 26568 16643
rect 26516 16600 26568 16609
rect 28632 16643 28684 16652
rect 28632 16609 28666 16643
rect 28666 16609 28684 16643
rect 30932 16643 30984 16652
rect 28632 16600 28684 16609
rect 30932 16609 30941 16643
rect 30941 16609 30975 16643
rect 30975 16609 30984 16643
rect 30932 16600 30984 16609
rect 31852 16600 31904 16652
rect 32312 16600 32364 16652
rect 32772 16600 32824 16652
rect 34612 16643 34664 16652
rect 11152 16532 11204 16584
rect 11336 16575 11388 16584
rect 11336 16541 11345 16575
rect 11345 16541 11379 16575
rect 11379 16541 11388 16575
rect 11336 16532 11388 16541
rect 24216 16532 24268 16584
rect 27528 16532 27580 16584
rect 28356 16575 28408 16584
rect 28356 16541 28365 16575
rect 28365 16541 28399 16575
rect 28399 16541 28408 16575
rect 28356 16532 28408 16541
rect 32864 16532 32916 16584
rect 34612 16609 34621 16643
rect 34621 16609 34655 16643
rect 34655 16609 34664 16643
rect 34612 16600 34664 16609
rect 33876 16532 33928 16584
rect 34336 16532 34388 16584
rect 35808 16643 35860 16652
rect 35808 16609 35817 16643
rect 35817 16609 35851 16643
rect 35851 16609 35860 16643
rect 35808 16600 35860 16609
rect 35624 16532 35676 16584
rect 24492 16464 24544 16516
rect 7840 16439 7892 16448
rect 7840 16405 7849 16439
rect 7849 16405 7883 16439
rect 7883 16405 7892 16439
rect 7840 16396 7892 16405
rect 9680 16439 9732 16448
rect 9680 16405 9689 16439
rect 9689 16405 9723 16439
rect 9723 16405 9732 16439
rect 9680 16396 9732 16405
rect 21456 16439 21508 16448
rect 21456 16405 21465 16439
rect 21465 16405 21499 16439
rect 21499 16405 21508 16439
rect 21456 16396 21508 16405
rect 26700 16439 26752 16448
rect 26700 16405 26709 16439
rect 26709 16405 26743 16439
rect 26743 16405 26752 16439
rect 26700 16396 26752 16405
rect 36176 16396 36228 16448
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 34966 16294 35018 16346
rect 35030 16294 35082 16346
rect 35094 16294 35146 16346
rect 35158 16294 35210 16346
rect 7104 16235 7156 16244
rect 7104 16201 7113 16235
rect 7113 16201 7147 16235
rect 7147 16201 7156 16235
rect 7104 16192 7156 16201
rect 11152 16235 11204 16244
rect 11152 16201 11161 16235
rect 11161 16201 11195 16235
rect 11195 16201 11204 16235
rect 11152 16192 11204 16201
rect 23664 16192 23716 16244
rect 24768 16192 24820 16244
rect 28632 16192 28684 16244
rect 29276 16192 29328 16244
rect 31852 16235 31904 16244
rect 22192 16056 22244 16108
rect 24216 16056 24268 16108
rect 7472 16031 7524 16040
rect 7472 15997 7506 16031
rect 7506 15997 7524 16031
rect 7472 15988 7524 15997
rect 11336 15988 11388 16040
rect 11888 15988 11940 16040
rect 12532 15988 12584 16040
rect 22100 15988 22152 16040
rect 24492 16031 24544 16040
rect 24492 15997 24501 16031
rect 24501 15997 24535 16031
rect 24535 15997 24544 16031
rect 24492 15988 24544 15997
rect 27528 16099 27580 16108
rect 27528 16065 27537 16099
rect 27537 16065 27571 16099
rect 27571 16065 27580 16099
rect 27528 16056 27580 16065
rect 31852 16201 31861 16235
rect 31861 16201 31895 16235
rect 31895 16201 31904 16235
rect 31852 16192 31904 16201
rect 32220 16235 32272 16244
rect 32220 16201 32229 16235
rect 32229 16201 32263 16235
rect 32263 16201 32272 16235
rect 32220 16192 32272 16201
rect 33048 16192 33100 16244
rect 34336 16235 34388 16244
rect 34336 16201 34345 16235
rect 34345 16201 34379 16235
rect 34379 16201 34388 16235
rect 34336 16192 34388 16201
rect 34612 16235 34664 16244
rect 34612 16201 34621 16235
rect 34621 16201 34655 16235
rect 34655 16201 34664 16235
rect 34612 16192 34664 16201
rect 35624 16235 35676 16244
rect 35624 16201 35633 16235
rect 35633 16201 35667 16235
rect 35667 16201 35676 16235
rect 35624 16192 35676 16201
rect 35900 16192 35952 16244
rect 30932 16124 30984 16176
rect 30380 16056 30432 16108
rect 33968 16124 34020 16176
rect 35532 16124 35584 16176
rect 9496 15920 9548 15972
rect 10140 15920 10192 15972
rect 24676 15920 24728 15972
rect 8576 15895 8628 15904
rect 8576 15861 8585 15895
rect 8585 15861 8619 15895
rect 8619 15861 8628 15895
rect 8576 15852 8628 15861
rect 13820 15895 13872 15904
rect 13820 15861 13829 15895
rect 13829 15861 13863 15895
rect 13863 15861 13872 15895
rect 13820 15852 13872 15861
rect 20904 15852 20956 15904
rect 21456 15852 21508 15904
rect 22744 15852 22796 15904
rect 26240 15852 26292 15904
rect 26884 15852 26936 15904
rect 28356 15852 28408 15904
rect 29184 15852 29236 15904
rect 29828 15852 29880 15904
rect 34428 15852 34480 15904
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 8300 15691 8352 15700
rect 8300 15657 8309 15691
rect 8309 15657 8343 15691
rect 8343 15657 8352 15691
rect 8300 15648 8352 15657
rect 9128 15691 9180 15700
rect 9128 15657 9137 15691
rect 9137 15657 9171 15691
rect 9171 15657 9180 15691
rect 9128 15648 9180 15657
rect 9496 15691 9548 15700
rect 9496 15657 9505 15691
rect 9505 15657 9539 15691
rect 9539 15657 9548 15691
rect 9496 15648 9548 15657
rect 10048 15691 10100 15700
rect 10048 15657 10057 15691
rect 10057 15657 10091 15691
rect 10091 15657 10100 15691
rect 10048 15648 10100 15657
rect 11244 15691 11296 15700
rect 11244 15657 11253 15691
rect 11253 15657 11287 15691
rect 11287 15657 11296 15691
rect 11244 15648 11296 15657
rect 12532 15648 12584 15700
rect 22100 15648 22152 15700
rect 22744 15648 22796 15700
rect 24308 15691 24360 15700
rect 24308 15657 24317 15691
rect 24317 15657 24351 15691
rect 24351 15657 24360 15691
rect 24308 15648 24360 15657
rect 24584 15648 24636 15700
rect 30564 15691 30616 15700
rect 30564 15657 30573 15691
rect 30573 15657 30607 15691
rect 30607 15657 30616 15691
rect 30564 15648 30616 15657
rect 34612 15648 34664 15700
rect 8208 15580 8260 15632
rect 8576 15580 8628 15632
rect 11612 15623 11664 15632
rect 11612 15589 11646 15623
rect 11646 15589 11664 15623
rect 11612 15580 11664 15589
rect 23388 15580 23440 15632
rect 32956 15580 33008 15632
rect 7104 15512 7156 15564
rect 11336 15555 11388 15564
rect 11336 15521 11345 15555
rect 11345 15521 11379 15555
rect 11379 15521 11388 15555
rect 11336 15512 11388 15521
rect 22192 15512 22244 15564
rect 23480 15512 23532 15564
rect 24676 15512 24728 15564
rect 26884 15555 26936 15564
rect 26884 15521 26893 15555
rect 26893 15521 26927 15555
rect 26927 15521 26936 15555
rect 26884 15512 26936 15521
rect 27528 15512 27580 15564
rect 29184 15555 29236 15564
rect 29184 15521 29193 15555
rect 29193 15521 29227 15555
rect 29227 15521 29236 15555
rect 29184 15512 29236 15521
rect 29460 15555 29512 15564
rect 29460 15521 29494 15555
rect 29494 15521 29512 15555
rect 29460 15512 29512 15521
rect 34060 15555 34112 15564
rect 34060 15521 34069 15555
rect 34069 15521 34103 15555
rect 34103 15521 34112 15555
rect 34060 15512 34112 15521
rect 34612 15512 34664 15564
rect 6368 15487 6420 15496
rect 6368 15453 6377 15487
rect 6377 15453 6411 15487
rect 6411 15453 6420 15487
rect 6368 15444 6420 15453
rect 9680 15444 9732 15496
rect 10232 15487 10284 15496
rect 10232 15453 10241 15487
rect 10241 15453 10275 15487
rect 10275 15453 10284 15487
rect 10232 15444 10284 15453
rect 22928 15444 22980 15496
rect 24216 15444 24268 15496
rect 25964 15444 26016 15496
rect 26424 15444 26476 15496
rect 22836 15419 22888 15428
rect 22836 15385 22845 15419
rect 22845 15385 22879 15419
rect 22879 15385 22888 15419
rect 22836 15376 22888 15385
rect 24768 15376 24820 15428
rect 26792 15376 26844 15428
rect 32404 15444 32456 15496
rect 35624 15487 35676 15496
rect 32864 15376 32916 15428
rect 35624 15453 35633 15487
rect 35633 15453 35667 15487
rect 35667 15453 35676 15487
rect 35624 15444 35676 15453
rect 35348 15376 35400 15428
rect 5264 15351 5316 15360
rect 5264 15317 5273 15351
rect 5273 15317 5307 15351
rect 5307 15317 5316 15351
rect 5264 15308 5316 15317
rect 7748 15351 7800 15360
rect 7748 15317 7757 15351
rect 7757 15317 7791 15351
rect 7791 15317 7800 15351
rect 7748 15308 7800 15317
rect 9496 15308 9548 15360
rect 19248 15351 19300 15360
rect 19248 15317 19257 15351
rect 19257 15317 19291 15351
rect 19291 15317 19300 15351
rect 19248 15308 19300 15317
rect 24400 15351 24452 15360
rect 24400 15317 24409 15351
rect 24409 15317 24443 15351
rect 24443 15317 24452 15351
rect 24400 15308 24452 15317
rect 26332 15351 26384 15360
rect 26332 15317 26341 15351
rect 26341 15317 26375 15351
rect 26375 15317 26384 15351
rect 26332 15308 26384 15317
rect 26516 15351 26568 15360
rect 26516 15317 26525 15351
rect 26525 15317 26559 15351
rect 26559 15317 26568 15351
rect 26516 15308 26568 15317
rect 27528 15308 27580 15360
rect 33048 15308 33100 15360
rect 33416 15308 33468 15360
rect 33968 15351 34020 15360
rect 33968 15317 33977 15351
rect 33977 15317 34011 15351
rect 34011 15317 34020 15351
rect 33968 15308 34020 15317
rect 35256 15308 35308 15360
rect 35992 15308 36044 15360
rect 36176 15351 36228 15360
rect 36176 15317 36185 15351
rect 36185 15317 36219 15351
rect 36219 15317 36228 15351
rect 36176 15308 36228 15317
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 34966 15206 35018 15258
rect 35030 15206 35082 15258
rect 35094 15206 35146 15258
rect 35158 15206 35210 15258
rect 9588 15104 9640 15156
rect 11336 15147 11388 15156
rect 11336 15113 11345 15147
rect 11345 15113 11379 15147
rect 11379 15113 11388 15147
rect 11336 15104 11388 15113
rect 11612 15104 11664 15156
rect 18880 15104 18932 15156
rect 5264 14968 5316 15020
rect 5816 15011 5868 15020
rect 5816 14977 5825 15011
rect 5825 14977 5859 15011
rect 5859 14977 5868 15011
rect 5816 14968 5868 14977
rect 9864 14968 9916 15020
rect 10232 14968 10284 15020
rect 17960 14968 18012 15020
rect 22744 15104 22796 15156
rect 23480 15147 23532 15156
rect 23480 15113 23489 15147
rect 23489 15113 23523 15147
rect 23523 15113 23532 15147
rect 23480 15104 23532 15113
rect 24492 15104 24544 15156
rect 26424 15104 26476 15156
rect 27620 15147 27672 15156
rect 27620 15113 27629 15147
rect 27629 15113 27663 15147
rect 27663 15113 27672 15147
rect 27620 15104 27672 15113
rect 29184 15104 29236 15156
rect 23388 15036 23440 15088
rect 24308 15079 24360 15088
rect 24308 15045 24317 15079
rect 24317 15045 24351 15079
rect 24351 15045 24360 15079
rect 24308 15036 24360 15045
rect 34428 15104 34480 15156
rect 37096 15147 37148 15156
rect 37096 15113 37105 15147
rect 37105 15113 37139 15147
rect 37139 15113 37148 15147
rect 37096 15104 37148 15113
rect 34060 15036 34112 15088
rect 33416 15011 33468 15020
rect 6368 14900 6420 14952
rect 10692 14900 10744 14952
rect 19248 14900 19300 14952
rect 24768 14943 24820 14952
rect 24768 14909 24802 14943
rect 24802 14909 24820 14943
rect 24768 14900 24820 14909
rect 26516 14900 26568 14952
rect 29460 14900 29512 14952
rect 30288 14900 30340 14952
rect 33416 14977 33425 15011
rect 33425 14977 33459 15011
rect 33459 14977 33468 15011
rect 33416 14968 33468 14977
rect 33968 14968 34020 15020
rect 35532 15011 35584 15020
rect 35532 14977 35541 15011
rect 35541 14977 35575 15011
rect 35575 14977 35584 15011
rect 35532 14968 35584 14977
rect 32128 14900 32180 14952
rect 33140 14900 33192 14952
rect 35256 14943 35308 14952
rect 35256 14909 35265 14943
rect 35265 14909 35299 14943
rect 35299 14909 35308 14943
rect 35256 14900 35308 14909
rect 37096 14900 37148 14952
rect 7748 14832 7800 14884
rect 7840 14832 7892 14884
rect 9864 14832 9916 14884
rect 5172 14807 5224 14816
rect 5172 14773 5181 14807
rect 5181 14773 5215 14807
rect 5215 14773 5224 14807
rect 5172 14764 5224 14773
rect 5540 14807 5592 14816
rect 5540 14773 5549 14807
rect 5549 14773 5583 14807
rect 5583 14773 5592 14807
rect 5540 14764 5592 14773
rect 5724 14764 5776 14816
rect 6644 14764 6696 14816
rect 10232 14807 10284 14816
rect 10232 14773 10241 14807
rect 10241 14773 10275 14807
rect 10275 14773 10284 14807
rect 10232 14764 10284 14773
rect 26792 14832 26844 14884
rect 28448 14832 28500 14884
rect 30748 14875 30800 14884
rect 30748 14841 30782 14875
rect 30782 14841 30800 14875
rect 30748 14832 30800 14841
rect 10784 14764 10836 14816
rect 20536 14807 20588 14816
rect 20536 14773 20545 14807
rect 20545 14773 20579 14807
rect 20579 14773 20588 14807
rect 20536 14764 20588 14773
rect 25872 14807 25924 14816
rect 25872 14773 25881 14807
rect 25881 14773 25915 14807
rect 25915 14773 25924 14807
rect 25872 14764 25924 14773
rect 26240 14764 26292 14816
rect 27068 14764 27120 14816
rect 31852 14807 31904 14816
rect 31852 14773 31861 14807
rect 31861 14773 31895 14807
rect 31895 14773 31904 14807
rect 31852 14764 31904 14773
rect 32404 14764 32456 14816
rect 32956 14764 33008 14816
rect 33600 14764 33652 14816
rect 34612 14807 34664 14816
rect 34612 14773 34621 14807
rect 34621 14773 34655 14807
rect 34655 14773 34664 14807
rect 34612 14764 34664 14773
rect 35256 14764 35308 14816
rect 35624 14764 35676 14816
rect 36636 14807 36688 14816
rect 36636 14773 36645 14807
rect 36645 14773 36679 14807
rect 36679 14773 36688 14807
rect 36636 14764 36688 14773
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 7748 14603 7800 14612
rect 7748 14569 7757 14603
rect 7757 14569 7791 14603
rect 7791 14569 7800 14603
rect 7748 14560 7800 14569
rect 10048 14560 10100 14612
rect 19248 14560 19300 14612
rect 22928 14603 22980 14612
rect 22928 14569 22937 14603
rect 22937 14569 22971 14603
rect 22971 14569 22980 14603
rect 22928 14560 22980 14569
rect 24308 14560 24360 14612
rect 26700 14560 26752 14612
rect 28080 14560 28132 14612
rect 28448 14603 28500 14612
rect 28448 14569 28457 14603
rect 28457 14569 28491 14603
rect 28491 14569 28500 14603
rect 28448 14560 28500 14569
rect 29828 14603 29880 14612
rect 29828 14569 29837 14603
rect 29837 14569 29871 14603
rect 29871 14569 29880 14603
rect 29828 14560 29880 14569
rect 30288 14603 30340 14612
rect 30288 14569 30297 14603
rect 30297 14569 30331 14603
rect 30331 14569 30340 14603
rect 30288 14560 30340 14569
rect 33416 14560 33468 14612
rect 34060 14603 34112 14612
rect 34060 14569 34069 14603
rect 34069 14569 34103 14603
rect 34103 14569 34112 14603
rect 34060 14560 34112 14569
rect 35532 14560 35584 14612
rect 36452 14603 36504 14612
rect 36452 14569 36461 14603
rect 36461 14569 36495 14603
rect 36495 14569 36504 14603
rect 36452 14560 36504 14569
rect 5540 14424 5592 14476
rect 6644 14424 6696 14476
rect 8760 14492 8812 14544
rect 9496 14492 9548 14544
rect 9864 14492 9916 14544
rect 16948 14492 17000 14544
rect 30196 14535 30248 14544
rect 30196 14501 30205 14535
rect 30205 14501 30239 14535
rect 30239 14501 30248 14535
rect 30196 14492 30248 14501
rect 31852 14492 31904 14544
rect 32864 14492 32916 14544
rect 9220 14424 9272 14476
rect 10232 14424 10284 14476
rect 11060 14424 11112 14476
rect 18052 14424 18104 14476
rect 23572 14424 23624 14476
rect 27068 14467 27120 14476
rect 27068 14433 27077 14467
rect 27077 14433 27111 14467
rect 27111 14433 27120 14467
rect 27068 14424 27120 14433
rect 32588 14424 32640 14476
rect 5724 14356 5776 14408
rect 17960 14399 18012 14408
rect 16580 14288 16632 14340
rect 17960 14365 17969 14399
rect 17969 14365 18003 14399
rect 18003 14365 18012 14399
rect 17960 14356 18012 14365
rect 27528 14356 27580 14408
rect 29920 14356 29972 14408
rect 30472 14399 30524 14408
rect 30472 14365 30481 14399
rect 30481 14365 30515 14399
rect 30515 14365 30524 14399
rect 30472 14356 30524 14365
rect 34612 14424 34664 14476
rect 6828 14220 6880 14272
rect 9496 14220 9548 14272
rect 9956 14220 10008 14272
rect 11244 14220 11296 14272
rect 15752 14220 15804 14272
rect 16396 14263 16448 14272
rect 16396 14229 16405 14263
rect 16405 14229 16439 14263
rect 16439 14229 16448 14263
rect 16396 14220 16448 14229
rect 18972 14220 19024 14272
rect 25412 14263 25464 14272
rect 25412 14229 25421 14263
rect 25421 14229 25455 14263
rect 25455 14229 25464 14263
rect 25412 14220 25464 14229
rect 26332 14263 26384 14272
rect 26332 14229 26341 14263
rect 26341 14229 26375 14263
rect 26375 14229 26384 14263
rect 26332 14220 26384 14229
rect 26700 14263 26752 14272
rect 26700 14229 26709 14263
rect 26709 14229 26743 14263
rect 26743 14229 26752 14263
rect 26700 14220 26752 14229
rect 27620 14220 27672 14272
rect 27804 14220 27856 14272
rect 32588 14220 32640 14272
rect 32956 14220 33008 14272
rect 33692 14356 33744 14408
rect 34428 14356 34480 14408
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 34966 14118 35018 14170
rect 35030 14118 35082 14170
rect 35094 14118 35146 14170
rect 35158 14118 35210 14170
rect 6644 14059 6696 14068
rect 6644 14025 6653 14059
rect 6653 14025 6687 14059
rect 6687 14025 6696 14059
rect 6644 14016 6696 14025
rect 8760 14059 8812 14068
rect 8760 14025 8769 14059
rect 8769 14025 8803 14059
rect 8803 14025 8812 14059
rect 8760 14016 8812 14025
rect 9220 14059 9272 14068
rect 9220 14025 9229 14059
rect 9229 14025 9263 14059
rect 9263 14025 9272 14059
rect 9220 14016 9272 14025
rect 9496 14059 9548 14068
rect 9496 14025 9505 14059
rect 9505 14025 9539 14059
rect 9539 14025 9548 14059
rect 9496 14016 9548 14025
rect 9956 14059 10008 14068
rect 9956 14025 9965 14059
rect 9965 14025 9999 14059
rect 9999 14025 10008 14059
rect 9956 14016 10008 14025
rect 17960 14016 18012 14068
rect 27068 14016 27120 14068
rect 30288 14016 30340 14068
rect 30472 14016 30524 14068
rect 31852 14059 31904 14068
rect 31852 14025 31861 14059
rect 31861 14025 31895 14059
rect 31895 14025 31904 14059
rect 31852 14016 31904 14025
rect 32128 14059 32180 14068
rect 32128 14025 32137 14059
rect 32137 14025 32171 14059
rect 32171 14025 32180 14059
rect 32128 14016 32180 14025
rect 32496 14016 32548 14068
rect 34612 14016 34664 14068
rect 5172 13991 5224 14000
rect 5172 13957 5181 13991
rect 5181 13957 5215 13991
rect 5215 13957 5224 13991
rect 5172 13948 5224 13957
rect 5816 13923 5868 13932
rect 5816 13889 5825 13923
rect 5825 13889 5859 13923
rect 5859 13889 5868 13923
rect 5816 13880 5868 13889
rect 6552 13880 6604 13932
rect 7380 13923 7432 13932
rect 7380 13889 7389 13923
rect 7389 13889 7423 13923
rect 7423 13889 7432 13923
rect 7380 13880 7432 13889
rect 7748 13880 7800 13932
rect 10324 13948 10376 14000
rect 28080 13991 28132 14000
rect 28080 13957 28089 13991
rect 28089 13957 28123 13991
rect 28123 13957 28132 13991
rect 28080 13948 28132 13957
rect 30196 13991 30248 14000
rect 30196 13957 30205 13991
rect 30205 13957 30239 13991
rect 30239 13957 30248 13991
rect 30196 13948 30248 13957
rect 18972 13880 19024 13932
rect 19064 13880 19116 13932
rect 6000 13744 6052 13796
rect 6828 13744 6880 13796
rect 7288 13787 7340 13796
rect 7288 13753 7297 13787
rect 7297 13753 7331 13787
rect 7331 13753 7340 13787
rect 9496 13812 9548 13864
rect 11060 13812 11112 13864
rect 7288 13744 7340 13753
rect 5540 13719 5592 13728
rect 5540 13685 5549 13719
rect 5549 13685 5583 13719
rect 5583 13685 5592 13719
rect 5540 13676 5592 13685
rect 5724 13676 5776 13728
rect 8208 13676 8260 13728
rect 10048 13719 10100 13728
rect 10048 13685 10057 13719
rect 10057 13685 10091 13719
rect 10091 13685 10100 13719
rect 10048 13676 10100 13685
rect 15200 13676 15252 13728
rect 15752 13855 15804 13864
rect 15752 13821 15786 13855
rect 15786 13821 15804 13855
rect 15752 13812 15804 13821
rect 18052 13812 18104 13864
rect 18604 13855 18656 13864
rect 18604 13821 18613 13855
rect 18613 13821 18647 13855
rect 18647 13821 18656 13855
rect 18604 13812 18656 13821
rect 19248 13812 19300 13864
rect 25964 13923 26016 13932
rect 19064 13744 19116 13796
rect 16948 13676 17000 13728
rect 18144 13719 18196 13728
rect 18144 13685 18153 13719
rect 18153 13685 18187 13719
rect 18187 13685 18196 13719
rect 18144 13676 18196 13685
rect 20536 13812 20588 13864
rect 23572 13812 23624 13864
rect 25964 13889 25973 13923
rect 25973 13889 26007 13923
rect 26007 13889 26016 13923
rect 25964 13880 26016 13889
rect 26332 13880 26384 13932
rect 26792 13923 26844 13932
rect 26792 13889 26801 13923
rect 26801 13889 26835 13923
rect 26835 13889 26844 13923
rect 26792 13880 26844 13889
rect 25872 13812 25924 13864
rect 26608 13812 26660 13864
rect 34428 13812 34480 13864
rect 24216 13744 24268 13796
rect 20904 13676 20956 13728
rect 21088 13719 21140 13728
rect 21088 13685 21097 13719
rect 21097 13685 21131 13719
rect 21131 13685 21140 13719
rect 21088 13676 21140 13685
rect 24308 13676 24360 13728
rect 25780 13719 25832 13728
rect 25780 13685 25789 13719
rect 25789 13685 25823 13719
rect 25823 13685 25832 13719
rect 25780 13676 25832 13685
rect 25872 13719 25924 13728
rect 25872 13685 25881 13719
rect 25881 13685 25915 13719
rect 25915 13685 25924 13719
rect 26240 13719 26292 13728
rect 25872 13676 25924 13685
rect 26240 13685 26249 13719
rect 26249 13685 26283 13719
rect 26283 13685 26292 13719
rect 26240 13676 26292 13685
rect 26516 13676 26568 13728
rect 27068 13719 27120 13728
rect 27068 13685 27077 13719
rect 27077 13685 27111 13719
rect 27111 13685 27120 13719
rect 27068 13676 27120 13685
rect 27804 13744 27856 13796
rect 32588 13787 32640 13796
rect 32588 13753 32622 13787
rect 32622 13753 32640 13787
rect 32588 13744 32640 13753
rect 35624 13787 35676 13796
rect 35624 13753 35658 13787
rect 35658 13753 35676 13787
rect 35624 13744 35676 13753
rect 27528 13676 27580 13728
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 5540 13472 5592 13524
rect 7104 13515 7156 13524
rect 7104 13481 7113 13515
rect 7113 13481 7147 13515
rect 7147 13481 7156 13515
rect 7104 13472 7156 13481
rect 18052 13515 18104 13524
rect 18052 13481 18061 13515
rect 18061 13481 18095 13515
rect 18095 13481 18104 13515
rect 18052 13472 18104 13481
rect 18604 13515 18656 13524
rect 18604 13481 18613 13515
rect 18613 13481 18647 13515
rect 18647 13481 18656 13515
rect 18604 13472 18656 13481
rect 19064 13515 19116 13524
rect 19064 13481 19073 13515
rect 19073 13481 19107 13515
rect 19107 13481 19116 13515
rect 19064 13472 19116 13481
rect 25872 13472 25924 13524
rect 26608 13515 26660 13524
rect 6000 13447 6052 13456
rect 6000 13413 6034 13447
rect 6034 13413 6052 13447
rect 6000 13404 6052 13413
rect 20076 13404 20128 13456
rect 21088 13404 21140 13456
rect 8208 13379 8260 13388
rect 8208 13345 8217 13379
rect 8217 13345 8251 13379
rect 8251 13345 8260 13379
rect 8208 13336 8260 13345
rect 9956 13336 10008 13388
rect 11704 13379 11756 13388
rect 11704 13345 11713 13379
rect 11713 13345 11747 13379
rect 11747 13345 11756 13379
rect 11704 13336 11756 13345
rect 12348 13336 12400 13388
rect 16948 13379 17000 13388
rect 16948 13345 16982 13379
rect 16982 13345 17000 13379
rect 16948 13336 17000 13345
rect 17776 13336 17828 13388
rect 20628 13336 20680 13388
rect 24216 13404 24268 13456
rect 26608 13481 26617 13515
rect 26617 13481 26651 13515
rect 26651 13481 26660 13515
rect 26608 13472 26660 13481
rect 27804 13472 27856 13524
rect 32588 13472 32640 13524
rect 34612 13515 34664 13524
rect 34612 13481 34621 13515
rect 34621 13481 34655 13515
rect 34655 13481 34664 13515
rect 34612 13472 34664 13481
rect 35624 13472 35676 13524
rect 26792 13404 26844 13456
rect 32956 13447 33008 13456
rect 32956 13413 32990 13447
rect 32990 13413 33008 13447
rect 32956 13404 33008 13413
rect 35348 13404 35400 13456
rect 24308 13336 24360 13388
rect 25872 13336 25924 13388
rect 26976 13379 27028 13388
rect 26976 13345 26985 13379
rect 26985 13345 27019 13379
rect 27019 13345 27028 13379
rect 26976 13336 27028 13345
rect 28080 13379 28132 13388
rect 28080 13345 28089 13379
rect 28089 13345 28123 13379
rect 28123 13345 28132 13379
rect 28080 13336 28132 13345
rect 30564 13336 30616 13388
rect 32128 13336 32180 13388
rect 36820 13336 36872 13388
rect 5724 13311 5776 13320
rect 5724 13277 5733 13311
rect 5733 13277 5767 13311
rect 5767 13277 5776 13311
rect 5724 13268 5776 13277
rect 11980 13311 12032 13320
rect 11980 13277 11989 13311
rect 11989 13277 12023 13311
rect 12023 13277 12032 13311
rect 11980 13268 12032 13277
rect 15200 13268 15252 13320
rect 16304 13200 16356 13252
rect 16580 13200 16632 13252
rect 7748 13132 7800 13184
rect 8392 13175 8444 13184
rect 8392 13141 8401 13175
rect 8401 13141 8435 13175
rect 8435 13141 8444 13175
rect 8392 13132 8444 13141
rect 10324 13132 10376 13184
rect 10692 13175 10744 13184
rect 10692 13141 10701 13175
rect 10701 13141 10735 13175
rect 10735 13141 10744 13175
rect 10692 13132 10744 13141
rect 12256 13132 12308 13184
rect 14464 13132 14516 13184
rect 15568 13175 15620 13184
rect 15568 13141 15577 13175
rect 15577 13141 15611 13175
rect 15611 13141 15620 13175
rect 15568 13132 15620 13141
rect 18972 13268 19024 13320
rect 19892 13311 19944 13320
rect 19892 13277 19901 13311
rect 19901 13277 19935 13311
rect 19935 13277 19944 13311
rect 19892 13268 19944 13277
rect 20904 13311 20956 13320
rect 20904 13277 20913 13311
rect 20913 13277 20947 13311
rect 20947 13277 20956 13311
rect 20904 13268 20956 13277
rect 26792 13268 26844 13320
rect 28172 13311 28224 13320
rect 25964 13200 26016 13252
rect 28172 13277 28181 13311
rect 28181 13277 28215 13311
rect 28215 13277 28224 13311
rect 28172 13268 28224 13277
rect 17868 13132 17920 13184
rect 19248 13175 19300 13184
rect 19248 13141 19257 13175
rect 19257 13141 19291 13175
rect 19291 13141 19300 13175
rect 19248 13132 19300 13141
rect 22284 13175 22336 13184
rect 22284 13141 22293 13175
rect 22293 13141 22327 13175
rect 22327 13141 22336 13175
rect 22284 13132 22336 13141
rect 24860 13175 24912 13184
rect 24860 13141 24869 13175
rect 24869 13141 24903 13175
rect 24903 13141 24912 13175
rect 25780 13175 25832 13184
rect 24860 13132 24912 13141
rect 25780 13141 25789 13175
rect 25789 13141 25823 13175
rect 25823 13141 25832 13175
rect 25780 13132 25832 13141
rect 28264 13132 28316 13184
rect 34428 13268 34480 13320
rect 29368 13175 29420 13184
rect 29368 13141 29377 13175
rect 29377 13141 29411 13175
rect 29411 13141 29420 13175
rect 29368 13132 29420 13141
rect 29644 13175 29696 13184
rect 29644 13141 29653 13175
rect 29653 13141 29687 13175
rect 29687 13141 29696 13175
rect 29644 13132 29696 13141
rect 30196 13132 30248 13184
rect 30564 13175 30616 13184
rect 30564 13141 30573 13175
rect 30573 13141 30607 13175
rect 30607 13141 30616 13175
rect 30564 13132 30616 13141
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 34966 13030 35018 13082
rect 35030 13030 35082 13082
rect 35094 13030 35146 13082
rect 35158 13030 35210 13082
rect 6000 12928 6052 12980
rect 8208 12928 8260 12980
rect 10048 12928 10100 12980
rect 11704 12971 11756 12980
rect 7104 12767 7156 12776
rect 7104 12733 7138 12767
rect 7138 12733 7156 12767
rect 7104 12724 7156 12733
rect 7840 12656 7892 12708
rect 11704 12937 11713 12971
rect 11713 12937 11747 12971
rect 11747 12937 11756 12971
rect 11704 12928 11756 12937
rect 17776 12971 17828 12980
rect 17776 12937 17785 12971
rect 17785 12937 17819 12971
rect 17819 12937 17828 12971
rect 17776 12928 17828 12937
rect 18144 12928 18196 12980
rect 20076 12971 20128 12980
rect 17868 12860 17920 12912
rect 10784 12792 10836 12844
rect 11244 12835 11296 12844
rect 11244 12801 11253 12835
rect 11253 12801 11287 12835
rect 11287 12801 11296 12835
rect 11244 12792 11296 12801
rect 14464 12835 14516 12844
rect 14464 12801 14473 12835
rect 14473 12801 14507 12835
rect 14507 12801 14516 12835
rect 14464 12792 14516 12801
rect 20076 12937 20085 12971
rect 20085 12937 20119 12971
rect 20119 12937 20128 12971
rect 20076 12928 20128 12937
rect 24308 12971 24360 12980
rect 24308 12937 24317 12971
rect 24317 12937 24351 12971
rect 24351 12937 24360 12971
rect 24308 12928 24360 12937
rect 25044 12928 25096 12980
rect 25412 12928 25464 12980
rect 25964 12928 26016 12980
rect 27436 12971 27488 12980
rect 27436 12937 27445 12971
rect 27445 12937 27479 12971
rect 27479 12937 27488 12971
rect 27436 12928 27488 12937
rect 28172 12928 28224 12980
rect 28816 12928 28868 12980
rect 30564 12928 30616 12980
rect 31576 12971 31628 12980
rect 31576 12937 31585 12971
rect 31585 12937 31619 12971
rect 31619 12937 31628 12971
rect 31576 12928 31628 12937
rect 32128 12971 32180 12980
rect 32128 12937 32137 12971
rect 32137 12937 32171 12971
rect 32171 12937 32180 12971
rect 32128 12928 32180 12937
rect 33600 12971 33652 12980
rect 33600 12937 33609 12971
rect 33609 12937 33643 12971
rect 33643 12937 33652 12971
rect 33600 12928 33652 12937
rect 34428 12928 34480 12980
rect 36820 12971 36872 12980
rect 23480 12860 23532 12912
rect 24216 12860 24268 12912
rect 26976 12860 27028 12912
rect 27896 12860 27948 12912
rect 29000 12860 29052 12912
rect 19524 12835 19576 12844
rect 19524 12801 19533 12835
rect 19533 12801 19567 12835
rect 19567 12801 19576 12835
rect 19524 12792 19576 12801
rect 29368 12792 29420 12844
rect 29736 12835 29788 12844
rect 29736 12801 29745 12835
rect 29745 12801 29779 12835
rect 29779 12801 29788 12835
rect 29736 12792 29788 12801
rect 30380 12860 30432 12912
rect 36820 12937 36829 12971
rect 36829 12937 36863 12971
rect 36863 12937 36872 12971
rect 36820 12928 36872 12937
rect 10692 12724 10744 12776
rect 15200 12724 15252 12776
rect 19248 12724 19300 12776
rect 15568 12656 15620 12708
rect 16488 12656 16540 12708
rect 20076 12656 20128 12708
rect 5724 12588 5776 12640
rect 6736 12588 6788 12640
rect 6920 12588 6972 12640
rect 9588 12588 9640 12640
rect 9956 12631 10008 12640
rect 9956 12597 9965 12631
rect 9965 12597 9999 12631
rect 9999 12597 10008 12631
rect 9956 12588 10008 12597
rect 10968 12588 11020 12640
rect 12348 12588 12400 12640
rect 13912 12631 13964 12640
rect 13912 12597 13921 12631
rect 13921 12597 13955 12631
rect 13955 12597 13964 12631
rect 13912 12588 13964 12597
rect 14280 12631 14332 12640
rect 14280 12597 14289 12631
rect 14289 12597 14323 12631
rect 14323 12597 14332 12631
rect 14280 12588 14332 12597
rect 15200 12588 15252 12640
rect 16856 12631 16908 12640
rect 16856 12597 16865 12631
rect 16865 12597 16899 12631
rect 16899 12597 16908 12631
rect 16856 12588 16908 12597
rect 18972 12631 19024 12640
rect 18972 12597 18981 12631
rect 18981 12597 19015 12631
rect 19015 12597 19024 12631
rect 18972 12588 19024 12597
rect 20628 12724 20680 12776
rect 22284 12724 22336 12776
rect 25412 12724 25464 12776
rect 26792 12724 26844 12776
rect 29644 12767 29696 12776
rect 29644 12733 29653 12767
rect 29653 12733 29687 12767
rect 29687 12733 29696 12767
rect 29644 12724 29696 12733
rect 31576 12724 31628 12776
rect 35348 12724 35400 12776
rect 25872 12699 25924 12708
rect 25872 12665 25881 12699
rect 25881 12665 25915 12699
rect 25915 12665 25924 12699
rect 25872 12656 25924 12665
rect 20904 12588 20956 12640
rect 21916 12631 21968 12640
rect 21916 12597 21925 12631
rect 21925 12597 21959 12631
rect 21959 12597 21968 12631
rect 21916 12588 21968 12597
rect 29276 12631 29328 12640
rect 29276 12597 29285 12631
rect 29285 12597 29319 12631
rect 29319 12597 29328 12631
rect 29276 12588 29328 12597
rect 30380 12588 30432 12640
rect 32404 12656 32456 12708
rect 35716 12699 35768 12708
rect 35716 12665 35750 12699
rect 35750 12665 35768 12699
rect 35716 12656 35768 12665
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 9956 12384 10008 12436
rect 10600 12384 10652 12436
rect 10784 12427 10836 12436
rect 10784 12393 10793 12427
rect 10793 12393 10827 12427
rect 10827 12393 10836 12427
rect 10784 12384 10836 12393
rect 14280 12384 14332 12436
rect 16580 12384 16632 12436
rect 18328 12427 18380 12436
rect 18328 12393 18337 12427
rect 18337 12393 18371 12427
rect 18371 12393 18380 12427
rect 18328 12384 18380 12393
rect 19340 12384 19392 12436
rect 20628 12427 20680 12436
rect 20628 12393 20637 12427
rect 20637 12393 20671 12427
rect 20671 12393 20680 12427
rect 20628 12384 20680 12393
rect 25964 12384 26016 12436
rect 27896 12427 27948 12436
rect 27896 12393 27905 12427
rect 27905 12393 27939 12427
rect 27939 12393 27948 12427
rect 27896 12384 27948 12393
rect 28080 12384 28132 12436
rect 30380 12427 30432 12436
rect 7012 12316 7064 12368
rect 8392 12316 8444 12368
rect 6736 12248 6788 12300
rect 9680 12248 9732 12300
rect 10048 12291 10100 12300
rect 10048 12257 10057 12291
rect 10057 12257 10091 12291
rect 10091 12257 10100 12291
rect 10048 12248 10100 12257
rect 11980 12248 12032 12300
rect 12440 12248 12492 12300
rect 14832 12248 14884 12300
rect 16212 12248 16264 12300
rect 18236 12291 18288 12300
rect 18236 12257 18245 12291
rect 18245 12257 18279 12291
rect 18279 12257 18288 12291
rect 18236 12248 18288 12257
rect 26792 12359 26844 12368
rect 26792 12325 26826 12359
rect 26826 12325 26844 12359
rect 26792 12316 26844 12325
rect 30380 12393 30389 12427
rect 30389 12393 30423 12427
rect 30423 12393 30432 12427
rect 30380 12384 30432 12393
rect 32404 12427 32456 12436
rect 32404 12393 32413 12427
rect 32413 12393 32447 12427
rect 32447 12393 32456 12427
rect 32404 12384 32456 12393
rect 32956 12384 33008 12436
rect 35256 12427 35308 12436
rect 35256 12393 35265 12427
rect 35265 12393 35299 12427
rect 35299 12393 35308 12427
rect 35256 12384 35308 12393
rect 35348 12384 35400 12436
rect 29092 12316 29144 12368
rect 32128 12316 32180 12368
rect 23664 12248 23716 12300
rect 24768 12248 24820 12300
rect 29000 12291 29052 12300
rect 29000 12257 29009 12291
rect 29009 12257 29043 12291
rect 29043 12257 29052 12291
rect 29000 12248 29052 12257
rect 10324 12223 10376 12232
rect 10324 12189 10333 12223
rect 10333 12189 10367 12223
rect 10367 12189 10376 12223
rect 10324 12180 10376 12189
rect 11244 12180 11296 12232
rect 11336 12180 11388 12232
rect 11888 12223 11940 12232
rect 11888 12189 11897 12223
rect 11897 12189 11931 12223
rect 11931 12189 11940 12223
rect 11888 12180 11940 12189
rect 15200 12180 15252 12232
rect 18144 12180 18196 12232
rect 19432 12180 19484 12232
rect 23480 12180 23532 12232
rect 25688 12180 25740 12232
rect 35716 12223 35768 12232
rect 35716 12189 35725 12223
rect 35725 12189 35759 12223
rect 35759 12189 35768 12223
rect 35716 12180 35768 12189
rect 35992 12180 36044 12232
rect 8024 12087 8076 12096
rect 8024 12053 8033 12087
rect 8033 12053 8067 12087
rect 8067 12053 8076 12087
rect 8024 12044 8076 12053
rect 13268 12087 13320 12096
rect 13268 12053 13277 12087
rect 13277 12053 13311 12087
rect 13311 12053 13320 12087
rect 13268 12044 13320 12053
rect 17868 12087 17920 12096
rect 17868 12053 17877 12087
rect 17877 12053 17911 12087
rect 17911 12053 17920 12087
rect 17868 12044 17920 12053
rect 19892 12044 19944 12096
rect 20904 12044 20956 12096
rect 25136 12087 25188 12096
rect 25136 12053 25145 12087
rect 25145 12053 25179 12087
rect 25179 12053 25188 12087
rect 25136 12044 25188 12053
rect 25320 12044 25372 12096
rect 28816 12087 28868 12096
rect 28816 12053 28825 12087
rect 28825 12053 28859 12087
rect 28859 12053 28868 12087
rect 28816 12044 28868 12053
rect 36820 12044 36872 12096
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 34966 11942 35018 11994
rect 35030 11942 35082 11994
rect 35094 11942 35146 11994
rect 35158 11942 35210 11994
rect 7012 11840 7064 11892
rect 8392 11840 8444 11892
rect 11244 11883 11296 11892
rect 11244 11849 11253 11883
rect 11253 11849 11287 11883
rect 11287 11849 11296 11883
rect 11244 11840 11296 11849
rect 11888 11883 11940 11892
rect 11888 11849 11897 11883
rect 11897 11849 11931 11883
rect 11931 11849 11940 11883
rect 11888 11840 11940 11849
rect 14832 11883 14884 11892
rect 14832 11849 14841 11883
rect 14841 11849 14875 11883
rect 14875 11849 14884 11883
rect 14832 11840 14884 11849
rect 16580 11840 16632 11892
rect 18236 11840 18288 11892
rect 18328 11840 18380 11892
rect 20904 11840 20956 11892
rect 23480 11840 23532 11892
rect 25320 11883 25372 11892
rect 25320 11849 25329 11883
rect 25329 11849 25363 11883
rect 25363 11849 25372 11883
rect 25320 11840 25372 11849
rect 26792 11840 26844 11892
rect 28264 11883 28316 11892
rect 28264 11849 28273 11883
rect 28273 11849 28307 11883
rect 28307 11849 28316 11883
rect 28264 11840 28316 11849
rect 28724 11883 28776 11892
rect 28724 11849 28733 11883
rect 28733 11849 28767 11883
rect 28767 11849 28776 11883
rect 28724 11840 28776 11849
rect 29000 11883 29052 11892
rect 29000 11849 29009 11883
rect 29009 11849 29043 11883
rect 29043 11849 29052 11883
rect 29000 11840 29052 11849
rect 35348 11840 35400 11892
rect 35992 11883 36044 11892
rect 35992 11849 36001 11883
rect 36001 11849 36035 11883
rect 36035 11849 36044 11883
rect 35992 11840 36044 11849
rect 16304 11772 16356 11824
rect 16672 11704 16724 11756
rect 6828 11679 6880 11688
rect 6828 11645 6837 11679
rect 6837 11645 6871 11679
rect 6871 11645 6880 11679
rect 6828 11636 6880 11645
rect 7932 11636 7984 11688
rect 13820 11636 13872 11688
rect 16212 11636 16264 11688
rect 6644 11568 6696 11620
rect 6920 11568 6972 11620
rect 9404 11568 9456 11620
rect 13268 11568 13320 11620
rect 17868 11636 17920 11688
rect 20260 11679 20312 11688
rect 20260 11645 20269 11679
rect 20269 11645 20303 11679
rect 20303 11645 20312 11679
rect 20260 11636 20312 11645
rect 21180 11636 21232 11688
rect 21916 11636 21968 11688
rect 23480 11679 23532 11688
rect 23480 11645 23489 11679
rect 23489 11645 23523 11679
rect 23523 11645 23532 11679
rect 23480 11636 23532 11645
rect 25688 11679 25740 11688
rect 25688 11645 25697 11679
rect 25697 11645 25731 11679
rect 25731 11645 25740 11679
rect 25688 11636 25740 11645
rect 35716 11704 35768 11756
rect 28724 11636 28776 11688
rect 19892 11611 19944 11620
rect 19892 11577 19901 11611
rect 19901 11577 19935 11611
rect 19935 11577 19944 11611
rect 19892 11568 19944 11577
rect 25136 11568 25188 11620
rect 28816 11568 28868 11620
rect 10692 11543 10744 11552
rect 10692 11509 10701 11543
rect 10701 11509 10735 11543
rect 10735 11509 10744 11543
rect 10692 11500 10744 11509
rect 13912 11500 13964 11552
rect 15200 11500 15252 11552
rect 15752 11543 15804 11552
rect 15752 11509 15761 11543
rect 15761 11509 15795 11543
rect 15795 11509 15804 11543
rect 15752 11500 15804 11509
rect 15936 11543 15988 11552
rect 15936 11509 15945 11543
rect 15945 11509 15979 11543
rect 15979 11509 15988 11543
rect 15936 11500 15988 11509
rect 16856 11500 16908 11552
rect 18236 11543 18288 11552
rect 18236 11509 18245 11543
rect 18245 11509 18279 11543
rect 18279 11509 18288 11543
rect 18236 11500 18288 11509
rect 20352 11543 20404 11552
rect 20352 11509 20361 11543
rect 20361 11509 20395 11543
rect 20395 11509 20404 11543
rect 20352 11500 20404 11509
rect 20444 11500 20496 11552
rect 20812 11500 20864 11552
rect 21364 11543 21416 11552
rect 21364 11509 21373 11543
rect 21373 11509 21407 11543
rect 21407 11509 21416 11543
rect 21364 11500 21416 11509
rect 29092 11500 29144 11552
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 8760 11296 8812 11348
rect 9404 11339 9456 11348
rect 9404 11305 9413 11339
rect 9413 11305 9447 11339
rect 9447 11305 9456 11339
rect 9404 11296 9456 11305
rect 10048 11296 10100 11348
rect 12440 11339 12492 11348
rect 12440 11305 12449 11339
rect 12449 11305 12483 11339
rect 12483 11305 12492 11339
rect 12440 11296 12492 11305
rect 13268 11296 13320 11348
rect 16856 11339 16908 11348
rect 16856 11305 16865 11339
rect 16865 11305 16899 11339
rect 16899 11305 16908 11339
rect 16856 11296 16908 11305
rect 17868 11296 17920 11348
rect 20352 11296 20404 11348
rect 20444 11296 20496 11348
rect 23664 11339 23716 11348
rect 23664 11305 23673 11339
rect 23673 11305 23707 11339
rect 23707 11305 23716 11339
rect 23664 11296 23716 11305
rect 24400 11339 24452 11348
rect 24400 11305 24409 11339
rect 24409 11305 24443 11339
rect 24443 11305 24452 11339
rect 24400 11296 24452 11305
rect 24860 11296 24912 11348
rect 25320 11296 25372 11348
rect 28816 11296 28868 11348
rect 29000 11296 29052 11348
rect 29368 11296 29420 11348
rect 30104 11339 30156 11348
rect 30104 11305 30113 11339
rect 30113 11305 30147 11339
rect 30147 11305 30156 11339
rect 30104 11296 30156 11305
rect 31760 11296 31812 11348
rect 6920 11228 6972 11280
rect 8024 11228 8076 11280
rect 10692 11228 10744 11280
rect 19708 11228 19760 11280
rect 21180 11271 21232 11280
rect 21180 11237 21214 11271
rect 21214 11237 21232 11271
rect 21180 11228 21232 11237
rect 23480 11228 23532 11280
rect 27896 11228 27948 11280
rect 6828 11135 6880 11144
rect 6828 11101 6837 11135
rect 6837 11101 6871 11135
rect 6871 11101 6880 11135
rect 7932 11160 7984 11212
rect 9956 11203 10008 11212
rect 9956 11169 9965 11203
rect 9965 11169 9999 11203
rect 9999 11169 10008 11203
rect 9956 11160 10008 11169
rect 11888 11160 11940 11212
rect 13544 11203 13596 11212
rect 13544 11169 13553 11203
rect 13553 11169 13587 11203
rect 13587 11169 13596 11203
rect 13544 11160 13596 11169
rect 15752 11203 15804 11212
rect 15752 11169 15786 11203
rect 15786 11169 15804 11203
rect 15752 11160 15804 11169
rect 18972 11160 19024 11212
rect 24492 11160 24544 11212
rect 25136 11160 25188 11212
rect 25688 11160 25740 11212
rect 27252 11160 27304 11212
rect 30012 11203 30064 11212
rect 30012 11169 30021 11203
rect 30021 11169 30055 11203
rect 30055 11169 30064 11203
rect 30012 11160 30064 11169
rect 32128 11203 32180 11212
rect 32128 11169 32137 11203
rect 32137 11169 32171 11203
rect 32171 11169 32180 11203
rect 32128 11160 32180 11169
rect 6828 11092 6880 11101
rect 15200 11092 15252 11144
rect 20904 11135 20956 11144
rect 20904 11101 20913 11135
rect 20913 11101 20947 11135
rect 20947 11101 20956 11135
rect 20904 11092 20956 11101
rect 25228 11092 25280 11144
rect 25964 11092 26016 11144
rect 29000 11092 29052 11144
rect 30196 11135 30248 11144
rect 30196 11101 30205 11135
rect 30205 11101 30239 11135
rect 30239 11101 30248 11135
rect 30196 11092 30248 11101
rect 10968 11024 11020 11076
rect 12532 11024 12584 11076
rect 18788 11024 18840 11076
rect 20352 11067 20404 11076
rect 20352 11033 20361 11067
rect 20361 11033 20395 11067
rect 20395 11033 20404 11067
rect 20352 11024 20404 11033
rect 32128 11024 32180 11076
rect 18144 10956 18196 11008
rect 19616 10999 19668 11008
rect 19616 10965 19625 10999
rect 19625 10965 19659 10999
rect 19659 10965 19668 10999
rect 19616 10956 19668 10965
rect 19984 10999 20036 11008
rect 19984 10965 19993 10999
rect 19993 10965 20027 10999
rect 20027 10965 20036 10999
rect 19984 10956 20036 10965
rect 35532 10999 35584 11008
rect 35532 10965 35541 10999
rect 35541 10965 35575 10999
rect 35575 10965 35584 10999
rect 35532 10956 35584 10965
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 34966 10854 35018 10906
rect 35030 10854 35082 10906
rect 35094 10854 35146 10906
rect 35158 10854 35210 10906
rect 6644 10795 6696 10804
rect 6644 10761 6653 10795
rect 6653 10761 6687 10795
rect 6687 10761 6696 10795
rect 7932 10795 7984 10804
rect 6644 10752 6696 10761
rect 6920 10684 6972 10736
rect 7932 10761 7941 10795
rect 7941 10761 7975 10795
rect 7975 10761 7984 10795
rect 7932 10752 7984 10761
rect 8300 10795 8352 10804
rect 8300 10761 8309 10795
rect 8309 10761 8343 10795
rect 8343 10761 8352 10795
rect 9956 10795 10008 10804
rect 8300 10752 8352 10761
rect 7380 10659 7432 10668
rect 7380 10625 7389 10659
rect 7389 10625 7423 10659
rect 7423 10625 7432 10659
rect 9956 10761 9965 10795
rect 9965 10761 9999 10795
rect 9999 10761 10008 10795
rect 9956 10752 10008 10761
rect 10692 10752 10744 10804
rect 11060 10752 11112 10804
rect 11704 10795 11756 10804
rect 11704 10761 11713 10795
rect 11713 10761 11747 10795
rect 11747 10761 11756 10795
rect 11704 10752 11756 10761
rect 11888 10752 11940 10804
rect 13544 10795 13596 10804
rect 13544 10761 13553 10795
rect 13553 10761 13587 10795
rect 13587 10761 13596 10795
rect 13544 10752 13596 10761
rect 15752 10752 15804 10804
rect 18972 10795 19024 10804
rect 18972 10761 18981 10795
rect 18981 10761 19015 10795
rect 19015 10761 19024 10795
rect 18972 10752 19024 10761
rect 20260 10795 20312 10804
rect 20260 10761 20269 10795
rect 20269 10761 20303 10795
rect 20303 10761 20312 10795
rect 20260 10752 20312 10761
rect 24492 10795 24544 10804
rect 24492 10761 24501 10795
rect 24501 10761 24535 10795
rect 24535 10761 24544 10795
rect 24492 10752 24544 10761
rect 24860 10795 24912 10804
rect 24860 10761 24869 10795
rect 24869 10761 24903 10795
rect 24903 10761 24912 10795
rect 24860 10752 24912 10761
rect 25228 10795 25280 10804
rect 25228 10761 25237 10795
rect 25237 10761 25271 10795
rect 25271 10761 25280 10795
rect 25228 10752 25280 10761
rect 25872 10795 25924 10804
rect 25872 10761 25881 10795
rect 25881 10761 25915 10795
rect 25915 10761 25924 10795
rect 25872 10752 25924 10761
rect 26240 10795 26292 10804
rect 26240 10761 26249 10795
rect 26249 10761 26283 10795
rect 26283 10761 26292 10795
rect 26240 10752 26292 10761
rect 18144 10684 18196 10736
rect 7380 10616 7432 10625
rect 8944 10659 8996 10668
rect 8944 10625 8953 10659
rect 8953 10625 8987 10659
rect 8987 10625 8996 10659
rect 8944 10616 8996 10625
rect 12440 10616 12492 10668
rect 12992 10616 13044 10668
rect 13268 10616 13320 10668
rect 15200 10616 15252 10668
rect 19708 10659 19760 10668
rect 19708 10625 19717 10659
rect 19717 10625 19751 10659
rect 19751 10625 19760 10659
rect 19708 10616 19760 10625
rect 19984 10684 20036 10736
rect 8760 10591 8812 10600
rect 8760 10557 8769 10591
rect 8769 10557 8803 10591
rect 8803 10557 8812 10591
rect 8760 10548 8812 10557
rect 10692 10548 10744 10600
rect 13728 10548 13780 10600
rect 19616 10591 19668 10600
rect 6552 10480 6604 10532
rect 6828 10455 6880 10464
rect 6828 10421 6837 10455
rect 6837 10421 6871 10455
rect 6871 10421 6880 10455
rect 6828 10412 6880 10421
rect 7012 10480 7064 10532
rect 7380 10412 7432 10464
rect 7656 10412 7708 10464
rect 16304 10480 16356 10532
rect 19616 10557 19625 10591
rect 19625 10557 19659 10591
rect 19659 10557 19668 10591
rect 19616 10548 19668 10557
rect 20076 10548 20128 10600
rect 20812 10591 20864 10600
rect 20812 10557 20821 10591
rect 20821 10557 20855 10591
rect 20855 10557 20864 10591
rect 20812 10548 20864 10557
rect 26240 10548 26292 10600
rect 27068 10752 27120 10804
rect 27160 10795 27212 10804
rect 27160 10761 27169 10795
rect 27169 10761 27203 10795
rect 27203 10761 27212 10795
rect 27896 10795 27948 10804
rect 27160 10752 27212 10761
rect 27896 10761 27905 10795
rect 27905 10761 27939 10795
rect 27939 10761 27948 10795
rect 27896 10752 27948 10761
rect 28908 10752 28960 10804
rect 29092 10795 29144 10804
rect 29092 10761 29101 10795
rect 29101 10761 29135 10795
rect 29135 10761 29144 10795
rect 29092 10752 29144 10761
rect 29368 10752 29420 10804
rect 32128 10795 32180 10804
rect 27252 10684 27304 10736
rect 28724 10727 28776 10736
rect 28724 10693 28733 10727
rect 28733 10693 28767 10727
rect 28767 10693 28776 10727
rect 28724 10684 28776 10693
rect 32128 10761 32137 10795
rect 32137 10761 32171 10795
rect 32171 10761 32180 10795
rect 32128 10752 32180 10761
rect 36820 10795 36872 10804
rect 36820 10761 36829 10795
rect 36829 10761 36863 10795
rect 36863 10761 36872 10795
rect 36820 10752 36872 10761
rect 29920 10548 29972 10600
rect 32312 10591 32364 10600
rect 32312 10557 32321 10591
rect 32321 10557 32355 10591
rect 32355 10557 32364 10591
rect 32312 10548 32364 10557
rect 30288 10480 30340 10532
rect 11336 10455 11388 10464
rect 11336 10421 11345 10455
rect 11345 10421 11379 10455
rect 11379 10421 11388 10455
rect 11336 10412 11388 10421
rect 12532 10412 12584 10464
rect 15200 10412 15252 10464
rect 18144 10412 18196 10464
rect 18696 10455 18748 10464
rect 18696 10421 18705 10455
rect 18705 10421 18739 10455
rect 18739 10421 18748 10455
rect 18696 10412 18748 10421
rect 19248 10455 19300 10464
rect 19248 10421 19257 10455
rect 19257 10421 19291 10455
rect 19291 10421 19300 10455
rect 19248 10412 19300 10421
rect 20904 10412 20956 10464
rect 21916 10412 21968 10464
rect 31208 10455 31260 10464
rect 31208 10421 31217 10455
rect 31217 10421 31251 10455
rect 31251 10421 31260 10455
rect 31208 10412 31260 10421
rect 32496 10455 32548 10464
rect 32496 10421 32505 10455
rect 32505 10421 32539 10455
rect 32539 10421 32548 10455
rect 32496 10412 32548 10421
rect 33324 10455 33376 10464
rect 33324 10421 33333 10455
rect 33333 10421 33367 10455
rect 33367 10421 33376 10455
rect 33324 10412 33376 10421
rect 35164 10412 35216 10464
rect 35532 10548 35584 10600
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 6552 10251 6604 10260
rect 6552 10217 6561 10251
rect 6561 10217 6595 10251
rect 6595 10217 6604 10251
rect 6552 10208 6604 10217
rect 6828 10208 6880 10260
rect 7104 10208 7156 10260
rect 7656 10251 7708 10260
rect 7656 10217 7665 10251
rect 7665 10217 7699 10251
rect 7699 10217 7708 10251
rect 7656 10208 7708 10217
rect 8760 10208 8812 10260
rect 10692 10208 10744 10260
rect 13268 10208 13320 10260
rect 15200 10208 15252 10260
rect 15752 10208 15804 10260
rect 15936 10208 15988 10260
rect 16580 10208 16632 10260
rect 18236 10208 18288 10260
rect 29460 10251 29512 10260
rect 29460 10217 29469 10251
rect 29469 10217 29503 10251
rect 29503 10217 29512 10251
rect 29460 10208 29512 10217
rect 30288 10208 30340 10260
rect 30380 10208 30432 10260
rect 31668 10208 31720 10260
rect 33232 10208 33284 10260
rect 33784 10208 33836 10260
rect 35532 10208 35584 10260
rect 11888 10140 11940 10192
rect 12992 10140 13044 10192
rect 20352 10140 20404 10192
rect 6828 10072 6880 10124
rect 7656 10072 7708 10124
rect 10416 10072 10468 10124
rect 14188 10072 14240 10124
rect 7012 10004 7064 10056
rect 7748 10004 7800 10056
rect 8300 10004 8352 10056
rect 10784 10047 10836 10056
rect 10784 10013 10793 10047
rect 10793 10013 10827 10047
rect 10827 10013 10836 10047
rect 10784 10004 10836 10013
rect 12164 10004 12216 10056
rect 7472 9936 7524 9988
rect 8944 9936 8996 9988
rect 14280 9979 14332 9988
rect 14280 9945 14289 9979
rect 14289 9945 14323 9979
rect 14323 9945 14332 9979
rect 14280 9936 14332 9945
rect 19248 10072 19300 10124
rect 28908 10115 28960 10124
rect 28908 10081 28917 10115
rect 28917 10081 28951 10115
rect 28951 10081 28960 10115
rect 28908 10072 28960 10081
rect 29828 10072 29880 10124
rect 32496 10072 32548 10124
rect 33048 10072 33100 10124
rect 34612 10072 34664 10124
rect 35164 10115 35216 10124
rect 35164 10081 35173 10115
rect 35173 10081 35207 10115
rect 35207 10081 35216 10115
rect 35164 10072 35216 10081
rect 35808 10072 35860 10124
rect 16488 10047 16540 10056
rect 16488 10013 16497 10047
rect 16497 10013 16531 10047
rect 16531 10013 16540 10047
rect 16488 10004 16540 10013
rect 18052 10047 18104 10056
rect 16120 9936 16172 9988
rect 18052 10013 18061 10047
rect 18061 10013 18095 10047
rect 18095 10013 18104 10047
rect 18052 10004 18104 10013
rect 18144 10047 18196 10056
rect 18144 10013 18153 10047
rect 18153 10013 18187 10047
rect 18187 10013 18196 10047
rect 18144 10004 18196 10013
rect 30564 10047 30616 10056
rect 30564 10013 30573 10047
rect 30573 10013 30607 10047
rect 30607 10013 30616 10047
rect 30564 10004 30616 10013
rect 31208 10004 31260 10056
rect 33324 10004 33376 10056
rect 34796 10004 34848 10056
rect 33232 9979 33284 9988
rect 33232 9945 33241 9979
rect 33241 9945 33275 9979
rect 33275 9945 33284 9979
rect 33232 9936 33284 9945
rect 7840 9868 7892 9920
rect 9680 9868 9732 9920
rect 12348 9868 12400 9920
rect 12900 9868 12952 9920
rect 17868 9868 17920 9920
rect 19248 9868 19300 9920
rect 19800 9911 19852 9920
rect 19800 9877 19809 9911
rect 19809 9877 19843 9911
rect 19843 9877 19852 9911
rect 19800 9868 19852 9877
rect 20168 9911 20220 9920
rect 20168 9877 20177 9911
rect 20177 9877 20211 9911
rect 20211 9877 20220 9911
rect 20168 9868 20220 9877
rect 20904 9868 20956 9920
rect 22008 9868 22060 9920
rect 25412 9911 25464 9920
rect 25412 9877 25421 9911
rect 25421 9877 25455 9911
rect 25455 9877 25464 9911
rect 25412 9868 25464 9877
rect 30012 9911 30064 9920
rect 30012 9877 30021 9911
rect 30021 9877 30055 9911
rect 30055 9877 30064 9911
rect 30012 9868 30064 9877
rect 32864 9911 32916 9920
rect 32864 9877 32873 9911
rect 32873 9877 32907 9911
rect 32907 9877 32916 9911
rect 32864 9868 32916 9877
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 34966 9766 35018 9818
rect 35030 9766 35082 9818
rect 35094 9766 35146 9818
rect 35158 9766 35210 9818
rect 7104 9664 7156 9716
rect 7472 9664 7524 9716
rect 10784 9707 10836 9716
rect 10784 9673 10793 9707
rect 10793 9673 10827 9707
rect 10827 9673 10836 9707
rect 10784 9664 10836 9673
rect 14188 9707 14240 9716
rect 14188 9673 14197 9707
rect 14197 9673 14231 9707
rect 14231 9673 14240 9707
rect 14188 9664 14240 9673
rect 6828 9596 6880 9648
rect 8300 9596 8352 9648
rect 9588 9596 9640 9648
rect 13912 9639 13964 9648
rect 13912 9605 13921 9639
rect 13921 9605 13955 9639
rect 13955 9605 13964 9639
rect 13912 9596 13964 9605
rect 16120 9664 16172 9716
rect 18236 9707 18288 9716
rect 18236 9673 18245 9707
rect 18245 9673 18279 9707
rect 18279 9673 18288 9707
rect 18236 9664 18288 9673
rect 20076 9707 20128 9716
rect 20076 9673 20085 9707
rect 20085 9673 20119 9707
rect 20119 9673 20128 9707
rect 20076 9664 20128 9673
rect 28908 9707 28960 9716
rect 28908 9673 28917 9707
rect 28917 9673 28951 9707
rect 28951 9673 28960 9707
rect 28908 9664 28960 9673
rect 29828 9707 29880 9716
rect 29828 9673 29837 9707
rect 29837 9673 29871 9707
rect 29871 9673 29880 9707
rect 29828 9664 29880 9673
rect 32496 9664 32548 9716
rect 33784 9707 33836 9716
rect 33784 9673 33793 9707
rect 33793 9673 33827 9707
rect 33827 9673 33836 9707
rect 33784 9664 33836 9673
rect 17592 9639 17644 9648
rect 17592 9605 17601 9639
rect 17601 9605 17635 9639
rect 17635 9605 17644 9639
rect 17592 9596 17644 9605
rect 18788 9639 18840 9648
rect 18788 9605 18797 9639
rect 18797 9605 18831 9639
rect 18831 9605 18840 9639
rect 18788 9596 18840 9605
rect 20352 9596 20404 9648
rect 11428 9571 11480 9580
rect 11428 9537 11437 9571
rect 11437 9537 11471 9571
rect 11471 9537 11480 9571
rect 11428 9528 11480 9537
rect 12624 9528 12676 9580
rect 12900 9571 12952 9580
rect 12900 9537 12909 9571
rect 12909 9537 12943 9571
rect 12943 9537 12952 9571
rect 12900 9528 12952 9537
rect 13084 9571 13136 9580
rect 13084 9537 13093 9571
rect 13093 9537 13127 9571
rect 13127 9537 13136 9571
rect 13084 9528 13136 9537
rect 12256 9460 12308 9512
rect 9404 9392 9456 9444
rect 10876 9392 10928 9444
rect 12532 9392 12584 9444
rect 10416 9324 10468 9376
rect 11244 9367 11296 9376
rect 11244 9333 11253 9367
rect 11253 9333 11287 9367
rect 11287 9333 11296 9367
rect 11888 9367 11940 9376
rect 11244 9324 11296 9333
rect 11888 9333 11897 9367
rect 11897 9333 11931 9367
rect 11931 9333 11940 9367
rect 11888 9324 11940 9333
rect 12164 9367 12216 9376
rect 12164 9333 12173 9367
rect 12173 9333 12207 9367
rect 12207 9333 12216 9367
rect 12164 9324 12216 9333
rect 12716 9324 12768 9376
rect 15016 9367 15068 9376
rect 15016 9333 15025 9367
rect 15025 9333 15059 9367
rect 15059 9333 15068 9367
rect 15016 9324 15068 9333
rect 15200 9324 15252 9376
rect 19248 9503 19300 9512
rect 19248 9469 19257 9503
rect 19257 9469 19291 9503
rect 19291 9469 19300 9503
rect 19248 9460 19300 9469
rect 19800 9528 19852 9580
rect 32496 9528 32548 9580
rect 20904 9503 20956 9512
rect 15752 9435 15804 9444
rect 15752 9401 15786 9435
rect 15786 9401 15804 9435
rect 15752 9392 15804 9401
rect 18144 9392 18196 9444
rect 20904 9469 20913 9503
rect 20913 9469 20947 9503
rect 20947 9469 20956 9503
rect 20904 9460 20956 9469
rect 20168 9392 20220 9444
rect 22008 9460 22060 9512
rect 16304 9324 16356 9376
rect 18880 9367 18932 9376
rect 18880 9333 18889 9367
rect 18889 9333 18923 9367
rect 18923 9333 18932 9367
rect 18880 9324 18932 9333
rect 20444 9367 20496 9376
rect 20444 9333 20453 9367
rect 20453 9333 20487 9367
rect 20487 9333 20496 9367
rect 20444 9324 20496 9333
rect 22284 9367 22336 9376
rect 22284 9333 22293 9367
rect 22293 9333 22327 9367
rect 22327 9333 22336 9367
rect 22284 9324 22336 9333
rect 25412 9460 25464 9512
rect 29920 9460 29972 9512
rect 32312 9503 32364 9512
rect 29736 9392 29788 9444
rect 30564 9435 30616 9444
rect 30564 9401 30576 9435
rect 30576 9401 30616 9435
rect 30564 9392 30616 9401
rect 26516 9324 26568 9376
rect 26700 9367 26752 9376
rect 26700 9333 26709 9367
rect 26709 9333 26743 9367
rect 26743 9333 26752 9367
rect 26700 9324 26752 9333
rect 32312 9469 32321 9503
rect 32321 9469 32355 9503
rect 32355 9469 32364 9503
rect 32312 9460 32364 9469
rect 34520 9460 34572 9512
rect 34888 9503 34940 9512
rect 34888 9469 34897 9503
rect 34897 9469 34931 9503
rect 34931 9469 34940 9503
rect 34888 9460 34940 9469
rect 32864 9392 32916 9444
rect 31024 9324 31076 9376
rect 31116 9324 31168 9376
rect 32956 9324 33008 9376
rect 34428 9392 34480 9444
rect 34796 9392 34848 9444
rect 33324 9324 33376 9376
rect 34612 9324 34664 9376
rect 34888 9324 34940 9376
rect 36268 9367 36320 9376
rect 36268 9333 36277 9367
rect 36277 9333 36311 9367
rect 36311 9333 36320 9367
rect 36268 9324 36320 9333
rect 36820 9367 36872 9376
rect 36820 9333 36829 9367
rect 36829 9333 36863 9367
rect 36863 9333 36872 9367
rect 36820 9324 36872 9333
rect 37096 9324 37148 9376
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 11244 9120 11296 9172
rect 12440 9120 12492 9172
rect 13176 9120 13228 9172
rect 14188 9163 14240 9172
rect 14188 9129 14197 9163
rect 14197 9129 14231 9163
rect 14231 9129 14240 9163
rect 14188 9120 14240 9129
rect 15016 9120 15068 9172
rect 16488 9120 16540 9172
rect 16580 9120 16632 9172
rect 17960 9120 18012 9172
rect 18328 9120 18380 9172
rect 19340 9163 19392 9172
rect 13084 9052 13136 9104
rect 16304 9095 16356 9104
rect 16304 9061 16313 9095
rect 16313 9061 16347 9095
rect 16347 9061 16356 9095
rect 16304 9052 16356 9061
rect 19340 9129 19349 9163
rect 19349 9129 19383 9163
rect 19383 9129 19392 9163
rect 19340 9120 19392 9129
rect 20168 9120 20220 9172
rect 25412 9120 25464 9172
rect 29736 9163 29788 9172
rect 29736 9129 29745 9163
rect 29745 9129 29779 9163
rect 29779 9129 29788 9163
rect 29736 9120 29788 9129
rect 30288 9120 30340 9172
rect 32312 9120 32364 9172
rect 32680 9120 32732 9172
rect 33140 9120 33192 9172
rect 33784 9120 33836 9172
rect 35992 9163 36044 9172
rect 35992 9129 36001 9163
rect 36001 9129 36035 9163
rect 36035 9129 36044 9163
rect 35992 9120 36044 9129
rect 19432 9052 19484 9104
rect 20444 9052 20496 9104
rect 21364 9052 21416 9104
rect 22284 9052 22336 9104
rect 26700 9052 26752 9104
rect 30012 9052 30064 9104
rect 6920 9027 6972 9036
rect 6920 8993 6929 9027
rect 6929 8993 6963 9027
rect 6963 8993 6972 9027
rect 7196 9027 7248 9036
rect 6920 8984 6972 8993
rect 7196 8993 7230 9027
rect 7230 8993 7248 9027
rect 7196 8984 7248 8993
rect 11704 9027 11756 9036
rect 11704 8993 11713 9027
rect 11713 8993 11747 9027
rect 11747 8993 11756 9027
rect 11704 8984 11756 8993
rect 17960 8984 18012 9036
rect 18880 8984 18932 9036
rect 30840 9027 30892 9036
rect 30840 8993 30849 9027
rect 30849 8993 30883 9027
rect 30883 8993 30892 9027
rect 30840 8984 30892 8993
rect 32404 9027 32456 9036
rect 32404 8993 32413 9027
rect 32413 8993 32447 9027
rect 32447 8993 32456 9027
rect 32404 8984 32456 8993
rect 37096 8984 37148 9036
rect 10140 8916 10192 8968
rect 15752 8916 15804 8968
rect 16488 8916 16540 8968
rect 16672 8916 16724 8968
rect 18788 8959 18840 8968
rect 18788 8925 18797 8959
rect 18797 8925 18831 8959
rect 18831 8925 18840 8959
rect 18788 8916 18840 8925
rect 20904 8959 20956 8968
rect 20904 8925 20913 8959
rect 20913 8925 20947 8959
rect 20947 8925 20956 8959
rect 20904 8916 20956 8925
rect 17868 8848 17920 8900
rect 26516 8959 26568 8968
rect 26516 8925 26525 8959
rect 26525 8925 26559 8959
rect 26559 8925 26568 8959
rect 26516 8916 26568 8925
rect 31116 8959 31168 8968
rect 31116 8925 31125 8959
rect 31125 8925 31159 8959
rect 31159 8925 31168 8959
rect 31116 8916 31168 8925
rect 33048 8959 33100 8968
rect 33048 8925 33057 8959
rect 33057 8925 33091 8959
rect 33091 8925 33100 8959
rect 33048 8916 33100 8925
rect 33324 8959 33376 8968
rect 33324 8925 33333 8959
rect 33333 8925 33367 8959
rect 33367 8925 33376 8959
rect 33324 8916 33376 8925
rect 34612 8916 34664 8968
rect 35716 8916 35768 8968
rect 36268 8916 36320 8968
rect 8300 8823 8352 8832
rect 8300 8789 8309 8823
rect 8309 8789 8343 8823
rect 8343 8789 8352 8823
rect 8300 8780 8352 8789
rect 11428 8780 11480 8832
rect 13728 8780 13780 8832
rect 18144 8823 18196 8832
rect 18144 8789 18153 8823
rect 18153 8789 18187 8823
rect 18187 8789 18196 8823
rect 18144 8780 18196 8789
rect 22284 8823 22336 8832
rect 22284 8789 22293 8823
rect 22293 8789 22327 8823
rect 22327 8789 22336 8823
rect 22284 8780 22336 8789
rect 24308 8823 24360 8832
rect 24308 8789 24317 8823
rect 24317 8789 24351 8823
rect 24351 8789 24360 8823
rect 24308 8780 24360 8789
rect 24768 8823 24820 8832
rect 24768 8789 24777 8823
rect 24777 8789 24811 8823
rect 24811 8789 24820 8823
rect 24768 8780 24820 8789
rect 25320 8780 25372 8832
rect 26884 8780 26936 8832
rect 34796 8780 34848 8832
rect 35440 8780 35492 8832
rect 35716 8780 35768 8832
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 34966 8678 35018 8730
rect 35030 8678 35082 8730
rect 35094 8678 35146 8730
rect 35158 8678 35210 8730
rect 7196 8576 7248 8628
rect 11244 8619 11296 8628
rect 11244 8585 11253 8619
rect 11253 8585 11287 8619
rect 11287 8585 11296 8619
rect 11244 8576 11296 8585
rect 12164 8576 12216 8628
rect 12624 8576 12676 8628
rect 16304 8619 16356 8628
rect 16304 8585 16313 8619
rect 16313 8585 16347 8619
rect 16347 8585 16356 8619
rect 16304 8576 16356 8585
rect 18328 8619 18380 8628
rect 18328 8585 18337 8619
rect 18337 8585 18371 8619
rect 18371 8585 18380 8619
rect 18328 8576 18380 8585
rect 19340 8576 19392 8628
rect 21364 8619 21416 8628
rect 21364 8585 21373 8619
rect 21373 8585 21407 8619
rect 21407 8585 21416 8619
rect 21364 8576 21416 8585
rect 25412 8576 25464 8628
rect 27620 8576 27672 8628
rect 30012 8619 30064 8628
rect 30012 8585 30021 8619
rect 30021 8585 30055 8619
rect 30055 8585 30064 8619
rect 30012 8576 30064 8585
rect 12256 8551 12308 8560
rect 12256 8517 12265 8551
rect 12265 8517 12299 8551
rect 12299 8517 12308 8551
rect 12256 8508 12308 8517
rect 16672 8508 16724 8560
rect 4712 8483 4764 8492
rect 4712 8449 4721 8483
rect 4721 8449 4755 8483
rect 4755 8449 4764 8483
rect 4712 8440 4764 8449
rect 12900 8440 12952 8492
rect 13176 8483 13228 8492
rect 13176 8449 13185 8483
rect 13185 8449 13219 8483
rect 13219 8449 13228 8483
rect 13176 8440 13228 8449
rect 13452 8483 13504 8492
rect 13452 8449 13461 8483
rect 13461 8449 13495 8483
rect 13495 8449 13504 8483
rect 13452 8440 13504 8449
rect 30840 8576 30892 8628
rect 32496 8619 32548 8628
rect 32496 8585 32505 8619
rect 32505 8585 32539 8619
rect 32539 8585 32548 8619
rect 32496 8576 32548 8585
rect 33048 8576 33100 8628
rect 35808 8576 35860 8628
rect 36820 8576 36872 8628
rect 37096 8619 37148 8628
rect 37096 8585 37105 8619
rect 37105 8585 37139 8619
rect 37139 8585 37148 8619
rect 37096 8576 37148 8585
rect 31024 8483 31076 8492
rect 31024 8449 31033 8483
rect 31033 8449 31067 8483
rect 31067 8449 31076 8483
rect 31024 8440 31076 8449
rect 5356 8372 5408 8424
rect 3056 8304 3108 8356
rect 5448 8304 5500 8356
rect 4068 8279 4120 8288
rect 4068 8245 4077 8279
rect 4077 8245 4111 8279
rect 4111 8245 4120 8279
rect 4068 8236 4120 8245
rect 6920 8372 6972 8424
rect 10508 8372 10560 8424
rect 11704 8372 11756 8424
rect 12808 8372 12860 8424
rect 7288 8304 7340 8356
rect 9956 8304 10008 8356
rect 11428 8304 11480 8356
rect 16488 8304 16540 8356
rect 17960 8372 18012 8424
rect 18052 8372 18104 8424
rect 18328 8304 18380 8356
rect 19340 8347 19392 8356
rect 19340 8313 19374 8347
rect 19374 8313 19392 8347
rect 19340 8304 19392 8313
rect 20904 8304 20956 8356
rect 6368 8236 6420 8288
rect 6552 8279 6604 8288
rect 6552 8245 6561 8279
rect 6561 8245 6595 8279
rect 6595 8245 6604 8279
rect 6552 8236 6604 8245
rect 7932 8236 7984 8288
rect 23480 8304 23532 8356
rect 24308 8372 24360 8424
rect 16672 8236 16724 8288
rect 22100 8236 22152 8288
rect 26884 8304 26936 8356
rect 33140 8347 33192 8356
rect 33140 8313 33149 8347
rect 33149 8313 33183 8347
rect 33183 8313 33192 8347
rect 33140 8304 33192 8313
rect 34336 8304 34388 8356
rect 26516 8279 26568 8288
rect 26516 8245 26525 8279
rect 26525 8245 26559 8279
rect 26559 8245 26568 8279
rect 26516 8236 26568 8245
rect 31116 8236 31168 8288
rect 33600 8279 33652 8288
rect 33600 8245 33609 8279
rect 33609 8245 33643 8279
rect 33643 8245 33652 8279
rect 33600 8236 33652 8245
rect 33968 8236 34020 8288
rect 34796 8304 34848 8356
rect 35164 8372 35216 8424
rect 36268 8372 36320 8424
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 6368 8075 6420 8084
rect 6368 8041 6377 8075
rect 6377 8041 6411 8075
rect 6411 8041 6420 8075
rect 6368 8032 6420 8041
rect 7932 8075 7984 8084
rect 7932 8041 7941 8075
rect 7941 8041 7975 8075
rect 7975 8041 7984 8075
rect 7932 8032 7984 8041
rect 9956 8075 10008 8084
rect 9956 8041 9965 8075
rect 9965 8041 9999 8075
rect 9999 8041 10008 8075
rect 9956 8032 10008 8041
rect 12808 8075 12860 8084
rect 12808 8041 12817 8075
rect 12817 8041 12851 8075
rect 12851 8041 12860 8075
rect 12808 8032 12860 8041
rect 16672 8075 16724 8084
rect 16672 8041 16681 8075
rect 16681 8041 16715 8075
rect 16715 8041 16724 8075
rect 16672 8032 16724 8041
rect 21088 8075 21140 8084
rect 21088 8041 21097 8075
rect 21097 8041 21131 8075
rect 21131 8041 21140 8075
rect 21088 8032 21140 8041
rect 24308 8032 24360 8084
rect 24676 8032 24728 8084
rect 25412 8075 25464 8084
rect 25412 8041 25421 8075
rect 25421 8041 25455 8075
rect 25455 8041 25464 8075
rect 25412 8032 25464 8041
rect 26700 8032 26752 8084
rect 26884 8032 26936 8084
rect 31116 8075 31168 8084
rect 31116 8041 31125 8075
rect 31125 8041 31159 8075
rect 31159 8041 31168 8075
rect 31116 8032 31168 8041
rect 34428 8032 34480 8084
rect 35164 8032 35216 8084
rect 12716 7964 12768 8016
rect 13452 8007 13504 8016
rect 13452 7973 13461 8007
rect 13461 7973 13495 8007
rect 13495 7973 13504 8007
rect 13452 7964 13504 7973
rect 15476 7964 15528 8016
rect 17408 8007 17460 8016
rect 17408 7973 17417 8007
rect 17417 7973 17451 8007
rect 17451 7973 17460 8007
rect 17408 7964 17460 7973
rect 19340 7964 19392 8016
rect 20444 7964 20496 8016
rect 23572 7964 23624 8016
rect 26976 8007 27028 8016
rect 26976 7973 26985 8007
rect 26985 7973 27019 8007
rect 27019 7973 27028 8007
rect 26976 7964 27028 7973
rect 27528 7964 27580 8016
rect 34520 7964 34572 8016
rect 35992 8032 36044 8084
rect 5264 7939 5316 7948
rect 5264 7905 5298 7939
rect 5298 7905 5316 7939
rect 5264 7896 5316 7905
rect 8208 7896 8260 7948
rect 4988 7871 5040 7880
rect 4988 7837 4997 7871
rect 4997 7837 5031 7871
rect 5031 7837 5040 7871
rect 4988 7828 5040 7837
rect 10508 7871 10560 7880
rect 7380 7760 7432 7812
rect 10508 7837 10517 7871
rect 10517 7837 10551 7871
rect 10551 7837 10560 7871
rect 10508 7828 10560 7837
rect 12164 7896 12216 7948
rect 18236 7939 18288 7948
rect 18236 7905 18245 7939
rect 18245 7905 18279 7939
rect 18279 7905 18288 7939
rect 18236 7896 18288 7905
rect 19524 7939 19576 7948
rect 19524 7905 19533 7939
rect 19533 7905 19567 7939
rect 19567 7905 19576 7939
rect 19524 7896 19576 7905
rect 21456 7896 21508 7948
rect 23480 7896 23532 7948
rect 28540 7939 28592 7948
rect 28540 7905 28574 7939
rect 28574 7905 28592 7939
rect 28540 7896 28592 7905
rect 33508 7896 33560 7948
rect 35256 7896 35308 7948
rect 13728 7828 13780 7880
rect 15200 7828 15252 7880
rect 17040 7828 17092 7880
rect 18512 7871 18564 7880
rect 18512 7837 18521 7871
rect 18521 7837 18555 7871
rect 18555 7837 18564 7871
rect 18512 7828 18564 7837
rect 19248 7828 19300 7880
rect 27160 7871 27212 7880
rect 27160 7837 27169 7871
rect 27169 7837 27203 7871
rect 27203 7837 27212 7871
rect 27160 7828 27212 7837
rect 28080 7828 28132 7880
rect 32680 7871 32732 7880
rect 32680 7837 32689 7871
rect 32689 7837 32723 7871
rect 32723 7837 32732 7871
rect 32680 7828 32732 7837
rect 12900 7760 12952 7812
rect 3056 7735 3108 7744
rect 3056 7701 3065 7735
rect 3065 7701 3099 7735
rect 3099 7701 3108 7735
rect 3056 7692 3108 7701
rect 4712 7692 4764 7744
rect 5172 7692 5224 7744
rect 6552 7692 6604 7744
rect 7288 7735 7340 7744
rect 7288 7701 7297 7735
rect 7297 7701 7331 7735
rect 7331 7701 7340 7735
rect 7288 7692 7340 7701
rect 7472 7735 7524 7744
rect 7472 7701 7481 7735
rect 7481 7701 7515 7735
rect 7515 7701 7524 7735
rect 7472 7692 7524 7701
rect 12348 7692 12400 7744
rect 12992 7735 13044 7744
rect 12992 7701 13001 7735
rect 13001 7701 13035 7735
rect 13035 7701 13044 7735
rect 12992 7692 13044 7701
rect 17776 7692 17828 7744
rect 26608 7735 26660 7744
rect 26608 7701 26617 7735
rect 26617 7701 26651 7735
rect 26651 7701 26660 7735
rect 26608 7692 26660 7701
rect 29644 7735 29696 7744
rect 29644 7701 29653 7735
rect 29653 7701 29687 7735
rect 29687 7701 29696 7735
rect 29644 7692 29696 7701
rect 32128 7692 32180 7744
rect 34796 7760 34848 7812
rect 35808 7760 35860 7812
rect 33968 7692 34020 7744
rect 35440 7735 35492 7744
rect 35440 7701 35449 7735
rect 35449 7701 35483 7735
rect 35483 7701 35492 7735
rect 35440 7692 35492 7701
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 34966 7590 35018 7642
rect 35030 7590 35082 7642
rect 35094 7590 35146 7642
rect 35158 7590 35210 7642
rect 5264 7488 5316 7540
rect 7932 7488 7984 7540
rect 10048 7488 10100 7540
rect 10508 7488 10560 7540
rect 10876 7488 10928 7540
rect 12164 7531 12216 7540
rect 12164 7497 12173 7531
rect 12173 7497 12207 7531
rect 12207 7497 12216 7531
rect 12164 7488 12216 7497
rect 12808 7531 12860 7540
rect 12808 7497 12817 7531
rect 12817 7497 12851 7531
rect 12851 7497 12860 7531
rect 12808 7488 12860 7497
rect 17040 7531 17092 7540
rect 17040 7497 17049 7531
rect 17049 7497 17083 7531
rect 17083 7497 17092 7531
rect 17040 7488 17092 7497
rect 18236 7488 18288 7540
rect 19524 7488 19576 7540
rect 20076 7488 20128 7540
rect 20444 7531 20496 7540
rect 20444 7497 20453 7531
rect 20453 7497 20487 7531
rect 20487 7497 20496 7531
rect 20444 7488 20496 7497
rect 20720 7531 20772 7540
rect 20720 7497 20729 7531
rect 20729 7497 20763 7531
rect 20763 7497 20772 7531
rect 20720 7488 20772 7497
rect 21456 7531 21508 7540
rect 21456 7497 21465 7531
rect 21465 7497 21499 7531
rect 21499 7497 21508 7531
rect 21456 7488 21508 7497
rect 22100 7488 22152 7540
rect 23480 7531 23532 7540
rect 23480 7497 23489 7531
rect 23489 7497 23523 7531
rect 23523 7497 23532 7531
rect 23480 7488 23532 7497
rect 26884 7488 26936 7540
rect 33508 7531 33560 7540
rect 33508 7497 33517 7531
rect 33517 7497 33551 7531
rect 33551 7497 33560 7531
rect 33508 7488 33560 7497
rect 37280 7531 37332 7540
rect 37280 7497 37289 7531
rect 37289 7497 37323 7531
rect 37323 7497 37332 7531
rect 37280 7488 37332 7497
rect 11704 7463 11756 7472
rect 11704 7429 11713 7463
rect 11713 7429 11747 7463
rect 11747 7429 11756 7463
rect 11704 7420 11756 7429
rect 11980 7420 12032 7472
rect 13360 7395 13412 7404
rect 13360 7361 13369 7395
rect 13369 7361 13403 7395
rect 13403 7361 13412 7395
rect 13360 7352 13412 7361
rect 3056 7284 3108 7336
rect 5540 7284 5592 7336
rect 6552 7284 6604 7336
rect 3976 7216 4028 7268
rect 4988 7259 5040 7268
rect 4988 7225 4997 7259
rect 4997 7225 5031 7259
rect 5031 7225 5040 7259
rect 4988 7216 5040 7225
rect 7932 7216 7984 7268
rect 12348 7284 12400 7336
rect 12900 7327 12952 7336
rect 12900 7293 12909 7327
rect 12909 7293 12943 7327
rect 12943 7293 12952 7327
rect 12900 7284 12952 7293
rect 17868 7420 17920 7472
rect 18052 7395 18104 7404
rect 12624 7216 12676 7268
rect 15200 7216 15252 7268
rect 18052 7361 18061 7395
rect 18061 7361 18095 7395
rect 18095 7361 18104 7395
rect 18052 7352 18104 7361
rect 19432 7284 19484 7336
rect 32128 7395 32180 7404
rect 32128 7361 32137 7395
rect 32137 7361 32171 7395
rect 32171 7361 32180 7395
rect 32128 7352 32180 7361
rect 34244 7352 34296 7404
rect 35164 7352 35216 7404
rect 35808 7352 35860 7404
rect 26976 7327 27028 7336
rect 26976 7293 27010 7327
rect 27010 7293 27028 7327
rect 17868 7216 17920 7268
rect 18512 7216 18564 7268
rect 23940 7259 23992 7268
rect 23940 7225 23974 7259
rect 23974 7225 23992 7259
rect 23940 7216 23992 7225
rect 26516 7216 26568 7268
rect 26976 7284 27028 7293
rect 28080 7284 28132 7336
rect 35256 7284 35308 7336
rect 36176 7327 36228 7336
rect 36176 7293 36185 7327
rect 36185 7293 36219 7327
rect 36219 7293 36228 7327
rect 36176 7284 36228 7293
rect 2504 7191 2556 7200
rect 2504 7157 2513 7191
rect 2513 7157 2547 7191
rect 2547 7157 2556 7191
rect 2504 7148 2556 7157
rect 2780 7191 2832 7200
rect 2780 7157 2789 7191
rect 2789 7157 2823 7191
rect 2823 7157 2832 7191
rect 2780 7148 2832 7157
rect 4160 7148 4212 7200
rect 5816 7191 5868 7200
rect 5816 7157 5825 7191
rect 5825 7157 5859 7191
rect 5859 7157 5868 7191
rect 5816 7148 5868 7157
rect 6552 7191 6604 7200
rect 6552 7157 6561 7191
rect 6561 7157 6595 7191
rect 6595 7157 6604 7191
rect 6552 7148 6604 7157
rect 8208 7191 8260 7200
rect 8208 7157 8217 7191
rect 8217 7157 8251 7191
rect 8251 7157 8260 7191
rect 8208 7148 8260 7157
rect 11152 7191 11204 7200
rect 11152 7157 11161 7191
rect 11161 7157 11195 7191
rect 11195 7157 11204 7191
rect 11152 7148 11204 7157
rect 14740 7191 14792 7200
rect 14740 7157 14749 7191
rect 14749 7157 14783 7191
rect 14783 7157 14792 7191
rect 14740 7148 14792 7157
rect 15476 7148 15528 7200
rect 19432 7191 19484 7200
rect 19432 7157 19441 7191
rect 19441 7157 19475 7191
rect 19475 7157 19484 7191
rect 19432 7148 19484 7157
rect 22468 7148 22520 7200
rect 22652 7191 22704 7200
rect 22652 7157 22661 7191
rect 22661 7157 22695 7191
rect 22695 7157 22704 7191
rect 22652 7148 22704 7157
rect 23572 7148 23624 7200
rect 27988 7148 28040 7200
rect 28540 7216 28592 7268
rect 32496 7216 32548 7268
rect 28908 7148 28960 7200
rect 33968 7148 34020 7200
rect 34520 7148 34572 7200
rect 35072 7148 35124 7200
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 2504 6944 2556 6996
rect 5448 6987 5500 6996
rect 5448 6953 5457 6987
rect 5457 6953 5491 6987
rect 5491 6953 5500 6987
rect 5448 6944 5500 6953
rect 11428 6987 11480 6996
rect 11428 6953 11437 6987
rect 11437 6953 11471 6987
rect 11471 6953 11480 6987
rect 11428 6944 11480 6953
rect 12624 6944 12676 6996
rect 13176 6944 13228 6996
rect 14740 6944 14792 6996
rect 15200 6944 15252 6996
rect 25504 6944 25556 6996
rect 26608 6944 26660 6996
rect 26976 6944 27028 6996
rect 33048 6944 33100 6996
rect 33600 6944 33652 6996
rect 34796 6987 34848 6996
rect 34796 6953 34805 6987
rect 34805 6953 34839 6987
rect 34839 6953 34848 6987
rect 34796 6944 34848 6953
rect 35440 6944 35492 6996
rect 2596 6808 2648 6860
rect 4160 6876 4212 6928
rect 4712 6808 4764 6860
rect 5356 6808 5408 6860
rect 6644 6808 6696 6860
rect 8300 6808 8352 6860
rect 10048 6851 10100 6860
rect 10048 6817 10057 6851
rect 10057 6817 10091 6851
rect 10091 6817 10100 6851
rect 10048 6808 10100 6817
rect 10692 6808 10744 6860
rect 11152 6876 11204 6928
rect 11980 6876 12032 6928
rect 11796 6808 11848 6860
rect 13360 6808 13412 6860
rect 13820 6808 13872 6860
rect 17500 6808 17552 6860
rect 35164 6876 35216 6928
rect 17960 6808 18012 6860
rect 19984 6808 20036 6860
rect 22376 6851 22428 6860
rect 22376 6817 22410 6851
rect 22410 6817 22428 6851
rect 22376 6808 22428 6817
rect 25320 6851 25372 6860
rect 25320 6817 25329 6851
rect 25329 6817 25363 6851
rect 25363 6817 25372 6851
rect 25320 6808 25372 6817
rect 26976 6808 27028 6860
rect 29000 6808 29052 6860
rect 29644 6808 29696 6860
rect 32956 6808 33008 6860
rect 33600 6808 33652 6860
rect 35624 6851 35676 6860
rect 35624 6817 35633 6851
rect 35633 6817 35667 6851
rect 35667 6817 35676 6851
rect 35624 6808 35676 6817
rect 3976 6740 4028 6792
rect 6552 6783 6604 6792
rect 6552 6749 6561 6783
rect 6561 6749 6595 6783
rect 6595 6749 6604 6783
rect 6552 6740 6604 6749
rect 12440 6740 12492 6792
rect 12808 6740 12860 6792
rect 13728 6740 13780 6792
rect 15292 6783 15344 6792
rect 15292 6749 15301 6783
rect 15301 6749 15335 6783
rect 15335 6749 15344 6783
rect 15292 6740 15344 6749
rect 17868 6740 17920 6792
rect 5080 6672 5132 6724
rect 6368 6715 6420 6724
rect 6368 6681 6377 6715
rect 6377 6681 6411 6715
rect 6411 6681 6420 6715
rect 6368 6672 6420 6681
rect 17776 6672 17828 6724
rect 17960 6672 18012 6724
rect 18420 6740 18472 6792
rect 19432 6740 19484 6792
rect 21916 6740 21968 6792
rect 22100 6783 22152 6792
rect 22100 6749 22109 6783
rect 22109 6749 22143 6783
rect 22143 6749 22152 6783
rect 25412 6783 25464 6792
rect 22100 6740 22152 6749
rect 25412 6749 25421 6783
rect 25421 6749 25455 6783
rect 25455 6749 25464 6783
rect 25412 6740 25464 6749
rect 28080 6740 28132 6792
rect 33508 6783 33560 6792
rect 33508 6749 33517 6783
rect 33517 6749 33551 6783
rect 33551 6749 33560 6783
rect 33508 6740 33560 6749
rect 35532 6740 35584 6792
rect 2412 6647 2464 6656
rect 2412 6613 2421 6647
rect 2421 6613 2455 6647
rect 2455 6613 2464 6647
rect 2412 6604 2464 6613
rect 3516 6647 3568 6656
rect 3516 6613 3525 6647
rect 3525 6613 3559 6647
rect 3559 6613 3568 6647
rect 3516 6604 3568 6613
rect 5540 6604 5592 6656
rect 7288 6604 7340 6656
rect 8392 6604 8444 6656
rect 12072 6647 12124 6656
rect 12072 6613 12081 6647
rect 12081 6613 12115 6647
rect 12115 6613 12124 6647
rect 12072 6604 12124 6613
rect 12532 6647 12584 6656
rect 12532 6613 12541 6647
rect 12541 6613 12575 6647
rect 12575 6613 12584 6647
rect 12532 6604 12584 6613
rect 16948 6604 17000 6656
rect 19432 6647 19484 6656
rect 19432 6613 19441 6647
rect 19441 6613 19475 6647
rect 19475 6613 19484 6647
rect 19432 6604 19484 6613
rect 22008 6647 22060 6656
rect 22008 6613 22017 6647
rect 22017 6613 22051 6647
rect 22051 6613 22060 6647
rect 22008 6604 22060 6613
rect 23480 6647 23532 6656
rect 23480 6613 23489 6647
rect 23489 6613 23523 6647
rect 23523 6613 23532 6647
rect 23480 6604 23532 6613
rect 23940 6604 23992 6656
rect 24124 6604 24176 6656
rect 24768 6672 24820 6724
rect 27160 6672 27212 6724
rect 27896 6672 27948 6724
rect 24860 6647 24912 6656
rect 24860 6613 24869 6647
rect 24869 6613 24903 6647
rect 24903 6613 24912 6647
rect 24860 6604 24912 6613
rect 26608 6604 26660 6656
rect 29644 6647 29696 6656
rect 29644 6613 29653 6647
rect 29653 6613 29687 6647
rect 29687 6613 29696 6647
rect 29644 6604 29696 6613
rect 32864 6647 32916 6656
rect 32864 6613 32873 6647
rect 32873 6613 32907 6647
rect 32907 6613 32916 6647
rect 32864 6604 32916 6613
rect 35808 6604 35860 6656
rect 35900 6604 35952 6656
rect 36176 6604 36228 6656
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 34966 6502 35018 6554
rect 35030 6502 35082 6554
rect 35094 6502 35146 6554
rect 35158 6502 35210 6554
rect 2228 6443 2280 6452
rect 2228 6409 2237 6443
rect 2237 6409 2271 6443
rect 2271 6409 2280 6443
rect 2228 6400 2280 6409
rect 2504 6400 2556 6452
rect 3240 6400 3292 6452
rect 3976 6400 4028 6452
rect 4712 6443 4764 6452
rect 4712 6409 4721 6443
rect 4721 6409 4755 6443
rect 4755 6409 4764 6443
rect 4712 6400 4764 6409
rect 8208 6400 8260 6452
rect 10048 6443 10100 6452
rect 10048 6409 10057 6443
rect 10057 6409 10091 6443
rect 10091 6409 10100 6443
rect 10048 6400 10100 6409
rect 11796 6443 11848 6452
rect 11796 6409 11805 6443
rect 11805 6409 11839 6443
rect 11839 6409 11848 6443
rect 11796 6400 11848 6409
rect 13452 6443 13504 6452
rect 13452 6409 13461 6443
rect 13461 6409 13495 6443
rect 13495 6409 13504 6443
rect 13452 6400 13504 6409
rect 6552 6375 6604 6384
rect 6552 6341 6561 6375
rect 6561 6341 6595 6375
rect 6595 6341 6604 6375
rect 6552 6332 6604 6341
rect 2228 6196 2280 6248
rect 6368 6264 6420 6316
rect 8300 6264 8352 6316
rect 10600 6307 10652 6316
rect 10600 6273 10609 6307
rect 10609 6273 10643 6307
rect 10643 6273 10652 6307
rect 10600 6264 10652 6273
rect 10692 6307 10744 6316
rect 10692 6273 10701 6307
rect 10701 6273 10735 6307
rect 10735 6273 10744 6307
rect 10692 6264 10744 6273
rect 11704 6264 11756 6316
rect 15108 6400 15160 6452
rect 17500 6443 17552 6452
rect 17500 6409 17509 6443
rect 17509 6409 17543 6443
rect 17543 6409 17552 6443
rect 17500 6400 17552 6409
rect 19984 6443 20036 6452
rect 19984 6409 19993 6443
rect 19993 6409 20027 6443
rect 20027 6409 20036 6443
rect 19984 6400 20036 6409
rect 21916 6443 21968 6452
rect 21916 6409 21925 6443
rect 21925 6409 21959 6443
rect 21959 6409 21968 6443
rect 21916 6400 21968 6409
rect 23572 6400 23624 6452
rect 24676 6443 24728 6452
rect 22008 6332 22060 6384
rect 24032 6332 24084 6384
rect 17316 6264 17368 6316
rect 18052 6307 18104 6316
rect 18052 6273 18061 6307
rect 18061 6273 18095 6307
rect 18095 6273 18104 6307
rect 18052 6264 18104 6273
rect 22376 6264 22428 6316
rect 22560 6307 22612 6316
rect 22560 6273 22569 6307
rect 22569 6273 22603 6307
rect 22603 6273 22612 6307
rect 24676 6409 24685 6443
rect 24685 6409 24719 6443
rect 24719 6409 24728 6443
rect 24676 6400 24728 6409
rect 25320 6400 25372 6452
rect 25504 6443 25556 6452
rect 25504 6409 25513 6443
rect 25513 6409 25547 6443
rect 25547 6409 25556 6443
rect 25504 6400 25556 6409
rect 29000 6443 29052 6452
rect 29000 6409 29009 6443
rect 29009 6409 29043 6443
rect 29043 6409 29052 6443
rect 29000 6400 29052 6409
rect 33048 6400 33100 6452
rect 33508 6400 33560 6452
rect 33600 6443 33652 6452
rect 33600 6409 33609 6443
rect 33609 6409 33643 6443
rect 33643 6409 33652 6443
rect 33600 6400 33652 6409
rect 22560 6264 22612 6273
rect 24216 6307 24268 6316
rect 24216 6273 24225 6307
rect 24225 6273 24259 6307
rect 24259 6273 24268 6307
rect 27896 6332 27948 6384
rect 24216 6264 24268 6273
rect 27988 6307 28040 6316
rect 2596 6239 2648 6248
rect 2596 6205 2630 6239
rect 2630 6205 2648 6239
rect 2596 6196 2648 6205
rect 3976 6196 4028 6248
rect 7472 6196 7524 6248
rect 8392 6239 8444 6248
rect 8392 6205 8401 6239
rect 8401 6205 8435 6239
rect 8435 6205 8444 6239
rect 8392 6196 8444 6205
rect 10784 6196 10836 6248
rect 13176 6196 13228 6248
rect 19156 6196 19208 6248
rect 24676 6196 24728 6248
rect 25412 6196 25464 6248
rect 27988 6273 27997 6307
rect 27997 6273 28031 6307
rect 28031 6273 28040 6307
rect 27988 6264 28040 6273
rect 35624 6400 35676 6452
rect 35532 6332 35584 6384
rect 27620 6196 27672 6248
rect 29000 6196 29052 6248
rect 29276 6239 29328 6248
rect 29276 6205 29285 6239
rect 29285 6205 29319 6239
rect 29319 6205 29328 6239
rect 29276 6196 29328 6205
rect 6644 6128 6696 6180
rect 12072 6128 12124 6180
rect 13912 6128 13964 6180
rect 14372 6128 14424 6180
rect 18420 6128 18472 6180
rect 23480 6128 23532 6180
rect 29736 6128 29788 6180
rect 5080 6103 5132 6112
rect 5080 6069 5089 6103
rect 5089 6069 5123 6103
rect 5123 6069 5132 6103
rect 5080 6060 5132 6069
rect 5448 6103 5500 6112
rect 5448 6069 5457 6103
rect 5457 6069 5491 6103
rect 5491 6069 5500 6103
rect 5448 6060 5500 6069
rect 6828 6103 6880 6112
rect 6828 6069 6837 6103
rect 6837 6069 6871 6103
rect 6871 6069 6880 6103
rect 6828 6060 6880 6069
rect 7288 6103 7340 6112
rect 7288 6069 7297 6103
rect 7297 6069 7331 6103
rect 7331 6069 7340 6103
rect 7288 6060 7340 6069
rect 8576 6103 8628 6112
rect 8576 6069 8585 6103
rect 8585 6069 8619 6103
rect 8619 6069 8628 6103
rect 8576 6060 8628 6069
rect 9772 6060 9824 6112
rect 10968 6060 11020 6112
rect 12164 6060 12216 6112
rect 12440 6103 12492 6112
rect 12440 6069 12449 6103
rect 12449 6069 12483 6103
rect 12483 6069 12492 6103
rect 12440 6060 12492 6069
rect 12532 6060 12584 6112
rect 14004 6060 14056 6112
rect 15476 6060 15528 6112
rect 16212 6060 16264 6112
rect 19340 6060 19392 6112
rect 22008 6103 22060 6112
rect 22008 6069 22017 6103
rect 22017 6069 22051 6103
rect 22051 6069 22060 6103
rect 22008 6060 22060 6069
rect 23664 6103 23716 6112
rect 23664 6069 23673 6103
rect 23673 6069 23707 6103
rect 23707 6069 23716 6103
rect 23664 6060 23716 6069
rect 25964 6103 26016 6112
rect 25964 6069 25973 6103
rect 25973 6069 26007 6103
rect 26007 6069 26016 6103
rect 25964 6060 26016 6069
rect 26240 6060 26292 6112
rect 26976 6103 27028 6112
rect 26976 6069 26985 6103
rect 26985 6069 27019 6103
rect 27019 6069 27028 6103
rect 26976 6060 27028 6069
rect 28080 6060 28132 6112
rect 29460 6103 29512 6112
rect 29460 6069 29469 6103
rect 29469 6069 29503 6103
rect 29503 6069 29512 6103
rect 29460 6060 29512 6069
rect 30288 6103 30340 6112
rect 30288 6069 30297 6103
rect 30297 6069 30331 6103
rect 30331 6069 30340 6103
rect 30288 6060 30340 6069
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 3976 5856 4028 5908
rect 4160 5856 4212 5908
rect 4620 5856 4672 5908
rect 6000 5899 6052 5908
rect 6000 5865 6009 5899
rect 6009 5865 6043 5899
rect 6043 5865 6052 5899
rect 6000 5856 6052 5865
rect 7288 5856 7340 5908
rect 7564 5899 7616 5908
rect 7564 5865 7573 5899
rect 7573 5865 7607 5899
rect 7607 5865 7616 5899
rect 7564 5856 7616 5865
rect 8300 5899 8352 5908
rect 8300 5865 8309 5899
rect 8309 5865 8343 5899
rect 8343 5865 8352 5899
rect 8300 5856 8352 5865
rect 10600 5899 10652 5908
rect 10600 5865 10609 5899
rect 10609 5865 10643 5899
rect 10643 5865 10652 5899
rect 10600 5856 10652 5865
rect 11704 5899 11756 5908
rect 11704 5865 11713 5899
rect 11713 5865 11747 5899
rect 11747 5865 11756 5899
rect 11704 5856 11756 5865
rect 12808 5899 12860 5908
rect 12808 5865 12817 5899
rect 12817 5865 12851 5899
rect 12851 5865 12860 5899
rect 12808 5856 12860 5865
rect 13176 5899 13228 5908
rect 13176 5865 13185 5899
rect 13185 5865 13219 5899
rect 13219 5865 13228 5899
rect 13176 5856 13228 5865
rect 13820 5856 13872 5908
rect 14372 5899 14424 5908
rect 14372 5865 14381 5899
rect 14381 5865 14415 5899
rect 14415 5865 14424 5899
rect 14372 5856 14424 5865
rect 16948 5856 17000 5908
rect 17960 5856 18012 5908
rect 22376 5856 22428 5908
rect 23664 5856 23716 5908
rect 23848 5899 23900 5908
rect 23848 5865 23857 5899
rect 23857 5865 23891 5899
rect 23891 5865 23900 5899
rect 23848 5856 23900 5865
rect 26516 5899 26568 5908
rect 2504 5788 2556 5840
rect 4436 5831 4488 5840
rect 4436 5797 4445 5831
rect 4445 5797 4479 5831
rect 4479 5797 4488 5831
rect 4436 5788 4488 5797
rect 5540 5788 5592 5840
rect 7472 5788 7524 5840
rect 10692 5788 10744 5840
rect 11520 5788 11572 5840
rect 12440 5788 12492 5840
rect 16856 5831 16908 5840
rect 16856 5797 16865 5831
rect 16865 5797 16899 5831
rect 16899 5797 16908 5831
rect 16856 5788 16908 5797
rect 26516 5865 26525 5899
rect 26525 5865 26559 5899
rect 26559 5865 26568 5899
rect 26516 5856 26568 5865
rect 27620 5899 27672 5908
rect 27620 5865 27629 5899
rect 27629 5865 27663 5899
rect 27663 5865 27672 5899
rect 27620 5856 27672 5865
rect 27896 5899 27948 5908
rect 27896 5865 27905 5899
rect 27905 5865 27939 5899
rect 27939 5865 27948 5899
rect 27896 5856 27948 5865
rect 30288 5856 30340 5908
rect 30748 5899 30800 5908
rect 30748 5865 30757 5899
rect 30757 5865 30791 5899
rect 30791 5865 30800 5899
rect 30748 5856 30800 5865
rect 35440 5856 35492 5908
rect 1492 5720 1544 5772
rect 2228 5720 2280 5772
rect 6920 5763 6972 5772
rect 6920 5729 6929 5763
rect 6929 5729 6963 5763
rect 6963 5729 6972 5763
rect 6920 5720 6972 5729
rect 7196 5720 7248 5772
rect 8116 5763 8168 5772
rect 8116 5729 8125 5763
rect 8125 5729 8159 5763
rect 8159 5729 8168 5763
rect 8116 5720 8168 5729
rect 9680 5763 9732 5772
rect 9680 5729 9689 5763
rect 9689 5729 9723 5763
rect 9723 5729 9732 5763
rect 9680 5720 9732 5729
rect 11796 5720 11848 5772
rect 13728 5763 13780 5772
rect 13728 5729 13737 5763
rect 13737 5729 13771 5763
rect 13771 5729 13780 5763
rect 13728 5720 13780 5729
rect 15936 5720 15988 5772
rect 3056 5584 3108 5636
rect 3516 5584 3568 5636
rect 6644 5652 6696 5704
rect 6000 5584 6052 5636
rect 7380 5652 7432 5704
rect 8208 5652 8260 5704
rect 12348 5695 12400 5704
rect 12348 5661 12357 5695
rect 12357 5661 12391 5695
rect 12391 5661 12400 5695
rect 12348 5652 12400 5661
rect 13176 5652 13228 5704
rect 14004 5695 14056 5704
rect 9864 5627 9916 5636
rect 9864 5593 9873 5627
rect 9873 5593 9907 5627
rect 9907 5593 9916 5627
rect 9864 5584 9916 5593
rect 14004 5661 14013 5695
rect 14013 5661 14047 5695
rect 14047 5661 14056 5695
rect 14004 5652 14056 5661
rect 15752 5695 15804 5704
rect 15752 5661 15761 5695
rect 15761 5661 15795 5695
rect 15795 5661 15804 5695
rect 15752 5652 15804 5661
rect 15476 5584 15528 5636
rect 16488 5584 16540 5636
rect 18052 5720 18104 5772
rect 18880 5763 18932 5772
rect 18880 5729 18889 5763
rect 18889 5729 18923 5763
rect 18923 5729 18932 5763
rect 18880 5720 18932 5729
rect 20720 5720 20772 5772
rect 26332 5720 26384 5772
rect 26700 5720 26752 5772
rect 28724 5788 28776 5840
rect 29644 5788 29696 5840
rect 30840 5720 30892 5772
rect 17960 5584 18012 5636
rect 20536 5652 20588 5704
rect 20904 5695 20956 5704
rect 20904 5661 20913 5695
rect 20913 5661 20947 5695
rect 20947 5661 20956 5695
rect 20904 5652 20956 5661
rect 24216 5652 24268 5704
rect 25412 5652 25464 5704
rect 26976 5695 27028 5704
rect 26976 5661 26985 5695
rect 26985 5661 27019 5695
rect 27019 5661 27028 5695
rect 26976 5652 27028 5661
rect 27160 5695 27212 5704
rect 27160 5661 27169 5695
rect 27169 5661 27203 5695
rect 27203 5661 27212 5695
rect 28080 5695 28132 5704
rect 27160 5652 27212 5661
rect 28080 5661 28089 5695
rect 28089 5661 28123 5695
rect 28123 5661 28132 5695
rect 28080 5652 28132 5661
rect 32036 5652 32088 5704
rect 22468 5584 22520 5636
rect 2780 5559 2832 5568
rect 2780 5525 2789 5559
rect 2789 5525 2823 5559
rect 2823 5525 2832 5559
rect 2780 5516 2832 5525
rect 3332 5559 3384 5568
rect 3332 5525 3341 5559
rect 3341 5525 3375 5559
rect 3375 5525 3384 5559
rect 3332 5516 3384 5525
rect 5080 5559 5132 5568
rect 5080 5525 5089 5559
rect 5089 5525 5123 5559
rect 5123 5525 5132 5559
rect 5080 5516 5132 5525
rect 7472 5516 7524 5568
rect 11612 5516 11664 5568
rect 13360 5559 13412 5568
rect 13360 5525 13369 5559
rect 13369 5525 13403 5559
rect 13403 5525 13412 5559
rect 13360 5516 13412 5525
rect 15292 5559 15344 5568
rect 15292 5525 15301 5559
rect 15301 5525 15335 5559
rect 15335 5525 15344 5559
rect 15292 5516 15344 5525
rect 17868 5516 17920 5568
rect 19892 5559 19944 5568
rect 19892 5525 19901 5559
rect 19901 5525 19935 5559
rect 19935 5525 19944 5559
rect 19892 5516 19944 5525
rect 22836 5559 22888 5568
rect 22836 5525 22845 5559
rect 22845 5525 22879 5559
rect 22879 5525 22888 5559
rect 22836 5516 22888 5525
rect 24124 5516 24176 5568
rect 24860 5559 24912 5568
rect 24860 5525 24869 5559
rect 24869 5525 24903 5559
rect 24903 5525 24912 5559
rect 24860 5516 24912 5525
rect 26240 5516 26292 5568
rect 29000 5516 29052 5568
rect 30104 5559 30156 5568
rect 30104 5525 30113 5559
rect 30113 5525 30147 5559
rect 30147 5525 30156 5559
rect 30104 5516 30156 5525
rect 31208 5559 31260 5568
rect 31208 5525 31217 5559
rect 31217 5525 31251 5559
rect 31251 5525 31260 5559
rect 31208 5516 31260 5525
rect 31760 5559 31812 5568
rect 31760 5525 31769 5559
rect 31769 5525 31803 5559
rect 31803 5525 31812 5559
rect 31760 5516 31812 5525
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 34966 5414 35018 5466
rect 35030 5414 35082 5466
rect 35094 5414 35146 5466
rect 35158 5414 35210 5466
rect 1492 5312 1544 5364
rect 3240 5355 3292 5364
rect 3240 5321 3249 5355
rect 3249 5321 3283 5355
rect 3283 5321 3292 5355
rect 3240 5312 3292 5321
rect 4620 5355 4672 5364
rect 4620 5321 4629 5355
rect 4629 5321 4663 5355
rect 4663 5321 4672 5355
rect 4620 5312 4672 5321
rect 5540 5312 5592 5364
rect 6736 5312 6788 5364
rect 9680 5312 9732 5364
rect 11796 5355 11848 5364
rect 11796 5321 11805 5355
rect 11805 5321 11839 5355
rect 11839 5321 11848 5355
rect 11796 5312 11848 5321
rect 13728 5312 13780 5364
rect 13912 5312 13964 5364
rect 14556 5312 14608 5364
rect 15752 5312 15804 5364
rect 15936 5355 15988 5364
rect 15936 5321 15945 5355
rect 15945 5321 15979 5355
rect 15979 5321 15988 5355
rect 15936 5312 15988 5321
rect 17776 5312 17828 5364
rect 18144 5312 18196 5364
rect 19156 5355 19208 5364
rect 19156 5321 19165 5355
rect 19165 5321 19199 5355
rect 19199 5321 19208 5355
rect 19156 5312 19208 5321
rect 20720 5355 20772 5364
rect 20720 5321 20729 5355
rect 20729 5321 20763 5355
rect 20763 5321 20772 5355
rect 20720 5312 20772 5321
rect 23848 5312 23900 5364
rect 25044 5355 25096 5364
rect 25044 5321 25053 5355
rect 25053 5321 25087 5355
rect 25087 5321 25096 5355
rect 25044 5312 25096 5321
rect 26240 5312 26292 5364
rect 28724 5355 28776 5364
rect 6644 5287 6696 5296
rect 6644 5253 6653 5287
rect 6653 5253 6687 5287
rect 6687 5253 6696 5287
rect 6644 5244 6696 5253
rect 15108 5244 15160 5296
rect 3056 5176 3108 5228
rect 5448 5219 5500 5228
rect 2596 5108 2648 5160
rect 2780 5108 2832 5160
rect 5448 5185 5457 5219
rect 5457 5185 5491 5219
rect 5491 5185 5500 5219
rect 5448 5176 5500 5185
rect 7288 5219 7340 5228
rect 7288 5185 7297 5219
rect 7297 5185 7331 5219
rect 7331 5185 7340 5219
rect 7288 5176 7340 5185
rect 7472 5219 7524 5228
rect 7472 5185 7481 5219
rect 7481 5185 7515 5219
rect 7515 5185 7524 5219
rect 7472 5176 7524 5185
rect 13360 5176 13412 5228
rect 13820 5176 13872 5228
rect 16856 5176 16908 5228
rect 18972 5176 19024 5228
rect 22008 5287 22060 5296
rect 22008 5253 22017 5287
rect 22017 5253 22051 5287
rect 22051 5253 22060 5287
rect 22008 5244 22060 5253
rect 24768 5244 24820 5296
rect 26976 5244 27028 5296
rect 28724 5321 28733 5355
rect 28733 5321 28767 5355
rect 28767 5321 28776 5355
rect 28724 5312 28776 5321
rect 31208 5312 31260 5364
rect 22560 5219 22612 5228
rect 3332 5040 3384 5092
rect 7564 5108 7616 5160
rect 4344 5083 4396 5092
rect 4344 5049 4353 5083
rect 4353 5049 4387 5083
rect 4387 5049 4396 5083
rect 4344 5040 4396 5049
rect 10600 5151 10652 5160
rect 10600 5117 10609 5151
rect 10609 5117 10643 5151
rect 10643 5117 10652 5151
rect 10600 5108 10652 5117
rect 12900 5108 12952 5160
rect 13452 5108 13504 5160
rect 22560 5185 22569 5219
rect 22569 5185 22603 5219
rect 22603 5185 22612 5219
rect 22560 5176 22612 5185
rect 24124 5219 24176 5228
rect 24124 5185 24133 5219
rect 24133 5185 24167 5219
rect 24167 5185 24176 5219
rect 24124 5176 24176 5185
rect 24216 5219 24268 5228
rect 24216 5185 24225 5219
rect 24225 5185 24259 5219
rect 24259 5185 24268 5219
rect 24216 5176 24268 5185
rect 25596 5176 25648 5228
rect 27896 5219 27948 5228
rect 27896 5185 27905 5219
rect 27905 5185 27939 5219
rect 27939 5185 27948 5219
rect 27896 5176 27948 5185
rect 31760 5176 31812 5228
rect 32128 5219 32180 5228
rect 32128 5185 32137 5219
rect 32137 5185 32171 5219
rect 32171 5185 32180 5219
rect 32128 5176 32180 5185
rect 32312 5219 32364 5228
rect 32312 5185 32321 5219
rect 32321 5185 32355 5219
rect 32355 5185 32364 5219
rect 32312 5176 32364 5185
rect 10876 5040 10928 5092
rect 16948 5040 17000 5092
rect 20904 5108 20956 5160
rect 22836 5108 22888 5160
rect 23388 5108 23440 5160
rect 25044 5108 25096 5160
rect 26884 5151 26936 5160
rect 26884 5117 26893 5151
rect 26893 5117 26927 5151
rect 26927 5117 26936 5151
rect 26884 5108 26936 5117
rect 29000 5108 29052 5160
rect 29276 5151 29328 5160
rect 29276 5117 29285 5151
rect 29285 5117 29319 5151
rect 29319 5117 29328 5151
rect 29276 5108 29328 5117
rect 19892 5040 19944 5092
rect 20628 5040 20680 5092
rect 25780 5040 25832 5092
rect 32036 5151 32088 5160
rect 32036 5117 32045 5151
rect 32045 5117 32079 5151
rect 32079 5117 32088 5151
rect 32036 5108 32088 5117
rect 2412 4972 2464 5024
rect 2596 5015 2648 5024
rect 2596 4981 2605 5015
rect 2605 4981 2639 5015
rect 2639 4981 2648 5015
rect 2596 4972 2648 4981
rect 2688 4972 2740 5024
rect 4620 4972 4672 5024
rect 7932 4972 7984 5024
rect 8116 5015 8168 5024
rect 8116 4981 8125 5015
rect 8125 4981 8159 5015
rect 8159 4981 8168 5015
rect 8116 4972 8168 4981
rect 8392 4972 8444 5024
rect 9036 5015 9088 5024
rect 9036 4981 9045 5015
rect 9045 4981 9079 5015
rect 9079 4981 9088 5015
rect 9036 4972 9088 4981
rect 9312 5015 9364 5024
rect 9312 4981 9321 5015
rect 9321 4981 9355 5015
rect 9355 4981 9364 5015
rect 9312 4972 9364 4981
rect 9496 4972 9548 5024
rect 10784 5015 10836 5024
rect 10784 4981 10793 5015
rect 10793 4981 10827 5015
rect 10827 4981 10836 5015
rect 10784 4972 10836 4981
rect 12716 4972 12768 5024
rect 14280 4972 14332 5024
rect 16396 5015 16448 5024
rect 16396 4981 16405 5015
rect 16405 4981 16439 5015
rect 16439 4981 16448 5015
rect 16396 4972 16448 4981
rect 16580 4972 16632 5024
rect 17776 5015 17828 5024
rect 17776 4981 17785 5015
rect 17785 4981 17819 5015
rect 17819 4981 17828 5015
rect 17776 4972 17828 4981
rect 18880 5015 18932 5024
rect 18880 4981 18889 5015
rect 18889 4981 18923 5015
rect 18923 4981 18932 5015
rect 18880 4972 18932 4981
rect 23112 5015 23164 5024
rect 23112 4981 23121 5015
rect 23121 4981 23155 5015
rect 23155 4981 23164 5015
rect 23112 4972 23164 4981
rect 24032 5015 24084 5024
rect 24032 4981 24041 5015
rect 24041 4981 24075 5015
rect 24075 4981 24084 5015
rect 24032 4972 24084 4981
rect 28080 4972 28132 5024
rect 29276 4972 29328 5024
rect 29460 5015 29512 5024
rect 29460 4981 29469 5015
rect 29469 4981 29503 5015
rect 29503 4981 29512 5015
rect 29460 4972 29512 4981
rect 30196 5015 30248 5024
rect 30196 4981 30205 5015
rect 30205 4981 30239 5015
rect 30239 4981 30248 5015
rect 30196 4972 30248 4981
rect 30564 5015 30616 5024
rect 30564 4981 30573 5015
rect 30573 4981 30607 5015
rect 30607 4981 30616 5015
rect 30564 4972 30616 4981
rect 30840 4972 30892 5024
rect 31668 4972 31720 5024
rect 32772 5015 32824 5024
rect 32772 4981 32781 5015
rect 32781 4981 32815 5015
rect 32815 4981 32824 5015
rect 32772 4972 32824 4981
rect 34520 4972 34572 5024
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 3332 4811 3384 4820
rect 3332 4777 3341 4811
rect 3341 4777 3375 4811
rect 3375 4777 3384 4811
rect 3332 4768 3384 4777
rect 5816 4768 5868 4820
rect 6736 4768 6788 4820
rect 7288 4768 7340 4820
rect 8024 4811 8076 4820
rect 8024 4777 8033 4811
rect 8033 4777 8067 4811
rect 8067 4777 8076 4811
rect 8024 4768 8076 4777
rect 9496 4811 9548 4820
rect 9496 4777 9505 4811
rect 9505 4777 9539 4811
rect 9539 4777 9548 4811
rect 9496 4768 9548 4777
rect 10232 4768 10284 4820
rect 10784 4768 10836 4820
rect 11520 4811 11572 4820
rect 11520 4777 11529 4811
rect 11529 4777 11563 4811
rect 11563 4777 11572 4811
rect 11520 4768 11572 4777
rect 14004 4811 14056 4820
rect 14004 4777 14013 4811
rect 14013 4777 14047 4811
rect 14047 4777 14056 4811
rect 14004 4768 14056 4777
rect 15292 4768 15344 4820
rect 16948 4768 17000 4820
rect 17224 4811 17276 4820
rect 17224 4777 17233 4811
rect 17233 4777 17267 4811
rect 17267 4777 17276 4811
rect 17224 4768 17276 4777
rect 19340 4768 19392 4820
rect 4804 4700 4856 4752
rect 7932 4743 7984 4752
rect 7932 4709 7941 4743
rect 7941 4709 7975 4743
rect 7975 4709 7984 4743
rect 7932 4700 7984 4709
rect 11704 4700 11756 4752
rect 12072 4700 12124 4752
rect 16580 4700 16632 4752
rect 17776 4700 17828 4752
rect 19432 4700 19484 4752
rect 19616 4700 19668 4752
rect 20444 4768 20496 4820
rect 21824 4811 21876 4820
rect 21824 4777 21833 4811
rect 21833 4777 21867 4811
rect 21867 4777 21876 4811
rect 21824 4768 21876 4777
rect 24216 4768 24268 4820
rect 27160 4811 27212 4820
rect 27160 4777 27169 4811
rect 27169 4777 27203 4811
rect 27203 4777 27212 4811
rect 27160 4768 27212 4777
rect 30288 4768 30340 4820
rect 32128 4811 32180 4820
rect 32128 4777 32137 4811
rect 32137 4777 32171 4811
rect 32171 4777 32180 4811
rect 32128 4768 32180 4777
rect 32772 4768 32824 4820
rect 34244 4768 34296 4820
rect 34612 4768 34664 4820
rect 23296 4700 23348 4752
rect 23664 4743 23716 4752
rect 23664 4709 23698 4743
rect 23698 4709 23716 4743
rect 23664 4700 23716 4709
rect 32036 4700 32088 4752
rect 1492 4632 1544 4684
rect 5172 4632 5224 4684
rect 6184 4632 6236 4684
rect 6828 4675 6880 4684
rect 6828 4641 6837 4675
rect 6837 4641 6871 4675
rect 6871 4641 6880 4675
rect 6828 4632 6880 4641
rect 7012 4632 7064 4684
rect 2780 4471 2832 4480
rect 2780 4437 2789 4471
rect 2789 4437 2823 4471
rect 2823 4437 2832 4471
rect 2780 4428 2832 4437
rect 3056 4428 3108 4480
rect 8484 4675 8536 4684
rect 8484 4641 8493 4675
rect 8493 4641 8527 4675
rect 8527 4641 8536 4675
rect 8484 4632 8536 4641
rect 10600 4632 10652 4684
rect 11980 4675 12032 4684
rect 11980 4641 11989 4675
rect 11989 4641 12023 4675
rect 12023 4641 12032 4675
rect 11980 4632 12032 4641
rect 15660 4675 15712 4684
rect 15660 4641 15669 4675
rect 15669 4641 15703 4675
rect 15703 4641 15712 4675
rect 15660 4632 15712 4641
rect 16856 4632 16908 4684
rect 17592 4675 17644 4684
rect 17592 4641 17615 4675
rect 17615 4641 17644 4675
rect 22192 4675 22244 4684
rect 17592 4632 17644 4641
rect 22192 4641 22201 4675
rect 22201 4641 22235 4675
rect 22235 4641 22244 4675
rect 22192 4632 22244 4641
rect 27804 4675 27856 4684
rect 27804 4641 27813 4675
rect 27813 4641 27847 4675
rect 27847 4641 27856 4675
rect 27804 4632 27856 4641
rect 28356 4632 28408 4684
rect 29368 4632 29420 4684
rect 32496 4675 32548 4684
rect 32496 4641 32505 4675
rect 32505 4641 32539 4675
rect 32539 4641 32548 4675
rect 32496 4632 32548 4641
rect 9496 4564 9548 4616
rect 9956 4564 10008 4616
rect 14096 4564 14148 4616
rect 15844 4607 15896 4616
rect 15844 4573 15853 4607
rect 15853 4573 15887 4607
rect 15887 4573 15896 4607
rect 15844 4564 15896 4573
rect 17316 4607 17368 4616
rect 17316 4573 17325 4607
rect 17325 4573 17359 4607
rect 17359 4573 17368 4607
rect 17316 4564 17368 4573
rect 22284 4607 22336 4616
rect 22284 4573 22293 4607
rect 22293 4573 22327 4607
rect 22327 4573 22336 4607
rect 22284 4564 22336 4573
rect 6000 4539 6052 4548
rect 6000 4505 6009 4539
rect 6009 4505 6043 4539
rect 6043 4505 6052 4539
rect 6000 4496 6052 4505
rect 8484 4496 8536 4548
rect 15200 4496 15252 4548
rect 22560 4564 22612 4616
rect 23204 4564 23256 4616
rect 27988 4607 28040 4616
rect 27988 4573 27997 4607
rect 27997 4573 28031 4607
rect 28031 4573 28040 4607
rect 29276 4607 29328 4616
rect 27988 4564 28040 4573
rect 29276 4573 29285 4607
rect 29285 4573 29319 4607
rect 29319 4573 29328 4607
rect 29276 4564 29328 4573
rect 5540 4428 5592 4480
rect 5632 4471 5684 4480
rect 5632 4437 5641 4471
rect 5641 4437 5675 4471
rect 5675 4437 5684 4471
rect 7104 4471 7156 4480
rect 5632 4428 5684 4437
rect 7104 4437 7113 4471
rect 7113 4437 7147 4471
rect 7147 4437 7156 4471
rect 7104 4428 7156 4437
rect 7564 4428 7616 4480
rect 9128 4471 9180 4480
rect 9128 4437 9137 4471
rect 9137 4437 9171 4471
rect 9171 4437 9180 4471
rect 9128 4428 9180 4437
rect 10324 4428 10376 4480
rect 12348 4428 12400 4480
rect 13636 4428 13688 4480
rect 13820 4428 13872 4480
rect 15476 4428 15528 4480
rect 19156 4428 19208 4480
rect 21272 4471 21324 4480
rect 21272 4437 21281 4471
rect 21281 4437 21315 4471
rect 21315 4437 21324 4471
rect 23112 4496 23164 4548
rect 21272 4428 21324 4437
rect 23204 4471 23256 4480
rect 23204 4437 23213 4471
rect 23213 4437 23247 4471
rect 23247 4437 23256 4471
rect 23204 4428 23256 4437
rect 25596 4496 25648 4548
rect 27620 4496 27672 4548
rect 24768 4471 24820 4480
rect 24768 4437 24777 4471
rect 24777 4437 24811 4471
rect 24811 4437 24820 4471
rect 24768 4428 24820 4437
rect 26700 4471 26752 4480
rect 26700 4437 26709 4471
rect 26709 4437 26743 4471
rect 26743 4437 26752 4471
rect 26700 4428 26752 4437
rect 27528 4428 27580 4480
rect 28448 4471 28500 4480
rect 28448 4437 28457 4471
rect 28457 4437 28491 4471
rect 28491 4437 28500 4471
rect 28448 4428 28500 4437
rect 30380 4428 30432 4480
rect 33048 4632 33100 4684
rect 34244 4675 34296 4684
rect 34244 4641 34278 4675
rect 34278 4641 34296 4675
rect 34244 4632 34296 4641
rect 33968 4607 34020 4616
rect 33968 4573 33977 4607
rect 33977 4573 34011 4607
rect 34011 4573 34020 4607
rect 33968 4564 34020 4573
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 34966 4326 35018 4378
rect 35030 4326 35082 4378
rect 35094 4326 35146 4378
rect 35158 4326 35210 4378
rect 3332 4224 3384 4276
rect 6184 4267 6236 4276
rect 6184 4233 6193 4267
rect 6193 4233 6227 4267
rect 6227 4233 6236 4267
rect 6184 4224 6236 4233
rect 11980 4267 12032 4276
rect 11980 4233 11989 4267
rect 11989 4233 12023 4267
rect 12023 4233 12032 4267
rect 11980 4224 12032 4233
rect 15752 4224 15804 4276
rect 2872 4088 2924 4140
rect 4620 4156 4672 4208
rect 6736 4156 6788 4208
rect 7564 4156 7616 4208
rect 5540 4131 5592 4140
rect 5540 4097 5549 4131
rect 5549 4097 5583 4131
rect 5583 4097 5592 4131
rect 5540 4088 5592 4097
rect 1492 4020 1544 4072
rect 2596 4020 2648 4072
rect 3792 3927 3844 3936
rect 3792 3893 3801 3927
rect 3801 3893 3835 3927
rect 3835 3893 3844 3927
rect 3792 3884 3844 3893
rect 4068 3927 4120 3936
rect 4068 3893 4077 3927
rect 4077 3893 4111 3927
rect 4111 3893 4120 3927
rect 4068 3884 4120 3893
rect 4712 4020 4764 4072
rect 5080 4020 5132 4072
rect 7104 4020 7156 4072
rect 9588 4020 9640 4072
rect 12440 4063 12492 4072
rect 4620 3884 4672 3936
rect 4804 3927 4856 3936
rect 4804 3893 4813 3927
rect 4813 3893 4847 3927
rect 4847 3893 4856 3927
rect 4804 3884 4856 3893
rect 5356 3952 5408 4004
rect 6920 3952 6972 4004
rect 8300 3952 8352 4004
rect 12440 4029 12449 4063
rect 12449 4029 12483 4063
rect 12483 4029 12492 4063
rect 12440 4020 12492 4029
rect 14096 4063 14148 4072
rect 14096 4029 14130 4063
rect 14130 4029 14148 4063
rect 11980 3952 12032 4004
rect 14096 4020 14148 4029
rect 17316 4224 17368 4276
rect 17592 4224 17644 4276
rect 18604 4267 18656 4276
rect 18604 4233 18613 4267
rect 18613 4233 18647 4267
rect 18647 4233 18656 4267
rect 18604 4224 18656 4233
rect 19984 4224 20036 4276
rect 20168 4224 20220 4276
rect 22192 4224 22244 4276
rect 23204 4224 23256 4276
rect 26700 4224 26752 4276
rect 27804 4224 27856 4276
rect 17224 4156 17276 4208
rect 17408 4088 17460 4140
rect 19432 4088 19484 4140
rect 20628 4088 20680 4140
rect 22284 4156 22336 4208
rect 25596 4199 25648 4208
rect 25596 4165 25605 4199
rect 25605 4165 25639 4199
rect 25639 4165 25648 4199
rect 25596 4156 25648 4165
rect 23572 4088 23624 4140
rect 26976 4156 27028 4208
rect 16948 3952 17000 4004
rect 19616 4020 19668 4072
rect 20168 4020 20220 4072
rect 23204 4020 23256 4072
rect 24768 4020 24820 4072
rect 26608 4020 26660 4072
rect 28448 4156 28500 4208
rect 29276 4088 29328 4140
rect 29644 4088 29696 4140
rect 30288 4088 30340 4140
rect 31208 4088 31260 4140
rect 33048 4088 33100 4140
rect 28264 4020 28316 4072
rect 30380 4020 30432 4072
rect 31116 4020 31168 4072
rect 31668 4020 31720 4072
rect 32496 4020 32548 4072
rect 5540 3884 5592 3936
rect 6828 3927 6880 3936
rect 6828 3893 6837 3927
rect 6837 3893 6871 3927
rect 6871 3893 6880 3927
rect 6828 3884 6880 3893
rect 9956 3927 10008 3936
rect 9956 3893 9965 3927
rect 9965 3893 9999 3927
rect 9999 3893 10008 3927
rect 9956 3884 10008 3893
rect 10600 3927 10652 3936
rect 10600 3893 10609 3927
rect 10609 3893 10643 3927
rect 10643 3893 10652 3927
rect 10600 3884 10652 3893
rect 11244 3927 11296 3936
rect 11244 3893 11253 3927
rect 11253 3893 11287 3927
rect 11287 3893 11296 3927
rect 11244 3884 11296 3893
rect 11704 3927 11756 3936
rect 11704 3893 11713 3927
rect 11713 3893 11747 3927
rect 11747 3893 11756 3927
rect 11704 3884 11756 3893
rect 12716 3884 12768 3936
rect 14372 3884 14424 3936
rect 14924 3884 14976 3936
rect 15660 3884 15712 3936
rect 16488 3884 16540 3936
rect 19064 3927 19116 3936
rect 19064 3893 19073 3927
rect 19073 3893 19107 3927
rect 19107 3893 19116 3927
rect 19064 3884 19116 3893
rect 19432 3927 19484 3936
rect 19432 3893 19441 3927
rect 19441 3893 19475 3927
rect 19475 3893 19484 3927
rect 19984 3927 20036 3936
rect 19432 3884 19484 3893
rect 19984 3893 19995 3927
rect 19995 3893 20029 3927
rect 20029 3893 20036 3927
rect 21364 3927 21416 3936
rect 19984 3884 20036 3893
rect 21364 3893 21373 3927
rect 21373 3893 21407 3927
rect 21407 3893 21416 3927
rect 21364 3884 21416 3893
rect 22652 3927 22704 3936
rect 22652 3893 22661 3927
rect 22661 3893 22695 3927
rect 22695 3893 22704 3927
rect 22652 3884 22704 3893
rect 23112 3927 23164 3936
rect 23112 3893 23121 3927
rect 23121 3893 23155 3927
rect 23155 3893 23164 3927
rect 23112 3884 23164 3893
rect 25044 3927 25096 3936
rect 25044 3893 25053 3927
rect 25053 3893 25087 3927
rect 25087 3893 25096 3927
rect 25044 3884 25096 3893
rect 26700 3884 26752 3936
rect 28356 3927 28408 3936
rect 28356 3893 28365 3927
rect 28365 3893 28399 3927
rect 28399 3893 28408 3927
rect 28356 3884 28408 3893
rect 29736 3884 29788 3936
rect 29920 3927 29972 3936
rect 29920 3893 29929 3927
rect 29929 3893 29963 3927
rect 29963 3893 29972 3927
rect 30472 3927 30524 3936
rect 29920 3884 29972 3893
rect 30472 3893 30481 3927
rect 30481 3893 30515 3927
rect 30515 3893 30524 3927
rect 30472 3884 30524 3893
rect 31024 3884 31076 3936
rect 32036 3884 32088 3936
rect 33600 3884 33652 3936
rect 33968 3927 34020 3936
rect 33968 3893 33977 3927
rect 33977 3893 34011 3927
rect 34011 3893 34020 3927
rect 33968 3884 34020 3893
rect 34244 3884 34296 3936
rect 34612 3884 34664 3936
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 2412 3680 2464 3732
rect 8484 3680 8536 3732
rect 9496 3723 9548 3732
rect 9496 3689 9505 3723
rect 9505 3689 9539 3723
rect 9539 3689 9548 3723
rect 9496 3680 9548 3689
rect 9680 3723 9732 3732
rect 9680 3689 9689 3723
rect 9689 3689 9723 3723
rect 9723 3689 9732 3723
rect 9680 3680 9732 3689
rect 10232 3723 10284 3732
rect 10232 3689 10241 3723
rect 10241 3689 10275 3723
rect 10275 3689 10284 3723
rect 10232 3680 10284 3689
rect 12072 3723 12124 3732
rect 12072 3689 12081 3723
rect 12081 3689 12115 3723
rect 12115 3689 12124 3723
rect 12072 3680 12124 3689
rect 13176 3723 13228 3732
rect 13176 3689 13185 3723
rect 13185 3689 13219 3723
rect 13219 3689 13228 3723
rect 13176 3680 13228 3689
rect 13728 3680 13780 3732
rect 14556 3723 14608 3732
rect 14556 3689 14565 3723
rect 14565 3689 14599 3723
rect 14599 3689 14608 3723
rect 14556 3680 14608 3689
rect 14924 3723 14976 3732
rect 14924 3689 14933 3723
rect 14933 3689 14967 3723
rect 14967 3689 14976 3723
rect 14924 3680 14976 3689
rect 15844 3680 15896 3732
rect 16212 3723 16264 3732
rect 16212 3689 16221 3723
rect 16221 3689 16255 3723
rect 16255 3689 16264 3723
rect 16212 3680 16264 3689
rect 16396 3680 16448 3732
rect 17776 3680 17828 3732
rect 20168 3680 20220 3732
rect 20628 3723 20680 3732
rect 20628 3689 20637 3723
rect 20637 3689 20671 3723
rect 20671 3689 20680 3723
rect 20628 3680 20680 3689
rect 23296 3680 23348 3732
rect 26608 3680 26660 3732
rect 28264 3680 28316 3732
rect 28632 3680 28684 3732
rect 28908 3680 28960 3732
rect 29368 3723 29420 3732
rect 29368 3689 29377 3723
rect 29377 3689 29411 3723
rect 29411 3689 29420 3723
rect 29368 3680 29420 3689
rect 30564 3680 30616 3732
rect 31576 3680 31628 3732
rect 32036 3680 32088 3732
rect 32312 3723 32364 3732
rect 32312 3689 32321 3723
rect 32321 3689 32355 3723
rect 32355 3689 32364 3723
rect 32312 3680 32364 3689
rect 32496 3680 32548 3732
rect 34612 3723 34664 3732
rect 34612 3689 34621 3723
rect 34621 3689 34655 3723
rect 34655 3689 34664 3723
rect 34612 3680 34664 3689
rect 2780 3612 2832 3664
rect 8208 3612 8260 3664
rect 9956 3612 10008 3664
rect 1492 3587 1544 3596
rect 1492 3553 1501 3587
rect 1501 3553 1535 3587
rect 1535 3553 1544 3587
rect 1492 3544 1544 3553
rect 4436 3587 4488 3596
rect 4436 3553 4445 3587
rect 4445 3553 4479 3587
rect 4479 3553 4488 3587
rect 4436 3544 4488 3553
rect 5632 3544 5684 3596
rect 6828 3544 6880 3596
rect 8944 3544 8996 3596
rect 9496 3544 9548 3596
rect 11980 3612 12032 3664
rect 12716 3612 12768 3664
rect 14464 3612 14516 3664
rect 15108 3612 15160 3664
rect 10784 3544 10836 3596
rect 4712 3519 4764 3528
rect 4712 3485 4721 3519
rect 4721 3485 4755 3519
rect 4755 3485 4764 3519
rect 4712 3476 4764 3485
rect 6000 3519 6052 3528
rect 6000 3485 6009 3519
rect 6009 3485 6043 3519
rect 6043 3485 6052 3519
rect 6000 3476 6052 3485
rect 3976 3408 4028 3460
rect 2964 3340 3016 3392
rect 5172 3383 5224 3392
rect 5172 3349 5181 3383
rect 5181 3349 5215 3383
rect 5215 3349 5224 3383
rect 5172 3340 5224 3349
rect 5448 3340 5500 3392
rect 7196 3340 7248 3392
rect 8668 3383 8720 3392
rect 8668 3349 8677 3383
rect 8677 3349 8711 3383
rect 8711 3349 8720 3383
rect 8668 3340 8720 3349
rect 10968 3340 11020 3392
rect 14372 3476 14424 3528
rect 17316 3612 17368 3664
rect 23480 3612 23532 3664
rect 25044 3612 25096 3664
rect 30288 3612 30340 3664
rect 30472 3612 30524 3664
rect 33140 3655 33192 3664
rect 33140 3621 33149 3655
rect 33149 3621 33183 3655
rect 33183 3621 33192 3655
rect 33140 3612 33192 3621
rect 17408 3587 17460 3596
rect 17408 3553 17417 3587
rect 17417 3553 17451 3587
rect 17451 3553 17460 3587
rect 17408 3544 17460 3553
rect 17684 3544 17736 3596
rect 21364 3587 21416 3596
rect 21364 3553 21373 3587
rect 21373 3553 21407 3587
rect 21407 3553 21416 3587
rect 21364 3544 21416 3553
rect 23204 3544 23256 3596
rect 26516 3587 26568 3596
rect 26516 3553 26525 3587
rect 26525 3553 26559 3587
rect 26559 3553 26568 3587
rect 26516 3544 26568 3553
rect 26884 3544 26936 3596
rect 17868 3519 17920 3528
rect 17868 3485 17877 3519
rect 17877 3485 17911 3519
rect 17911 3485 17920 3519
rect 17868 3476 17920 3485
rect 18144 3519 18196 3528
rect 18144 3485 18153 3519
rect 18153 3485 18187 3519
rect 18187 3485 18196 3519
rect 18144 3476 18196 3485
rect 21456 3519 21508 3528
rect 21456 3485 21465 3519
rect 21465 3485 21499 3519
rect 21499 3485 21508 3519
rect 21456 3476 21508 3485
rect 22560 3476 22612 3528
rect 27528 3476 27580 3528
rect 28448 3519 28500 3528
rect 28448 3485 28457 3519
rect 28457 3485 28491 3519
rect 28491 3485 28500 3519
rect 28448 3476 28500 3485
rect 29644 3544 29696 3596
rect 31944 3544 31996 3596
rect 34060 3544 34112 3596
rect 35440 3544 35492 3596
rect 28724 3476 28776 3528
rect 29368 3476 29420 3528
rect 19984 3408 20036 3460
rect 22468 3408 22520 3460
rect 26332 3408 26384 3460
rect 27436 3408 27488 3460
rect 15844 3383 15896 3392
rect 15844 3349 15853 3383
rect 15853 3349 15887 3383
rect 15887 3349 15896 3383
rect 15844 3340 15896 3349
rect 20904 3383 20956 3392
rect 20904 3349 20913 3383
rect 20913 3349 20947 3383
rect 20947 3349 20956 3383
rect 20904 3340 20956 3349
rect 22652 3383 22704 3392
rect 22652 3349 22661 3383
rect 22661 3349 22695 3383
rect 22695 3349 22704 3383
rect 22652 3340 22704 3349
rect 23572 3340 23624 3392
rect 30196 3340 30248 3392
rect 30932 3383 30984 3392
rect 30932 3349 30941 3383
rect 30941 3349 30975 3383
rect 30975 3349 30984 3383
rect 30932 3340 30984 3349
rect 33600 3340 33652 3392
rect 35348 3340 35400 3392
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 34966 3238 35018 3290
rect 35030 3238 35082 3290
rect 35094 3238 35146 3290
rect 35158 3238 35210 3290
rect 1492 3136 1544 3188
rect 5632 3179 5684 3188
rect 4160 3068 4212 3120
rect 5632 3145 5641 3179
rect 5641 3145 5675 3179
rect 5675 3145 5684 3179
rect 5632 3136 5684 3145
rect 8300 3179 8352 3188
rect 8300 3145 8309 3179
rect 8309 3145 8343 3179
rect 8343 3145 8352 3179
rect 8300 3136 8352 3145
rect 10784 3179 10836 3188
rect 10784 3145 10793 3179
rect 10793 3145 10827 3179
rect 10827 3145 10836 3179
rect 10784 3136 10836 3145
rect 11980 3136 12032 3188
rect 12624 3179 12676 3188
rect 12624 3145 12633 3179
rect 12633 3145 12667 3179
rect 12667 3145 12676 3179
rect 12624 3136 12676 3145
rect 13728 3136 13780 3188
rect 15752 3179 15804 3188
rect 15752 3145 15761 3179
rect 15761 3145 15795 3179
rect 15795 3145 15804 3179
rect 15752 3136 15804 3145
rect 16212 3136 16264 3188
rect 16672 3179 16724 3188
rect 16672 3145 16681 3179
rect 16681 3145 16715 3179
rect 16715 3145 16724 3179
rect 16672 3136 16724 3145
rect 17040 3179 17092 3188
rect 17040 3145 17049 3179
rect 17049 3145 17083 3179
rect 17083 3145 17092 3179
rect 17040 3136 17092 3145
rect 17684 3136 17736 3188
rect 6000 3068 6052 3120
rect 1768 3043 1820 3052
rect 1768 3009 1777 3043
rect 1777 3009 1811 3043
rect 1811 3009 1820 3043
rect 1768 3000 1820 3009
rect 3792 3000 3844 3052
rect 4160 2975 4212 2984
rect 4160 2941 4169 2975
rect 4169 2941 4203 2975
rect 4203 2941 4212 2975
rect 4160 2932 4212 2941
rect 5448 2932 5500 2984
rect 12532 3068 12584 3120
rect 18144 3136 18196 3188
rect 18420 3179 18472 3188
rect 18420 3145 18429 3179
rect 18429 3145 18463 3179
rect 18463 3145 18472 3179
rect 18420 3136 18472 3145
rect 18972 3136 19024 3188
rect 14280 3000 14332 3052
rect 14464 3000 14516 3052
rect 14556 3000 14608 3052
rect 18880 3043 18932 3052
rect 7196 2975 7248 2984
rect 7196 2941 7230 2975
rect 7230 2941 7248 2975
rect 2964 2864 3016 2916
rect 1676 2796 1728 2848
rect 2688 2796 2740 2848
rect 4804 2864 4856 2916
rect 7196 2932 7248 2941
rect 8944 2975 8996 2984
rect 8944 2941 8953 2975
rect 8953 2941 8987 2975
rect 8987 2941 8996 2975
rect 8944 2932 8996 2941
rect 9496 2932 9548 2984
rect 9956 2932 10008 2984
rect 10324 2864 10376 2916
rect 14004 2932 14056 2984
rect 16672 2932 16724 2984
rect 18880 3009 18889 3043
rect 18889 3009 18923 3043
rect 18923 3009 18932 3043
rect 18880 3000 18932 3009
rect 20720 3136 20772 3188
rect 24584 3136 24636 3188
rect 21364 3111 21416 3120
rect 21364 3077 21373 3111
rect 21373 3077 21407 3111
rect 21407 3077 21416 3111
rect 21364 3068 21416 3077
rect 26056 3136 26108 3188
rect 26516 3179 26568 3188
rect 26516 3145 26525 3179
rect 26525 3145 26559 3179
rect 26559 3145 26568 3179
rect 26516 3136 26568 3145
rect 27620 3136 27672 3188
rect 27988 3179 28040 3188
rect 27988 3145 27997 3179
rect 27997 3145 28031 3179
rect 28031 3145 28040 3179
rect 27988 3136 28040 3145
rect 28908 3136 28960 3188
rect 31024 3179 31076 3188
rect 31024 3145 31033 3179
rect 31033 3145 31067 3179
rect 31067 3145 31076 3179
rect 31024 3136 31076 3145
rect 31944 3136 31996 3188
rect 34244 3179 34296 3188
rect 34244 3145 34253 3179
rect 34253 3145 34287 3179
rect 34287 3145 34296 3179
rect 34244 3136 34296 3145
rect 34520 3136 34572 3188
rect 26240 3068 26292 3120
rect 28632 3111 28684 3120
rect 28632 3077 28641 3111
rect 28641 3077 28675 3111
rect 28675 3077 28684 3111
rect 28632 3068 28684 3077
rect 20904 3000 20956 3052
rect 22468 3043 22520 3052
rect 19984 2932 20036 2984
rect 22468 3009 22477 3043
rect 22477 3009 22511 3043
rect 22511 3009 22520 3043
rect 22468 3000 22520 3009
rect 29736 3000 29788 3052
rect 30104 3043 30156 3052
rect 30104 3009 30113 3043
rect 30113 3009 30147 3043
rect 30147 3009 30156 3043
rect 30104 3000 30156 3009
rect 22652 2932 22704 2984
rect 20628 2864 20680 2916
rect 22100 2864 22152 2916
rect 23204 2932 23256 2984
rect 23756 2932 23808 2984
rect 26608 2975 26660 2984
rect 26608 2941 26624 2975
rect 26624 2941 26658 2975
rect 26658 2941 26660 2975
rect 26884 2975 26936 2984
rect 26608 2932 26660 2941
rect 23572 2864 23624 2916
rect 25688 2864 25740 2916
rect 26884 2941 26918 2975
rect 26918 2941 26936 2975
rect 26884 2932 26936 2941
rect 31116 2975 31168 2984
rect 31116 2941 31125 2975
rect 31125 2941 31159 2975
rect 31159 2941 31168 2975
rect 31116 2932 31168 2941
rect 3700 2839 3752 2848
rect 3700 2805 3709 2839
rect 3709 2805 3743 2839
rect 3743 2805 3752 2839
rect 3700 2796 3752 2805
rect 12440 2796 12492 2848
rect 13084 2839 13136 2848
rect 13084 2805 13093 2839
rect 13093 2805 13127 2839
rect 13127 2805 13136 2839
rect 13084 2796 13136 2805
rect 20812 2796 20864 2848
rect 21824 2839 21876 2848
rect 21824 2805 21833 2839
rect 21833 2805 21867 2839
rect 21867 2805 21876 2839
rect 21824 2796 21876 2805
rect 26608 2796 26660 2848
rect 29644 2864 29696 2916
rect 30656 2864 30708 2916
rect 29552 2839 29604 2848
rect 29552 2805 29561 2839
rect 29561 2805 29595 2839
rect 29595 2805 29604 2839
rect 29552 2796 29604 2805
rect 31576 3043 31628 3052
rect 31576 3009 31585 3043
rect 31585 3009 31619 3043
rect 31619 3009 31628 3043
rect 31576 3000 31628 3009
rect 32036 3000 32088 3052
rect 32956 3043 33008 3052
rect 32956 3009 32965 3043
rect 32965 3009 32999 3043
rect 32999 3009 33008 3043
rect 32956 3000 33008 3009
rect 35348 3043 35400 3052
rect 35348 3009 35357 3043
rect 35357 3009 35391 3043
rect 35391 3009 35400 3043
rect 35348 3000 35400 3009
rect 35440 3043 35492 3052
rect 35440 3009 35449 3043
rect 35449 3009 35483 3043
rect 35483 3009 35492 3043
rect 35440 3000 35492 3009
rect 37280 2864 37332 2916
rect 38292 2864 38344 2916
rect 33600 2839 33652 2848
rect 33600 2805 33609 2839
rect 33609 2805 33643 2839
rect 33643 2805 33652 2839
rect 33600 2796 33652 2805
rect 34888 2839 34940 2848
rect 34888 2805 34897 2839
rect 34897 2805 34931 2839
rect 34931 2805 34940 2839
rect 34888 2796 34940 2805
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 1768 2635 1820 2644
rect 1768 2601 1777 2635
rect 1777 2601 1811 2635
rect 1811 2601 1820 2635
rect 1768 2592 1820 2601
rect 2412 2635 2464 2644
rect 2412 2601 2421 2635
rect 2421 2601 2455 2635
rect 2455 2601 2464 2635
rect 2412 2592 2464 2601
rect 2780 2592 2832 2644
rect 3700 2592 3752 2644
rect 5448 2635 5500 2644
rect 5448 2601 5457 2635
rect 5457 2601 5491 2635
rect 5491 2601 5500 2635
rect 5448 2592 5500 2601
rect 7012 2592 7064 2644
rect 7196 2592 7248 2644
rect 8300 2635 8352 2644
rect 8300 2601 8309 2635
rect 8309 2601 8343 2635
rect 8343 2601 8352 2635
rect 8300 2592 8352 2601
rect 2964 2524 3016 2576
rect 9312 2592 9364 2644
rect 10324 2635 10376 2644
rect 10324 2601 10333 2635
rect 10333 2601 10367 2635
rect 10367 2601 10376 2635
rect 10324 2592 10376 2601
rect 10784 2592 10836 2644
rect 14096 2592 14148 2644
rect 16856 2635 16908 2644
rect 16856 2601 16865 2635
rect 16865 2601 16899 2635
rect 16899 2601 16908 2635
rect 16856 2592 16908 2601
rect 17868 2592 17920 2644
rect 10140 2524 10192 2576
rect 12440 2524 12492 2576
rect 13728 2524 13780 2576
rect 4804 2456 4856 2508
rect 6920 2456 6972 2508
rect 12072 2499 12124 2508
rect 3056 2431 3108 2440
rect 3056 2397 3065 2431
rect 3065 2397 3099 2431
rect 3099 2397 3108 2431
rect 3056 2388 3108 2397
rect 4068 2431 4120 2440
rect 4068 2397 4077 2431
rect 4077 2397 4111 2431
rect 4111 2397 4120 2431
rect 4068 2388 4120 2397
rect 8208 2388 8260 2440
rect 12072 2465 12081 2499
rect 12081 2465 12115 2499
rect 12115 2465 12124 2499
rect 12072 2456 12124 2465
rect 13636 2456 13688 2508
rect 9220 2431 9272 2440
rect 9220 2397 9229 2431
rect 9229 2397 9263 2431
rect 9263 2397 9272 2431
rect 9220 2388 9272 2397
rect 10784 2388 10836 2440
rect 12532 2388 12584 2440
rect 18972 2592 19024 2644
rect 19156 2592 19208 2644
rect 19984 2635 20036 2644
rect 19248 2524 19300 2576
rect 19984 2601 19993 2635
rect 19993 2601 20027 2635
rect 20027 2601 20036 2635
rect 19984 2592 20036 2601
rect 20720 2592 20772 2644
rect 22560 2635 22612 2644
rect 22560 2601 22569 2635
rect 22569 2601 22603 2635
rect 22603 2601 22612 2635
rect 22560 2592 22612 2601
rect 23756 2635 23808 2644
rect 23756 2601 23765 2635
rect 23765 2601 23799 2635
rect 23799 2601 23808 2635
rect 23756 2592 23808 2601
rect 25688 2635 25740 2644
rect 25688 2601 25697 2635
rect 25697 2601 25731 2635
rect 25731 2601 25740 2635
rect 25688 2592 25740 2601
rect 26240 2635 26292 2644
rect 26240 2601 26249 2635
rect 26249 2601 26283 2635
rect 26283 2601 26292 2635
rect 26608 2635 26660 2644
rect 26240 2592 26292 2601
rect 26608 2601 26617 2635
rect 26617 2601 26651 2635
rect 26651 2601 26660 2635
rect 26608 2592 26660 2601
rect 28632 2592 28684 2644
rect 20720 2456 20772 2508
rect 22008 2456 22060 2508
rect 24584 2567 24636 2576
rect 24584 2533 24618 2567
rect 24618 2533 24636 2567
rect 24584 2524 24636 2533
rect 27528 2524 27580 2576
rect 30196 2524 30248 2576
rect 34060 2592 34112 2644
rect 34796 2635 34848 2644
rect 34796 2601 34805 2635
rect 34805 2601 34839 2635
rect 34839 2601 34848 2635
rect 34796 2592 34848 2601
rect 35164 2635 35216 2644
rect 35164 2601 35173 2635
rect 35173 2601 35207 2635
rect 35207 2601 35216 2635
rect 35164 2592 35216 2601
rect 35348 2592 35400 2644
rect 37004 2635 37056 2644
rect 37004 2601 37013 2635
rect 37013 2601 37047 2635
rect 37047 2601 37056 2635
rect 37004 2592 37056 2601
rect 29644 2456 29696 2508
rect 33600 2456 33652 2508
rect 34796 2456 34848 2508
rect 35164 2388 35216 2440
rect 10968 2320 11020 2372
rect 28908 2320 28960 2372
rect 11060 2252 11112 2304
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 34966 2150 35018 2202
rect 35030 2150 35082 2202
rect 35094 2150 35146 2202
rect 35158 2150 35210 2202
<< metal2 >>
rect 36174 39400 36230 39409
rect 36174 39335 36230 39344
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 35622 37088 35678 37097
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 34940 37020 35236 37040
rect 35622 37023 35678 37032
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19580 36400 19876 36420
rect 33874 36136 33930 36145
rect 33874 36071 33930 36080
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 30472 35556 30524 35562
rect 30472 35498 30524 35504
rect 30012 35488 30064 35494
rect 30012 35430 30064 35436
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 29092 35080 29144 35086
rect 29092 35022 29144 35028
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 29104 34746 29132 35022
rect 29092 34740 29144 34746
rect 29092 34682 29144 34688
rect 29104 34626 29132 34682
rect 29012 34598 29132 34626
rect 29012 34490 29040 34598
rect 30024 34542 30052 35430
rect 30288 35284 30340 35290
rect 30288 35226 30340 35232
rect 30300 34542 30328 35226
rect 30484 35154 30512 35498
rect 30840 35488 30892 35494
rect 30840 35430 30892 35436
rect 30852 35290 30880 35430
rect 30840 35284 30892 35290
rect 30840 35226 30892 35232
rect 30472 35148 30524 35154
rect 30472 35090 30524 35096
rect 32036 35148 32088 35154
rect 32036 35090 32088 35096
rect 31668 34944 31720 34950
rect 31668 34886 31720 34892
rect 30380 34740 30432 34746
rect 30380 34682 30432 34688
rect 28920 34462 29040 34490
rect 30012 34536 30064 34542
rect 30012 34478 30064 34484
rect 30288 34536 30340 34542
rect 30288 34478 30340 34484
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 27712 34196 27764 34202
rect 27712 34138 27764 34144
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 27724 33658 27752 34138
rect 28724 34060 28776 34066
rect 28724 34002 28776 34008
rect 27988 33856 28040 33862
rect 27988 33798 28040 33804
rect 27712 33652 27764 33658
rect 27712 33594 27764 33600
rect 28000 33289 28028 33798
rect 28736 33658 28764 34002
rect 28920 33998 28948 34462
rect 29368 34400 29420 34406
rect 29368 34342 29420 34348
rect 29380 33998 29408 34342
rect 29736 34196 29788 34202
rect 29736 34138 29788 34144
rect 28908 33992 28960 33998
rect 28908 33934 28960 33940
rect 29368 33992 29420 33998
rect 29368 33934 29420 33940
rect 28724 33652 28776 33658
rect 28724 33594 28776 33600
rect 27986 33280 28042 33289
rect 19580 33212 19876 33232
rect 27986 33215 28042 33224
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 28920 33114 28948 33934
rect 29380 33318 29408 33934
rect 29748 33454 29776 34138
rect 30392 34082 30420 34682
rect 30300 34066 30420 34082
rect 30288 34060 30420 34066
rect 30340 34054 30420 34060
rect 31576 34060 31628 34066
rect 30288 34002 30340 34008
rect 31576 34002 31628 34008
rect 30932 33856 30984 33862
rect 30932 33798 30984 33804
rect 30944 33454 30972 33798
rect 29736 33448 29788 33454
rect 29736 33390 29788 33396
rect 30932 33448 30984 33454
rect 30932 33390 30984 33396
rect 29368 33312 29420 33318
rect 29368 33254 29420 33260
rect 28908 33108 28960 33114
rect 28908 33050 28960 33056
rect 29380 32910 29408 33254
rect 29748 33114 29776 33390
rect 31588 33318 31616 34002
rect 31680 33538 31708 34886
rect 32048 34678 32076 35090
rect 32772 35080 32824 35086
rect 32772 35022 32824 35028
rect 32784 34746 32812 35022
rect 33324 34944 33376 34950
rect 33324 34886 33376 34892
rect 33692 34944 33744 34950
rect 33692 34886 33744 34892
rect 32772 34740 32824 34746
rect 32772 34682 32824 34688
rect 33140 34740 33192 34746
rect 33140 34682 33192 34688
rect 32036 34672 32088 34678
rect 32034 34640 32036 34649
rect 32088 34640 32090 34649
rect 32034 34575 32090 34584
rect 32128 33992 32180 33998
rect 32128 33934 32180 33940
rect 32140 33658 32168 33934
rect 32772 33856 32824 33862
rect 32772 33798 32824 33804
rect 32128 33652 32180 33658
rect 32128 33594 32180 33600
rect 31680 33522 31800 33538
rect 32784 33522 32812 33798
rect 31680 33516 31812 33522
rect 31680 33510 31760 33516
rect 31760 33458 31812 33464
rect 32772 33516 32824 33522
rect 32772 33458 32824 33464
rect 31852 33380 31904 33386
rect 31852 33322 31904 33328
rect 30472 33312 30524 33318
rect 30472 33254 30524 33260
rect 31576 33312 31628 33318
rect 31864 33289 31892 33322
rect 32128 33312 32180 33318
rect 31576 33254 31628 33260
rect 31850 33280 31906 33289
rect 29826 33144 29882 33153
rect 29736 33108 29788 33114
rect 29826 33079 29882 33088
rect 29736 33050 29788 33056
rect 29840 33046 29868 33079
rect 29828 33040 29880 33046
rect 29828 32982 29880 32988
rect 29368 32904 29420 32910
rect 29368 32846 29420 32852
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 29380 32366 29408 32846
rect 29840 32570 29868 32982
rect 29828 32564 29880 32570
rect 29828 32506 29880 32512
rect 29368 32360 29420 32366
rect 29368 32302 29420 32308
rect 29380 32230 29408 32302
rect 29368 32224 29420 32230
rect 29368 32166 29420 32172
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 28908 31884 28960 31890
rect 28908 31826 28960 31832
rect 28920 31770 28948 31826
rect 28920 31742 29040 31770
rect 29380 31754 29408 32166
rect 29840 31890 29868 32506
rect 30104 32224 30156 32230
rect 30104 32166 30156 32172
rect 29828 31884 29880 31890
rect 29828 31826 29880 31832
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 29012 31482 29040 31742
rect 29368 31748 29420 31754
rect 29368 31690 29420 31696
rect 29000 31476 29052 31482
rect 29000 31418 29052 31424
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 29380 30802 29408 31690
rect 29840 31482 29868 31826
rect 29920 31748 29972 31754
rect 29920 31690 29972 31696
rect 29932 31482 29960 31690
rect 29828 31476 29880 31482
rect 29828 31418 29880 31424
rect 29920 31476 29972 31482
rect 29920 31418 29972 31424
rect 30116 30870 30144 32166
rect 30380 32020 30432 32026
rect 30380 31962 30432 31968
rect 30288 31952 30340 31958
rect 30288 31894 30340 31900
rect 30300 30920 30328 31894
rect 30392 31346 30420 31962
rect 30484 31822 30512 33254
rect 32128 33254 32180 33260
rect 31850 33215 31906 33224
rect 31864 33114 31892 33215
rect 31852 33108 31904 33114
rect 31852 33050 31904 33056
rect 32036 32972 32088 32978
rect 32036 32914 32088 32920
rect 31760 32836 31812 32842
rect 31760 32778 31812 32784
rect 30932 32768 30984 32774
rect 30932 32710 30984 32716
rect 30944 32298 30972 32710
rect 30932 32292 30984 32298
rect 30932 32234 30984 32240
rect 30472 31816 30524 31822
rect 30472 31758 30524 31764
rect 30562 31376 30618 31385
rect 30380 31340 30432 31346
rect 31772 31362 31800 32778
rect 32048 32570 32076 32914
rect 32036 32564 32088 32570
rect 32036 32506 32088 32512
rect 32140 32366 32168 33254
rect 32588 32904 32640 32910
rect 32588 32846 32640 32852
rect 32600 32570 32628 32846
rect 32588 32564 32640 32570
rect 32588 32506 32640 32512
rect 32128 32360 32180 32366
rect 32128 32302 32180 32308
rect 32600 32298 32628 32506
rect 32784 32502 32812 33458
rect 33152 32910 33180 34682
rect 33336 34542 33364 34886
rect 33324 34536 33376 34542
rect 33324 34478 33376 34484
rect 33232 34400 33284 34406
rect 33232 34342 33284 34348
rect 33244 33114 33272 34342
rect 33508 33856 33560 33862
rect 33508 33798 33560 33804
rect 33520 33153 33548 33798
rect 33506 33144 33562 33153
rect 33232 33108 33284 33114
rect 33506 33079 33562 33088
rect 33232 33050 33284 33056
rect 33140 32904 33192 32910
rect 33140 32846 33192 32852
rect 32772 32496 32824 32502
rect 32772 32438 32824 32444
rect 32588 32292 32640 32298
rect 32588 32234 32640 32240
rect 32036 32224 32088 32230
rect 32036 32166 32088 32172
rect 30562 31311 30564 31320
rect 30380 31282 30432 31288
rect 30616 31311 30618 31320
rect 31680 31334 31800 31362
rect 32048 31346 32076 32166
rect 33152 31958 33180 32846
rect 33244 32366 33272 33050
rect 33416 32496 33468 32502
rect 33416 32438 33468 32444
rect 33232 32360 33284 32366
rect 33232 32302 33284 32308
rect 33232 32224 33284 32230
rect 33232 32166 33284 32172
rect 33140 31952 33192 31958
rect 33140 31894 33192 31900
rect 33244 31890 33272 32166
rect 33428 32026 33456 32438
rect 33704 32434 33732 34886
rect 33888 33658 33916 36071
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 35636 35834 35664 37023
rect 35624 35828 35676 35834
rect 35624 35770 35676 35776
rect 35440 35624 35492 35630
rect 35440 35566 35492 35572
rect 34704 35148 34756 35154
rect 34704 35090 34756 35096
rect 34520 34944 34572 34950
rect 34520 34886 34572 34892
rect 34152 34740 34204 34746
rect 34152 34682 34204 34688
rect 34164 34610 34192 34682
rect 34428 34672 34480 34678
rect 34428 34614 34480 34620
rect 34152 34604 34204 34610
rect 34152 34546 34204 34552
rect 34164 34202 34192 34546
rect 34440 34218 34468 34614
rect 34532 34610 34560 34886
rect 34520 34604 34572 34610
rect 34520 34546 34572 34552
rect 34612 34400 34664 34406
rect 34612 34342 34664 34348
rect 34152 34196 34204 34202
rect 34152 34138 34204 34144
rect 34348 34190 34560 34218
rect 33876 33652 33928 33658
rect 33876 33594 33928 33600
rect 34244 33584 34296 33590
rect 34244 33526 34296 33532
rect 34256 32910 34284 33526
rect 34348 33114 34376 34190
rect 34532 34134 34560 34190
rect 34520 34128 34572 34134
rect 34520 34070 34572 34076
rect 34624 33998 34652 34342
rect 34612 33992 34664 33998
rect 34612 33934 34664 33940
rect 34624 33590 34652 33934
rect 34716 33862 34744 35090
rect 34796 35012 34848 35018
rect 34796 34954 34848 34960
rect 34808 34746 34836 34954
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34940 34768 35236 34788
rect 34796 34740 34848 34746
rect 34796 34682 34848 34688
rect 34704 33856 34756 33862
rect 34704 33798 34756 33804
rect 34612 33584 34664 33590
rect 34612 33526 34664 33532
rect 34716 33386 34744 33798
rect 34808 33538 34836 34682
rect 34940 33756 35236 33776
rect 34996 33754 35020 33756
rect 35076 33754 35100 33756
rect 35156 33754 35180 33756
rect 35018 33702 35020 33754
rect 35082 33702 35094 33754
rect 35156 33702 35158 33754
rect 34996 33700 35020 33702
rect 35076 33700 35100 33702
rect 35156 33700 35180 33702
rect 34940 33680 35236 33700
rect 34808 33510 34928 33538
rect 34704 33380 34756 33386
rect 34704 33322 34756 33328
rect 34796 33312 34848 33318
rect 34796 33254 34848 33260
rect 34336 33108 34388 33114
rect 34336 33050 34388 33056
rect 34244 32904 34296 32910
rect 34244 32846 34296 32852
rect 34256 32570 34284 32846
rect 34244 32564 34296 32570
rect 34244 32506 34296 32512
rect 34428 32564 34480 32570
rect 34428 32506 34480 32512
rect 33692 32428 33744 32434
rect 33692 32370 33744 32376
rect 33416 32020 33468 32026
rect 33416 31962 33468 31968
rect 33784 32020 33836 32026
rect 33784 31962 33836 31968
rect 32956 31884 33008 31890
rect 32956 31826 33008 31832
rect 33232 31884 33284 31890
rect 33232 31826 33284 31832
rect 32128 31680 32180 31686
rect 32128 31622 32180 31628
rect 32140 31346 32168 31622
rect 32968 31482 32996 31826
rect 33048 31680 33100 31686
rect 33048 31622 33100 31628
rect 32956 31476 33008 31482
rect 32956 31418 33008 31424
rect 32036 31340 32088 31346
rect 30564 31282 30616 31288
rect 31680 31210 31708 31334
rect 32036 31282 32088 31288
rect 32128 31340 32180 31346
rect 32128 31282 32180 31288
rect 31668 31204 31720 31210
rect 31668 31146 31720 31152
rect 31576 31136 31628 31142
rect 31576 31078 31628 31084
rect 31944 31136 31996 31142
rect 31944 31078 31996 31084
rect 30380 30932 30432 30938
rect 30300 30892 30380 30920
rect 30380 30874 30432 30880
rect 30104 30864 30156 30870
rect 30104 30806 30156 30812
rect 29368 30796 29420 30802
rect 29368 30738 29420 30744
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 28816 30320 28868 30326
rect 28816 30262 28868 30268
rect 28724 30252 28776 30258
rect 28724 30194 28776 30200
rect 27988 30048 28040 30054
rect 27988 29990 28040 29996
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 27712 29504 27764 29510
rect 27712 29446 27764 29452
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 27724 29102 27752 29446
rect 28000 29306 28028 29990
rect 28736 29714 28764 30194
rect 28724 29708 28776 29714
rect 28724 29650 28776 29656
rect 28448 29504 28500 29510
rect 28448 29446 28500 29452
rect 27988 29300 28040 29306
rect 27988 29242 28040 29248
rect 28460 29170 28488 29446
rect 28736 29238 28764 29650
rect 28724 29232 28776 29238
rect 28724 29174 28776 29180
rect 28448 29164 28500 29170
rect 28448 29106 28500 29112
rect 27712 29096 27764 29102
rect 27712 29038 27764 29044
rect 28172 29028 28224 29034
rect 28172 28970 28224 28976
rect 27620 28960 27672 28966
rect 27620 28902 27672 28908
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19580 27696 19876 27716
rect 23112 27532 23164 27538
rect 23112 27474 23164 27480
rect 24308 27532 24360 27538
rect 24308 27474 24360 27480
rect 21916 27328 21968 27334
rect 21916 27270 21968 27276
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 21824 26988 21876 26994
rect 21824 26930 21876 26936
rect 19580 26684 19876 26704
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 20904 26376 20956 26382
rect 20904 26318 20956 26324
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 20916 26042 20944 26318
rect 21180 26240 21232 26246
rect 21180 26182 21232 26188
rect 20904 26036 20956 26042
rect 20904 25978 20956 25984
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 20916 25362 20944 25978
rect 21192 25770 21220 26182
rect 21180 25764 21232 25770
rect 21180 25706 21232 25712
rect 21548 25764 21600 25770
rect 21548 25706 21600 25712
rect 20904 25356 20956 25362
rect 20904 25298 20956 25304
rect 21180 25356 21232 25362
rect 21180 25298 21232 25304
rect 20628 25152 20680 25158
rect 20628 25094 20680 25100
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 20536 24812 20588 24818
rect 20536 24754 20588 24760
rect 20260 24608 20312 24614
rect 20260 24550 20312 24556
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 20272 24342 20300 24550
rect 20548 24410 20576 24754
rect 20640 24698 20668 25094
rect 20916 24954 20944 25298
rect 20904 24948 20956 24954
rect 20904 24890 20956 24896
rect 20640 24682 20760 24698
rect 20640 24676 20772 24682
rect 20640 24670 20720 24676
rect 20720 24618 20772 24624
rect 20536 24404 20588 24410
rect 20536 24346 20588 24352
rect 20260 24336 20312 24342
rect 20260 24278 20312 24284
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 20272 23866 20300 24278
rect 20732 23866 20760 24618
rect 21192 24342 21220 25298
rect 21560 25158 21588 25706
rect 21548 25152 21600 25158
rect 21548 25094 21600 25100
rect 21180 24336 21232 24342
rect 21180 24278 21232 24284
rect 21560 24274 21588 25094
rect 21548 24268 21600 24274
rect 21548 24210 21600 24216
rect 21560 23866 21588 24210
rect 21836 24206 21864 26930
rect 21928 26926 21956 27270
rect 21916 26920 21968 26926
rect 21916 26862 21968 26868
rect 21928 26586 21956 26862
rect 23124 26790 23152 27474
rect 23296 27328 23348 27334
rect 23296 27270 23348 27276
rect 22008 26784 22060 26790
rect 22008 26726 22060 26732
rect 22284 26784 22336 26790
rect 22284 26726 22336 26732
rect 22744 26784 22796 26790
rect 22744 26726 22796 26732
rect 23112 26784 23164 26790
rect 23112 26726 23164 26732
rect 21916 26580 21968 26586
rect 21916 26522 21968 26528
rect 21916 24608 21968 24614
rect 21916 24550 21968 24556
rect 21928 24342 21956 24550
rect 22020 24426 22048 26726
rect 22296 26518 22324 26726
rect 22284 26512 22336 26518
rect 22284 26454 22336 26460
rect 22296 26042 22324 26454
rect 22284 26036 22336 26042
rect 22284 25978 22336 25984
rect 22020 24398 22140 24426
rect 22756 24410 22784 26726
rect 23308 26353 23336 27270
rect 23294 26344 23350 26353
rect 23294 26279 23350 26288
rect 24032 25832 24084 25838
rect 24032 25774 24084 25780
rect 24044 25498 24072 25774
rect 24032 25492 24084 25498
rect 24032 25434 24084 25440
rect 24124 25288 24176 25294
rect 24124 25230 24176 25236
rect 23480 24608 23532 24614
rect 23400 24568 23480 24596
rect 22112 24342 22140 24398
rect 22744 24404 22796 24410
rect 22744 24346 22796 24352
rect 21916 24336 21968 24342
rect 21916 24278 21968 24284
rect 22100 24336 22152 24342
rect 22100 24278 22152 24284
rect 23112 24336 23164 24342
rect 23112 24278 23164 24284
rect 21824 24200 21876 24206
rect 21824 24142 21876 24148
rect 22836 24200 22888 24206
rect 22836 24142 22888 24148
rect 21836 24041 21864 24142
rect 22848 24070 22876 24142
rect 22836 24064 22888 24070
rect 21822 24032 21878 24041
rect 22836 24006 22888 24012
rect 21822 23967 21878 23976
rect 20260 23860 20312 23866
rect 20260 23802 20312 23808
rect 20720 23860 20772 23866
rect 20720 23802 20772 23808
rect 21548 23860 21600 23866
rect 21548 23802 21600 23808
rect 20732 23662 20760 23802
rect 21836 23730 21864 23967
rect 22848 23866 22876 24006
rect 23124 23866 23152 24278
rect 22836 23860 22888 23866
rect 22836 23802 22888 23808
rect 23112 23860 23164 23866
rect 23112 23802 23164 23808
rect 21824 23724 21876 23730
rect 21824 23666 21876 23672
rect 20720 23656 20772 23662
rect 20720 23598 20772 23604
rect 19984 23520 20036 23526
rect 19984 23462 20036 23468
rect 20996 23520 21048 23526
rect 20996 23462 21048 23468
rect 21180 23520 21232 23526
rect 21180 23462 21232 23468
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 19996 23322 20024 23462
rect 19984 23316 20036 23322
rect 19984 23258 20036 23264
rect 21008 23186 21036 23462
rect 21192 23361 21220 23462
rect 21178 23352 21234 23361
rect 21836 23322 21864 23666
rect 22100 23656 22152 23662
rect 22100 23598 22152 23604
rect 22112 23322 22140 23598
rect 23400 23322 23428 24568
rect 23480 24550 23532 24556
rect 23848 24608 23900 24614
rect 23848 24550 23900 24556
rect 23860 23662 23888 24550
rect 24136 24070 24164 25230
rect 24320 24410 24348 27474
rect 24768 27328 24820 27334
rect 24768 27270 24820 27276
rect 24676 26920 24728 26926
rect 24676 26862 24728 26868
rect 24688 26450 24716 26862
rect 24676 26444 24728 26450
rect 24676 26386 24728 26392
rect 24584 26240 24636 26246
rect 24584 26182 24636 26188
rect 24596 25770 24624 26182
rect 24688 25838 24716 26386
rect 24676 25832 24728 25838
rect 24676 25774 24728 25780
rect 24584 25764 24636 25770
rect 24584 25706 24636 25712
rect 24596 25430 24624 25706
rect 24676 25492 24728 25498
rect 24676 25434 24728 25440
rect 24584 25424 24636 25430
rect 24584 25366 24636 25372
rect 24398 25256 24454 25265
rect 24398 25191 24454 25200
rect 24308 24404 24360 24410
rect 24308 24346 24360 24352
rect 24124 24064 24176 24070
rect 24122 24032 24124 24041
rect 24176 24032 24178 24041
rect 24122 23967 24178 23976
rect 24412 23798 24440 25191
rect 24596 24886 24624 25366
rect 24688 24954 24716 25434
rect 24780 25242 24808 27270
rect 25320 26852 25372 26858
rect 25320 26794 25372 26800
rect 25332 26042 25360 26794
rect 26056 26784 26108 26790
rect 26056 26726 26108 26732
rect 27528 26784 27580 26790
rect 27528 26726 27580 26732
rect 25320 26036 25372 26042
rect 25320 25978 25372 25984
rect 25332 25498 25360 25978
rect 26068 25770 26096 26726
rect 26516 26444 26568 26450
rect 26516 26386 26568 26392
rect 26792 26444 26844 26450
rect 26792 26386 26844 26392
rect 26422 26344 26478 26353
rect 26422 26279 26478 26288
rect 26056 25764 26108 25770
rect 26056 25706 26108 25712
rect 26068 25498 26096 25706
rect 25320 25492 25372 25498
rect 25320 25434 25372 25440
rect 26056 25492 26108 25498
rect 26056 25434 26108 25440
rect 25504 25424 25556 25430
rect 25504 25366 25556 25372
rect 24780 25214 24900 25242
rect 24768 25152 24820 25158
rect 24768 25094 24820 25100
rect 24676 24948 24728 24954
rect 24676 24890 24728 24896
rect 24584 24880 24636 24886
rect 24584 24822 24636 24828
rect 24780 24342 24808 25094
rect 24872 24750 24900 25214
rect 24860 24744 24912 24750
rect 24860 24686 24912 24692
rect 25516 24614 25544 25366
rect 25596 25288 25648 25294
rect 25596 25230 25648 25236
rect 25608 24818 25636 25230
rect 26240 25152 26292 25158
rect 26160 25100 26240 25106
rect 26160 25094 26292 25100
rect 26160 25078 26280 25094
rect 25596 24812 25648 24818
rect 25596 24754 25648 24760
rect 26160 24682 26188 25078
rect 26436 24818 26464 26279
rect 26528 25838 26556 26386
rect 26516 25832 26568 25838
rect 26516 25774 26568 25780
rect 26700 25356 26752 25362
rect 26700 25298 26752 25304
rect 26712 25265 26740 25298
rect 26698 25256 26754 25265
rect 26698 25191 26754 25200
rect 26712 24954 26740 25191
rect 26804 25158 26832 26386
rect 27436 26240 27488 26246
rect 27436 26182 27488 26188
rect 27448 25498 27476 26182
rect 27436 25492 27488 25498
rect 27436 25434 27488 25440
rect 26792 25152 26844 25158
rect 26792 25094 26844 25100
rect 26700 24948 26752 24954
rect 26700 24890 26752 24896
rect 26424 24812 26476 24818
rect 26424 24754 26476 24760
rect 27160 24812 27212 24818
rect 27160 24754 27212 24760
rect 26884 24744 26936 24750
rect 26884 24686 26936 24692
rect 26148 24676 26200 24682
rect 26148 24618 26200 24624
rect 26896 24614 26924 24686
rect 25044 24608 25096 24614
rect 25044 24550 25096 24556
rect 25412 24608 25464 24614
rect 25412 24550 25464 24556
rect 25504 24608 25556 24614
rect 26884 24608 26936 24614
rect 25504 24550 25556 24556
rect 26606 24576 26662 24585
rect 25056 24410 25084 24550
rect 25424 24410 25452 24550
rect 26884 24550 26936 24556
rect 26606 24511 26662 24520
rect 25044 24404 25096 24410
rect 25044 24346 25096 24352
rect 25412 24404 25464 24410
rect 25412 24346 25464 24352
rect 26148 24404 26200 24410
rect 26148 24346 26200 24352
rect 24768 24336 24820 24342
rect 24768 24278 24820 24284
rect 24780 23866 24808 24278
rect 24768 23860 24820 23866
rect 24768 23802 24820 23808
rect 24400 23792 24452 23798
rect 24400 23734 24452 23740
rect 23848 23656 23900 23662
rect 23848 23598 23900 23604
rect 23754 23352 23810 23361
rect 21178 23287 21234 23296
rect 21824 23316 21876 23322
rect 21824 23258 21876 23264
rect 22100 23316 22152 23322
rect 22100 23258 22152 23264
rect 23388 23316 23440 23322
rect 23860 23322 23888 23598
rect 24860 23588 24912 23594
rect 24860 23530 24912 23536
rect 24872 23322 24900 23530
rect 23754 23287 23756 23296
rect 23388 23258 23440 23264
rect 23808 23287 23810 23296
rect 23848 23316 23900 23322
rect 23756 23258 23808 23264
rect 23848 23258 23900 23264
rect 24860 23316 24912 23322
rect 24860 23258 24912 23264
rect 20628 23180 20680 23186
rect 20628 23122 20680 23128
rect 20996 23180 21048 23186
rect 20996 23122 21048 23128
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 20640 22438 20668 23122
rect 20904 23112 20956 23118
rect 20904 23054 20956 23060
rect 21546 23080 21602 23089
rect 20916 22778 20944 23054
rect 21546 23015 21602 23024
rect 21560 22778 21588 23015
rect 20904 22772 20956 22778
rect 20904 22714 20956 22720
rect 21548 22772 21600 22778
rect 21548 22714 21600 22720
rect 20628 22432 20680 22438
rect 20628 22374 20680 22380
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 20640 22234 20668 22374
rect 20628 22228 20680 22234
rect 20628 22170 20680 22176
rect 20720 22092 20772 22098
rect 20720 22034 20772 22040
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 20732 21146 20760 22034
rect 20916 22030 20944 22714
rect 21836 22642 21864 23258
rect 21824 22636 21876 22642
rect 21824 22578 21876 22584
rect 21364 22432 21416 22438
rect 21364 22374 21416 22380
rect 20904 22024 20956 22030
rect 20904 21966 20956 21972
rect 20916 21690 20944 21966
rect 20904 21684 20956 21690
rect 20904 21626 20956 21632
rect 20720 21140 20772 21146
rect 20720 21082 20772 21088
rect 20916 21010 20944 21626
rect 21376 21418 21404 22374
rect 21836 22166 21864 22578
rect 23664 22568 23716 22574
rect 23664 22510 23716 22516
rect 21916 22432 21968 22438
rect 21916 22374 21968 22380
rect 23112 22432 23164 22438
rect 23112 22374 23164 22380
rect 21824 22160 21876 22166
rect 21824 22102 21876 22108
rect 21928 22098 21956 22374
rect 23124 22234 23152 22374
rect 23112 22228 23164 22234
rect 23112 22170 23164 22176
rect 21916 22092 21968 22098
rect 21916 22034 21968 22040
rect 23204 22092 23256 22098
rect 23204 22034 23256 22040
rect 21928 21690 21956 22034
rect 21916 21684 21968 21690
rect 21916 21626 21968 21632
rect 21364 21412 21416 21418
rect 21364 21354 21416 21360
rect 22284 21412 22336 21418
rect 22284 21354 22336 21360
rect 22296 21146 22324 21354
rect 23216 21146 23244 22034
rect 23676 21690 23704 22510
rect 23768 22438 23796 23258
rect 24952 23180 25004 23186
rect 24952 23122 25004 23128
rect 23848 23112 23900 23118
rect 23846 23080 23848 23089
rect 24032 23112 24084 23118
rect 23900 23080 23902 23089
rect 24032 23054 24084 23060
rect 23846 23015 23902 23024
rect 23860 22778 23888 23015
rect 23848 22772 23900 22778
rect 23848 22714 23900 22720
rect 24044 22642 24072 23054
rect 24964 22710 24992 23122
rect 25056 23118 25084 24346
rect 25412 24200 25464 24206
rect 25412 24142 25464 24148
rect 25424 23526 25452 24142
rect 26160 23866 26188 24346
rect 26620 23866 26648 24511
rect 27172 24410 27200 24754
rect 27160 24404 27212 24410
rect 27160 24346 27212 24352
rect 27540 24274 27568 26726
rect 27528 24268 27580 24274
rect 27528 24210 27580 24216
rect 27540 23866 27568 24210
rect 26148 23860 26200 23866
rect 26148 23802 26200 23808
rect 26608 23860 26660 23866
rect 26608 23802 26660 23808
rect 27528 23860 27580 23866
rect 27528 23802 27580 23808
rect 26620 23662 26648 23802
rect 27632 23662 27660 28902
rect 27988 28620 28040 28626
rect 27988 28562 28040 28568
rect 28000 28218 28028 28562
rect 27988 28212 28040 28218
rect 27988 28154 28040 28160
rect 28184 28082 28212 28970
rect 28460 28694 28488 29106
rect 28448 28688 28500 28694
rect 28448 28630 28500 28636
rect 28460 28218 28488 28630
rect 28736 28626 28764 29174
rect 28724 28620 28776 28626
rect 28724 28562 28776 28568
rect 28632 28416 28684 28422
rect 28632 28358 28684 28364
rect 28448 28212 28500 28218
rect 28448 28154 28500 28160
rect 28172 28076 28224 28082
rect 28172 28018 28224 28024
rect 27896 26852 27948 26858
rect 27896 26794 27948 26800
rect 27908 26586 27936 26794
rect 27896 26580 27948 26586
rect 27896 26522 27948 26528
rect 27908 26042 27936 26522
rect 28448 26444 28500 26450
rect 28448 26386 28500 26392
rect 27896 26036 27948 26042
rect 27896 25978 27948 25984
rect 27804 25696 27856 25702
rect 27804 25638 27856 25644
rect 27816 25158 27844 25638
rect 28264 25356 28316 25362
rect 28264 25298 28316 25304
rect 27804 25152 27856 25158
rect 27804 25094 27856 25100
rect 28276 24682 28304 25298
rect 28356 25288 28408 25294
rect 28356 25230 28408 25236
rect 28368 24954 28396 25230
rect 28356 24948 28408 24954
rect 28356 24890 28408 24896
rect 28264 24676 28316 24682
rect 28264 24618 28316 24624
rect 28264 24336 28316 24342
rect 28264 24278 28316 24284
rect 28276 23730 28304 24278
rect 28460 24274 28488 26386
rect 28644 24342 28672 28358
rect 28736 27130 28764 28562
rect 28828 28098 28856 30262
rect 29380 30258 29408 30738
rect 29552 30592 29604 30598
rect 29552 30534 29604 30540
rect 29368 30252 29420 30258
rect 29368 30194 29420 30200
rect 29564 30122 29592 30534
rect 29552 30116 29604 30122
rect 29552 30058 29604 30064
rect 29092 30048 29144 30054
rect 29092 29990 29144 29996
rect 29104 29782 29132 29990
rect 30116 29850 30144 30806
rect 30840 30592 30892 30598
rect 30840 30534 30892 30540
rect 30654 30288 30710 30297
rect 30654 30223 30710 30232
rect 30104 29844 30156 29850
rect 30104 29786 30156 29792
rect 30668 29782 30696 30223
rect 29092 29776 29144 29782
rect 29092 29718 29144 29724
rect 30656 29776 30708 29782
rect 30656 29718 30708 29724
rect 29104 29238 29132 29718
rect 30668 29306 30696 29718
rect 30852 29714 30880 30534
rect 30840 29708 30892 29714
rect 30840 29650 30892 29656
rect 30748 29504 30800 29510
rect 30748 29446 30800 29452
rect 30656 29300 30708 29306
rect 30656 29242 30708 29248
rect 29092 29232 29144 29238
rect 29092 29174 29144 29180
rect 29828 29232 29880 29238
rect 29828 29174 29880 29180
rect 28908 29096 28960 29102
rect 28960 29044 29040 29050
rect 28908 29038 29040 29044
rect 28920 29022 29040 29038
rect 29012 28218 29040 29022
rect 29092 28756 29144 28762
rect 29092 28698 29144 28704
rect 29000 28212 29052 28218
rect 29000 28154 29052 28160
rect 28828 28082 29040 28098
rect 28828 28076 29052 28082
rect 28828 28070 29000 28076
rect 29000 28018 29052 28024
rect 28908 27532 28960 27538
rect 28908 27474 28960 27480
rect 28816 27328 28868 27334
rect 28816 27270 28868 27276
rect 28724 27124 28776 27130
rect 28724 27066 28776 27072
rect 28724 26784 28776 26790
rect 28722 26752 28724 26761
rect 28776 26752 28778 26761
rect 28722 26687 28778 26696
rect 28828 25514 28856 27270
rect 28920 26314 28948 27474
rect 29000 27464 29052 27470
rect 29000 27406 29052 27412
rect 28908 26308 28960 26314
rect 28908 26250 28960 26256
rect 29012 26042 29040 27406
rect 29000 26036 29052 26042
rect 29000 25978 29052 25984
rect 28828 25486 29040 25514
rect 29012 25430 29040 25486
rect 29000 25424 29052 25430
rect 29000 25366 29052 25372
rect 28724 25288 28776 25294
rect 28724 25230 28776 25236
rect 28736 24614 28764 25230
rect 28724 24608 28776 24614
rect 28724 24550 28776 24556
rect 28736 24410 28764 24550
rect 28724 24404 28776 24410
rect 28724 24346 28776 24352
rect 28632 24336 28684 24342
rect 28632 24278 28684 24284
rect 28448 24268 28500 24274
rect 28448 24210 28500 24216
rect 28460 23866 28488 24210
rect 28448 23860 28500 23866
rect 28448 23802 28500 23808
rect 28264 23724 28316 23730
rect 28264 23666 28316 23672
rect 26608 23656 26660 23662
rect 26608 23598 26660 23604
rect 26976 23656 27028 23662
rect 26976 23598 27028 23604
rect 27620 23656 27672 23662
rect 27620 23598 27672 23604
rect 25412 23520 25464 23526
rect 25412 23462 25464 23468
rect 25044 23112 25096 23118
rect 25044 23054 25096 23060
rect 25424 22778 25452 23462
rect 26988 23322 27016 23598
rect 28172 23520 28224 23526
rect 28172 23462 28224 23468
rect 27158 23352 27214 23361
rect 26976 23316 27028 23322
rect 27158 23287 27214 23296
rect 26976 23258 27028 23264
rect 25412 22772 25464 22778
rect 25412 22714 25464 22720
rect 24952 22704 25004 22710
rect 24952 22646 25004 22652
rect 25870 22672 25926 22681
rect 24032 22636 24084 22642
rect 24032 22578 24084 22584
rect 23756 22432 23808 22438
rect 23756 22374 23808 22380
rect 24044 22234 24072 22578
rect 24964 22234 24992 22646
rect 25870 22607 25872 22616
rect 25924 22607 25926 22616
rect 26240 22636 26292 22642
rect 25872 22578 25924 22584
rect 26240 22578 26292 22584
rect 25778 22264 25834 22273
rect 24032 22228 24084 22234
rect 24032 22170 24084 22176
rect 24952 22228 25004 22234
rect 25778 22199 25834 22208
rect 24952 22170 25004 22176
rect 23756 22160 23808 22166
rect 23756 22102 23808 22108
rect 24768 22160 24820 22166
rect 24768 22102 24820 22108
rect 23664 21684 23716 21690
rect 23664 21626 23716 21632
rect 23664 21344 23716 21350
rect 23664 21286 23716 21292
rect 22284 21140 22336 21146
rect 22284 21082 22336 21088
rect 23204 21140 23256 21146
rect 23204 21082 23256 21088
rect 23676 21078 23704 21286
rect 21364 21072 21416 21078
rect 21364 21014 21416 21020
rect 23480 21072 23532 21078
rect 23480 21014 23532 21020
rect 23664 21072 23716 21078
rect 23664 21014 23716 21020
rect 20904 21004 20956 21010
rect 20904 20946 20956 20952
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 20916 20602 20944 20946
rect 21376 20777 21404 21014
rect 23296 20936 23348 20942
rect 23296 20878 23348 20884
rect 21362 20768 21418 20777
rect 21362 20703 21418 20712
rect 21376 20602 21404 20703
rect 20904 20596 20956 20602
rect 20904 20538 20956 20544
rect 21364 20596 21416 20602
rect 21364 20538 21416 20544
rect 22468 20528 22520 20534
rect 22468 20470 22520 20476
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 3422 20088 3478 20097
rect 19580 20080 19876 20100
rect 3422 20023 3478 20032
rect 3436 18193 3464 20023
rect 22480 19854 22508 20470
rect 23308 20330 23336 20878
rect 23492 20618 23520 21014
rect 23768 20777 23796 22102
rect 24216 22024 24268 22030
rect 24216 21966 24268 21972
rect 24228 21554 24256 21966
rect 24676 21888 24728 21894
rect 24676 21830 24728 21836
rect 24216 21548 24268 21554
rect 24216 21490 24268 21496
rect 23940 21412 23992 21418
rect 23940 21354 23992 21360
rect 23754 20768 23810 20777
rect 23754 20703 23810 20712
rect 23400 20602 23520 20618
rect 23388 20596 23520 20602
rect 23440 20590 23520 20596
rect 23388 20538 23440 20544
rect 23296 20324 23348 20330
rect 23296 20266 23348 20272
rect 22742 20224 22798 20233
rect 22742 20159 22798 20168
rect 22756 19922 22784 20159
rect 22744 19916 22796 19922
rect 22744 19858 22796 19864
rect 22468 19848 22520 19854
rect 22468 19790 22520 19796
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 22480 19446 22508 19790
rect 22756 19514 22784 19858
rect 22744 19508 22796 19514
rect 22744 19450 22796 19456
rect 23308 19446 23336 20266
rect 23768 20058 23796 20703
rect 23952 20398 23980 21354
rect 24688 21350 24716 21830
rect 24780 21690 24808 22102
rect 25792 22098 25820 22199
rect 25320 22092 25372 22098
rect 25320 22034 25372 22040
rect 25780 22092 25832 22098
rect 25780 22034 25832 22040
rect 25332 21690 25360 22034
rect 26054 21992 26110 22001
rect 26054 21927 26110 21936
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 25320 21684 25372 21690
rect 25320 21626 25372 21632
rect 24768 21412 24820 21418
rect 24768 21354 24820 21360
rect 24124 21344 24176 21350
rect 24122 21312 24124 21321
rect 24676 21344 24728 21350
rect 24176 21312 24178 21321
rect 24676 21286 24728 21292
rect 24122 21247 24178 21256
rect 23940 20392 23992 20398
rect 23940 20334 23992 20340
rect 23952 20058 23980 20334
rect 24688 20233 24716 21286
rect 24780 21146 24808 21354
rect 26068 21350 26096 21927
rect 25228 21344 25280 21350
rect 25228 21286 25280 21292
rect 26056 21344 26108 21350
rect 26056 21286 26108 21292
rect 24768 21140 24820 21146
rect 24768 21082 24820 21088
rect 25240 21010 25268 21286
rect 25228 21004 25280 21010
rect 25228 20946 25280 20952
rect 25872 20596 25924 20602
rect 25872 20538 25924 20544
rect 25044 20256 25096 20262
rect 24674 20224 24730 20233
rect 24674 20159 24730 20168
rect 25042 20224 25044 20233
rect 25096 20224 25098 20233
rect 25042 20159 25098 20168
rect 23756 20052 23808 20058
rect 23756 19994 23808 20000
rect 23940 20052 23992 20058
rect 23940 19994 23992 20000
rect 22468 19440 22520 19446
rect 22468 19382 22520 19388
rect 23296 19440 23348 19446
rect 23296 19382 23348 19388
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 25884 18970 25912 20538
rect 25872 18964 25924 18970
rect 25872 18906 25924 18912
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 24492 18284 24544 18290
rect 24492 18226 24544 18232
rect 18880 18216 18932 18222
rect 3422 18184 3478 18193
rect 3422 18119 3478 18128
rect 18694 18184 18750 18193
rect 18880 18158 18932 18164
rect 18694 18119 18696 18128
rect 18748 18119 18750 18128
rect 18696 18090 18748 18096
rect 11612 17740 11664 17746
rect 11612 17682 11664 17688
rect 11336 17672 11388 17678
rect 11336 17614 11388 17620
rect 8024 17536 8076 17542
rect 8024 17478 8076 17484
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 8036 17134 8064 17478
rect 10888 17202 10916 17478
rect 11348 17338 11376 17614
rect 11336 17332 11388 17338
rect 11336 17274 11388 17280
rect 10876 17196 10928 17202
rect 10876 17138 10928 17144
rect 8024 17128 8076 17134
rect 8024 17070 8076 17076
rect 7104 16992 7156 16998
rect 7104 16934 7156 16940
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 7116 16250 7144 16934
rect 7472 16788 7524 16794
rect 7472 16730 7524 16736
rect 7104 16244 7156 16250
rect 7104 16186 7156 16192
rect 5814 15736 5870 15745
rect 5814 15671 5870 15680
rect 5264 15360 5316 15366
rect 5264 15302 5316 15308
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 5276 15026 5304 15302
rect 5828 15026 5856 15671
rect 7116 15570 7144 16186
rect 7484 16046 7512 16730
rect 8036 16726 8064 17070
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 8312 16794 8340 16934
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 8024 16720 8076 16726
rect 8024 16662 8076 16668
rect 7748 16652 7800 16658
rect 7748 16594 7800 16600
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 7472 16040 7524 16046
rect 7472 15982 7524 15988
rect 7760 15745 7788 16594
rect 7840 16448 7892 16454
rect 7840 16390 7892 16396
rect 7852 15881 7880 16390
rect 7838 15872 7894 15881
rect 7838 15807 7894 15816
rect 7746 15736 7802 15745
rect 7746 15671 7802 15680
rect 8220 15638 8248 16594
rect 8312 15706 8340 16730
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 9128 16516 9180 16522
rect 9128 16458 9180 16464
rect 8576 15904 8628 15910
rect 8576 15846 8628 15852
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 8588 15638 8616 15846
rect 9140 15706 9168 16458
rect 9680 16448 9732 16454
rect 9680 16390 9732 16396
rect 9496 15972 9548 15978
rect 9496 15914 9548 15920
rect 9508 15706 9536 15914
rect 9128 15700 9180 15706
rect 9128 15642 9180 15648
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 8208 15632 8260 15638
rect 8208 15574 8260 15580
rect 8576 15632 8628 15638
rect 8576 15574 8628 15580
rect 7104 15564 7156 15570
rect 7104 15506 7156 15512
rect 9692 15502 9720 16390
rect 10152 16017 10180 16526
rect 10138 16008 10194 16017
rect 10138 15943 10140 15952
rect 10192 15943 10194 15952
rect 10140 15914 10192 15920
rect 10046 15872 10102 15881
rect 10046 15807 10102 15816
rect 10060 15706 10088 15807
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 6368 15496 6420 15502
rect 9680 15496 9732 15502
rect 6368 15438 6420 15444
rect 9600 15444 9680 15450
rect 9600 15438 9732 15444
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 5816 15020 5868 15026
rect 5816 14962 5868 14968
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5540 14816 5592 14822
rect 5540 14758 5592 14764
rect 5724 14816 5776 14822
rect 5724 14758 5776 14764
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 5184 14113 5212 14758
rect 5552 14482 5580 14758
rect 5540 14476 5592 14482
rect 5540 14418 5592 14424
rect 5736 14414 5764 14758
rect 5724 14408 5776 14414
rect 5724 14350 5776 14356
rect 5170 14104 5226 14113
rect 5170 14039 5226 14048
rect 5172 14000 5224 14006
rect 5170 13968 5172 13977
rect 5224 13968 5226 13977
rect 5170 13903 5226 13912
rect 5736 13734 5764 14350
rect 5828 13938 5856 14962
rect 6380 14958 6408 15438
rect 9600 15422 9720 15438
rect 7748 15360 7800 15366
rect 7748 15302 7800 15308
rect 9496 15360 9548 15366
rect 9496 15302 9548 15308
rect 6368 14952 6420 14958
rect 6368 14894 6420 14900
rect 7760 14890 7788 15302
rect 7748 14884 7800 14890
rect 7748 14826 7800 14832
rect 7840 14884 7892 14890
rect 7840 14826 7892 14832
rect 6644 14816 6696 14822
rect 6644 14758 6696 14764
rect 6656 14482 6684 14758
rect 7760 14618 7788 14826
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 6644 14476 6696 14482
rect 6644 14418 6696 14424
rect 6656 14074 6684 14418
rect 6828 14272 6880 14278
rect 6828 14214 6880 14220
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 5816 13932 5868 13938
rect 5816 13874 5868 13880
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 6000 13796 6052 13802
rect 6000 13738 6052 13744
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5724 13728 5776 13734
rect 5724 13670 5776 13676
rect 5552 13530 5580 13670
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5736 13326 5764 13670
rect 6012 13462 6040 13738
rect 6000 13456 6052 13462
rect 6000 13398 6052 13404
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 5736 12646 5764 13262
rect 6012 12986 6040 13398
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 6564 10538 6592 13874
rect 6840 13802 6868 14214
rect 7378 14104 7434 14113
rect 7378 14039 7434 14048
rect 7286 13968 7342 13977
rect 7392 13938 7420 14039
rect 7286 13903 7342 13912
rect 7380 13932 7432 13938
rect 7300 13802 7328 13903
rect 7380 13874 7432 13880
rect 7748 13932 7800 13938
rect 7852 13920 7880 14826
rect 9508 14550 9536 15302
rect 9600 15162 9628 15422
rect 9588 15156 9640 15162
rect 9588 15098 9640 15104
rect 9864 15020 9916 15026
rect 9864 14962 9916 14968
rect 9876 14890 9904 14962
rect 9864 14884 9916 14890
rect 9864 14826 9916 14832
rect 9876 14550 9904 14826
rect 10060 14618 10088 15642
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 10244 15026 10272 15438
rect 10232 15020 10284 15026
rect 10232 14962 10284 14968
rect 10704 14958 10732 16934
rect 10888 16590 10916 17138
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 11164 16726 11192 16934
rect 11152 16720 11204 16726
rect 11152 16662 11204 16668
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 10876 16584 10928 16590
rect 10876 16526 10928 16532
rect 11152 16584 11204 16590
rect 11152 16526 11204 16532
rect 11164 16250 11192 16526
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11256 15706 11284 16594
rect 11348 16590 11376 17274
rect 11624 17134 11652 17682
rect 18892 17542 18920 18158
rect 20260 18080 20312 18086
rect 20260 18022 20312 18028
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 12808 17536 12860 17542
rect 12808 17478 12860 17484
rect 13268 17536 13320 17542
rect 13268 17478 13320 17484
rect 18880 17536 18932 17542
rect 18880 17478 18932 17484
rect 11888 17332 11940 17338
rect 11888 17274 11940 17280
rect 11520 17128 11572 17134
rect 11520 17070 11572 17076
rect 11612 17128 11664 17134
rect 11612 17070 11664 17076
rect 11532 16810 11560 17070
rect 11532 16794 11652 16810
rect 11532 16788 11664 16794
rect 11532 16782 11612 16788
rect 11612 16730 11664 16736
rect 11336 16584 11388 16590
rect 11336 16526 11388 16532
rect 11336 16040 11388 16046
rect 11336 15982 11388 15988
rect 11244 15700 11296 15706
rect 11244 15642 11296 15648
rect 11348 15570 11376 15982
rect 11624 15638 11652 16730
rect 11900 16046 11928 17274
rect 12820 16998 12848 17478
rect 13280 17202 13308 17478
rect 13268 17196 13320 17202
rect 13268 17138 13320 17144
rect 13544 17128 13596 17134
rect 13542 17096 13544 17105
rect 13596 17096 13598 17105
rect 13542 17031 13598 17040
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11612 15632 11664 15638
rect 11612 15574 11664 15580
rect 11336 15564 11388 15570
rect 11336 15506 11388 15512
rect 11348 15162 11376 15506
rect 11624 15162 11652 15574
rect 11336 15156 11388 15162
rect 11336 15098 11388 15104
rect 11612 15156 11664 15162
rect 11612 15098 11664 15104
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 10782 14920 10838 14929
rect 10782 14855 10838 14864
rect 10796 14822 10824 14855
rect 10232 14816 10284 14822
rect 10232 14758 10284 14764
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 8760 14544 8812 14550
rect 8760 14486 8812 14492
rect 9496 14544 9548 14550
rect 9496 14486 9548 14492
rect 9864 14544 9916 14550
rect 9864 14486 9916 14492
rect 8772 14074 8800 14486
rect 10244 14482 10272 14758
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 9232 14074 9260 14418
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9956 14272 10008 14278
rect 9956 14214 10008 14220
rect 9508 14074 9536 14214
rect 9968 14074 9996 14214
rect 8760 14068 8812 14074
rect 8760 14010 8812 14016
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 7800 13892 7880 13920
rect 7748 13874 7800 13880
rect 6828 13796 6880 13802
rect 6828 13738 6880 13744
rect 7288 13796 7340 13802
rect 7288 13738 7340 13744
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 7116 12782 7144 13466
rect 7760 13190 7788 13874
rect 9508 13870 9536 14010
rect 10324 14000 10376 14006
rect 10324 13942 10376 13948
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 10048 13728 10100 13734
rect 10048 13670 10100 13676
rect 8220 13394 8248 13670
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 6736 12640 6788 12646
rect 6736 12582 6788 12588
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6748 12306 6776 12582
rect 6736 12300 6788 12306
rect 6788 12260 6868 12288
rect 6736 12242 6788 12248
rect 6840 11694 6868 12260
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6644 11620 6696 11626
rect 6644 11562 6696 11568
rect 6656 10810 6684 11562
rect 6840 11150 6868 11630
rect 6932 11626 6960 12582
rect 7012 12368 7064 12374
rect 7012 12310 7064 12316
rect 7024 11898 7052 12310
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 6920 11280 6972 11286
rect 6920 11222 6972 11228
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6840 10554 6868 11086
rect 6932 10742 6960 11222
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 6552 10532 6604 10538
rect 6840 10526 6960 10554
rect 7024 10538 7052 11834
rect 7380 10668 7432 10674
rect 7380 10610 7432 10616
rect 6552 10474 6604 10480
rect 6564 10266 6592 10474
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6840 10266 6868 10406
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 6840 9654 6868 10066
rect 6828 9648 6880 9654
rect 6828 9590 6880 9596
rect 6932 9042 6960 10526
rect 7012 10532 7064 10538
rect 7012 10474 7064 10480
rect 7024 10062 7052 10474
rect 7392 10470 7420 10610
rect 7380 10464 7432 10470
rect 7656 10464 7708 10470
rect 7432 10424 7512 10452
rect 7380 10406 7432 10412
rect 7104 10260 7156 10266
rect 7104 10202 7156 10208
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 7116 9722 7144 10202
rect 7484 9994 7512 10424
rect 7656 10406 7708 10412
rect 7668 10266 7696 10406
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7668 10130 7696 10202
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7760 10062 7788 13126
rect 8220 12986 8248 13330
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 8208 12980 8260 12986
rect 8208 12922 8260 12928
rect 7840 12708 7892 12714
rect 7840 12650 7892 12656
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 7472 9988 7524 9994
rect 7472 9930 7524 9936
rect 7484 9722 7512 9930
rect 7852 9926 7880 12650
rect 8404 12374 8432 13126
rect 9968 12646 9996 13330
rect 10060 12986 10088 13670
rect 10336 13190 10364 13942
rect 11072 13870 11100 14418
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 10324 13184 10376 13190
rect 10324 13126 10376 13132
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 9588 12640 9640 12646
rect 9956 12640 10008 12646
rect 9640 12600 9720 12628
rect 9588 12582 9640 12588
rect 8392 12368 8444 12374
rect 8392 12310 8444 12316
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 7932 11688 7984 11694
rect 7932 11630 7984 11636
rect 7944 11218 7972 11630
rect 8036 11286 8064 12038
rect 8404 11898 8432 12310
rect 9692 12306 9720 12600
rect 9954 12608 9956 12617
rect 10008 12608 10010 12617
rect 9954 12543 10010 12552
rect 9956 12436 10008 12442
rect 9956 12378 10008 12384
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 9404 11620 9456 11626
rect 9404 11562 9456 11568
rect 9416 11354 9444 11562
rect 8760 11348 8812 11354
rect 8760 11290 8812 11296
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 8024 11280 8076 11286
rect 8024 11222 8076 11228
rect 7932 11212 7984 11218
rect 7932 11154 7984 11160
rect 7944 10810 7972 11154
rect 8036 10962 8064 11222
rect 8036 10934 8340 10962
rect 8312 10810 8340 10934
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8772 10606 8800 11290
rect 9968 11218 9996 12378
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 10060 11354 10088 12242
rect 10336 12238 10364 13126
rect 10704 12782 10732 13126
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10692 12776 10744 12782
rect 10692 12718 10744 12724
rect 10600 12436 10652 12442
rect 10704 12424 10732 12718
rect 10796 12442 10824 12786
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 10652 12396 10732 12424
rect 10784 12436 10836 12442
rect 10600 12378 10652 12384
rect 10784 12378 10836 12384
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 10704 11286 10732 11494
rect 10692 11280 10744 11286
rect 10980 11257 11008 12582
rect 10692 11222 10744 11228
rect 10966 11248 11022 11257
rect 9956 11212 10008 11218
rect 9956 11154 10008 11160
rect 9968 10810 9996 11154
rect 10704 10810 10732 11222
rect 10966 11183 11022 11192
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8772 10266 8800 10542
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 7472 9716 7524 9722
rect 7472 9658 7524 9664
rect 8312 9654 8340 9998
rect 8956 9994 8984 10610
rect 10704 10606 10732 10746
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 10704 10266 10732 10542
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 8944 9988 8996 9994
rect 8944 9930 8996 9936
rect 9680 9920 9732 9926
rect 9600 9868 9680 9874
rect 9600 9862 9732 9868
rect 9600 9846 9720 9862
rect 9600 9654 9628 9846
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 9404 9444 9456 9450
rect 9404 9386 9456 9392
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 3056 8356 3108 8362
rect 3056 8298 3108 8304
rect 3068 7750 3096 8298
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 3056 7744 3108 7750
rect 3056 7686 3108 7692
rect 3068 7342 3096 7686
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 3976 7268 4028 7274
rect 3976 7210 4028 7216
rect 2504 7200 2556 7206
rect 2504 7142 2556 7148
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2516 7002 2544 7142
rect 2504 6996 2556 7002
rect 2504 6938 2556 6944
rect 2226 6760 2282 6769
rect 2226 6695 2282 6704
rect 2240 6458 2268 6695
rect 2412 6656 2464 6662
rect 2412 6598 2464 6604
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2240 6254 2268 6394
rect 2228 6248 2280 6254
rect 2228 6190 2280 6196
rect 2240 5778 2268 6190
rect 2424 5953 2452 6598
rect 2516 6458 2544 6938
rect 2596 6860 2648 6866
rect 2596 6802 2648 6808
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2410 5944 2466 5953
rect 2410 5879 2466 5888
rect 2516 5846 2544 6394
rect 2608 6254 2636 6802
rect 2792 6769 2820 7142
rect 3988 6905 4016 7210
rect 3974 6896 4030 6905
rect 3974 6831 4030 6840
rect 3988 6798 4016 6831
rect 3976 6792 4028 6798
rect 2778 6760 2834 6769
rect 2778 6695 2834 6704
rect 3514 6760 3570 6769
rect 3976 6734 4028 6740
rect 3514 6695 3570 6704
rect 3528 6662 3556 6695
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 2504 5840 2556 5846
rect 2504 5782 2556 5788
rect 1492 5772 1544 5778
rect 1492 5714 1544 5720
rect 2228 5772 2280 5778
rect 2228 5714 2280 5720
rect 1504 5370 1532 5714
rect 3056 5636 3108 5642
rect 3056 5578 3108 5584
rect 2780 5568 2832 5574
rect 2780 5510 2832 5516
rect 1492 5364 1544 5370
rect 1492 5306 1544 5312
rect 1504 4690 1532 5306
rect 2792 5166 2820 5510
rect 3068 5234 3096 5578
rect 3252 5370 3280 6394
rect 3528 5642 3556 6598
rect 3988 6458 4016 6734
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 3988 5914 4016 6190
rect 4080 5930 4108 8230
rect 4724 7750 4752 8434
rect 6932 8430 6960 8978
rect 7208 8673 7236 8978
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 7194 8664 7250 8673
rect 7194 8599 7196 8608
rect 7248 8599 7250 8608
rect 7196 8570 7248 8576
rect 7208 8539 7236 8570
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 5000 7274 5028 7822
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 4988 7268 5040 7274
rect 4988 7210 5040 7216
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 4172 6934 4200 7142
rect 4160 6928 4212 6934
rect 4160 6870 4212 6876
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 4724 6458 4752 6802
rect 5184 6769 5212 7686
rect 5276 7546 5304 7890
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5368 6866 5396 8366
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 7288 8356 7340 8362
rect 7288 8298 7340 8304
rect 5460 7002 5488 8298
rect 6368 8288 6420 8294
rect 6368 8230 6420 8236
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6380 8090 6408 8230
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 6564 7750 6592 8230
rect 7300 7750 7328 8298
rect 7932 8288 7984 8294
rect 7932 8230 7984 8236
rect 7944 8090 7972 8230
rect 7932 8084 7984 8090
rect 7932 8026 7984 8032
rect 7380 7812 7432 7818
rect 7380 7754 7432 7760
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 6564 7342 6592 7686
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 5170 6760 5226 6769
rect 5080 6724 5132 6730
rect 5170 6695 5226 6704
rect 5080 6666 5132 6672
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 5092 6118 5120 6666
rect 5552 6662 5580 7278
rect 6564 7206 6592 7278
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 5540 6656 5592 6662
rect 5368 6616 5540 6644
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 4434 5944 4490 5953
rect 4080 5914 4200 5930
rect 3976 5908 4028 5914
rect 4080 5908 4212 5914
rect 4080 5902 4160 5908
rect 3976 5850 4028 5856
rect 4434 5879 4490 5888
rect 4620 5908 4672 5914
rect 4160 5850 4212 5856
rect 4448 5846 4476 5879
rect 4620 5850 4672 5856
rect 4436 5840 4488 5846
rect 4436 5782 4488 5788
rect 3516 5636 3568 5642
rect 3516 5578 3568 5584
rect 3332 5568 3384 5574
rect 3332 5510 3384 5516
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 2596 5160 2648 5166
rect 2596 5102 2648 5108
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2608 5030 2636 5102
rect 2412 5024 2464 5030
rect 2412 4966 2464 4972
rect 2596 5024 2648 5030
rect 2596 4966 2648 4972
rect 2688 5024 2740 5030
rect 2688 4966 2740 4972
rect 1492 4684 1544 4690
rect 1492 4626 1544 4632
rect 1504 4078 1532 4626
rect 1492 4072 1544 4078
rect 1492 4014 1544 4020
rect 1504 3602 1532 4014
rect 2424 3738 2452 4966
rect 2608 4078 2636 4966
rect 2596 4072 2648 4078
rect 2596 4014 2648 4020
rect 2412 3732 2464 3738
rect 2412 3674 2464 3680
rect 1492 3596 1544 3602
rect 1492 3538 1544 3544
rect 1504 3194 1532 3538
rect 2410 3496 2466 3505
rect 2410 3431 2466 3440
rect 1492 3188 1544 3194
rect 1492 3130 1544 3136
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 1676 2848 1728 2854
rect 570 2816 626 2825
rect 1676 2790 1728 2796
rect 570 2751 626 2760
rect 584 480 612 2751
rect 1688 480 1716 2790
rect 1780 2650 1808 2994
rect 2424 2650 2452 3431
rect 2700 2854 2728 4966
rect 3068 4486 3096 5170
rect 3344 5098 3372 5510
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 4632 5370 4660 5850
rect 5092 5574 5120 6054
rect 5080 5568 5132 5574
rect 5080 5510 5132 5516
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4342 5128 4398 5137
rect 3332 5092 3384 5098
rect 4342 5063 4344 5072
rect 3332 5034 3384 5040
rect 4396 5063 4398 5072
rect 4344 5034 4396 5040
rect 3344 4826 3372 5034
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 2792 3670 2820 4422
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2780 3664 2832 3670
rect 2780 3606 2832 3612
rect 2688 2848 2740 2854
rect 2688 2790 2740 2796
rect 2792 2650 2820 3606
rect 1768 2644 1820 2650
rect 1768 2586 1820 2592
rect 2412 2644 2464 2650
rect 2412 2586 2464 2592
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 2884 2530 2912 4082
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 2976 2922 3004 3334
rect 2964 2916 3016 2922
rect 2964 2858 3016 2864
rect 2976 2582 3004 2858
rect 2792 2502 2912 2530
rect 2964 2576 3016 2582
rect 2964 2518 3016 2524
rect 2792 480 2820 2502
rect 3068 2446 3096 4422
rect 3344 4282 3372 4762
rect 3974 4720 4030 4729
rect 3974 4655 4030 4664
rect 3882 4584 3938 4593
rect 3882 4519 3938 4528
rect 3332 4276 3384 4282
rect 3332 4218 3384 4224
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3804 3058 3832 3878
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 3700 2848 3752 2854
rect 3700 2790 3752 2796
rect 3712 2650 3740 2790
rect 3700 2644 3752 2650
rect 3700 2586 3752 2592
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 3896 480 3924 4519
rect 3988 3466 4016 4655
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 4632 4214 4660 4966
rect 4804 4752 4856 4758
rect 4804 4694 4856 4700
rect 4620 4208 4672 4214
rect 4620 4150 4672 4156
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 3976 3460 4028 3466
rect 3976 3402 4028 3408
rect 4080 2825 4108 3878
rect 4436 3596 4488 3602
rect 4436 3538 4488 3544
rect 4448 3505 4476 3538
rect 4434 3496 4490 3505
rect 4434 3431 4490 3440
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 4160 3120 4212 3126
rect 4632 3097 4660 3878
rect 4724 3534 4752 4014
rect 4816 3942 4844 4694
rect 4986 4176 5042 4185
rect 4986 4111 5042 4120
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4712 3528 4764 3534
rect 4712 3470 4764 3476
rect 4160 3062 4212 3068
rect 4618 3088 4674 3097
rect 4172 2990 4200 3062
rect 4618 3023 4674 3032
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 4066 2816 4122 2825
rect 4066 2751 4122 2760
rect 4172 2666 4200 2926
rect 4816 2922 4844 3878
rect 4804 2916 4856 2922
rect 4804 2858 4856 2864
rect 4080 2638 4200 2666
rect 4080 2446 4108 2638
rect 4816 2514 4844 2858
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 5000 480 5028 4111
rect 5092 4078 5120 5510
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5080 4072 5132 4078
rect 5080 4014 5132 4020
rect 5184 3398 5212 4626
rect 5368 4010 5396 6616
rect 5540 6598 5592 6604
rect 5630 6216 5686 6225
rect 5630 6151 5686 6160
rect 5448 6112 5500 6118
rect 5446 6080 5448 6089
rect 5500 6080 5502 6089
rect 5446 6015 5502 6024
rect 5540 5840 5592 5846
rect 5540 5782 5592 5788
rect 5552 5370 5580 5782
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5446 5264 5502 5273
rect 5446 5199 5448 5208
rect 5500 5199 5502 5208
rect 5448 5170 5500 5176
rect 5644 4729 5672 6151
rect 5828 4826 5856 7142
rect 6564 6798 6592 7142
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6552 6792 6604 6798
rect 5998 6760 6054 6769
rect 6552 6734 6604 6740
rect 5998 6695 6054 6704
rect 6368 6724 6420 6730
rect 6012 5914 6040 6695
rect 6368 6666 6420 6672
rect 6380 6322 6408 6666
rect 6564 6390 6592 6734
rect 6552 6384 6604 6390
rect 6552 6326 6604 6332
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6656 6186 6684 6802
rect 7300 6662 7328 7686
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7300 6202 7328 6598
rect 6644 6180 6696 6186
rect 6644 6122 6696 6128
rect 7208 6174 7328 6202
rect 6000 5908 6052 5914
rect 6000 5850 6052 5856
rect 6012 5642 6040 5850
rect 6656 5710 6684 6122
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6840 5953 6868 6054
rect 6826 5944 6882 5953
rect 6826 5879 6882 5888
rect 7208 5778 7236 6174
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7300 5914 7328 6054
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 6644 5704 6696 5710
rect 6932 5658 6960 5714
rect 7392 5710 7420 7754
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7484 6254 7512 7686
rect 7944 7546 7972 8026
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 7944 7274 7972 7482
rect 7932 7268 7984 7274
rect 7932 7210 7984 7216
rect 8220 7206 8248 7890
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 8220 6458 8248 7142
rect 8312 6866 8340 8774
rect 8300 6860 8352 6866
rect 8300 6802 8352 6808
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7484 5846 7512 6190
rect 7562 6080 7618 6089
rect 7562 6015 7618 6024
rect 7576 5914 7604 6015
rect 8312 5914 8340 6258
rect 8404 6254 8432 6598
rect 8392 6248 8444 6254
rect 8390 6216 8392 6225
rect 8444 6216 8446 6225
rect 8390 6151 8446 6160
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 7472 5840 7524 5846
rect 7472 5782 7524 5788
rect 7380 5704 7432 5710
rect 6644 5646 6696 5652
rect 6000 5636 6052 5642
rect 6000 5578 6052 5584
rect 6656 5302 6684 5646
rect 6748 5630 6960 5658
rect 7286 5672 7342 5681
rect 6748 5370 6776 5630
rect 7380 5646 7432 5652
rect 7286 5607 7342 5616
rect 6826 5400 6882 5409
rect 6736 5364 6788 5370
rect 6826 5335 6882 5344
rect 6736 5306 6788 5312
rect 6644 5296 6696 5302
rect 6644 5238 6696 5244
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 5630 4720 5686 4729
rect 5630 4655 5686 4664
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 5998 4584 6054 4593
rect 5998 4519 6000 4528
rect 6052 4519 6054 4528
rect 6000 4490 6052 4496
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5552 4146 5580 4422
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5356 4004 5408 4010
rect 5356 3946 5408 3952
rect 5540 3936 5592 3942
rect 5644 3890 5672 4422
rect 6196 4321 6224 4626
rect 6182 4312 6238 4321
rect 6182 4247 6184 4256
rect 6236 4247 6238 4256
rect 6184 4218 6236 4224
rect 6748 4214 6776 4762
rect 6840 4690 6868 5335
rect 7300 5234 7328 5607
rect 7472 5568 7524 5574
rect 7472 5510 7524 5516
rect 7484 5234 7512 5510
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7300 4826 7328 5170
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 6736 4208 6788 4214
rect 6736 4150 6788 4156
rect 6840 4162 6868 4626
rect 6840 4134 6960 4162
rect 6932 4010 6960 4134
rect 7024 4026 7052 4626
rect 7484 4570 7512 5170
rect 7576 5166 7604 5850
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 7564 5160 7616 5166
rect 7564 5102 7616 5108
rect 8022 5128 8078 5137
rect 8022 5063 8078 5072
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 7944 4758 7972 4966
rect 8036 4826 8064 5063
rect 8128 5030 8156 5714
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8116 5024 8168 5030
rect 8116 4966 8168 4972
rect 8128 4865 8156 4966
rect 8114 4856 8170 4865
rect 8024 4820 8076 4826
rect 8114 4791 8170 4800
rect 8024 4762 8076 4768
rect 7932 4752 7984 4758
rect 7932 4694 7984 4700
rect 7484 4542 7604 4570
rect 7576 4486 7604 4542
rect 7104 4480 7156 4486
rect 7104 4422 7156 4428
rect 7564 4480 7616 4486
rect 7564 4422 7616 4428
rect 7116 4185 7144 4422
rect 7576 4214 7604 4422
rect 7564 4208 7616 4214
rect 7102 4176 7158 4185
rect 7564 4150 7616 4156
rect 7102 4111 7158 4120
rect 7104 4072 7156 4078
rect 7024 4020 7104 4026
rect 7024 4014 7156 4020
rect 6920 4004 6972 4010
rect 7024 3998 7144 4014
rect 6920 3946 6972 3952
rect 6828 3936 6880 3942
rect 5592 3884 5672 3890
rect 5540 3878 5672 3884
rect 5552 3862 5672 3878
rect 6826 3904 6828 3913
rect 6880 3904 6882 3913
rect 5552 3505 5580 3862
rect 6826 3839 6882 3848
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 5538 3496 5594 3505
rect 5538 3431 5594 3440
rect 5172 3392 5224 3398
rect 5172 3334 5224 3340
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5460 2990 5488 3334
rect 5644 3194 5672 3538
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 6012 3126 6040 3470
rect 6000 3120 6052 3126
rect 6000 3062 6052 3068
rect 6840 3074 6868 3538
rect 7010 3496 7066 3505
rect 7010 3431 7066 3440
rect 6840 3046 6960 3074
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5460 2650 5488 2926
rect 6090 2816 6146 2825
rect 6090 2751 6146 2760
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 6104 480 6132 2751
rect 6932 2514 6960 3046
rect 7024 2650 7052 3431
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 7116 1873 7144 3998
rect 8220 3670 8248 5646
rect 8588 5409 8616 6054
rect 8574 5400 8630 5409
rect 8574 5335 8630 5344
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 9036 5024 9088 5030
rect 9036 4966 9088 4972
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 8300 4004 8352 4010
rect 8300 3946 8352 3952
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 7208 2990 7236 3334
rect 7196 2984 7248 2990
rect 7196 2926 7248 2932
rect 7208 2650 7236 2926
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 8220 2446 8248 3606
rect 8312 3194 8340 3946
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8312 2650 8340 3130
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8404 2530 8432 4966
rect 8482 4720 8538 4729
rect 8482 4655 8484 4664
rect 8536 4655 8538 4664
rect 8484 4626 8536 4632
rect 8484 4548 8536 4554
rect 8484 4490 8536 4496
rect 8496 3913 8524 4490
rect 8482 3904 8538 3913
rect 8482 3839 8538 3848
rect 8496 3738 8524 3839
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8944 3596 8996 3602
rect 8944 3538 8996 3544
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8680 2825 8708 3334
rect 8956 2990 8984 3538
rect 9048 3097 9076 4966
rect 9128 4480 9180 4486
rect 9126 4448 9128 4457
rect 9180 4448 9182 4457
rect 9126 4383 9182 4392
rect 9034 3088 9090 3097
rect 9034 3023 9090 3032
rect 8944 2984 8996 2990
rect 8942 2952 8944 2961
rect 8996 2952 8998 2961
rect 8942 2887 8998 2896
rect 8666 2816 8722 2825
rect 8666 2751 8722 2760
rect 9324 2650 9352 4966
rect 9312 2644 9364 2650
rect 9312 2586 9364 2592
rect 8312 2502 8432 2530
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 7102 1864 7158 1873
rect 7102 1799 7158 1808
rect 7194 1456 7250 1465
rect 7194 1391 7250 1400
rect 7208 480 7236 1391
rect 8312 480 8340 2502
rect 9220 2440 9272 2446
rect 9218 2408 9220 2417
rect 9272 2408 9274 2417
rect 9218 2343 9274 2352
rect 9416 480 9444 9386
rect 10428 9382 10456 10066
rect 10784 10056 10836 10062
rect 10784 9998 10836 10004
rect 10796 9722 10824 9998
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 9956 8356 10008 8362
rect 9956 8298 10008 8304
rect 9968 8090 9996 8298
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 10060 6866 10088 7482
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10060 6458 10088 6802
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9678 5944 9734 5953
rect 9678 5879 9734 5888
rect 9692 5778 9720 5879
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9692 5370 9720 5714
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9508 4826 9536 4966
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9508 4622 9536 4762
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 9588 4072 9640 4078
rect 9494 4040 9550 4049
rect 9588 4014 9640 4020
rect 9494 3975 9550 3984
rect 9508 3738 9536 3975
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 9496 3596 9548 3602
rect 9600 3584 9628 4014
rect 9678 3768 9734 3777
rect 9678 3703 9680 3712
rect 9732 3703 9734 3712
rect 9680 3674 9732 3680
rect 9548 3556 9628 3584
rect 9496 3538 9548 3544
rect 9508 2990 9536 3538
rect 9784 3233 9812 6054
rect 9862 5672 9918 5681
rect 9862 5607 9864 5616
rect 9916 5607 9918 5616
rect 9864 5578 9916 5584
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 9968 3942 9996 4558
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 9968 3670 9996 3878
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 9770 3224 9826 3233
rect 9770 3159 9826 3168
rect 9968 2990 9996 3606
rect 9496 2984 9548 2990
rect 9496 2926 9548 2932
rect 9956 2984 10008 2990
rect 9956 2926 10008 2932
rect 10152 2582 10180 8910
rect 10428 6202 10456 9318
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10520 7886 10548 8366
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10520 7546 10548 7822
rect 10888 7546 10916 9386
rect 10980 8265 11008 11018
rect 11072 10810 11100 13806
rect 11256 12850 11284 14214
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 11150 12608 11206 12617
rect 11150 12543 11206 12552
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 11164 10690 11192 12543
rect 11348 12238 11376 15098
rect 12452 14929 12480 16934
rect 12532 16720 12584 16726
rect 12532 16662 12584 16668
rect 12544 16046 12572 16662
rect 12820 16658 12848 16934
rect 12808 16652 12860 16658
rect 12808 16594 12860 16600
rect 12532 16040 12584 16046
rect 12532 15982 12584 15988
rect 13818 16008 13874 16017
rect 12544 15706 12572 15982
rect 13818 15943 13874 15952
rect 13832 15910 13860 15943
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 18892 15162 18920 17478
rect 20272 17066 20300 18022
rect 22652 17740 22704 17746
rect 22652 17682 22704 17688
rect 23112 17740 23164 17746
rect 23112 17682 23164 17688
rect 21456 17672 21508 17678
rect 21456 17614 21508 17620
rect 21468 17134 21496 17614
rect 22664 17338 22692 17682
rect 23124 17338 23152 17682
rect 23756 17536 23808 17542
rect 23756 17478 23808 17484
rect 24308 17536 24360 17542
rect 24504 17524 24532 18226
rect 25884 18222 25912 18906
rect 25872 18216 25924 18222
rect 25872 18158 25924 18164
rect 24360 17496 24532 17524
rect 24308 17478 24360 17484
rect 22652 17332 22704 17338
rect 22652 17274 22704 17280
rect 23112 17332 23164 17338
rect 23112 17274 23164 17280
rect 21456 17128 21508 17134
rect 21456 17070 21508 17076
rect 20260 17060 20312 17066
rect 20260 17002 20312 17008
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 21468 16454 21496 17070
rect 22192 17060 22244 17066
rect 22192 17002 22244 17008
rect 22100 16992 22152 16998
rect 22100 16934 22152 16940
rect 22112 16726 22140 16934
rect 22100 16720 22152 16726
rect 22100 16662 22152 16668
rect 21456 16448 21508 16454
rect 21456 16390 21508 16396
rect 21468 15910 21496 16390
rect 22112 16046 22140 16662
rect 22204 16114 22232 17002
rect 22664 16794 22692 17274
rect 23768 17134 23796 17478
rect 23756 17128 23808 17134
rect 23756 17070 23808 17076
rect 22652 16788 22704 16794
rect 22652 16730 22704 16736
rect 23480 16788 23532 16794
rect 23480 16730 23532 16736
rect 22834 16552 22890 16561
rect 22834 16487 22890 16496
rect 22192 16108 22244 16114
rect 22192 16050 22244 16056
rect 22100 16040 22152 16046
rect 22100 15982 22152 15988
rect 20904 15904 20956 15910
rect 20904 15846 20956 15852
rect 21456 15904 21508 15910
rect 21456 15846 21508 15852
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 19248 15360 19300 15366
rect 19248 15302 19300 15308
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 12438 14920 12494 14929
rect 12438 14855 12494 14864
rect 16948 14544 17000 14550
rect 16948 14486 17000 14492
rect 16580 14340 16632 14346
rect 16580 14282 16632 14288
rect 15752 14272 15804 14278
rect 15752 14214 15804 14220
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 15764 13870 15792 14214
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15200 13728 15252 13734
rect 15200 13670 15252 13676
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 12348 13388 12400 13394
rect 12348 13330 12400 13336
rect 11716 12986 11744 13330
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11992 12306 12020 13262
rect 12256 13184 12308 13190
rect 12256 13126 12308 13132
rect 11980 12300 12032 12306
rect 11980 12242 12032 12248
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11256 11898 11284 12174
rect 11900 11898 11928 12174
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11900 11218 11928 11834
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 11900 10810 11928 11154
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11072 10662 11192 10690
rect 10966 8256 11022 8265
rect 10966 8191 11022 8200
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10598 6352 10654 6361
rect 10704 6322 10732 6802
rect 10782 6488 10838 6497
rect 10782 6423 10838 6432
rect 10598 6287 10600 6296
rect 10652 6287 10654 6296
rect 10692 6316 10744 6322
rect 10600 6258 10652 6264
rect 10692 6258 10744 6264
rect 10428 6174 10548 6202
rect 10232 4820 10284 4826
rect 10232 4762 10284 4768
rect 10244 3738 10272 4762
rect 10324 4480 10376 4486
rect 10324 4422 10376 4428
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 10230 3224 10286 3233
rect 10230 3159 10286 3168
rect 10140 2576 10192 2582
rect 10140 2518 10192 2524
rect 10244 2145 10272 3159
rect 10336 2922 10364 4422
rect 10324 2916 10376 2922
rect 10324 2858 10376 2864
rect 10336 2650 10364 2858
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 10230 2136 10286 2145
rect 10230 2071 10286 2080
rect 10520 480 10548 6174
rect 10612 5914 10640 6258
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10704 5846 10732 6258
rect 10796 6254 10824 6423
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10692 5840 10744 5846
rect 10692 5782 10744 5788
rect 10600 5160 10652 5166
rect 10598 5128 10600 5137
rect 10652 5128 10654 5137
rect 10598 5063 10654 5072
rect 10874 5128 10930 5137
rect 10874 5063 10876 5072
rect 10928 5063 10930 5072
rect 10876 5034 10928 5040
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 10796 4826 10824 4966
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10612 3942 10640 4626
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10612 3641 10640 3878
rect 10598 3632 10654 3641
rect 10598 3567 10654 3576
rect 10784 3596 10836 3602
rect 10784 3538 10836 3544
rect 10796 3194 10824 3538
rect 10980 3398 11008 6054
rect 11072 3482 11100 10662
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11348 10169 11376 10406
rect 11334 10160 11390 10169
rect 11334 10095 11390 10104
rect 11428 9580 11480 9586
rect 11428 9522 11480 9528
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11256 9178 11284 9318
rect 11244 9172 11296 9178
rect 11244 9114 11296 9120
rect 11440 8838 11468 9522
rect 11716 9042 11744 10746
rect 12268 10690 12296 13126
rect 12360 12646 12388 13330
rect 15212 13326 15240 13670
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 14464 13184 14516 13190
rect 14464 13126 14516 13132
rect 14476 12850 14504 13126
rect 14464 12844 14516 12850
rect 14464 12786 14516 12792
rect 15212 12782 15240 13262
rect 15568 13184 15620 13190
rect 15568 13126 15620 13132
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15212 12646 15240 12718
rect 15580 12714 15608 13126
rect 15568 12708 15620 12714
rect 15568 12650 15620 12656
rect 12348 12640 12400 12646
rect 13912 12640 13964 12646
rect 12400 12600 12572 12628
rect 12348 12582 12400 12588
rect 12440 12300 12492 12306
rect 12440 12242 12492 12248
rect 12452 11354 12480 12242
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12544 11082 12572 12600
rect 14280 12640 14332 12646
rect 13912 12582 13964 12588
rect 14278 12608 14280 12617
rect 15200 12640 15252 12646
rect 14332 12608 14334 12617
rect 13924 12481 13952 12582
rect 15764 12617 15792 13806
rect 16304 13252 16356 13258
rect 16304 13194 16356 13200
rect 15200 12582 15252 12588
rect 15750 12608 15806 12617
rect 14278 12543 14334 12552
rect 13910 12472 13966 12481
rect 14292 12442 14320 12543
rect 13910 12407 13966 12416
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 14832 12300 14884 12306
rect 14832 12242 14884 12248
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 13280 11626 13308 12038
rect 14844 11898 14872 12242
rect 15212 12238 15240 12582
rect 15750 12543 15806 12552
rect 16212 12300 16264 12306
rect 16212 12242 16264 12248
rect 15200 12232 15252 12238
rect 15200 12174 15252 12180
rect 14832 11892 14884 11898
rect 14832 11834 14884 11840
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 13268 11620 13320 11626
rect 13268 11562 13320 11568
rect 13280 11354 13308 11562
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 12532 11076 12584 11082
rect 12532 11018 12584 11024
rect 12268 10674 12480 10690
rect 13280 10674 13308 11290
rect 13542 11248 13598 11257
rect 13542 11183 13544 11192
rect 13596 11183 13598 11192
rect 13544 11154 13596 11160
rect 13556 10810 13584 11154
rect 13544 10804 13596 10810
rect 13544 10746 13596 10752
rect 13832 10690 13860 11630
rect 15212 11558 15240 12174
rect 16224 11694 16252 12242
rect 16316 11830 16344 13194
rect 16408 12322 16436 14214
rect 16592 13258 16620 14282
rect 16960 13734 16988 14486
rect 17972 14414 18000 14962
rect 19260 14958 19288 15302
rect 19248 14952 19300 14958
rect 19248 14894 19300 14900
rect 19260 14618 19288 14894
rect 20536 14816 20588 14822
rect 20536 14758 20588 14764
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 19248 14612 19300 14618
rect 19248 14554 19300 14560
rect 18052 14476 18104 14482
rect 18052 14418 18104 14424
rect 17960 14408 18012 14414
rect 17960 14350 18012 14356
rect 17972 14074 18000 14350
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 17972 13818 18000 14010
rect 18064 13870 18092 14418
rect 18972 14272 19024 14278
rect 18972 14214 19024 14220
rect 18984 13938 19012 14214
rect 18972 13932 19024 13938
rect 18972 13874 19024 13880
rect 19064 13932 19116 13938
rect 19064 13874 19116 13880
rect 17880 13790 18000 13818
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 18604 13864 18656 13870
rect 18604 13806 18656 13812
rect 16948 13728 17000 13734
rect 16948 13670 17000 13676
rect 16960 13394 16988 13670
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 17776 13388 17828 13394
rect 17776 13330 17828 13336
rect 16580 13252 16632 13258
rect 16580 13194 16632 13200
rect 17788 12986 17816 13330
rect 17880 13190 17908 13790
rect 18064 13530 18092 13806
rect 18144 13728 18196 13734
rect 18144 13670 18196 13676
rect 18052 13524 18104 13530
rect 18052 13466 18104 13472
rect 17868 13184 17920 13190
rect 17868 13126 17920 13132
rect 17776 12980 17828 12986
rect 17776 12922 17828 12928
rect 17880 12918 17908 13126
rect 18156 12986 18184 13670
rect 18616 13530 18644 13806
rect 18604 13524 18656 13530
rect 18604 13466 18656 13472
rect 18984 13326 19012 13874
rect 19076 13802 19104 13874
rect 19260 13870 19288 14554
rect 20548 13870 20576 14758
rect 19248 13864 19300 13870
rect 19248 13806 19300 13812
rect 20536 13864 20588 13870
rect 20536 13806 20588 13812
rect 19064 13796 19116 13802
rect 19064 13738 19116 13744
rect 19076 13530 19104 13738
rect 20916 13734 20944 15846
rect 22112 15706 22140 15982
rect 22100 15700 22152 15706
rect 22100 15642 22152 15648
rect 22204 15570 22232 16050
rect 22744 15904 22796 15910
rect 22744 15846 22796 15852
rect 22756 15706 22784 15846
rect 22744 15700 22796 15706
rect 22744 15642 22796 15648
rect 22192 15564 22244 15570
rect 22192 15506 22244 15512
rect 22756 15162 22784 15642
rect 22848 15434 22876 16487
rect 23492 15722 23520 16730
rect 23768 16726 23796 17070
rect 24504 17066 24532 17496
rect 25320 17536 25372 17542
rect 25320 17478 25372 17484
rect 24584 17332 24636 17338
rect 24584 17274 24636 17280
rect 24492 17060 24544 17066
rect 24492 17002 24544 17008
rect 23664 16720 23716 16726
rect 23664 16662 23716 16668
rect 23756 16720 23808 16726
rect 23756 16662 23808 16668
rect 24308 16720 24360 16726
rect 24308 16662 24360 16668
rect 23676 16250 23704 16662
rect 24216 16584 24268 16590
rect 24216 16526 24268 16532
rect 23664 16244 23716 16250
rect 23664 16186 23716 16192
rect 24228 16114 24256 16526
rect 24216 16108 24268 16114
rect 24216 16050 24268 16056
rect 23400 15694 23520 15722
rect 23400 15638 23428 15694
rect 23388 15632 23440 15638
rect 23388 15574 23440 15580
rect 22928 15496 22980 15502
rect 22928 15438 22980 15444
rect 22836 15428 22888 15434
rect 22836 15370 22888 15376
rect 22940 15201 22968 15438
rect 22926 15192 22982 15201
rect 22744 15156 22796 15162
rect 22926 15127 22982 15136
rect 22744 15098 22796 15104
rect 22940 14618 22968 15127
rect 23400 15094 23428 15574
rect 23480 15564 23532 15570
rect 23480 15506 23532 15512
rect 23492 15162 23520 15506
rect 24228 15502 24256 16050
rect 24320 15706 24348 16662
rect 24504 16522 24532 17002
rect 24492 16516 24544 16522
rect 24492 16458 24544 16464
rect 24504 16046 24532 16458
rect 24492 16040 24544 16046
rect 24492 15982 24544 15988
rect 24308 15700 24360 15706
rect 24308 15642 24360 15648
rect 24216 15496 24268 15502
rect 24504 15450 24532 15982
rect 24596 15706 24624 17274
rect 25332 16658 25360 17478
rect 24860 16652 24912 16658
rect 24860 16594 24912 16600
rect 25320 16652 25372 16658
rect 25320 16594 25372 16600
rect 24872 16402 24900 16594
rect 24688 16374 24900 16402
rect 24688 15978 24716 16374
rect 24768 16244 24820 16250
rect 24768 16186 24820 16192
rect 24676 15972 24728 15978
rect 24676 15914 24728 15920
rect 24584 15700 24636 15706
rect 24584 15642 24636 15648
rect 24216 15438 24268 15444
rect 24320 15422 24532 15450
rect 23480 15156 23532 15162
rect 23480 15098 23532 15104
rect 24320 15094 24348 15422
rect 24400 15360 24452 15366
rect 24398 15328 24400 15337
rect 24452 15328 24454 15337
rect 24398 15263 24454 15272
rect 24596 15178 24624 15642
rect 24688 15570 24716 15914
rect 24676 15564 24728 15570
rect 24676 15506 24728 15512
rect 24780 15434 24808 16186
rect 25964 15496 26016 15502
rect 25964 15438 26016 15444
rect 24768 15428 24820 15434
rect 24768 15370 24820 15376
rect 24504 15162 24624 15178
rect 24492 15156 24624 15162
rect 24544 15150 24624 15156
rect 24492 15098 24544 15104
rect 23388 15088 23440 15094
rect 23388 15030 23440 15036
rect 24308 15088 24360 15094
rect 24308 15030 24360 15036
rect 24320 14618 24348 15030
rect 24780 14958 24808 15370
rect 24768 14952 24820 14958
rect 24768 14894 24820 14900
rect 25872 14816 25924 14822
rect 25872 14758 25924 14764
rect 22928 14612 22980 14618
rect 22928 14554 22980 14560
rect 24308 14612 24360 14618
rect 24308 14554 24360 14560
rect 23572 14476 23624 14482
rect 23572 14418 23624 14424
rect 23584 13870 23612 14418
rect 23572 13864 23624 13870
rect 24320 13818 24348 14554
rect 25412 14272 25464 14278
rect 25412 14214 25464 14220
rect 23572 13806 23624 13812
rect 20904 13728 20956 13734
rect 20904 13670 20956 13676
rect 21088 13728 21140 13734
rect 21088 13670 21140 13676
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 19064 13524 19116 13530
rect 19064 13466 19116 13472
rect 20076 13456 20128 13462
rect 20076 13398 20128 13404
rect 18972 13320 19024 13326
rect 18972 13262 19024 13268
rect 19892 13320 19944 13326
rect 19892 13262 19944 13268
rect 19248 13184 19300 13190
rect 19248 13126 19300 13132
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 17868 12912 17920 12918
rect 17868 12854 17920 12860
rect 19260 12782 19288 13126
rect 19524 12844 19576 12850
rect 19524 12786 19576 12792
rect 19248 12776 19300 12782
rect 19248 12718 19300 12724
rect 16488 12708 16540 12714
rect 16540 12668 16620 12696
rect 16488 12650 16540 12656
rect 16592 12442 16620 12668
rect 16856 12640 16908 12646
rect 16854 12608 16856 12617
rect 18972 12640 19024 12646
rect 16908 12608 16910 12617
rect 18972 12582 19024 12588
rect 16854 12543 16910 12552
rect 18326 12472 18382 12481
rect 16580 12436 16632 12442
rect 18326 12407 18328 12416
rect 16580 12378 16632 12384
rect 18380 12407 18382 12416
rect 18328 12378 18380 12384
rect 16408 12294 16620 12322
rect 16592 11898 16620 12294
rect 18236 12300 18288 12306
rect 18236 12242 18288 12248
rect 18144 12232 18196 12238
rect 18144 12174 18196 12180
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 16580 11892 16632 11898
rect 16580 11834 16632 11840
rect 16304 11824 16356 11830
rect 16304 11766 16356 11772
rect 16672 11756 16724 11762
rect 16672 11698 16724 11704
rect 16212 11688 16264 11694
rect 16212 11630 16264 11636
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 15936 11552 15988 11558
rect 15936 11494 15988 11500
rect 12268 10668 12492 10674
rect 12268 10662 12440 10668
rect 12440 10610 12492 10616
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 13740 10662 13860 10690
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 11888 10192 11940 10198
rect 11888 10134 11940 10140
rect 11900 9382 11928 10134
rect 12164 10056 12216 10062
rect 12164 9998 12216 10004
rect 12176 9382 12204 9998
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 12360 9738 12388 9862
rect 12360 9710 12480 9738
rect 12256 9512 12308 9518
rect 12256 9454 12308 9460
rect 11888 9376 11940 9382
rect 11886 9344 11888 9353
rect 12164 9376 12216 9382
rect 11940 9344 11942 9353
rect 12164 9318 12216 9324
rect 11886 9279 11942 9288
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11428 8832 11480 8838
rect 11428 8774 11480 8780
rect 11242 8664 11298 8673
rect 11242 8599 11244 8608
rect 11296 8599 11298 8608
rect 11244 8570 11296 8576
rect 11440 8362 11468 8774
rect 11716 8430 11744 8978
rect 12176 8634 12204 9318
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12268 8566 12296 9454
rect 12452 9178 12480 9710
rect 12544 9450 12572 10406
rect 13004 10198 13032 10610
rect 13280 10266 13308 10610
rect 13740 10606 13768 10662
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 12992 10192 13044 10198
rect 12992 10134 13044 10140
rect 13266 10160 13322 10169
rect 13266 10095 13322 10104
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 12912 9586 12940 9862
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 12532 9444 12584 9450
rect 12532 9386 12584 9392
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 12636 8634 12664 9522
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12256 8560 12308 8566
rect 12254 8528 12256 8537
rect 12308 8528 12310 8537
rect 12254 8463 12310 8472
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 11428 8356 11480 8362
rect 11428 8298 11480 8304
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 11164 6934 11192 7142
rect 11440 7002 11468 8298
rect 11716 7478 11744 8366
rect 11794 8256 11850 8265
rect 11794 8191 11850 8200
rect 11704 7472 11756 7478
rect 11704 7414 11756 7420
rect 11428 6996 11480 7002
rect 11428 6938 11480 6944
rect 11152 6928 11204 6934
rect 11152 6870 11204 6876
rect 11808 6866 11836 8191
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 12176 7546 12204 7890
rect 12348 7744 12400 7750
rect 12400 7704 12480 7732
rect 12348 7686 12400 7692
rect 12164 7540 12216 7546
rect 12164 7482 12216 7488
rect 11980 7472 12032 7478
rect 11980 7414 12032 7420
rect 11992 6934 12020 7414
rect 12348 7336 12400 7342
rect 12452 7324 12480 7704
rect 12400 7296 12480 7324
rect 12348 7278 12400 7284
rect 11980 6928 12032 6934
rect 11980 6870 12032 6876
rect 11796 6860 11848 6866
rect 11796 6802 11848 6808
rect 11808 6458 11836 6802
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11716 5914 11744 6258
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11520 5840 11572 5846
rect 11520 5782 11572 5788
rect 11532 4826 11560 5782
rect 11612 5568 11664 5574
rect 11612 5510 11664 5516
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11624 4321 11652 5510
rect 11716 4758 11744 5850
rect 11796 5772 11848 5778
rect 11796 5714 11848 5720
rect 11808 5370 11836 5714
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11704 4752 11756 4758
rect 11704 4694 11756 4700
rect 11992 4690 12020 6870
rect 12452 6798 12480 7296
rect 12636 7274 12664 8570
rect 12728 8022 12756 9318
rect 13096 9110 13124 9522
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 13084 9104 13136 9110
rect 13084 9046 13136 9052
rect 13188 8498 13216 9114
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 12808 8424 12860 8430
rect 12808 8366 12860 8372
rect 12820 8090 12848 8366
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 12716 8016 12768 8022
rect 12716 7958 12768 7964
rect 12820 7546 12848 8026
rect 12912 7818 12940 8434
rect 12900 7812 12952 7818
rect 12900 7754 12952 7760
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 12624 7268 12676 7274
rect 12624 7210 12676 7216
rect 12636 7002 12664 7210
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12820 6882 12848 7482
rect 12912 7342 12940 7754
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12728 6854 12848 6882
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 12072 6656 12124 6662
rect 12072 6598 12124 6604
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12084 6186 12112 6598
rect 12544 6361 12572 6598
rect 12530 6352 12586 6361
rect 12530 6287 12586 6296
rect 12072 6180 12124 6186
rect 12072 6122 12124 6128
rect 12176 6174 12572 6202
rect 12176 6118 12204 6174
rect 12544 6118 12572 6174
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12452 5846 12480 6054
rect 12440 5840 12492 5846
rect 12440 5782 12492 5788
rect 12348 5704 12400 5710
rect 12348 5646 12400 5652
rect 12072 4752 12124 4758
rect 12072 4694 12124 4700
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 11610 4312 11666 4321
rect 11992 4282 12020 4626
rect 11610 4247 11666 4256
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 11242 4040 11298 4049
rect 11992 4010 12020 4218
rect 11242 3975 11298 3984
rect 11980 4004 12032 4010
rect 11256 3942 11284 3975
rect 11980 3946 12032 3952
rect 11244 3936 11296 3942
rect 11704 3936 11756 3942
rect 11244 3878 11296 3884
rect 11702 3904 11704 3913
rect 11756 3904 11758 3913
rect 11702 3839 11758 3848
rect 11992 3670 12020 3946
rect 12084 3738 12112 4694
rect 12360 4486 12388 5646
rect 12728 5030 12756 6854
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12820 5914 12848 6734
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12912 5166 12940 7278
rect 13004 5409 13032 7686
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 13188 6254 13216 6938
rect 13176 6248 13228 6254
rect 13176 6190 13228 6196
rect 13188 5914 13216 6190
rect 13176 5908 13228 5914
rect 13176 5850 13228 5856
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 12990 5400 13046 5409
rect 12990 5335 13046 5344
rect 12900 5160 12952 5166
rect 12898 5128 12900 5137
rect 12952 5128 12954 5137
rect 12898 5063 12954 5072
rect 12716 5024 12768 5030
rect 13004 5001 13032 5335
rect 12716 4966 12768 4972
rect 12990 4992 13046 5001
rect 12990 4927 13046 4936
rect 12348 4480 12400 4486
rect 12348 4422 12400 4428
rect 12622 4448 12678 4457
rect 12622 4383 12678 4392
rect 12440 4072 12492 4078
rect 12438 4040 12440 4049
rect 12492 4040 12494 4049
rect 12438 3975 12494 3984
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 11980 3664 12032 3670
rect 11980 3606 12032 3612
rect 11072 3454 11652 3482
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 10796 2650 10824 3130
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 10796 2446 10824 2586
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 10980 2378 11008 3334
rect 10968 2372 11020 2378
rect 10968 2314 11020 2320
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 11072 1465 11100 2246
rect 11058 1456 11114 1465
rect 11058 1391 11114 1400
rect 11624 480 11652 3454
rect 11992 3194 12020 3606
rect 12636 3194 12664 4383
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12728 3670 12756 3878
rect 13188 3738 13216 5646
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 12716 3664 12768 3670
rect 12716 3606 12768 3612
rect 13280 3482 13308 10095
rect 13924 9654 13952 11494
rect 15212 11150 15240 11494
rect 15764 11218 15792 11494
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15212 10674 15240 11086
rect 15764 10810 15792 11154
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 15212 10470 15240 10610
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15212 10266 15240 10406
rect 15764 10266 15792 10746
rect 15948 10266 15976 11494
rect 16304 10532 16356 10538
rect 16304 10474 16356 10480
rect 16118 10432 16174 10441
rect 16118 10367 16174 10376
rect 15200 10260 15252 10266
rect 15200 10202 15252 10208
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 14188 10124 14240 10130
rect 14188 10066 14240 10072
rect 14200 9722 14228 10066
rect 14278 10024 14334 10033
rect 14278 9959 14280 9968
rect 14332 9959 14334 9968
rect 14280 9930 14332 9936
rect 14188 9716 14240 9722
rect 14188 9658 14240 9664
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 15212 9382 15240 10202
rect 16132 9994 16160 10367
rect 16120 9988 16172 9994
rect 16120 9930 16172 9936
rect 16132 9722 16160 9930
rect 16120 9716 16172 9722
rect 16120 9658 16172 9664
rect 15752 9444 15804 9450
rect 15752 9386 15804 9392
rect 15016 9376 15068 9382
rect 14186 9344 14242 9353
rect 15016 9318 15068 9324
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 14186 9279 14242 9288
rect 14200 9178 14228 9279
rect 15028 9178 15056 9318
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 15016 9172 15068 9178
rect 15016 9114 15068 9120
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13450 8528 13506 8537
rect 13450 8463 13452 8472
rect 13504 8463 13506 8472
rect 13452 8434 13504 8440
rect 13452 8016 13504 8022
rect 13452 7958 13504 7964
rect 13360 7404 13412 7410
rect 13360 7346 13412 7352
rect 13372 6866 13400 7346
rect 13360 6860 13412 6866
rect 13360 6802 13412 6808
rect 13464 6458 13492 7958
rect 13740 7886 13768 8774
rect 15212 7886 15240 9318
rect 15764 8974 15792 9386
rect 16316 9382 16344 10474
rect 16580 10260 16632 10266
rect 16580 10202 16632 10208
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16316 9110 16344 9318
rect 16500 9178 16528 9998
rect 16592 9178 16620 10202
rect 16488 9172 16540 9178
rect 16488 9114 16540 9120
rect 16580 9172 16632 9178
rect 16580 9114 16632 9120
rect 16304 9104 16356 9110
rect 16304 9046 16356 9052
rect 15752 8968 15804 8974
rect 15752 8910 15804 8916
rect 16316 8634 16344 9046
rect 16684 8974 16712 11698
rect 17880 11694 17908 12038
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16868 11354 16896 11494
rect 17880 11354 17908 11630
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 17868 11348 17920 11354
rect 17868 11290 17920 11296
rect 18156 11014 18184 12174
rect 18248 11898 18276 12242
rect 18340 11898 18368 12378
rect 18236 11892 18288 11898
rect 18236 11834 18288 11840
rect 18328 11892 18380 11898
rect 18328 11834 18380 11840
rect 18236 11552 18288 11558
rect 18236 11494 18288 11500
rect 18144 11008 18196 11014
rect 18144 10950 18196 10956
rect 18156 10742 18184 10950
rect 18144 10736 18196 10742
rect 18144 10678 18196 10684
rect 18156 10470 18184 10678
rect 18144 10464 18196 10470
rect 18142 10432 18144 10441
rect 18196 10432 18198 10441
rect 18142 10367 18198 10376
rect 18248 10266 18276 11494
rect 18984 11218 19012 12582
rect 19260 12458 19288 12718
rect 19536 12696 19564 12786
rect 19444 12668 19564 12696
rect 19260 12442 19380 12458
rect 19260 12436 19392 12442
rect 19260 12430 19340 12436
rect 19340 12378 19392 12384
rect 19444 12238 19472 12668
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19904 12102 19932 13262
rect 20088 12986 20116 13398
rect 20628 13388 20680 13394
rect 20628 13330 20680 13336
rect 20076 12980 20128 12986
rect 20076 12922 20128 12928
rect 20088 12714 20116 12922
rect 20640 12782 20668 13330
rect 20916 13326 20944 13670
rect 21100 13462 21128 13670
rect 21088 13456 21140 13462
rect 21088 13398 21140 13404
rect 20904 13320 20956 13326
rect 20904 13262 20956 13268
rect 20628 12776 20680 12782
rect 20628 12718 20680 12724
rect 20076 12708 20128 12714
rect 20076 12650 20128 12656
rect 20640 12442 20668 12718
rect 20916 12646 20944 13262
rect 22284 13184 22336 13190
rect 22284 13126 22336 13132
rect 22296 12782 22324 13126
rect 23480 12912 23532 12918
rect 23480 12854 23532 12860
rect 22284 12776 22336 12782
rect 22284 12718 22336 12724
rect 20904 12640 20956 12646
rect 20904 12582 20956 12588
rect 21916 12640 21968 12646
rect 21916 12582 21968 12588
rect 20628 12436 20680 12442
rect 20628 12378 20680 12384
rect 20916 12102 20944 12582
rect 21362 12200 21418 12209
rect 21362 12135 21418 12144
rect 19892 12096 19944 12102
rect 19892 12038 19944 12044
rect 20904 12096 20956 12102
rect 20904 12038 20956 12044
rect 19904 11626 19932 12038
rect 20916 11898 20944 12038
rect 20904 11892 20956 11898
rect 20904 11834 20956 11840
rect 20260 11688 20312 11694
rect 20260 11630 20312 11636
rect 19892 11620 19944 11626
rect 19892 11562 19944 11568
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 19708 11280 19760 11286
rect 19708 11222 19760 11228
rect 18972 11212 19024 11218
rect 18972 11154 19024 11160
rect 18788 11076 18840 11082
rect 18788 11018 18840 11024
rect 18696 10464 18748 10470
rect 18696 10406 18748 10412
rect 18236 10260 18288 10266
rect 18236 10202 18288 10208
rect 18052 10056 18104 10062
rect 17590 10024 17646 10033
rect 17590 9959 17646 9968
rect 18050 10024 18052 10033
rect 18144 10056 18196 10062
rect 18104 10024 18106 10033
rect 18144 9998 18196 10004
rect 18050 9959 18106 9968
rect 17604 9654 17632 9959
rect 17868 9920 17920 9926
rect 17868 9862 17920 9868
rect 17592 9648 17644 9654
rect 17592 9590 17644 9596
rect 17880 9160 17908 9862
rect 18156 9450 18184 9998
rect 18248 9722 18276 10202
rect 18708 10169 18736 10406
rect 18694 10160 18750 10169
rect 18694 10095 18750 10104
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18800 9654 18828 11018
rect 18984 10810 19012 11154
rect 19616 11008 19668 11014
rect 19616 10950 19668 10956
rect 18972 10804 19024 10810
rect 18972 10746 19024 10752
rect 19628 10606 19656 10950
rect 19720 10674 19748 11222
rect 19708 10668 19760 10674
rect 19708 10610 19760 10616
rect 19616 10600 19668 10606
rect 19616 10542 19668 10548
rect 19248 10464 19300 10470
rect 19248 10406 19300 10412
rect 19260 10130 19288 10406
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 19904 10248 19932 11562
rect 19984 11008 20036 11014
rect 19984 10950 20036 10956
rect 19996 10742 20024 10950
rect 20272 10810 20300 11630
rect 20352 11552 20404 11558
rect 20352 11494 20404 11500
rect 20444 11552 20496 11558
rect 20444 11494 20496 11500
rect 20812 11552 20864 11558
rect 20812 11494 20864 11500
rect 20364 11354 20392 11494
rect 20456 11354 20484 11494
rect 20352 11348 20404 11354
rect 20352 11290 20404 11296
rect 20444 11348 20496 11354
rect 20444 11290 20496 11296
rect 20456 11234 20484 11290
rect 20364 11206 20484 11234
rect 20364 11082 20392 11206
rect 20352 11076 20404 11082
rect 20352 11018 20404 11024
rect 20260 10804 20312 10810
rect 20260 10746 20312 10752
rect 19984 10736 20036 10742
rect 19984 10678 20036 10684
rect 20076 10600 20128 10606
rect 20076 10542 20128 10548
rect 19982 10432 20038 10441
rect 19982 10367 20038 10376
rect 19812 10220 19932 10248
rect 19248 10124 19300 10130
rect 19248 10066 19300 10072
rect 19260 10010 19288 10066
rect 19260 9982 19380 10010
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 18788 9648 18840 9654
rect 18788 9590 18840 9596
rect 19260 9518 19288 9862
rect 19248 9512 19300 9518
rect 19248 9454 19300 9460
rect 18144 9444 18196 9450
rect 18144 9386 18196 9392
rect 17960 9172 18012 9178
rect 17880 9132 17960 9160
rect 17960 9114 18012 9120
rect 17960 9036 18012 9042
rect 17960 8978 18012 8984
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16672 8968 16724 8974
rect 16672 8910 16724 8916
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16500 8362 16528 8910
rect 16684 8566 16712 8910
rect 17868 8900 17920 8906
rect 17868 8842 17920 8848
rect 16672 8560 16724 8566
rect 16672 8502 16724 8508
rect 16488 8356 16540 8362
rect 16488 8298 16540 8304
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 16684 8090 16712 8230
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 15476 8016 15528 8022
rect 17408 8016 17460 8022
rect 15476 7958 15528 7964
rect 17406 7984 17408 7993
rect 17460 7984 17462 7993
rect 13728 7880 13780 7886
rect 15200 7880 15252 7886
rect 13780 7828 13860 7834
rect 13728 7822 13860 7828
rect 15200 7822 15252 7828
rect 13740 7806 13860 7822
rect 13832 6866 13860 7806
rect 15212 7274 15240 7822
rect 15200 7268 15252 7274
rect 15200 7210 15252 7216
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14752 7002 14780 7142
rect 15212 7002 15240 7210
rect 15488 7206 15516 7958
rect 17406 7919 17462 7928
rect 17040 7880 17092 7886
rect 17040 7822 17092 7828
rect 17052 7546 17080 7822
rect 17776 7744 17828 7750
rect 17776 7686 17828 7692
rect 17040 7540 17092 7546
rect 17040 7482 17092 7488
rect 15476 7200 15528 7206
rect 15476 7142 15528 7148
rect 14740 6996 14792 7002
rect 14740 6938 14792 6944
rect 15200 6996 15252 7002
rect 15200 6938 15252 6944
rect 15212 6882 15240 6938
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 15120 6854 15240 6882
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13740 5778 13768 6734
rect 15120 6458 15148 6854
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15304 6497 15332 6734
rect 15290 6488 15346 6497
rect 15108 6452 15160 6458
rect 15290 6423 15346 6432
rect 15108 6394 15160 6400
rect 13912 6180 13964 6186
rect 13912 6122 13964 6128
rect 14372 6180 14424 6186
rect 14372 6122 14424 6128
rect 13820 5908 13872 5914
rect 13820 5850 13872 5856
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 13360 5568 13412 5574
rect 13360 5510 13412 5516
rect 13372 5234 13400 5510
rect 13740 5370 13768 5714
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 13832 5234 13860 5850
rect 13924 5370 13952 6122
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 14016 5710 14044 6054
rect 14384 5914 14412 6122
rect 15488 6118 15516 7142
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 15476 6112 15528 6118
rect 15476 6054 15528 6060
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 14372 5908 14424 5914
rect 14372 5850 14424 5856
rect 14004 5704 14056 5710
rect 14004 5646 14056 5652
rect 13912 5364 13964 5370
rect 13912 5306 13964 5312
rect 13360 5228 13412 5234
rect 13820 5228 13872 5234
rect 13360 5170 13412 5176
rect 13740 5188 13820 5216
rect 13452 5160 13504 5166
rect 13452 5102 13504 5108
rect 13464 4593 13492 5102
rect 13450 4584 13506 4593
rect 13450 4519 13506 4528
rect 13636 4480 13688 4486
rect 13636 4422 13688 4428
rect 12728 3454 13308 3482
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 12624 3188 12676 3194
rect 12624 3130 12676 3136
rect 12532 3120 12584 3126
rect 12532 3062 12584 3068
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12452 2582 12480 2790
rect 12440 2576 12492 2582
rect 12070 2544 12126 2553
rect 12440 2518 12492 2524
rect 12070 2479 12072 2488
rect 12124 2479 12126 2488
rect 12072 2450 12124 2456
rect 12544 2446 12572 3062
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 12728 480 12756 3454
rect 13084 2848 13136 2854
rect 13082 2816 13084 2825
rect 13136 2816 13138 2825
rect 13082 2751 13138 2760
rect 13648 2514 13676 4422
rect 13740 3738 13768 5188
rect 13820 5170 13872 5176
rect 14016 4826 14044 5646
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 14004 4820 14056 4826
rect 14004 4762 14056 4768
rect 14096 4616 14148 4622
rect 14002 4584 14058 4593
rect 14096 4558 14148 4564
rect 14002 4519 14058 4528
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13740 3194 13768 3674
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13832 3074 13860 4422
rect 13910 3904 13966 3913
rect 13910 3839 13966 3848
rect 13740 3046 13860 3074
rect 13740 2582 13768 3046
rect 13728 2576 13780 2582
rect 13728 2518 13780 2524
rect 13636 2508 13688 2514
rect 13636 2450 13688 2456
rect 13924 480 13952 3839
rect 14016 3505 14044 4519
rect 14108 4078 14136 4558
rect 14096 4072 14148 4078
rect 14096 4014 14148 4020
rect 14002 3496 14058 3505
rect 14002 3431 14058 3440
rect 14016 2990 14044 3431
rect 14004 2984 14056 2990
rect 14004 2926 14056 2932
rect 14108 2650 14136 4014
rect 14292 3233 14320 4966
rect 14384 3942 14412 5850
rect 15936 5772 15988 5778
rect 15936 5714 15988 5720
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 15476 5636 15528 5642
rect 15476 5578 15528 5584
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 14384 3534 14412 3878
rect 14568 3738 14596 5306
rect 15108 5296 15160 5302
rect 15108 5238 15160 5244
rect 15198 5264 15254 5273
rect 15014 4856 15070 4865
rect 15014 4791 15070 4800
rect 14924 3936 14976 3942
rect 14924 3878 14976 3884
rect 14936 3738 14964 3878
rect 14556 3732 14608 3738
rect 14556 3674 14608 3680
rect 14924 3732 14976 3738
rect 14924 3674 14976 3680
rect 14464 3664 14516 3670
rect 14464 3606 14516 3612
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 14278 3224 14334 3233
rect 14278 3159 14334 3168
rect 14292 3058 14320 3159
rect 14476 3058 14504 3606
rect 14568 3058 14596 3674
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14096 2644 14148 2650
rect 14096 2586 14148 2592
rect 15028 480 15056 4791
rect 15120 3670 15148 5238
rect 15198 5199 15254 5208
rect 15212 4593 15240 5199
rect 15304 4826 15332 5510
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 15198 4584 15254 4593
rect 15198 4519 15200 4528
rect 15252 4519 15254 4528
rect 15200 4490 15252 4496
rect 15212 4459 15240 4490
rect 15488 4486 15516 5578
rect 15764 5370 15792 5646
rect 15948 5370 15976 5714
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15936 5364 15988 5370
rect 15936 5306 15988 5312
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15476 4480 15528 4486
rect 15474 4448 15476 4457
rect 15528 4448 15530 4457
rect 15474 4383 15530 4392
rect 15672 3942 15700 4626
rect 15764 4282 15792 5306
rect 15844 4616 15896 4622
rect 15844 4558 15896 4564
rect 15752 4276 15804 4282
rect 15752 4218 15804 4224
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 15672 3777 15700 3878
rect 15658 3768 15714 3777
rect 15658 3703 15714 3712
rect 15108 3664 15160 3670
rect 15108 3606 15160 3612
rect 15764 3194 15792 4218
rect 15856 3738 15884 4558
rect 16224 3738 16252 6054
rect 16854 5944 16910 5953
rect 16960 5914 16988 6598
rect 17512 6458 17540 6802
rect 17788 6730 17816 7686
rect 17880 7478 17908 8842
rect 17972 8430 18000 8978
rect 18156 8838 18184 9386
rect 18880 9376 18932 9382
rect 18880 9318 18932 9324
rect 18328 9172 18380 9178
rect 18328 9114 18380 9120
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 18052 8424 18104 8430
rect 18052 8366 18104 8372
rect 17868 7472 17920 7478
rect 17868 7414 17920 7420
rect 17868 7268 17920 7274
rect 17868 7210 17920 7216
rect 17880 6798 17908 7210
rect 17972 6866 18000 8366
rect 18064 7410 18092 8366
rect 18052 7404 18104 7410
rect 18052 7346 18104 7352
rect 17960 6860 18012 6866
rect 17960 6802 18012 6808
rect 17868 6792 17920 6798
rect 17868 6734 17920 6740
rect 17776 6724 17828 6730
rect 17776 6666 17828 6672
rect 17960 6724 18012 6730
rect 17960 6666 18012 6672
rect 17500 6452 17552 6458
rect 17500 6394 17552 6400
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 16854 5879 16910 5888
rect 16948 5908 17000 5914
rect 16868 5846 16896 5879
rect 16948 5850 17000 5856
rect 16856 5840 16908 5846
rect 16856 5782 16908 5788
rect 16488 5636 16540 5642
rect 16488 5578 16540 5584
rect 16396 5024 16448 5030
rect 16396 4966 16448 4972
rect 16408 3738 16436 4966
rect 16500 3942 16528 5578
rect 16868 5234 16896 5782
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 16580 5024 16632 5030
rect 16580 4966 16632 4972
rect 16592 4758 16620 4966
rect 16580 4752 16632 4758
rect 16580 4694 16632 4700
rect 16670 4720 16726 4729
rect 16868 4690 16896 5170
rect 16960 5098 16988 5850
rect 17222 5128 17278 5137
rect 16948 5092 17000 5098
rect 17222 5063 17278 5072
rect 16948 5034 17000 5040
rect 16960 4826 16988 5034
rect 17236 4826 17264 5063
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 16670 4655 16726 4664
rect 16856 4684 16908 4690
rect 16488 3936 16540 3942
rect 16488 3878 16540 3884
rect 15844 3732 15896 3738
rect 15844 3674 15896 3680
rect 16212 3732 16264 3738
rect 16212 3674 16264 3680
rect 16396 3732 16448 3738
rect 16396 3674 16448 3680
rect 15844 3392 15896 3398
rect 15844 3334 15896 3340
rect 15752 3188 15804 3194
rect 15752 3130 15804 3136
rect 15856 2961 15884 3334
rect 16224 3194 16252 3674
rect 16684 3194 16712 4655
rect 16856 4626 16908 4632
rect 16854 4448 16910 4457
rect 16854 4383 16910 4392
rect 16212 3188 16264 3194
rect 16212 3130 16264 3136
rect 16672 3188 16724 3194
rect 16672 3130 16724 3136
rect 16684 2990 16712 3130
rect 16672 2984 16724 2990
rect 15842 2952 15898 2961
rect 16672 2926 16724 2932
rect 15842 2887 15898 2896
rect 15856 2009 15884 2887
rect 16118 2816 16174 2825
rect 16118 2751 16174 2760
rect 15842 2000 15898 2009
rect 15842 1935 15898 1944
rect 16132 480 16160 2751
rect 16868 2650 16896 4383
rect 16960 4010 16988 4762
rect 17236 4214 17264 4762
rect 17328 4622 17356 6258
rect 17972 5914 18000 6666
rect 18064 6322 18092 7346
rect 18052 6316 18104 6322
rect 18052 6258 18104 6264
rect 17960 5908 18012 5914
rect 17960 5850 18012 5856
rect 18052 5772 18104 5778
rect 18052 5714 18104 5720
rect 17958 5672 18014 5681
rect 17788 5630 17958 5658
rect 17788 5370 17816 5630
rect 17958 5607 17960 5616
rect 18012 5607 18014 5616
rect 17960 5578 18012 5584
rect 17868 5568 17920 5574
rect 17972 5547 18000 5578
rect 17868 5510 17920 5516
rect 17776 5364 17828 5370
rect 17776 5306 17828 5312
rect 17776 5024 17828 5030
rect 17774 4992 17776 5001
rect 17828 4992 17830 5001
rect 17774 4927 17830 4936
rect 17776 4752 17828 4758
rect 17776 4694 17828 4700
rect 17592 4684 17644 4690
rect 17592 4626 17644 4632
rect 17316 4616 17368 4622
rect 17316 4558 17368 4564
rect 17328 4282 17356 4558
rect 17604 4282 17632 4626
rect 17316 4276 17368 4282
rect 17316 4218 17368 4224
rect 17592 4276 17644 4282
rect 17592 4218 17644 4224
rect 17224 4208 17276 4214
rect 17224 4150 17276 4156
rect 17408 4140 17460 4146
rect 17408 4082 17460 4088
rect 16948 4004 17000 4010
rect 16948 3946 17000 3952
rect 17316 3664 17368 3670
rect 17038 3632 17094 3641
rect 17038 3567 17094 3576
rect 17314 3632 17316 3641
rect 17368 3632 17370 3641
rect 17420 3602 17448 4082
rect 17682 3768 17738 3777
rect 17788 3738 17816 4694
rect 17682 3703 17738 3712
rect 17776 3732 17828 3738
rect 17696 3602 17724 3703
rect 17776 3674 17828 3680
rect 17314 3567 17370 3576
rect 17408 3596 17460 3602
rect 17052 3194 17080 3567
rect 17408 3538 17460 3544
rect 17684 3596 17736 3602
rect 17684 3538 17736 3544
rect 17420 3505 17448 3538
rect 17406 3496 17462 3505
rect 17406 3431 17462 3440
rect 17696 3233 17724 3538
rect 17880 3534 17908 5510
rect 18064 5001 18092 5714
rect 18156 5370 18184 8774
rect 18340 8634 18368 9114
rect 18892 9042 18920 9318
rect 19352 9178 19380 9982
rect 19812 9926 19840 10220
rect 19800 9920 19852 9926
rect 19800 9862 19852 9868
rect 19812 9586 19840 9862
rect 19800 9580 19852 9586
rect 19800 9522 19852 9528
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 19432 9104 19484 9110
rect 19432 9046 19484 9052
rect 19996 9058 20024 10367
rect 20088 9722 20116 10542
rect 20364 10198 20392 11018
rect 20824 10606 20852 11494
rect 20916 11150 20944 11834
rect 21180 11688 21232 11694
rect 21180 11630 21232 11636
rect 21192 11286 21220 11630
rect 21376 11558 21404 12135
rect 21928 11694 21956 12582
rect 23492 12238 23520 12854
rect 23480 12232 23532 12238
rect 23480 12174 23532 12180
rect 23492 11898 23520 12174
rect 23480 11892 23532 11898
rect 23480 11834 23532 11840
rect 23492 11694 23520 11834
rect 21916 11688 21968 11694
rect 21916 11630 21968 11636
rect 23480 11688 23532 11694
rect 23480 11630 23532 11636
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 23492 11286 23520 11630
rect 21180 11280 21232 11286
rect 21180 11222 21232 11228
rect 23480 11280 23532 11286
rect 23480 11222 23532 11228
rect 20904 11144 20956 11150
rect 20904 11086 20956 11092
rect 20812 10600 20864 10606
rect 20812 10542 20864 10548
rect 20916 10470 20944 11086
rect 20904 10464 20956 10470
rect 20904 10406 20956 10412
rect 21916 10464 21968 10470
rect 21916 10406 21968 10412
rect 20352 10192 20404 10198
rect 20258 10160 20314 10169
rect 20352 10134 20404 10140
rect 20258 10095 20314 10104
rect 20168 9920 20220 9926
rect 20168 9862 20220 9868
rect 20076 9716 20128 9722
rect 20076 9658 20128 9664
rect 20180 9450 20208 9862
rect 20168 9444 20220 9450
rect 20272 9432 20300 10095
rect 20364 9654 20392 10134
rect 20916 9926 20944 10406
rect 20904 9920 20956 9926
rect 20904 9862 20956 9868
rect 20352 9648 20404 9654
rect 20352 9590 20404 9596
rect 20916 9518 20944 9862
rect 20904 9512 20956 9518
rect 20904 9454 20956 9460
rect 20272 9404 20392 9432
rect 20168 9386 20220 9392
rect 20180 9178 20208 9386
rect 20168 9172 20220 9178
rect 20168 9114 20220 9120
rect 18880 9036 18932 9042
rect 18880 8978 18932 8984
rect 18788 8968 18840 8974
rect 18788 8910 18840 8916
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 18328 8356 18380 8362
rect 18328 8298 18380 8304
rect 18236 7948 18288 7954
rect 18236 7890 18288 7896
rect 18248 7857 18276 7890
rect 18234 7848 18290 7857
rect 18234 7783 18290 7792
rect 18248 7546 18276 7783
rect 18236 7540 18288 7546
rect 18236 7482 18288 7488
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 18050 4992 18106 5001
rect 18050 4927 18106 4936
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 17682 3224 17738 3233
rect 17040 3188 17092 3194
rect 17682 3159 17684 3168
rect 17040 3130 17092 3136
rect 17736 3159 17738 3168
rect 17684 3130 17736 3136
rect 17696 3099 17724 3130
rect 17880 2650 17908 3470
rect 18156 3194 18184 3470
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 16856 2644 16908 2650
rect 16856 2586 16908 2592
rect 17868 2644 17920 2650
rect 17868 2586 17920 2592
rect 17222 2408 17278 2417
rect 17222 2343 17278 2352
rect 17236 480 17264 2343
rect 18340 480 18368 8298
rect 18800 7993 18828 8910
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 19352 8514 19380 8570
rect 19260 8486 19380 8514
rect 18786 7984 18842 7993
rect 18786 7919 18842 7928
rect 19260 7886 19288 8486
rect 19340 8356 19392 8362
rect 19340 8298 19392 8304
rect 19352 8022 19380 8298
rect 19340 8016 19392 8022
rect 19340 7958 19392 7964
rect 18512 7880 18564 7886
rect 18512 7822 18564 7828
rect 19248 7880 19300 7886
rect 19248 7822 19300 7828
rect 18524 7274 18552 7822
rect 19444 7342 19472 9046
rect 19996 9030 20208 9058
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 19524 7948 19576 7954
rect 19524 7890 19576 7896
rect 19536 7546 19564 7890
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 20076 7540 20128 7546
rect 20076 7482 20128 7488
rect 19432 7336 19484 7342
rect 19432 7278 19484 7284
rect 18512 7268 18564 7274
rect 18512 7210 18564 7216
rect 19432 7200 19484 7206
rect 19432 7142 19484 7148
rect 19444 6798 19472 7142
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 19984 6860 20036 6866
rect 19984 6802 20036 6808
rect 18420 6792 18472 6798
rect 18420 6734 18472 6740
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 18432 6186 18460 6734
rect 19432 6656 19484 6662
rect 19432 6598 19484 6604
rect 19156 6248 19208 6254
rect 19156 6190 19208 6196
rect 18420 6180 18472 6186
rect 18420 6122 18472 6128
rect 18878 5808 18934 5817
rect 18878 5743 18880 5752
rect 18932 5743 18934 5752
rect 18880 5714 18932 5720
rect 19168 5370 19196 6190
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 19352 5953 19380 6054
rect 19338 5944 19394 5953
rect 19338 5879 19394 5888
rect 19156 5364 19208 5370
rect 19156 5306 19208 5312
rect 18418 5264 18474 5273
rect 18418 5199 18474 5208
rect 18972 5228 19024 5234
rect 18432 3194 18460 5199
rect 18972 5170 19024 5176
rect 18880 5024 18932 5030
rect 18880 4966 18932 4972
rect 18892 4729 18920 4966
rect 18878 4720 18934 4729
rect 18878 4655 18934 4664
rect 18602 4448 18658 4457
rect 18602 4383 18658 4392
rect 18616 4282 18644 4383
rect 18604 4276 18656 4282
rect 18604 4218 18656 4224
rect 18984 3194 19012 5170
rect 19338 4992 19394 5001
rect 19338 4927 19394 4936
rect 19352 4826 19380 4927
rect 19340 4820 19392 4826
rect 19340 4762 19392 4768
rect 19444 4758 19472 6598
rect 19996 6458 20024 6802
rect 19984 6452 20036 6458
rect 19984 6394 20036 6400
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 19892 5568 19944 5574
rect 19892 5510 19944 5516
rect 19904 5137 19932 5510
rect 19890 5128 19946 5137
rect 19890 5063 19892 5072
rect 19944 5063 19946 5072
rect 19892 5034 19944 5040
rect 19904 5003 19932 5034
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 19432 4752 19484 4758
rect 19432 4694 19484 4700
rect 19616 4752 19668 4758
rect 19616 4694 19668 4700
rect 19156 4480 19208 4486
rect 19156 4422 19208 4428
rect 19064 3936 19116 3942
rect 19064 3878 19116 3884
rect 19076 3369 19104 3878
rect 19168 3641 19196 4422
rect 19444 4146 19472 4694
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 19628 4078 19656 4694
rect 19984 4276 20036 4282
rect 19984 4218 20036 4224
rect 19616 4072 19668 4078
rect 19616 4014 19668 4020
rect 19996 3942 20024 4218
rect 19432 3936 19484 3942
rect 19432 3878 19484 3884
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 19444 3777 19472 3878
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19430 3768 19486 3777
rect 19580 3760 19876 3780
rect 20088 3777 20116 7482
rect 20180 4282 20208 9030
rect 20168 4276 20220 4282
rect 20168 4218 20220 4224
rect 20168 4072 20220 4078
rect 20168 4014 20220 4020
rect 20074 3768 20130 3777
rect 19430 3703 19486 3712
rect 20180 3738 20208 4014
rect 20074 3703 20130 3712
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 19154 3632 19210 3641
rect 20364 3618 20392 9404
rect 20444 9376 20496 9382
rect 20444 9318 20496 9324
rect 20456 9110 20484 9318
rect 20444 9104 20496 9110
rect 20444 9046 20496 9052
rect 20916 8974 20944 9454
rect 21364 9104 21416 9110
rect 21928 9081 21956 10406
rect 23584 10146 23612 13806
rect 24228 13802 24348 13818
rect 24216 13796 24348 13802
rect 24268 13790 24348 13796
rect 24216 13738 24268 13744
rect 24228 13462 24256 13738
rect 24308 13728 24360 13734
rect 24308 13670 24360 13676
rect 24216 13456 24268 13462
rect 24216 13398 24268 13404
rect 24228 12918 24256 13398
rect 24320 13394 24348 13670
rect 24308 13388 24360 13394
rect 24308 13330 24360 13336
rect 24320 12986 24348 13330
rect 24860 13184 24912 13190
rect 24780 13132 24860 13138
rect 24780 13126 24912 13132
rect 24780 13110 24900 13126
rect 24308 12980 24360 12986
rect 24308 12922 24360 12928
rect 24216 12912 24268 12918
rect 24216 12854 24268 12860
rect 24780 12306 24808 13110
rect 25424 12986 25452 14214
rect 25884 13870 25912 14758
rect 25976 13938 26004 15438
rect 25964 13932 26016 13938
rect 25964 13874 26016 13880
rect 25872 13864 25924 13870
rect 25872 13806 25924 13812
rect 25780 13728 25832 13734
rect 25780 13670 25832 13676
rect 25872 13728 25924 13734
rect 25872 13670 25924 13676
rect 25792 13190 25820 13670
rect 25884 13530 25912 13670
rect 25872 13524 25924 13530
rect 25872 13466 25924 13472
rect 25872 13388 25924 13394
rect 25872 13330 25924 13336
rect 25780 13184 25832 13190
rect 25780 13126 25832 13132
rect 25044 12980 25096 12986
rect 25044 12922 25096 12928
rect 25412 12980 25464 12986
rect 25412 12922 25464 12928
rect 23664 12300 23716 12306
rect 23664 12242 23716 12248
rect 24768 12300 24820 12306
rect 24768 12242 24820 12248
rect 23676 11354 23704 12242
rect 25056 12209 25084 12922
rect 25424 12782 25452 12922
rect 25412 12776 25464 12782
rect 25884 12753 25912 13330
rect 25976 13258 26004 13874
rect 25964 13252 26016 13258
rect 25964 13194 26016 13200
rect 25976 12986 26004 13194
rect 25964 12980 26016 12986
rect 25964 12922 26016 12928
rect 25412 12718 25464 12724
rect 25870 12744 25926 12753
rect 25870 12679 25872 12688
rect 25924 12679 25926 12688
rect 25872 12650 25924 12656
rect 25976 12442 26004 12922
rect 25964 12436 26016 12442
rect 25964 12378 26016 12384
rect 25688 12232 25740 12238
rect 25042 12200 25098 12209
rect 25688 12174 25740 12180
rect 25042 12135 25098 12144
rect 25136 12096 25188 12102
rect 25136 12038 25188 12044
rect 25320 12096 25372 12102
rect 25320 12038 25372 12044
rect 25148 11626 25176 12038
rect 25332 11898 25360 12038
rect 25320 11892 25372 11898
rect 25320 11834 25372 11840
rect 25136 11620 25188 11626
rect 25136 11562 25188 11568
rect 24398 11384 24454 11393
rect 23664 11348 23716 11354
rect 24398 11319 24400 11328
rect 23664 11290 23716 11296
rect 24452 11319 24454 11328
rect 24860 11348 24912 11354
rect 24400 11290 24452 11296
rect 24860 11290 24912 11296
rect 24492 11212 24544 11218
rect 24492 11154 24544 11160
rect 24504 10810 24532 11154
rect 24872 10810 24900 11290
rect 25148 11218 25176 11562
rect 25332 11354 25360 11834
rect 25700 11694 25728 12174
rect 25688 11688 25740 11694
rect 25688 11630 25740 11636
rect 25320 11348 25372 11354
rect 25320 11290 25372 11296
rect 25700 11218 25728 11630
rect 25136 11212 25188 11218
rect 25136 11154 25188 11160
rect 25688 11212 25740 11218
rect 25688 11154 25740 11160
rect 25976 11150 26004 12378
rect 25228 11144 25280 11150
rect 25228 11086 25280 11092
rect 25964 11144 26016 11150
rect 25964 11086 26016 11092
rect 25240 10810 25268 11086
rect 25870 10976 25926 10985
rect 25870 10911 25926 10920
rect 25884 10810 25912 10911
rect 24492 10804 24544 10810
rect 24492 10746 24544 10752
rect 24860 10804 24912 10810
rect 24860 10746 24912 10752
rect 25228 10804 25280 10810
rect 25228 10746 25280 10752
rect 25872 10804 25924 10810
rect 25872 10746 25924 10752
rect 26068 10441 26096 21286
rect 26148 21072 26200 21078
rect 26148 21014 26200 21020
rect 26160 20466 26188 21014
rect 26148 20460 26200 20466
rect 26148 20402 26200 20408
rect 26160 18426 26188 20402
rect 26252 20398 26280 22578
rect 26988 22574 27016 23258
rect 26976 22568 27028 22574
rect 26976 22510 27028 22516
rect 27172 22506 27200 23287
rect 27896 23180 27948 23186
rect 27896 23122 27948 23128
rect 27908 22778 27936 23122
rect 28184 23050 28212 23462
rect 28276 23322 28304 23666
rect 28264 23316 28316 23322
rect 28264 23258 28316 23264
rect 28356 23180 28408 23186
rect 28356 23122 28408 23128
rect 28172 23044 28224 23050
rect 28172 22986 28224 22992
rect 28080 22976 28132 22982
rect 28080 22918 28132 22924
rect 27896 22772 27948 22778
rect 27896 22714 27948 22720
rect 27528 22636 27580 22642
rect 27528 22578 27580 22584
rect 27160 22500 27212 22506
rect 27160 22442 27212 22448
rect 26884 22432 26936 22438
rect 26884 22374 26936 22380
rect 26792 22024 26844 22030
rect 26792 21966 26844 21972
rect 26516 21888 26568 21894
rect 26516 21830 26568 21836
rect 26332 21480 26384 21486
rect 26528 21457 26556 21830
rect 26804 21593 26832 21966
rect 26790 21584 26846 21593
rect 26790 21519 26846 21528
rect 26332 21422 26384 21428
rect 26514 21448 26570 21457
rect 26344 21078 26372 21422
rect 26514 21383 26516 21392
rect 26568 21383 26570 21392
rect 26516 21354 26568 21360
rect 26804 21146 26832 21519
rect 26896 21146 26924 22374
rect 27172 22098 27200 22442
rect 27436 22228 27488 22234
rect 27436 22170 27488 22176
rect 27160 22092 27212 22098
rect 27160 22034 27212 22040
rect 27252 22024 27304 22030
rect 27448 22001 27476 22170
rect 27252 21966 27304 21972
rect 27434 21992 27490 22001
rect 27264 21418 27292 21966
rect 27434 21927 27490 21936
rect 27540 21672 27568 22578
rect 27712 22024 27764 22030
rect 27712 21966 27764 21972
rect 27620 21684 27672 21690
rect 27540 21644 27620 21672
rect 27620 21626 27672 21632
rect 27252 21412 27304 21418
rect 27252 21354 27304 21360
rect 26792 21140 26844 21146
rect 26792 21082 26844 21088
rect 26884 21140 26936 21146
rect 26884 21082 26936 21088
rect 26332 21072 26384 21078
rect 26332 21014 26384 21020
rect 26700 21004 26752 21010
rect 26700 20946 26752 20952
rect 26240 20392 26292 20398
rect 26240 20334 26292 20340
rect 26252 20058 26280 20334
rect 26712 20058 26740 20946
rect 26896 20058 26924 21082
rect 27160 20936 27212 20942
rect 27160 20878 27212 20884
rect 27172 20602 27200 20878
rect 27264 20874 27292 21354
rect 27724 21146 27752 21966
rect 28092 21690 28120 22918
rect 28184 22030 28212 22986
rect 28368 22778 28396 23122
rect 28460 23118 28488 23802
rect 29104 23338 29132 28698
rect 29840 28082 29868 29174
rect 30760 29170 30788 29446
rect 30852 29238 30880 29650
rect 30840 29232 30892 29238
rect 30840 29174 30892 29180
rect 30748 29164 30800 29170
rect 30748 29106 30800 29112
rect 30472 29096 30524 29102
rect 30472 29038 30524 29044
rect 30380 29028 30432 29034
rect 30380 28970 30432 28976
rect 30392 28778 30420 28970
rect 30300 28762 30420 28778
rect 30288 28756 30420 28762
rect 30340 28750 30420 28756
rect 30288 28698 30340 28704
rect 30484 28626 30512 29038
rect 31588 29034 31616 31078
rect 31956 30938 31984 31078
rect 31944 30932 31996 30938
rect 31944 30874 31996 30880
rect 32140 30666 32168 31282
rect 33060 30938 33088 31622
rect 33796 31385 33824 31962
rect 34152 31952 34204 31958
rect 34152 31894 34204 31900
rect 34164 31822 34192 31894
rect 34152 31816 34204 31822
rect 34152 31758 34204 31764
rect 33782 31376 33838 31385
rect 33782 31311 33838 31320
rect 33796 30954 33824 31311
rect 33048 30932 33100 30938
rect 33048 30874 33100 30880
rect 33600 30932 33652 30938
rect 33796 30926 33916 30954
rect 33600 30874 33652 30880
rect 32680 30728 32732 30734
rect 32680 30670 32732 30676
rect 31668 30660 31720 30666
rect 31668 30602 31720 30608
rect 32128 30660 32180 30666
rect 32128 30602 32180 30608
rect 31680 30326 31708 30602
rect 31760 30592 31812 30598
rect 31760 30534 31812 30540
rect 31668 30320 31720 30326
rect 31668 30262 31720 30268
rect 31772 29186 31800 30534
rect 32692 30394 32720 30670
rect 33060 30394 33088 30874
rect 33140 30728 33192 30734
rect 33140 30670 33192 30676
rect 32680 30388 32732 30394
rect 32680 30330 32732 30336
rect 33048 30388 33100 30394
rect 33048 30330 33100 30336
rect 32128 29708 32180 29714
rect 32128 29650 32180 29656
rect 32140 29306 32168 29650
rect 32128 29300 32180 29306
rect 32128 29242 32180 29248
rect 33152 29238 33180 30670
rect 33612 30190 33640 30874
rect 33888 30258 33916 30926
rect 33876 30252 33928 30258
rect 33876 30194 33928 30200
rect 33600 30184 33652 30190
rect 33600 30126 33652 30132
rect 33692 30048 33744 30054
rect 33692 29990 33744 29996
rect 33704 29850 33732 29990
rect 33692 29844 33744 29850
rect 33692 29786 33744 29792
rect 33888 29510 33916 30194
rect 34164 29782 34192 31758
rect 34440 31686 34468 32506
rect 34520 31884 34572 31890
rect 34520 31826 34572 31832
rect 34244 31680 34296 31686
rect 34244 31622 34296 31628
rect 34428 31680 34480 31686
rect 34428 31622 34480 31628
rect 34256 30938 34284 31622
rect 34532 31498 34560 31826
rect 34704 31816 34756 31822
rect 34704 31758 34756 31764
rect 34612 31680 34664 31686
rect 34612 31622 34664 31628
rect 34440 31482 34560 31498
rect 34624 31482 34652 31622
rect 34428 31476 34560 31482
rect 34480 31470 34560 31476
rect 34612 31476 34664 31482
rect 34428 31418 34480 31424
rect 34612 31418 34664 31424
rect 34624 30954 34652 31418
rect 34716 31210 34744 31758
rect 34704 31204 34756 31210
rect 34704 31146 34756 31152
rect 34244 30932 34296 30938
rect 34244 30874 34296 30880
rect 34532 30926 34652 30954
rect 34532 30802 34560 30926
rect 34612 30864 34664 30870
rect 34612 30806 34664 30812
rect 34520 30796 34572 30802
rect 34520 30738 34572 30744
rect 34532 30394 34560 30738
rect 34624 30598 34652 30806
rect 34612 30592 34664 30598
rect 34612 30534 34664 30540
rect 34520 30388 34572 30394
rect 34520 30330 34572 30336
rect 34520 30116 34572 30122
rect 34520 30058 34572 30064
rect 34152 29776 34204 29782
rect 34152 29718 34204 29724
rect 34532 29646 34560 30058
rect 34624 30054 34652 30534
rect 34612 30048 34664 30054
rect 34612 29990 34664 29996
rect 34624 29714 34652 29990
rect 34808 29730 34836 33254
rect 34900 33046 34928 33510
rect 34888 33040 34940 33046
rect 34888 32982 34940 32988
rect 34940 32668 35236 32688
rect 34996 32666 35020 32668
rect 35076 32666 35100 32668
rect 35156 32666 35180 32668
rect 35018 32614 35020 32666
rect 35082 32614 35094 32666
rect 35156 32614 35158 32666
rect 34996 32612 35020 32614
rect 35076 32612 35100 32614
rect 35156 32612 35180 32614
rect 34940 32592 35236 32612
rect 35164 32292 35216 32298
rect 35164 32234 35216 32240
rect 35176 31890 35204 32234
rect 35164 31884 35216 31890
rect 35164 31826 35216 31832
rect 35348 31884 35400 31890
rect 35348 31826 35400 31832
rect 34940 31580 35236 31600
rect 34996 31578 35020 31580
rect 35076 31578 35100 31580
rect 35156 31578 35180 31580
rect 35018 31526 35020 31578
rect 35082 31526 35094 31578
rect 35156 31526 35158 31578
rect 34996 31524 35020 31526
rect 35076 31524 35100 31526
rect 35156 31524 35180 31526
rect 34940 31504 35236 31524
rect 35164 31204 35216 31210
rect 35164 31146 35216 31152
rect 35176 30938 35204 31146
rect 35164 30932 35216 30938
rect 35164 30874 35216 30880
rect 34940 30492 35236 30512
rect 34996 30490 35020 30492
rect 35076 30490 35100 30492
rect 35156 30490 35180 30492
rect 35018 30438 35020 30490
rect 35082 30438 35094 30490
rect 35156 30438 35158 30490
rect 34996 30436 35020 30438
rect 35076 30436 35100 30438
rect 35156 30436 35180 30438
rect 34940 30416 35236 30436
rect 34888 30252 34940 30258
rect 34888 30194 34940 30200
rect 34900 29850 34928 30194
rect 34888 29844 34940 29850
rect 34888 29786 34940 29792
rect 34612 29708 34664 29714
rect 34612 29650 34664 29656
rect 34716 29702 34836 29730
rect 34520 29640 34572 29646
rect 34440 29588 34520 29594
rect 34440 29582 34572 29588
rect 34440 29566 34560 29582
rect 33876 29504 33928 29510
rect 33876 29446 33928 29452
rect 31680 29158 31800 29186
rect 33140 29232 33192 29238
rect 33140 29174 33192 29180
rect 34334 29200 34390 29209
rect 31680 29102 31708 29158
rect 34334 29135 34336 29144
rect 34388 29135 34390 29144
rect 34336 29106 34388 29112
rect 31668 29096 31720 29102
rect 31668 29038 31720 29044
rect 31576 29028 31628 29034
rect 31576 28970 31628 28976
rect 32310 28792 32366 28801
rect 34440 28762 34468 29566
rect 34624 29306 34652 29650
rect 34612 29300 34664 29306
rect 34612 29242 34664 29248
rect 32310 28727 32366 28736
rect 34428 28756 34480 28762
rect 30472 28620 30524 28626
rect 30472 28562 30524 28568
rect 30484 28218 30512 28562
rect 32220 28552 32272 28558
rect 32220 28494 32272 28500
rect 30656 28416 30708 28422
rect 30656 28358 30708 28364
rect 30472 28212 30524 28218
rect 30472 28154 30524 28160
rect 29828 28076 29880 28082
rect 29828 28018 29880 28024
rect 29840 27674 29868 28018
rect 30668 28014 30696 28358
rect 32232 28218 32260 28494
rect 32324 28218 32352 28727
rect 34428 28698 34480 28704
rect 32220 28212 32272 28218
rect 32220 28154 32272 28160
rect 32312 28212 32364 28218
rect 32312 28154 32364 28160
rect 32232 28014 32260 28154
rect 34518 28112 34574 28121
rect 32864 28076 32916 28082
rect 34518 28047 34574 28056
rect 32864 28018 32916 28024
rect 30656 28008 30708 28014
rect 30656 27950 30708 27956
rect 32220 28008 32272 28014
rect 32220 27950 32272 27956
rect 31668 27940 31720 27946
rect 31668 27882 31720 27888
rect 31680 27674 31708 27882
rect 29828 27668 29880 27674
rect 29828 27610 29880 27616
rect 31668 27668 31720 27674
rect 31668 27610 31720 27616
rect 31852 27532 31904 27538
rect 31852 27474 31904 27480
rect 30104 27464 30156 27470
rect 30104 27406 30156 27412
rect 31300 27464 31352 27470
rect 31300 27406 31352 27412
rect 29552 27396 29604 27402
rect 29552 27338 29604 27344
rect 29184 26988 29236 26994
rect 29184 26930 29236 26936
rect 29196 26790 29224 26930
rect 29564 26926 29592 27338
rect 29552 26920 29604 26926
rect 29552 26862 29604 26868
rect 29184 26784 29236 26790
rect 29184 26726 29236 26732
rect 29196 26500 29224 26726
rect 29564 26586 29592 26862
rect 29552 26580 29604 26586
rect 29552 26522 29604 26528
rect 29368 26512 29420 26518
rect 29196 26472 29368 26500
rect 29196 25702 29224 26472
rect 29368 26454 29420 26460
rect 29276 25832 29328 25838
rect 29276 25774 29328 25780
rect 29184 25696 29236 25702
rect 29184 25638 29236 25644
rect 29288 25498 29316 25774
rect 29550 25528 29606 25537
rect 29276 25492 29328 25498
rect 30116 25498 30144 27406
rect 31312 27130 31340 27406
rect 31300 27124 31352 27130
rect 31300 27066 31352 27072
rect 30656 26784 30708 26790
rect 30656 26726 30708 26732
rect 30668 25838 30696 26726
rect 31864 26314 31892 27474
rect 32588 27464 32640 27470
rect 32588 27406 32640 27412
rect 32036 27396 32088 27402
rect 32036 27338 32088 27344
rect 32048 26926 32076 27338
rect 32036 26920 32088 26926
rect 32036 26862 32088 26868
rect 32048 26518 32076 26862
rect 32404 26852 32456 26858
rect 32404 26794 32456 26800
rect 32036 26512 32088 26518
rect 32036 26454 32088 26460
rect 31852 26308 31904 26314
rect 31852 26250 31904 26256
rect 30380 25832 30432 25838
rect 30380 25774 30432 25780
rect 30656 25832 30708 25838
rect 30656 25774 30708 25780
rect 30288 25764 30340 25770
rect 30288 25706 30340 25712
rect 29550 25463 29552 25472
rect 29276 25434 29328 25440
rect 29604 25463 29606 25472
rect 30104 25492 30156 25498
rect 29552 25434 29604 25440
rect 30104 25434 30156 25440
rect 30116 24954 30144 25434
rect 30300 25294 30328 25706
rect 30392 25702 30420 25774
rect 30380 25696 30432 25702
rect 30380 25638 30432 25644
rect 31864 25537 31892 26250
rect 32048 26042 32076 26454
rect 32416 26382 32444 26794
rect 32404 26376 32456 26382
rect 32404 26318 32456 26324
rect 32036 26036 32088 26042
rect 32036 25978 32088 25984
rect 32416 25838 32444 26318
rect 32404 25832 32456 25838
rect 32404 25774 32456 25780
rect 32128 25696 32180 25702
rect 32128 25638 32180 25644
rect 31850 25528 31906 25537
rect 31850 25463 31906 25472
rect 30472 25424 30524 25430
rect 30472 25366 30524 25372
rect 30288 25288 30340 25294
rect 30288 25230 30340 25236
rect 30104 24948 30156 24954
rect 30104 24890 30156 24896
rect 30300 24886 30328 25230
rect 30288 24880 30340 24886
rect 30288 24822 30340 24828
rect 30380 24608 30432 24614
rect 30380 24550 30432 24556
rect 30392 24410 30420 24550
rect 30380 24404 30432 24410
rect 30380 24346 30432 24352
rect 30484 24342 30512 25366
rect 31942 25256 31998 25265
rect 31942 25191 31944 25200
rect 31996 25191 31998 25200
rect 31944 25162 31996 25168
rect 30932 24676 30984 24682
rect 30932 24618 30984 24624
rect 30472 24336 30524 24342
rect 30472 24278 30524 24284
rect 29828 24064 29880 24070
rect 29828 24006 29880 24012
rect 29840 23730 29868 24006
rect 29828 23724 29880 23730
rect 29828 23666 29880 23672
rect 28920 23310 29132 23338
rect 28920 23254 28948 23310
rect 28908 23248 28960 23254
rect 28908 23190 28960 23196
rect 29840 23186 29868 23666
rect 29828 23180 29880 23186
rect 29828 23122 29880 23128
rect 28448 23112 28500 23118
rect 28448 23054 28500 23060
rect 28460 22778 28488 23054
rect 29368 22976 29420 22982
rect 29368 22918 29420 22924
rect 30656 22976 30708 22982
rect 30656 22918 30708 22924
rect 28356 22772 28408 22778
rect 28356 22714 28408 22720
rect 28448 22772 28500 22778
rect 28448 22714 28500 22720
rect 28632 22772 28684 22778
rect 28632 22714 28684 22720
rect 28644 22080 28672 22714
rect 29380 22574 29408 22918
rect 29368 22568 29420 22574
rect 29368 22510 29420 22516
rect 30472 22432 30524 22438
rect 30472 22374 30524 22380
rect 28460 22052 28672 22080
rect 29552 22092 29604 22098
rect 28172 22024 28224 22030
rect 28172 21966 28224 21972
rect 28080 21684 28132 21690
rect 28080 21626 28132 21632
rect 27712 21140 27764 21146
rect 27712 21082 27764 21088
rect 28460 21010 28488 22052
rect 29552 22034 29604 22040
rect 29090 21992 29146 22001
rect 29090 21927 29146 21936
rect 29276 21956 29328 21962
rect 29104 21350 29132 21927
rect 29276 21898 29328 21904
rect 29288 21593 29316 21898
rect 29564 21894 29592 22034
rect 30012 22024 30064 22030
rect 30012 21966 30064 21972
rect 30288 22024 30340 22030
rect 30340 21972 30420 21978
rect 30288 21966 30420 21972
rect 29552 21888 29604 21894
rect 29552 21830 29604 21836
rect 29736 21888 29788 21894
rect 29736 21830 29788 21836
rect 29564 21690 29592 21830
rect 29552 21684 29604 21690
rect 29552 21626 29604 21632
rect 29274 21584 29330 21593
rect 29564 21554 29592 21626
rect 29274 21519 29276 21528
rect 29328 21519 29330 21528
rect 29552 21548 29604 21554
rect 29276 21490 29328 21496
rect 29552 21490 29604 21496
rect 29092 21344 29144 21350
rect 28998 21312 29054 21321
rect 29092 21286 29144 21292
rect 28998 21247 29054 21256
rect 29012 21146 29040 21247
rect 29000 21140 29052 21146
rect 29000 21082 29052 21088
rect 28448 21004 28500 21010
rect 28448 20946 28500 20952
rect 28632 21004 28684 21010
rect 28632 20946 28684 20952
rect 27252 20868 27304 20874
rect 27252 20810 27304 20816
rect 27160 20596 27212 20602
rect 27160 20538 27212 20544
rect 28460 20262 28488 20946
rect 28644 20913 28672 20946
rect 28630 20904 28686 20913
rect 28630 20839 28686 20848
rect 28448 20256 28500 20262
rect 28448 20198 28500 20204
rect 28644 20058 28672 20839
rect 29644 20800 29696 20806
rect 29644 20742 29696 20748
rect 29368 20528 29420 20534
rect 29366 20496 29368 20505
rect 29420 20496 29422 20505
rect 29366 20431 29422 20440
rect 28816 20256 28868 20262
rect 28816 20198 28868 20204
rect 26240 20052 26292 20058
rect 26240 19994 26292 20000
rect 26700 20052 26752 20058
rect 26700 19994 26752 20000
rect 26884 20052 26936 20058
rect 26884 19994 26936 20000
rect 28632 20052 28684 20058
rect 28632 19994 28684 20000
rect 28828 19174 28856 20198
rect 28816 19168 28868 19174
rect 28816 19110 28868 19116
rect 28264 18896 28316 18902
rect 28264 18838 28316 18844
rect 28172 18828 28224 18834
rect 28172 18770 28224 18776
rect 26148 18420 26200 18426
rect 26148 18362 26200 18368
rect 28080 18148 28132 18154
rect 28080 18090 28132 18096
rect 27160 18080 27212 18086
rect 27160 18022 27212 18028
rect 27172 17105 27200 18022
rect 28092 17678 28120 18090
rect 28184 18086 28212 18770
rect 28172 18080 28224 18086
rect 28172 18022 28224 18028
rect 28080 17672 28132 17678
rect 28080 17614 28132 17620
rect 27988 17536 28040 17542
rect 27988 17478 28040 17484
rect 28000 17134 28028 17478
rect 27988 17128 28040 17134
rect 27158 17096 27214 17105
rect 27988 17070 28040 17076
rect 27158 17031 27214 17040
rect 28092 16998 28120 17614
rect 28184 17270 28212 18022
rect 28172 17264 28224 17270
rect 28172 17206 28224 17212
rect 28184 17134 28212 17206
rect 28276 17202 28304 18838
rect 28828 18766 28856 19110
rect 28816 18760 28868 18766
rect 28816 18702 28868 18708
rect 28540 18216 28592 18222
rect 28540 18158 28592 18164
rect 28552 17814 28580 18158
rect 28828 18154 28856 18702
rect 29000 18624 29052 18630
rect 28920 18572 29000 18578
rect 28920 18566 29052 18572
rect 28920 18550 29040 18566
rect 28816 18148 28868 18154
rect 28816 18090 28868 18096
rect 28540 17808 28592 17814
rect 28540 17750 28592 17756
rect 28920 17542 28948 18550
rect 29276 18080 29328 18086
rect 29276 18022 29328 18028
rect 28908 17536 28960 17542
rect 28908 17478 28960 17484
rect 28264 17196 28316 17202
rect 28264 17138 28316 17144
rect 28172 17128 28224 17134
rect 28170 17096 28172 17105
rect 28224 17096 28226 17105
rect 28170 17031 28226 17040
rect 28080 16992 28132 16998
rect 28080 16934 28132 16940
rect 28356 16992 28408 16998
rect 28356 16934 28408 16940
rect 26516 16652 26568 16658
rect 26516 16594 26568 16600
rect 26528 16561 26556 16594
rect 28368 16590 28396 16934
rect 28632 16652 28684 16658
rect 28632 16594 28684 16600
rect 27528 16584 27580 16590
rect 26514 16552 26570 16561
rect 27528 16526 27580 16532
rect 28356 16584 28408 16590
rect 28356 16526 28408 16532
rect 26514 16487 26570 16496
rect 26700 16448 26752 16454
rect 26700 16390 26752 16396
rect 26240 15904 26292 15910
rect 26240 15846 26292 15852
rect 26252 14822 26280 15846
rect 26424 15496 26476 15502
rect 26424 15438 26476 15444
rect 26332 15360 26384 15366
rect 26436 15337 26464 15438
rect 26516 15360 26568 15366
rect 26332 15302 26384 15308
rect 26422 15328 26478 15337
rect 26344 15201 26372 15302
rect 26516 15302 26568 15308
rect 26422 15263 26478 15272
rect 26330 15192 26386 15201
rect 26436 15162 26464 15263
rect 26330 15127 26386 15136
rect 26424 15156 26476 15162
rect 26424 15098 26476 15104
rect 26528 14958 26556 15302
rect 26516 14952 26568 14958
rect 26516 14894 26568 14900
rect 26240 14816 26292 14822
rect 26240 14758 26292 14764
rect 26712 14618 26740 16390
rect 27540 16114 27568 16526
rect 27528 16108 27580 16114
rect 27528 16050 27580 16056
rect 28368 15910 28396 16526
rect 28644 16250 28672 16594
rect 29288 16250 29316 18022
rect 29552 17876 29604 17882
rect 29552 17818 29604 17824
rect 29564 17134 29592 17818
rect 29552 17128 29604 17134
rect 29552 17070 29604 17076
rect 29656 16946 29684 20742
rect 29748 20466 29776 21830
rect 30024 21554 30052 21966
rect 30300 21950 30420 21966
rect 30012 21548 30064 21554
rect 30012 21490 30064 21496
rect 30392 21350 30420 21950
rect 30484 21457 30512 22374
rect 30668 22030 30696 22918
rect 30656 22024 30708 22030
rect 30656 21966 30708 21972
rect 30470 21448 30526 21457
rect 30470 21383 30526 21392
rect 29828 21344 29880 21350
rect 29828 21286 29880 21292
rect 30380 21344 30432 21350
rect 30380 21286 30432 21292
rect 29840 21078 29868 21286
rect 29828 21072 29880 21078
rect 29828 21014 29880 21020
rect 30288 20936 30340 20942
rect 30288 20878 30340 20884
rect 29736 20460 29788 20466
rect 29736 20402 29788 20408
rect 30012 20460 30064 20466
rect 30012 20402 30064 20408
rect 30024 20058 30052 20402
rect 30300 20330 30328 20878
rect 30392 20806 30420 21286
rect 30380 20800 30432 20806
rect 30380 20742 30432 20748
rect 30484 20466 30512 21383
rect 30668 21146 30696 21966
rect 30944 21962 30972 24618
rect 32140 22574 32168 25638
rect 32600 25265 32628 27406
rect 32876 27130 32904 28018
rect 34244 27600 34296 27606
rect 34244 27542 34296 27548
rect 33876 27464 33928 27470
rect 33876 27406 33928 27412
rect 32864 27124 32916 27130
rect 32864 27066 32916 27072
rect 32876 26518 32904 27066
rect 33888 26858 33916 27406
rect 33876 26852 33928 26858
rect 33876 26794 33928 26800
rect 34256 26790 34284 27542
rect 34244 26784 34296 26790
rect 34244 26726 34296 26732
rect 33876 26580 33928 26586
rect 33876 26522 33928 26528
rect 32864 26512 32916 26518
rect 32864 26454 32916 26460
rect 32678 26208 32734 26217
rect 32678 26143 32734 26152
rect 32692 25498 32720 26143
rect 32680 25492 32732 25498
rect 32680 25434 32732 25440
rect 32876 25430 32904 26454
rect 33416 26308 33468 26314
rect 33416 26250 33468 26256
rect 33428 26194 33456 26250
rect 33336 26166 33456 26194
rect 33232 25696 33284 25702
rect 33232 25638 33284 25644
rect 32864 25424 32916 25430
rect 32864 25366 32916 25372
rect 33048 25356 33100 25362
rect 33048 25298 33100 25304
rect 32680 25288 32732 25294
rect 32586 25256 32642 25265
rect 32680 25230 32732 25236
rect 32586 25191 32642 25200
rect 32600 24818 32628 25191
rect 32312 24812 32364 24818
rect 32312 24754 32364 24760
rect 32588 24812 32640 24818
rect 32588 24754 32640 24760
rect 32324 24410 32352 24754
rect 32692 24614 32720 25230
rect 32680 24608 32732 24614
rect 32680 24550 32732 24556
rect 32312 24404 32364 24410
rect 32312 24346 32364 24352
rect 32692 24070 32720 24550
rect 33060 24410 33088 25298
rect 33244 24886 33272 25638
rect 33336 25294 33364 26166
rect 33888 25906 33916 26522
rect 34256 26314 34284 26726
rect 34244 26308 34296 26314
rect 34244 26250 34296 26256
rect 33876 25900 33928 25906
rect 33876 25842 33928 25848
rect 33692 25696 33744 25702
rect 33692 25638 33744 25644
rect 33704 25537 33732 25638
rect 33690 25528 33746 25537
rect 33690 25463 33692 25472
rect 33744 25463 33746 25472
rect 33692 25434 33744 25440
rect 33704 25403 33732 25434
rect 33324 25288 33376 25294
rect 33324 25230 33376 25236
rect 34060 25288 34112 25294
rect 34060 25230 34112 25236
rect 33232 24880 33284 24886
rect 33232 24822 33284 24828
rect 33336 24410 33364 25230
rect 33048 24404 33100 24410
rect 33048 24346 33100 24352
rect 33324 24404 33376 24410
rect 33324 24346 33376 24352
rect 34072 24070 34100 25230
rect 32680 24064 32732 24070
rect 32680 24006 32732 24012
rect 34060 24064 34112 24070
rect 34060 24006 34112 24012
rect 32692 23497 32720 24006
rect 32678 23488 32734 23497
rect 32678 23423 32734 23432
rect 32956 22772 33008 22778
rect 32956 22714 33008 22720
rect 32128 22568 32180 22574
rect 32128 22510 32180 22516
rect 32140 22438 32168 22510
rect 32968 22506 32996 22714
rect 32956 22500 33008 22506
rect 32956 22442 33008 22448
rect 32128 22432 32180 22438
rect 32128 22374 32180 22380
rect 33600 22432 33652 22438
rect 33600 22374 33652 22380
rect 31760 22092 31812 22098
rect 31760 22034 31812 22040
rect 30932 21956 30984 21962
rect 30932 21898 30984 21904
rect 30656 21140 30708 21146
rect 30656 21082 30708 21088
rect 30944 21010 30972 21898
rect 31772 21690 31800 22034
rect 31760 21684 31812 21690
rect 31680 21644 31760 21672
rect 30932 21004 30984 21010
rect 30932 20946 30984 20952
rect 31680 20466 31708 21644
rect 31760 21626 31812 21632
rect 32140 21554 32168 22374
rect 32588 22024 32640 22030
rect 32588 21966 32640 21972
rect 32312 21956 32364 21962
rect 32312 21898 32364 21904
rect 32128 21548 32180 21554
rect 32128 21490 32180 21496
rect 31944 21480 31996 21486
rect 31944 21422 31996 21428
rect 31956 21146 31984 21422
rect 32140 21418 32168 21490
rect 32128 21412 32180 21418
rect 32128 21354 32180 21360
rect 32324 21350 32352 21898
rect 32312 21344 32364 21350
rect 32312 21286 32364 21292
rect 31944 21140 31996 21146
rect 31944 21082 31996 21088
rect 32324 20942 32352 21286
rect 32312 20936 32364 20942
rect 32310 20904 32312 20913
rect 32404 20936 32456 20942
rect 32364 20904 32366 20913
rect 32404 20878 32456 20884
rect 32310 20839 32366 20848
rect 30472 20460 30524 20466
rect 30472 20402 30524 20408
rect 31668 20460 31720 20466
rect 31668 20402 31720 20408
rect 30288 20324 30340 20330
rect 30288 20266 30340 20272
rect 30012 20052 30064 20058
rect 30012 19994 30064 20000
rect 30012 19712 30064 19718
rect 30012 19654 30064 19660
rect 30024 19242 30052 19654
rect 30012 19236 30064 19242
rect 30012 19178 30064 19184
rect 29920 18896 29972 18902
rect 29920 18838 29972 18844
rect 29932 18290 29960 18838
rect 30024 18630 30052 19178
rect 32416 19174 32444 20878
rect 32600 20602 32628 21966
rect 32956 21888 33008 21894
rect 32956 21830 33008 21836
rect 33140 21888 33192 21894
rect 33140 21830 33192 21836
rect 32772 21140 32824 21146
rect 32772 21082 32824 21088
rect 32588 20596 32640 20602
rect 32588 20538 32640 20544
rect 32784 20534 32812 21082
rect 32968 20942 32996 21830
rect 33152 21010 33180 21830
rect 33612 21486 33640 22374
rect 34072 21962 34100 24006
rect 34244 23656 34296 23662
rect 34244 23598 34296 23604
rect 34256 23322 34284 23598
rect 34426 23488 34482 23497
rect 34426 23423 34482 23432
rect 34244 23316 34296 23322
rect 34244 23258 34296 23264
rect 34440 22681 34468 23423
rect 34532 23338 34560 28047
rect 34612 26784 34664 26790
rect 34612 26726 34664 26732
rect 34624 26382 34652 26726
rect 34612 26376 34664 26382
rect 34612 26318 34664 26324
rect 34716 26330 34744 29702
rect 34900 29594 34928 29786
rect 34808 29566 34928 29594
rect 35256 29640 35308 29646
rect 35256 29582 35308 29588
rect 34808 29306 34836 29566
rect 34940 29404 35236 29424
rect 34996 29402 35020 29404
rect 35076 29402 35100 29404
rect 35156 29402 35180 29404
rect 35018 29350 35020 29402
rect 35082 29350 35094 29402
rect 35156 29350 35158 29402
rect 34996 29348 35020 29350
rect 35076 29348 35100 29350
rect 35156 29348 35180 29350
rect 34940 29328 35236 29348
rect 34796 29300 34848 29306
rect 34796 29242 34848 29248
rect 34980 29028 35032 29034
rect 34980 28970 35032 28976
rect 34992 28762 35020 28970
rect 34980 28756 35032 28762
rect 34980 28698 35032 28704
rect 34940 28316 35236 28336
rect 34996 28314 35020 28316
rect 35076 28314 35100 28316
rect 35156 28314 35180 28316
rect 35018 28262 35020 28314
rect 35082 28262 35094 28314
rect 35156 28262 35158 28314
rect 34996 28260 35020 28262
rect 35076 28260 35100 28262
rect 35156 28260 35180 28262
rect 34940 28240 35236 28260
rect 35268 28218 35296 29582
rect 35256 28212 35308 28218
rect 35256 28154 35308 28160
rect 35256 27328 35308 27334
rect 35256 27270 35308 27276
rect 34940 27228 35236 27248
rect 34996 27226 35020 27228
rect 35076 27226 35100 27228
rect 35156 27226 35180 27228
rect 35018 27174 35020 27226
rect 35082 27174 35094 27226
rect 35156 27174 35158 27226
rect 34996 27172 35020 27174
rect 35076 27172 35100 27174
rect 35156 27172 35180 27174
rect 34940 27152 35236 27172
rect 35268 26518 35296 27270
rect 35256 26512 35308 26518
rect 35256 26454 35308 26460
rect 34624 25838 34652 26318
rect 34716 26302 34836 26330
rect 34704 26240 34756 26246
rect 34702 26208 34704 26217
rect 34756 26208 34758 26217
rect 34702 26143 34758 26152
rect 34716 25838 34744 26143
rect 34808 25974 34836 26302
rect 34940 26140 35236 26160
rect 34996 26138 35020 26140
rect 35076 26138 35100 26140
rect 35156 26138 35180 26140
rect 35018 26086 35020 26138
rect 35082 26086 35094 26138
rect 35156 26086 35158 26138
rect 34996 26084 35020 26086
rect 35076 26084 35100 26086
rect 35156 26084 35180 26086
rect 34940 26064 35236 26084
rect 34796 25968 34848 25974
rect 34796 25910 34848 25916
rect 35268 25906 35296 26454
rect 35256 25900 35308 25906
rect 35256 25842 35308 25848
rect 34612 25832 34664 25838
rect 34612 25774 34664 25780
rect 34704 25832 34756 25838
rect 34704 25774 34756 25780
rect 35164 25696 35216 25702
rect 35164 25638 35216 25644
rect 35176 25294 35204 25638
rect 34612 25288 34664 25294
rect 34888 25288 34940 25294
rect 34612 25230 34664 25236
rect 34808 25236 34888 25242
rect 34808 25230 34940 25236
rect 35164 25288 35216 25294
rect 35164 25230 35216 25236
rect 34624 24954 34652 25230
rect 34808 25214 34928 25230
rect 34808 24954 34836 25214
rect 34940 25052 35236 25072
rect 34996 25050 35020 25052
rect 35076 25050 35100 25052
rect 35156 25050 35180 25052
rect 35018 24998 35020 25050
rect 35082 24998 35094 25050
rect 35156 24998 35158 25050
rect 34996 24996 35020 24998
rect 35076 24996 35100 24998
rect 35156 24996 35180 24998
rect 34940 24976 35236 24996
rect 34612 24948 34664 24954
rect 34796 24948 34848 24954
rect 34664 24908 34744 24936
rect 34612 24890 34664 24896
rect 34612 24064 34664 24070
rect 34612 24006 34664 24012
rect 34624 23526 34652 24006
rect 34612 23520 34664 23526
rect 34612 23462 34664 23468
rect 34532 23310 34652 23338
rect 34426 22672 34482 22681
rect 34426 22607 34482 22616
rect 34244 22432 34296 22438
rect 34244 22374 34296 22380
rect 34518 22400 34574 22409
rect 34060 21956 34112 21962
rect 34060 21898 34112 21904
rect 33876 21888 33928 21894
rect 33876 21830 33928 21836
rect 33232 21480 33284 21486
rect 33232 21422 33284 21428
rect 33600 21480 33652 21486
rect 33600 21422 33652 21428
rect 33140 21004 33192 21010
rect 33140 20946 33192 20952
rect 32956 20936 33008 20942
rect 32956 20878 33008 20884
rect 32968 20754 32996 20878
rect 32968 20726 33180 20754
rect 33152 20602 33180 20726
rect 33140 20596 33192 20602
rect 33140 20538 33192 20544
rect 32772 20528 32824 20534
rect 32772 20470 32824 20476
rect 33244 20466 33272 21422
rect 33324 20936 33376 20942
rect 33324 20878 33376 20884
rect 32588 20460 32640 20466
rect 32588 20402 32640 20408
rect 33232 20460 33284 20466
rect 33232 20402 33284 20408
rect 31024 19168 31076 19174
rect 31024 19110 31076 19116
rect 32404 19168 32456 19174
rect 32404 19110 32456 19116
rect 31036 18630 31064 19110
rect 30012 18624 30064 18630
rect 30012 18566 30064 18572
rect 31024 18624 31076 18630
rect 31024 18566 31076 18572
rect 29920 18284 29972 18290
rect 29920 18226 29972 18232
rect 29736 18216 29788 18222
rect 29736 18158 29788 18164
rect 29564 16918 29684 16946
rect 28632 16244 28684 16250
rect 28632 16186 28684 16192
rect 29276 16244 29328 16250
rect 29276 16186 29328 16192
rect 26884 15904 26936 15910
rect 26884 15846 26936 15852
rect 28356 15904 28408 15910
rect 28356 15846 28408 15852
rect 26896 15570 26924 15846
rect 28644 15745 28672 16186
rect 29184 15904 29236 15910
rect 29184 15846 29236 15852
rect 28630 15736 28686 15745
rect 28630 15671 28686 15680
rect 29196 15570 29224 15846
rect 26884 15564 26936 15570
rect 26884 15506 26936 15512
rect 27528 15564 27580 15570
rect 27528 15506 27580 15512
rect 29184 15564 29236 15570
rect 29184 15506 29236 15512
rect 29460 15564 29512 15570
rect 29460 15506 29512 15512
rect 27540 15450 27568 15506
rect 26792 15428 26844 15434
rect 27540 15422 27660 15450
rect 26792 15370 26844 15376
rect 26804 14890 26832 15370
rect 27528 15360 27580 15366
rect 27528 15302 27580 15308
rect 26792 14884 26844 14890
rect 26792 14826 26844 14832
rect 26700 14612 26752 14618
rect 26700 14554 26752 14560
rect 26332 14272 26384 14278
rect 26332 14214 26384 14220
rect 26700 14272 26752 14278
rect 26700 14214 26752 14220
rect 26344 13938 26372 14214
rect 26332 13932 26384 13938
rect 26332 13874 26384 13880
rect 26608 13864 26660 13870
rect 26608 13806 26660 13812
rect 26240 13728 26292 13734
rect 26240 13670 26292 13676
rect 26516 13728 26568 13734
rect 26516 13670 26568 13676
rect 26252 10810 26280 13670
rect 26528 11393 26556 13670
rect 26620 13530 26648 13806
rect 26608 13524 26660 13530
rect 26608 13466 26660 13472
rect 26712 11393 26740 14214
rect 26804 13938 26832 14826
rect 27068 14816 27120 14822
rect 27068 14758 27120 14764
rect 27080 14482 27108 14758
rect 27068 14476 27120 14482
rect 27068 14418 27120 14424
rect 27080 14074 27108 14418
rect 27540 14414 27568 15302
rect 27632 15162 27660 15422
rect 29196 15162 29224 15506
rect 27620 15156 27672 15162
rect 27620 15098 27672 15104
rect 29184 15156 29236 15162
rect 29184 15098 29236 15104
rect 29472 14958 29500 15506
rect 29460 14952 29512 14958
rect 29460 14894 29512 14900
rect 28448 14884 28500 14890
rect 28448 14826 28500 14832
rect 28460 14618 28488 14826
rect 28080 14612 28132 14618
rect 28080 14554 28132 14560
rect 28448 14612 28500 14618
rect 28448 14554 28500 14560
rect 27528 14408 27580 14414
rect 27528 14350 27580 14356
rect 27540 14113 27568 14350
rect 27620 14272 27672 14278
rect 27620 14214 27672 14220
rect 27804 14272 27856 14278
rect 27804 14214 27856 14220
rect 27526 14104 27582 14113
rect 27068 14068 27120 14074
rect 27526 14039 27582 14048
rect 27068 14010 27120 14016
rect 26792 13932 26844 13938
rect 26792 13874 26844 13880
rect 26804 13462 26832 13874
rect 27632 13818 27660 14214
rect 27540 13790 27660 13818
rect 27816 13802 27844 14214
rect 28092 14006 28120 14554
rect 28906 14104 28962 14113
rect 28906 14039 28962 14048
rect 28080 14000 28132 14006
rect 28080 13942 28132 13948
rect 28920 13818 28948 14039
rect 27804 13796 27856 13802
rect 27540 13734 27568 13790
rect 28920 13790 29040 13818
rect 27804 13738 27856 13744
rect 27068 13728 27120 13734
rect 27068 13670 27120 13676
rect 27528 13728 27580 13734
rect 27528 13670 27580 13676
rect 26792 13456 26844 13462
rect 26792 13398 26844 13404
rect 26976 13388 27028 13394
rect 26976 13330 27028 13336
rect 26792 13320 26844 13326
rect 26792 13262 26844 13268
rect 26804 12782 26832 13262
rect 26988 12918 27016 13330
rect 26976 12912 27028 12918
rect 26976 12854 27028 12860
rect 26792 12776 26844 12782
rect 26792 12718 26844 12724
rect 26804 12374 26832 12718
rect 26792 12368 26844 12374
rect 26792 12310 26844 12316
rect 26804 11898 26832 12310
rect 26792 11892 26844 11898
rect 26792 11834 26844 11840
rect 26514 11384 26570 11393
rect 26514 11319 26570 11328
rect 26698 11384 26754 11393
rect 26698 11319 26754 11328
rect 27080 10810 27108 13670
rect 27434 13560 27490 13569
rect 27816 13530 27844 13738
rect 27434 13495 27490 13504
rect 27804 13524 27856 13530
rect 27448 12986 27476 13495
rect 27804 13466 27856 13472
rect 28080 13388 28132 13394
rect 28080 13330 28132 13336
rect 27436 12980 27488 12986
rect 27436 12922 27488 12928
rect 27896 12912 27948 12918
rect 27896 12854 27948 12860
rect 27908 12442 27936 12854
rect 28092 12442 28120 13330
rect 28172 13320 28224 13326
rect 28172 13262 28224 13268
rect 28184 12986 28212 13262
rect 28264 13184 28316 13190
rect 28264 13126 28316 13132
rect 28172 12980 28224 12986
rect 28172 12922 28224 12928
rect 27896 12436 27948 12442
rect 27896 12378 27948 12384
rect 28080 12436 28132 12442
rect 28080 12378 28132 12384
rect 27908 11286 27936 12378
rect 28276 11898 28304 13126
rect 28816 12980 28868 12986
rect 28816 12922 28868 12928
rect 28722 12200 28778 12209
rect 28722 12135 28778 12144
rect 28736 11898 28764 12135
rect 28828 12102 28856 12922
rect 29012 12918 29040 13790
rect 29368 13184 29420 13190
rect 29368 13126 29420 13132
rect 29000 12912 29052 12918
rect 29000 12854 29052 12860
rect 29380 12850 29408 13126
rect 29368 12844 29420 12850
rect 29368 12786 29420 12792
rect 29276 12640 29328 12646
rect 29276 12582 29328 12588
rect 29092 12368 29144 12374
rect 29092 12310 29144 12316
rect 29000 12300 29052 12306
rect 29000 12242 29052 12248
rect 28816 12096 28868 12102
rect 28816 12038 28868 12044
rect 28264 11892 28316 11898
rect 28264 11834 28316 11840
rect 28724 11892 28776 11898
rect 28724 11834 28776 11840
rect 28736 11694 28764 11834
rect 28724 11688 28776 11694
rect 28724 11630 28776 11636
rect 28828 11626 28856 12038
rect 29012 11898 29040 12242
rect 29000 11892 29052 11898
rect 29000 11834 29052 11840
rect 28816 11620 28868 11626
rect 28816 11562 28868 11568
rect 28828 11354 28856 11562
rect 29012 11354 29040 11834
rect 29104 11558 29132 12310
rect 29092 11552 29144 11558
rect 29092 11494 29144 11500
rect 28816 11348 28868 11354
rect 28816 11290 28868 11296
rect 29000 11348 29052 11354
rect 29000 11290 29052 11296
rect 27896 11280 27948 11286
rect 27896 11222 27948 11228
rect 27252 11212 27304 11218
rect 27252 11154 27304 11160
rect 27158 10840 27214 10849
rect 26240 10804 26292 10810
rect 26240 10746 26292 10752
rect 27068 10804 27120 10810
rect 27158 10775 27160 10784
rect 27068 10746 27120 10752
rect 27212 10775 27214 10784
rect 27160 10746 27212 10752
rect 26252 10606 26280 10746
rect 27264 10742 27292 11154
rect 27908 10810 27936 11222
rect 29000 11144 29052 11150
rect 28920 11092 29000 11098
rect 28920 11086 29052 11092
rect 28920 11070 29040 11086
rect 28920 10810 28948 11070
rect 29104 10810 29132 11494
rect 27896 10804 27948 10810
rect 27896 10746 27948 10752
rect 28908 10804 28960 10810
rect 28908 10746 28960 10752
rect 29092 10804 29144 10810
rect 29092 10746 29144 10752
rect 27252 10736 27304 10742
rect 28724 10736 28776 10742
rect 27252 10678 27304 10684
rect 28722 10704 28724 10713
rect 29288 10713 29316 12582
rect 29458 11384 29514 11393
rect 29368 11348 29420 11354
rect 29458 11319 29514 11328
rect 29368 11290 29420 11296
rect 29380 10810 29408 11290
rect 29368 10804 29420 10810
rect 29368 10746 29420 10752
rect 28776 10704 28778 10713
rect 28722 10639 28778 10648
rect 29274 10704 29330 10713
rect 29274 10639 29330 10648
rect 26240 10600 26292 10606
rect 26240 10542 26292 10548
rect 26054 10432 26110 10441
rect 26054 10367 26110 10376
rect 29472 10266 29500 11319
rect 29460 10260 29512 10266
rect 29460 10202 29512 10208
rect 23584 10118 23704 10146
rect 22008 9920 22060 9926
rect 22008 9862 22060 9868
rect 22020 9518 22048 9862
rect 22008 9512 22060 9518
rect 22008 9454 22060 9460
rect 22284 9376 22336 9382
rect 22284 9318 22336 9324
rect 22296 9110 22324 9318
rect 22284 9104 22336 9110
rect 21364 9046 21416 9052
rect 21914 9072 21970 9081
rect 20904 8968 20956 8974
rect 20904 8910 20956 8916
rect 20916 8362 20944 8910
rect 21376 8634 21404 9046
rect 22284 9046 22336 9052
rect 21914 9007 21970 9016
rect 21364 8628 21416 8634
rect 21364 8570 21416 8576
rect 20904 8356 20956 8362
rect 20904 8298 20956 8304
rect 21088 8084 21140 8090
rect 21088 8026 21140 8032
rect 20444 8016 20496 8022
rect 21100 7993 21128 8026
rect 20444 7958 20496 7964
rect 21086 7984 21142 7993
rect 20456 7585 20484 7958
rect 21086 7919 21142 7928
rect 21456 7948 21508 7954
rect 21456 7890 21508 7896
rect 20718 7848 20774 7857
rect 20718 7783 20774 7792
rect 20442 7576 20498 7585
rect 20732 7546 20760 7783
rect 21468 7546 21496 7890
rect 20442 7511 20444 7520
rect 20496 7511 20498 7520
rect 20720 7540 20772 7546
rect 20444 7482 20496 7488
rect 20720 7482 20772 7488
rect 21456 7540 21508 7546
rect 21456 7482 21508 7488
rect 21928 6905 21956 9007
rect 22284 8832 22336 8838
rect 22284 8774 22336 8780
rect 22100 8288 22152 8294
rect 22100 8230 22152 8236
rect 22112 7546 22140 8230
rect 22296 7585 22324 8774
rect 23480 8356 23532 8362
rect 23480 8298 23532 8304
rect 23492 7954 23520 8298
rect 23572 8016 23624 8022
rect 23676 7993 23704 10118
rect 28908 10124 28960 10130
rect 28908 10066 28960 10072
rect 25412 9920 25464 9926
rect 25412 9862 25464 9868
rect 25424 9518 25452 9862
rect 28920 9722 28948 10066
rect 28908 9716 28960 9722
rect 28908 9658 28960 9664
rect 25412 9512 25464 9518
rect 25412 9454 25464 9460
rect 25424 9178 25452 9454
rect 26516 9376 26568 9382
rect 26516 9318 26568 9324
rect 26700 9376 26752 9382
rect 26700 9318 26752 9324
rect 25412 9172 25464 9178
rect 25412 9114 25464 9120
rect 24308 8832 24360 8838
rect 24308 8774 24360 8780
rect 24768 8832 24820 8838
rect 24768 8774 24820 8780
rect 25320 8832 25372 8838
rect 25320 8774 25372 8780
rect 24320 8430 24348 8774
rect 24308 8424 24360 8430
rect 24308 8366 24360 8372
rect 24320 8090 24348 8366
rect 24308 8084 24360 8090
rect 24308 8026 24360 8032
rect 24676 8084 24728 8090
rect 24676 8026 24728 8032
rect 23572 7958 23624 7964
rect 23662 7984 23718 7993
rect 23480 7948 23532 7954
rect 23480 7890 23532 7896
rect 22282 7576 22338 7585
rect 22100 7540 22152 7546
rect 23492 7546 23520 7890
rect 22282 7511 22338 7520
rect 23480 7540 23532 7546
rect 22100 7482 22152 7488
rect 23480 7482 23532 7488
rect 20442 6896 20498 6905
rect 20442 6831 20498 6840
rect 21914 6896 21970 6905
rect 21914 6831 21970 6840
rect 20456 5817 20484 6831
rect 22112 6798 22140 7482
rect 23584 7206 23612 7958
rect 23662 7919 23718 7928
rect 23940 7268 23992 7274
rect 23940 7210 23992 7216
rect 22468 7200 22520 7206
rect 22468 7142 22520 7148
rect 22652 7200 22704 7206
rect 22652 7142 22704 7148
rect 23572 7200 23624 7206
rect 23572 7142 23624 7148
rect 22376 6860 22428 6866
rect 22376 6802 22428 6808
rect 21916 6792 21968 6798
rect 21916 6734 21968 6740
rect 22100 6792 22152 6798
rect 22100 6734 22152 6740
rect 21928 6458 21956 6734
rect 22008 6656 22060 6662
rect 22008 6598 22060 6604
rect 21916 6452 21968 6458
rect 21916 6394 21968 6400
rect 22020 6390 22048 6598
rect 22008 6384 22060 6390
rect 22008 6326 22060 6332
rect 22388 6322 22416 6802
rect 22376 6316 22428 6322
rect 22376 6258 22428 6264
rect 22008 6112 22060 6118
rect 22008 6054 22060 6060
rect 22020 5953 22048 6054
rect 22006 5944 22062 5953
rect 22388 5914 22416 6258
rect 22006 5879 22062 5888
rect 22376 5908 22428 5914
rect 22376 5850 22428 5856
rect 20442 5808 20498 5817
rect 20442 5743 20498 5752
rect 20720 5772 20772 5778
rect 20456 4826 20484 5743
rect 20720 5714 20772 5720
rect 20536 5704 20588 5710
rect 20732 5681 20760 5714
rect 20904 5704 20956 5710
rect 20536 5646 20588 5652
rect 20718 5672 20774 5681
rect 20444 4820 20496 4826
rect 20444 4762 20496 4768
rect 20442 4720 20498 4729
rect 20442 4655 20498 4664
rect 19154 3567 19210 3576
rect 19444 3590 20392 3618
rect 19062 3360 19118 3369
rect 19062 3295 19118 3304
rect 18420 3188 18472 3194
rect 18420 3130 18472 3136
rect 18972 3188 19024 3194
rect 18972 3130 19024 3136
rect 18878 3088 18934 3097
rect 18878 3023 18880 3032
rect 18932 3023 18934 3032
rect 18880 2994 18932 3000
rect 18984 2650 19012 3130
rect 19168 2650 19196 3567
rect 19246 3496 19302 3505
rect 19246 3431 19302 3440
rect 18972 2644 19024 2650
rect 18972 2586 19024 2592
rect 19156 2644 19208 2650
rect 19156 2586 19208 2592
rect 19260 2582 19288 3431
rect 19248 2576 19300 2582
rect 19248 2518 19300 2524
rect 19444 480 19472 3590
rect 19984 3460 20036 3466
rect 19984 3402 20036 3408
rect 19996 2990 20024 3402
rect 20456 3074 20484 4655
rect 20548 3210 20576 5646
rect 20904 5646 20956 5652
rect 20718 5607 20774 5616
rect 20732 5370 20760 5607
rect 20720 5364 20772 5370
rect 20720 5306 20772 5312
rect 20916 5166 20944 5646
rect 22480 5642 22508 7142
rect 22664 7041 22692 7142
rect 22650 7032 22706 7041
rect 22650 6967 22706 6976
rect 23480 6656 23532 6662
rect 23480 6598 23532 6604
rect 22560 6316 22612 6322
rect 22560 6258 22612 6264
rect 22468 5636 22520 5642
rect 22468 5578 22520 5584
rect 22008 5296 22060 5302
rect 22006 5264 22008 5273
rect 22060 5264 22062 5273
rect 22572 5234 22600 6258
rect 23492 6186 23520 6598
rect 23584 6458 23612 7142
rect 23952 6662 23980 7210
rect 23940 6656 23992 6662
rect 23940 6598 23992 6604
rect 24124 6656 24176 6662
rect 24124 6598 24176 6604
rect 23572 6452 23624 6458
rect 23572 6394 23624 6400
rect 24032 6384 24084 6390
rect 24136 6372 24164 6598
rect 24688 6458 24716 8026
rect 24780 6730 24808 8774
rect 25042 7032 25098 7041
rect 25042 6967 25098 6976
rect 24768 6724 24820 6730
rect 24768 6666 24820 6672
rect 24860 6656 24912 6662
rect 24860 6598 24912 6604
rect 24676 6452 24728 6458
rect 24676 6394 24728 6400
rect 24084 6344 24164 6372
rect 24032 6326 24084 6332
rect 24136 6338 24164 6344
rect 24136 6322 24256 6338
rect 24136 6316 24268 6322
rect 24136 6310 24216 6316
rect 24216 6258 24268 6264
rect 24688 6254 24716 6394
rect 24872 6361 24900 6598
rect 24858 6352 24914 6361
rect 24858 6287 24914 6296
rect 24676 6248 24728 6254
rect 24676 6190 24728 6196
rect 23480 6180 23532 6186
rect 23480 6122 23532 6128
rect 23664 6112 23716 6118
rect 23664 6054 23716 6060
rect 24766 6080 24822 6089
rect 23676 5914 23704 6054
rect 24766 6015 24822 6024
rect 23846 5944 23902 5953
rect 23664 5908 23716 5914
rect 23846 5879 23848 5888
rect 23664 5850 23716 5856
rect 23900 5879 23902 5888
rect 23848 5850 23900 5856
rect 22836 5568 22888 5574
rect 22836 5510 22888 5516
rect 22006 5199 22062 5208
rect 22560 5228 22612 5234
rect 22560 5170 22612 5176
rect 20904 5160 20956 5166
rect 20904 5102 20956 5108
rect 20628 5092 20680 5098
rect 20628 5034 20680 5040
rect 20640 4978 20668 5034
rect 21822 4992 21878 5001
rect 20640 4950 20852 4978
rect 20628 4140 20680 4146
rect 20628 4082 20680 4088
rect 20640 3738 20668 4082
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 20548 3194 20760 3210
rect 20548 3188 20772 3194
rect 20548 3182 20720 3188
rect 20720 3130 20772 3136
rect 20456 3046 20576 3074
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 19996 2650 20024 2926
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 20548 480 20576 3046
rect 20628 2916 20680 2922
rect 20628 2858 20680 2864
rect 20640 2802 20668 2858
rect 20824 2854 20852 4950
rect 21822 4927 21878 4936
rect 21836 4826 21864 4927
rect 21824 4820 21876 4826
rect 21824 4762 21876 4768
rect 22192 4684 22244 4690
rect 22192 4626 22244 4632
rect 21272 4480 21324 4486
rect 21270 4448 21272 4457
rect 21324 4448 21326 4457
rect 21270 4383 21326 4392
rect 22204 4282 22232 4626
rect 22572 4622 22600 5170
rect 22848 5166 22876 5510
rect 23860 5370 23888 5850
rect 24216 5704 24268 5710
rect 24216 5646 24268 5652
rect 24124 5568 24176 5574
rect 24124 5510 24176 5516
rect 23848 5364 23900 5370
rect 23848 5306 23900 5312
rect 24136 5273 24164 5510
rect 24122 5264 24178 5273
rect 24228 5234 24256 5646
rect 24780 5302 24808 6015
rect 24860 5568 24912 5574
rect 24860 5510 24912 5516
rect 24768 5296 24820 5302
rect 24768 5238 24820 5244
rect 24122 5199 24124 5208
rect 24176 5199 24178 5208
rect 24216 5228 24268 5234
rect 24124 5170 24176 5176
rect 24216 5170 24268 5176
rect 22836 5160 22888 5166
rect 22836 5102 22888 5108
rect 23388 5160 23440 5166
rect 24228 5137 24256 5170
rect 23388 5102 23440 5108
rect 24214 5128 24270 5137
rect 23112 5024 23164 5030
rect 23112 4966 23164 4972
rect 22284 4616 22336 4622
rect 22284 4558 22336 4564
rect 22560 4616 22612 4622
rect 22560 4558 22612 4564
rect 22192 4276 22244 4282
rect 22192 4218 22244 4224
rect 21364 3936 21416 3942
rect 21364 3878 21416 3884
rect 21376 3641 21404 3878
rect 21638 3768 21694 3777
rect 21638 3703 21694 3712
rect 21362 3632 21418 3641
rect 21362 3567 21364 3576
rect 21416 3567 21418 3576
rect 21364 3538 21416 3544
rect 20904 3392 20956 3398
rect 20904 3334 20956 3340
rect 20916 3058 20944 3334
rect 21376 3126 21404 3538
rect 21456 3528 21508 3534
rect 21454 3496 21456 3505
rect 21508 3496 21510 3505
rect 21454 3431 21510 3440
rect 21364 3120 21416 3126
rect 21364 3062 21416 3068
rect 20904 3052 20956 3058
rect 20904 2994 20956 3000
rect 20812 2848 20864 2854
rect 20640 2774 20760 2802
rect 20812 2790 20864 2796
rect 20732 2650 20760 2774
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 20732 2514 20760 2586
rect 20720 2508 20772 2514
rect 20720 2450 20772 2456
rect 21652 480 21680 3703
rect 22204 3505 22232 4218
rect 22296 4214 22324 4558
rect 23124 4554 23152 4966
rect 23296 4752 23348 4758
rect 23296 4694 23348 4700
rect 23204 4616 23256 4622
rect 23204 4558 23256 4564
rect 23112 4548 23164 4554
rect 23112 4490 23164 4496
rect 23216 4486 23244 4558
rect 23204 4480 23256 4486
rect 23204 4422 23256 4428
rect 23216 4282 23244 4422
rect 23204 4276 23256 4282
rect 23204 4218 23256 4224
rect 22284 4208 22336 4214
rect 22284 4150 22336 4156
rect 22650 4176 22706 4185
rect 22650 4111 22706 4120
rect 22664 3942 22692 4111
rect 23216 4078 23244 4218
rect 23204 4072 23256 4078
rect 23204 4014 23256 4020
rect 22652 3936 22704 3942
rect 23112 3936 23164 3942
rect 22652 3878 22704 3884
rect 23110 3904 23112 3913
rect 23164 3904 23166 3913
rect 23110 3839 23166 3848
rect 23216 3602 23244 4014
rect 23308 3738 23336 4694
rect 23296 3732 23348 3738
rect 23296 3674 23348 3680
rect 23400 3618 23428 5102
rect 24214 5063 24270 5072
rect 24032 5024 24084 5030
rect 24030 4992 24032 5001
rect 24084 4992 24086 5001
rect 24030 4927 24086 4936
rect 23662 4856 23718 4865
rect 24228 4826 24256 5063
rect 24872 5001 24900 5510
rect 25056 5370 25084 6967
rect 25332 6866 25360 8774
rect 25424 8634 25452 9114
rect 26528 8974 26556 9318
rect 26712 9110 26740 9318
rect 26700 9104 26752 9110
rect 26700 9046 26752 9052
rect 26516 8968 26568 8974
rect 26516 8910 26568 8916
rect 25412 8628 25464 8634
rect 25412 8570 25464 8576
rect 25424 8090 25452 8570
rect 26528 8294 26556 8910
rect 26516 8288 26568 8294
rect 26516 8230 26568 8236
rect 25412 8084 25464 8090
rect 25412 8026 25464 8032
rect 26528 7274 26556 8230
rect 26712 8090 26740 9046
rect 26884 8832 26936 8838
rect 26884 8774 26936 8780
rect 26896 8362 26924 8774
rect 27620 8628 27672 8634
rect 27620 8570 27672 8576
rect 26884 8356 26936 8362
rect 26884 8298 26936 8304
rect 26896 8090 26924 8298
rect 27632 8106 27660 8570
rect 29564 8537 29592 16918
rect 29748 16794 29776 18158
rect 29736 16788 29788 16794
rect 29736 16730 29788 16736
rect 29828 15904 29880 15910
rect 29828 15846 29880 15852
rect 29840 14618 29868 15846
rect 29828 14612 29880 14618
rect 29828 14554 29880 14560
rect 29932 14414 29960 18226
rect 31036 18154 31064 18566
rect 31024 18148 31076 18154
rect 31024 18090 31076 18096
rect 31668 18148 31720 18154
rect 31668 18090 31720 18096
rect 30288 18080 30340 18086
rect 30288 18022 30340 18028
rect 31680 18034 31708 18090
rect 32312 18080 32364 18086
rect 30300 17882 30328 18022
rect 31680 18006 31800 18034
rect 32312 18022 32364 18028
rect 30288 17876 30340 17882
rect 30288 17818 30340 17824
rect 30932 17740 30984 17746
rect 30932 17682 30984 17688
rect 30380 17536 30432 17542
rect 30380 17478 30432 17484
rect 30392 16794 30420 17478
rect 30944 17338 30972 17682
rect 30932 17332 30984 17338
rect 30932 17274 30984 17280
rect 31116 17128 31168 17134
rect 30654 17096 30710 17105
rect 31116 17070 31168 17076
rect 30654 17031 30710 17040
rect 30668 16998 30696 17031
rect 30656 16992 30708 16998
rect 30656 16934 30708 16940
rect 31128 16794 31156 17070
rect 30380 16788 30432 16794
rect 30380 16730 30432 16736
rect 31116 16788 31168 16794
rect 31116 16730 31168 16736
rect 30392 16114 30420 16730
rect 31772 16726 31800 18006
rect 31852 17536 31904 17542
rect 31852 17478 31904 17484
rect 31864 17202 31892 17478
rect 31852 17196 31904 17202
rect 31852 17138 31904 17144
rect 32128 16992 32180 16998
rect 32128 16934 32180 16940
rect 32140 16794 32168 16934
rect 32128 16788 32180 16794
rect 32128 16730 32180 16736
rect 31760 16720 31812 16726
rect 31760 16662 31812 16668
rect 32220 16720 32272 16726
rect 32220 16662 32272 16668
rect 30932 16652 30984 16658
rect 30932 16594 30984 16600
rect 31852 16652 31904 16658
rect 31852 16594 31904 16600
rect 30944 16182 30972 16594
rect 31574 16552 31630 16561
rect 31574 16487 31630 16496
rect 30932 16176 30984 16182
rect 30932 16118 30984 16124
rect 30380 16108 30432 16114
rect 30380 16050 30432 16056
rect 30194 15736 30250 15745
rect 30194 15671 30250 15680
rect 30562 15736 30618 15745
rect 30562 15671 30564 15680
rect 30208 14550 30236 15671
rect 30616 15671 30618 15680
rect 30564 15642 30616 15648
rect 30288 14952 30340 14958
rect 30288 14894 30340 14900
rect 30746 14920 30802 14929
rect 30300 14657 30328 14894
rect 30746 14855 30748 14864
rect 30800 14855 30802 14864
rect 30748 14826 30800 14832
rect 30286 14648 30342 14657
rect 30286 14583 30288 14592
rect 30340 14583 30342 14592
rect 30288 14554 30340 14560
rect 30196 14544 30248 14550
rect 30196 14486 30248 14492
rect 29920 14408 29972 14414
rect 29920 14350 29972 14356
rect 30208 14006 30236 14486
rect 30300 14074 30328 14554
rect 30472 14408 30524 14414
rect 30472 14350 30524 14356
rect 30484 14074 30512 14350
rect 30288 14068 30340 14074
rect 30288 14010 30340 14016
rect 30472 14068 30524 14074
rect 30472 14010 30524 14016
rect 30196 14000 30248 14006
rect 30196 13942 30248 13948
rect 30378 13832 30434 13841
rect 30378 13767 30434 13776
rect 29644 13184 29696 13190
rect 29644 13126 29696 13132
rect 30196 13184 30248 13190
rect 30196 13126 30248 13132
rect 29656 12782 29684 13126
rect 29736 12844 29788 12850
rect 29736 12786 29788 12792
rect 29644 12776 29696 12782
rect 29644 12718 29696 12724
rect 29656 10849 29684 12718
rect 29748 10985 29776 12786
rect 30102 11384 30158 11393
rect 30102 11319 30104 11328
rect 30156 11319 30158 11328
rect 30104 11290 30156 11296
rect 30012 11212 30064 11218
rect 30012 11154 30064 11160
rect 29734 10976 29790 10985
rect 29734 10911 29790 10920
rect 29642 10840 29698 10849
rect 29642 10775 29698 10784
rect 30024 10713 30052 11154
rect 30208 11150 30236 13126
rect 30392 12918 30420 13767
rect 30564 13388 30616 13394
rect 30564 13330 30616 13336
rect 30576 13190 30604 13330
rect 30564 13184 30616 13190
rect 30564 13126 30616 13132
rect 30576 12986 30604 13126
rect 31588 12986 31616 16487
rect 31864 16250 31892 16594
rect 32232 16250 32260 16662
rect 32324 16658 32352 18022
rect 32312 16652 32364 16658
rect 32312 16594 32364 16600
rect 32416 16538 32444 19110
rect 32600 18306 32628 20402
rect 32956 20256 33008 20262
rect 32956 20198 33008 20204
rect 33048 20256 33100 20262
rect 33048 20198 33100 20204
rect 32968 19802 32996 20198
rect 33060 20058 33088 20198
rect 33244 20058 33272 20402
rect 33336 20330 33364 20878
rect 33324 20324 33376 20330
rect 33324 20266 33376 20272
rect 33048 20052 33100 20058
rect 33048 19994 33100 20000
rect 33232 20052 33284 20058
rect 33232 19994 33284 20000
rect 32968 19774 33088 19802
rect 33060 19718 33088 19774
rect 33048 19712 33100 19718
rect 33048 19654 33100 19660
rect 33060 19394 33088 19654
rect 33888 19514 33916 21830
rect 34256 21486 34284 22374
rect 34518 22335 34574 22344
rect 34336 22228 34388 22234
rect 34336 22170 34388 22176
rect 34348 21690 34376 22170
rect 34428 22092 34480 22098
rect 34428 22034 34480 22040
rect 34336 21684 34388 21690
rect 34336 21626 34388 21632
rect 34244 21480 34296 21486
rect 34244 21422 34296 21428
rect 34244 21140 34296 21146
rect 34348 21128 34376 21626
rect 34440 21146 34468 22034
rect 34296 21100 34376 21128
rect 34428 21140 34480 21146
rect 34244 21082 34296 21088
rect 34428 21082 34480 21088
rect 34428 20256 34480 20262
rect 34428 20198 34480 20204
rect 34440 19514 34468 20198
rect 33876 19508 33928 19514
rect 33876 19450 33928 19456
rect 34428 19508 34480 19514
rect 34428 19450 34480 19456
rect 33060 19366 33272 19394
rect 32772 18828 32824 18834
rect 32772 18770 32824 18776
rect 32956 18828 33008 18834
rect 32956 18770 33008 18776
rect 32600 18278 32720 18306
rect 32324 16510 32444 16538
rect 31852 16244 31904 16250
rect 31852 16186 31904 16192
rect 32220 16244 32272 16250
rect 32220 16186 32272 16192
rect 32128 14952 32180 14958
rect 32128 14894 32180 14900
rect 31852 14816 31904 14822
rect 31852 14758 31904 14764
rect 31864 14657 31892 14758
rect 31850 14648 31906 14657
rect 31850 14583 31906 14592
rect 31852 14544 31904 14550
rect 31852 14486 31904 14492
rect 31864 14074 31892 14486
rect 32140 14074 32168 14894
rect 31852 14068 31904 14074
rect 31852 14010 31904 14016
rect 32128 14068 32180 14074
rect 32128 14010 32180 14016
rect 32140 13394 32168 14010
rect 32324 13569 32352 16510
rect 32404 15496 32456 15502
rect 32404 15438 32456 15444
rect 32416 14822 32444 15438
rect 32404 14816 32456 14822
rect 32404 14758 32456 14764
rect 32416 14090 32444 14758
rect 32588 14476 32640 14482
rect 32588 14418 32640 14424
rect 32600 14278 32628 14418
rect 32588 14272 32640 14278
rect 32588 14214 32640 14220
rect 32416 14074 32536 14090
rect 32416 14068 32548 14074
rect 32416 14062 32496 14068
rect 32310 13560 32366 13569
rect 32310 13495 32366 13504
rect 32128 13388 32180 13394
rect 32128 13330 32180 13336
rect 32140 12986 32168 13330
rect 30564 12980 30616 12986
rect 30564 12922 30616 12928
rect 31576 12980 31628 12986
rect 31576 12922 31628 12928
rect 32128 12980 32180 12986
rect 32128 12922 32180 12928
rect 30380 12912 30432 12918
rect 30380 12854 30432 12860
rect 31588 12782 31616 12922
rect 31576 12776 31628 12782
rect 31576 12718 31628 12724
rect 30380 12640 30432 12646
rect 30380 12582 30432 12588
rect 30392 12442 30420 12582
rect 30380 12436 30432 12442
rect 30380 12378 30432 12384
rect 30196 11144 30248 11150
rect 30392 11098 30420 12378
rect 32140 12374 32168 12922
rect 32416 12714 32444 14062
rect 32496 14010 32548 14016
rect 32600 13802 32628 14214
rect 32588 13796 32640 13802
rect 32588 13738 32640 13744
rect 32600 13530 32628 13738
rect 32588 13524 32640 13530
rect 32588 13466 32640 13472
rect 32404 12708 32456 12714
rect 32404 12650 32456 12656
rect 32416 12442 32444 12650
rect 32404 12436 32456 12442
rect 32404 12378 32456 12384
rect 32128 12368 32180 12374
rect 32128 12310 32180 12316
rect 31760 11348 31812 11354
rect 31760 11290 31812 11296
rect 30196 11086 30248 11092
rect 30300 11070 30420 11098
rect 30010 10704 30066 10713
rect 30010 10639 30066 10648
rect 29920 10600 29972 10606
rect 29920 10542 29972 10548
rect 29828 10124 29880 10130
rect 29828 10066 29880 10072
rect 29840 9722 29868 10066
rect 29828 9716 29880 9722
rect 29828 9658 29880 9664
rect 29932 9518 29960 10542
rect 30300 10538 30328 11070
rect 30288 10532 30340 10538
rect 30288 10474 30340 10480
rect 30300 10266 30328 10474
rect 31208 10464 31260 10470
rect 31208 10406 31260 10412
rect 30288 10260 30340 10266
rect 30288 10202 30340 10208
rect 30380 10260 30432 10266
rect 30380 10202 30432 10208
rect 30012 9920 30064 9926
rect 30012 9862 30064 9868
rect 29920 9512 29972 9518
rect 29920 9454 29972 9460
rect 29736 9444 29788 9450
rect 29736 9386 29788 9392
rect 29748 9178 29776 9386
rect 29736 9172 29788 9178
rect 29736 9114 29788 9120
rect 30024 9110 30052 9862
rect 30392 9738 30420 10202
rect 31220 10062 31248 10406
rect 31772 10282 31800 11290
rect 32128 11212 32180 11218
rect 32128 11154 32180 11160
rect 32140 11082 32168 11154
rect 32128 11076 32180 11082
rect 32128 11018 32180 11024
rect 32140 10810 32168 11018
rect 32128 10804 32180 10810
rect 32128 10746 32180 10752
rect 32310 10704 32366 10713
rect 32310 10639 32366 10648
rect 32324 10606 32352 10639
rect 32312 10600 32364 10606
rect 32312 10542 32364 10548
rect 32496 10464 32548 10470
rect 32496 10406 32548 10412
rect 31680 10266 31800 10282
rect 31668 10260 31800 10266
rect 31720 10254 31800 10260
rect 31668 10202 31720 10208
rect 32508 10130 32536 10406
rect 32496 10124 32548 10130
rect 32496 10066 32548 10072
rect 30564 10056 30616 10062
rect 30564 9998 30616 10004
rect 31208 10056 31260 10062
rect 31208 9998 31260 10004
rect 30300 9710 30420 9738
rect 30300 9178 30328 9710
rect 30576 9450 30604 9998
rect 32508 9722 32536 10066
rect 32496 9716 32548 9722
rect 32496 9658 32548 9664
rect 32496 9580 32548 9586
rect 32496 9522 32548 9528
rect 32312 9512 32364 9518
rect 32312 9454 32364 9460
rect 30564 9444 30616 9450
rect 30564 9386 30616 9392
rect 31024 9376 31076 9382
rect 31024 9318 31076 9324
rect 31116 9376 31168 9382
rect 31116 9318 31168 9324
rect 30288 9172 30340 9178
rect 30288 9114 30340 9120
rect 30012 9104 30064 9110
rect 30012 9046 30064 9052
rect 30024 8634 30052 9046
rect 30840 9036 30892 9042
rect 30840 8978 30892 8984
rect 30852 8634 30880 8978
rect 30012 8628 30064 8634
rect 30012 8570 30064 8576
rect 30840 8628 30892 8634
rect 30840 8570 30892 8576
rect 29550 8528 29606 8537
rect 31036 8498 31064 9318
rect 31128 8974 31156 9318
rect 32324 9178 32352 9454
rect 32312 9172 32364 9178
rect 32312 9114 32364 9120
rect 32402 9072 32458 9081
rect 32402 9007 32404 9016
rect 32456 9007 32458 9016
rect 32404 8978 32456 8984
rect 31116 8968 31168 8974
rect 31116 8910 31168 8916
rect 29550 8463 29606 8472
rect 31024 8492 31076 8498
rect 31024 8434 31076 8440
rect 31128 8294 31156 8910
rect 32508 8634 32536 9522
rect 32692 9178 32720 18278
rect 32784 18222 32812 18770
rect 32772 18216 32824 18222
rect 32772 18158 32824 18164
rect 32968 18154 32996 18770
rect 32956 18148 33008 18154
rect 32956 18090 33008 18096
rect 33140 18080 33192 18086
rect 33060 18028 33140 18034
rect 33060 18022 33192 18028
rect 33060 18006 33180 18022
rect 32864 17536 32916 17542
rect 32864 17478 32916 17484
rect 32876 17241 32904 17478
rect 32862 17232 32918 17241
rect 32772 17196 32824 17202
rect 32862 17167 32918 17176
rect 32772 17138 32824 17144
rect 32784 16658 32812 17138
rect 32772 16652 32824 16658
rect 32772 16594 32824 16600
rect 32864 16584 32916 16590
rect 32864 16526 32916 16532
rect 32876 15434 32904 16526
rect 33060 16250 33088 18006
rect 33140 17876 33192 17882
rect 33140 17818 33192 17824
rect 33152 16794 33180 17818
rect 33140 16788 33192 16794
rect 33140 16730 33192 16736
rect 33048 16244 33100 16250
rect 33048 16186 33100 16192
rect 32956 15632 33008 15638
rect 32956 15574 33008 15580
rect 32864 15428 32916 15434
rect 32864 15370 32916 15376
rect 32876 14550 32904 15370
rect 32968 14929 32996 15574
rect 33048 15360 33100 15366
rect 33100 15308 33180 15314
rect 33048 15302 33180 15308
rect 33060 15286 33180 15302
rect 33152 14958 33180 15286
rect 33140 14952 33192 14958
rect 32954 14920 33010 14929
rect 33140 14894 33192 14900
rect 32954 14855 33010 14864
rect 32968 14822 32996 14855
rect 32956 14816 33008 14822
rect 32956 14758 33008 14764
rect 32864 14544 32916 14550
rect 32864 14486 32916 14492
rect 32956 14272 33008 14278
rect 32956 14214 33008 14220
rect 32968 13462 32996 14214
rect 32956 13456 33008 13462
rect 32956 13398 33008 13404
rect 32968 12442 32996 13398
rect 32956 12436 33008 12442
rect 32956 12378 33008 12384
rect 33244 10266 33272 19366
rect 33508 19168 33560 19174
rect 34336 19168 34388 19174
rect 33508 19110 33560 19116
rect 34058 19136 34114 19145
rect 33324 17672 33376 17678
rect 33324 17614 33376 17620
rect 33336 17338 33364 17614
rect 33324 17332 33376 17338
rect 33324 17274 33376 17280
rect 33520 17241 33548 19110
rect 34336 19110 34388 19116
rect 34058 19071 34114 19080
rect 33690 18864 33746 18873
rect 33690 18799 33746 18808
rect 33704 18222 33732 18799
rect 34072 18630 34100 19071
rect 34244 18828 34296 18834
rect 34244 18770 34296 18776
rect 34060 18624 34112 18630
rect 34060 18566 34112 18572
rect 33692 18216 33744 18222
rect 33692 18158 33744 18164
rect 33704 17882 33732 18158
rect 33692 17876 33744 17882
rect 33692 17818 33744 17824
rect 34072 17746 34100 18566
rect 34256 18086 34284 18770
rect 34348 18154 34376 19110
rect 34428 18760 34480 18766
rect 34428 18702 34480 18708
rect 34336 18148 34388 18154
rect 34336 18090 34388 18096
rect 34244 18080 34296 18086
rect 34244 18022 34296 18028
rect 33600 17740 33652 17746
rect 33600 17682 33652 17688
rect 34060 17740 34112 17746
rect 34060 17682 34112 17688
rect 33612 17338 33640 17682
rect 34348 17678 34376 18090
rect 34336 17672 34388 17678
rect 34336 17614 34388 17620
rect 34060 17604 34112 17610
rect 34060 17546 34112 17552
rect 33600 17332 33652 17338
rect 33600 17274 33652 17280
rect 33506 17232 33562 17241
rect 33506 17167 33562 17176
rect 33784 17128 33836 17134
rect 33784 17070 33836 17076
rect 33796 16794 33824 17070
rect 33784 16788 33836 16794
rect 33784 16730 33836 16736
rect 33968 16788 34020 16794
rect 33968 16730 34020 16736
rect 33876 16584 33928 16590
rect 33876 16526 33928 16532
rect 33888 15994 33916 16526
rect 33980 16182 34008 16730
rect 34072 16726 34100 17546
rect 34348 17202 34376 17614
rect 34440 17338 34468 18702
rect 34428 17332 34480 17338
rect 34428 17274 34480 17280
rect 34336 17196 34388 17202
rect 34336 17138 34388 17144
rect 34060 16720 34112 16726
rect 34060 16662 34112 16668
rect 34336 16584 34388 16590
rect 34336 16526 34388 16532
rect 34348 16250 34376 16526
rect 34336 16244 34388 16250
rect 34336 16186 34388 16192
rect 33968 16176 34020 16182
rect 33968 16118 34020 16124
rect 33888 15966 34008 15994
rect 33980 15366 34008 15966
rect 34428 15904 34480 15910
rect 34428 15846 34480 15852
rect 34060 15564 34112 15570
rect 34060 15506 34112 15512
rect 33416 15360 33468 15366
rect 33416 15302 33468 15308
rect 33968 15360 34020 15366
rect 33968 15302 34020 15308
rect 33428 15026 33456 15302
rect 33980 15026 34008 15302
rect 34072 15094 34100 15506
rect 34440 15162 34468 15846
rect 34428 15156 34480 15162
rect 34428 15098 34480 15104
rect 34060 15088 34112 15094
rect 34060 15030 34112 15036
rect 33416 15020 33468 15026
rect 33416 14962 33468 14968
rect 33968 15020 34020 15026
rect 33968 14962 34020 14968
rect 33428 14618 33456 14962
rect 33600 14816 33652 14822
rect 33600 14758 33652 14764
rect 33416 14612 33468 14618
rect 33416 14554 33468 14560
rect 33612 12986 33640 14758
rect 34072 14618 34100 15030
rect 34060 14612 34112 14618
rect 34060 14554 34112 14560
rect 33692 14408 33744 14414
rect 33690 14376 33692 14385
rect 34428 14408 34480 14414
rect 33744 14376 33746 14385
rect 34428 14350 34480 14356
rect 33690 14311 33746 14320
rect 34440 13870 34468 14350
rect 34428 13864 34480 13870
rect 34428 13806 34480 13812
rect 34242 13560 34298 13569
rect 34242 13495 34298 13504
rect 33600 12980 33652 12986
rect 33600 12922 33652 12928
rect 33324 10464 33376 10470
rect 33324 10406 33376 10412
rect 33232 10260 33284 10266
rect 33232 10202 33284 10208
rect 33048 10124 33100 10130
rect 33048 10066 33100 10072
rect 32864 9920 32916 9926
rect 32864 9862 32916 9868
rect 32876 9450 32904 9862
rect 32864 9444 32916 9450
rect 32864 9386 32916 9392
rect 32956 9376 33008 9382
rect 32956 9318 33008 9324
rect 32680 9172 32732 9178
rect 32680 9114 32732 9120
rect 32496 8628 32548 8634
rect 32496 8570 32548 8576
rect 31116 8288 31168 8294
rect 31116 8230 31168 8236
rect 26700 8084 26752 8090
rect 26700 8026 26752 8032
rect 26884 8084 26936 8090
rect 26884 8026 26936 8032
rect 27540 8078 27660 8106
rect 31128 8090 31156 8230
rect 31116 8084 31168 8090
rect 26608 7744 26660 7750
rect 26608 7686 26660 7692
rect 26516 7268 26568 7274
rect 26516 7210 26568 7216
rect 26620 7002 26648 7686
rect 26896 7546 26924 8026
rect 27540 8022 27568 8078
rect 31116 8026 31168 8032
rect 26976 8016 27028 8022
rect 26976 7958 27028 7964
rect 27528 8016 27580 8022
rect 27528 7958 27580 7964
rect 26884 7540 26936 7546
rect 26884 7482 26936 7488
rect 26988 7342 27016 7958
rect 28540 7948 28592 7954
rect 28540 7890 28592 7896
rect 27160 7880 27212 7886
rect 27160 7822 27212 7828
rect 28080 7880 28132 7886
rect 28080 7822 28132 7828
rect 26976 7336 27028 7342
rect 26976 7278 27028 7284
rect 26988 7002 27016 7278
rect 25504 6996 25556 7002
rect 25504 6938 25556 6944
rect 26608 6996 26660 7002
rect 26608 6938 26660 6944
rect 26976 6996 27028 7002
rect 26976 6938 27028 6944
rect 25320 6860 25372 6866
rect 25320 6802 25372 6808
rect 25332 6458 25360 6802
rect 25412 6792 25464 6798
rect 25412 6734 25464 6740
rect 25320 6452 25372 6458
rect 25320 6394 25372 6400
rect 25424 6254 25452 6734
rect 25516 6458 25544 6938
rect 26976 6860 27028 6866
rect 26976 6802 27028 6808
rect 26608 6656 26660 6662
rect 26608 6598 26660 6604
rect 25504 6452 25556 6458
rect 25504 6394 25556 6400
rect 25412 6248 25464 6254
rect 25412 6190 25464 6196
rect 25424 5710 25452 6190
rect 25964 6112 26016 6118
rect 25964 6054 26016 6060
rect 26240 6112 26292 6118
rect 26240 6054 26292 6060
rect 25412 5704 25464 5710
rect 25976 5681 26004 6054
rect 25412 5646 25464 5652
rect 25962 5672 26018 5681
rect 25962 5607 26018 5616
rect 26252 5574 26280 6054
rect 26516 5908 26568 5914
rect 26516 5850 26568 5856
rect 26528 5817 26556 5850
rect 26514 5808 26570 5817
rect 26332 5772 26384 5778
rect 26514 5743 26570 5752
rect 26332 5714 26384 5720
rect 26240 5568 26292 5574
rect 26240 5510 26292 5516
rect 26252 5370 26280 5510
rect 25044 5364 25096 5370
rect 25044 5306 25096 5312
rect 26240 5364 26292 5370
rect 26240 5306 26292 5312
rect 25056 5166 25084 5306
rect 25778 5264 25834 5273
rect 25596 5228 25648 5234
rect 25778 5199 25834 5208
rect 25596 5170 25648 5176
rect 25044 5160 25096 5166
rect 25044 5102 25096 5108
rect 24858 4992 24914 5001
rect 24858 4927 24914 4936
rect 23662 4791 23718 4800
rect 24216 4820 24268 4826
rect 23676 4758 23704 4791
rect 24216 4762 24268 4768
rect 23664 4752 23716 4758
rect 23664 4694 23716 4700
rect 25608 4554 25636 5170
rect 25792 5098 25820 5199
rect 25780 5092 25832 5098
rect 25780 5034 25832 5040
rect 25596 4548 25648 4554
rect 25596 4490 25648 4496
rect 24768 4480 24820 4486
rect 24768 4422 24820 4428
rect 23572 4140 23624 4146
rect 23572 4082 23624 4088
rect 23480 3664 23532 3670
rect 23400 3612 23480 3618
rect 23400 3606 23532 3612
rect 23204 3596 23256 3602
rect 23400 3590 23520 3606
rect 23204 3538 23256 3544
rect 22560 3528 22612 3534
rect 22190 3496 22246 3505
rect 22560 3470 22612 3476
rect 22190 3431 22246 3440
rect 22468 3460 22520 3466
rect 22468 3402 22520 3408
rect 22480 3058 22508 3402
rect 22468 3052 22520 3058
rect 22468 2994 22520 3000
rect 22100 2916 22152 2922
rect 22100 2858 22152 2864
rect 21824 2848 21876 2854
rect 22112 2802 22140 2858
rect 21824 2790 21876 2796
rect 21836 1873 21864 2790
rect 22020 2774 22140 2802
rect 22020 2514 22048 2774
rect 22572 2650 22600 3470
rect 22652 3392 22704 3398
rect 22652 3334 22704 3340
rect 22742 3360 22798 3369
rect 22664 2990 22692 3334
rect 22742 3295 22798 3304
rect 22652 2984 22704 2990
rect 22652 2926 22704 2932
rect 22560 2644 22612 2650
rect 22560 2586 22612 2592
rect 22008 2508 22060 2514
rect 22008 2450 22060 2456
rect 21822 1864 21878 1873
rect 21822 1799 21878 1808
rect 22756 480 22784 3295
rect 23216 2990 23244 3538
rect 23584 3398 23612 4082
rect 24780 4078 24808 4422
rect 25608 4214 25636 4490
rect 25596 4208 25648 4214
rect 25594 4176 25596 4185
rect 25648 4176 25650 4185
rect 25594 4111 25650 4120
rect 24768 4072 24820 4078
rect 24768 4014 24820 4020
rect 25044 3936 25096 3942
rect 24950 3904 25006 3913
rect 25044 3878 25096 3884
rect 24950 3839 25006 3848
rect 24582 3496 24638 3505
rect 24582 3431 24638 3440
rect 23572 3392 23624 3398
rect 23572 3334 23624 3340
rect 23204 2984 23256 2990
rect 23204 2926 23256 2932
rect 23584 2922 23612 3334
rect 24596 3194 24624 3431
rect 24584 3188 24636 3194
rect 24584 3130 24636 3136
rect 23846 3088 23902 3097
rect 23846 3023 23902 3032
rect 23756 2984 23808 2990
rect 23756 2926 23808 2932
rect 23572 2916 23624 2922
rect 23572 2858 23624 2864
rect 23768 2650 23796 2926
rect 23756 2644 23808 2650
rect 23756 2586 23808 2592
rect 23860 480 23888 3023
rect 24596 2582 24624 3130
rect 24584 2576 24636 2582
rect 24584 2518 24636 2524
rect 24964 480 24992 3839
rect 25056 3670 25084 3878
rect 25044 3664 25096 3670
rect 25044 3606 25096 3612
rect 26344 3466 26372 5714
rect 26620 4078 26648 6598
rect 26988 6118 27016 6802
rect 27172 6730 27200 7822
rect 28092 7342 28120 7822
rect 28080 7336 28132 7342
rect 28080 7278 28132 7284
rect 27988 7200 28040 7206
rect 27988 7142 28040 7148
rect 27160 6724 27212 6730
rect 27160 6666 27212 6672
rect 27896 6724 27948 6730
rect 27896 6666 27948 6672
rect 27908 6390 27936 6666
rect 27896 6384 27948 6390
rect 27896 6326 27948 6332
rect 27620 6248 27672 6254
rect 27620 6190 27672 6196
rect 26976 6112 27028 6118
rect 26974 6080 26976 6089
rect 27028 6080 27030 6089
rect 26974 6015 27030 6024
rect 27632 5914 27660 6190
rect 27908 5914 27936 6326
rect 28000 6322 28028 7142
rect 28092 6798 28120 7278
rect 28552 7274 28580 7890
rect 29644 7744 29696 7750
rect 29644 7686 29696 7692
rect 32128 7744 32180 7750
rect 32128 7686 32180 7692
rect 28540 7268 28592 7274
rect 28540 7210 28592 7216
rect 28908 7200 28960 7206
rect 28908 7142 28960 7148
rect 28080 6792 28132 6798
rect 28080 6734 28132 6740
rect 27988 6316 28040 6322
rect 27988 6258 28040 6264
rect 28092 6118 28120 6734
rect 28080 6112 28132 6118
rect 28080 6054 28132 6060
rect 27620 5908 27672 5914
rect 27620 5850 27672 5856
rect 27896 5908 27948 5914
rect 27896 5850 27948 5856
rect 26700 5772 26752 5778
rect 26700 5714 26752 5720
rect 26712 5001 26740 5714
rect 26976 5704 27028 5710
rect 26976 5646 27028 5652
rect 27160 5704 27212 5710
rect 27160 5646 27212 5652
rect 26988 5302 27016 5646
rect 26976 5296 27028 5302
rect 26976 5238 27028 5244
rect 26884 5160 26936 5166
rect 26884 5102 26936 5108
rect 26698 4992 26754 5001
rect 26698 4927 26754 4936
rect 26712 4486 26740 4927
rect 26896 4865 26924 5102
rect 26882 4856 26938 4865
rect 26882 4791 26938 4800
rect 26700 4480 26752 4486
rect 26700 4422 26752 4428
rect 26712 4282 26740 4422
rect 26700 4276 26752 4282
rect 26700 4218 26752 4224
rect 26988 4214 27016 5238
rect 27172 4826 27200 5646
rect 27908 5234 27936 5850
rect 28092 5710 28120 6054
rect 28538 5944 28594 5953
rect 28538 5879 28594 5888
rect 28080 5704 28132 5710
rect 28080 5646 28132 5652
rect 27896 5228 27948 5234
rect 27896 5170 27948 5176
rect 28092 5030 28120 5646
rect 28080 5024 28132 5030
rect 28080 4966 28132 4972
rect 27160 4820 27212 4826
rect 27160 4762 27212 4768
rect 27804 4684 27856 4690
rect 27804 4626 27856 4632
rect 28356 4684 28408 4690
rect 28356 4626 28408 4632
rect 27448 4554 27660 4570
rect 27448 4548 27672 4554
rect 27448 4542 27620 4548
rect 26976 4208 27028 4214
rect 26976 4150 27028 4156
rect 26608 4072 26660 4078
rect 26608 4014 26660 4020
rect 26698 4040 26754 4049
rect 26620 3738 26648 4014
rect 26698 3975 26754 3984
rect 26712 3942 26740 3975
rect 26700 3936 26752 3942
rect 26700 3878 26752 3884
rect 26608 3732 26660 3738
rect 26608 3674 26660 3680
rect 26516 3596 26568 3602
rect 26516 3538 26568 3544
rect 26884 3596 26936 3602
rect 26884 3538 26936 3544
rect 26332 3460 26384 3466
rect 26332 3402 26384 3408
rect 26528 3194 26556 3538
rect 26056 3188 26108 3194
rect 26056 3130 26108 3136
rect 26516 3188 26568 3194
rect 26516 3130 26568 3136
rect 25688 2916 25740 2922
rect 25688 2858 25740 2864
rect 25700 2650 25728 2858
rect 25688 2644 25740 2650
rect 25688 2586 25740 2592
rect 26068 480 26096 3130
rect 26240 3120 26292 3126
rect 26240 3062 26292 3068
rect 26252 2650 26280 3062
rect 26896 2990 26924 3538
rect 27448 3466 27476 4542
rect 27620 4490 27672 4496
rect 27528 4480 27580 4486
rect 27528 4422 27580 4428
rect 27540 3534 27568 4422
rect 27816 4282 27844 4626
rect 27988 4616 28040 4622
rect 27988 4558 28040 4564
rect 27804 4276 27856 4282
rect 27804 4218 27856 4224
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 27436 3460 27488 3466
rect 27436 3402 27488 3408
rect 28000 3194 28028 4558
rect 28264 4072 28316 4078
rect 28264 4014 28316 4020
rect 28276 3738 28304 4014
rect 28368 3942 28396 4626
rect 28448 4480 28500 4486
rect 28448 4422 28500 4428
rect 28460 4214 28488 4422
rect 28448 4208 28500 4214
rect 28448 4150 28500 4156
rect 28356 3936 28408 3942
rect 28354 3904 28356 3913
rect 28408 3904 28410 3913
rect 28354 3839 28410 3848
rect 28552 3754 28580 5879
rect 28724 5840 28776 5846
rect 28724 5782 28776 5788
rect 28736 5370 28764 5782
rect 28724 5364 28776 5370
rect 28724 5306 28776 5312
rect 28264 3732 28316 3738
rect 28264 3674 28316 3680
rect 28368 3726 28580 3754
rect 28920 3738 28948 7142
rect 29656 6866 29684 7686
rect 32140 7410 32168 7686
rect 32128 7404 32180 7410
rect 32128 7346 32180 7352
rect 32508 7274 32536 8570
rect 32680 7880 32732 7886
rect 32678 7848 32680 7857
rect 32732 7848 32734 7857
rect 32678 7783 32734 7792
rect 32496 7268 32548 7274
rect 32496 7210 32548 7216
rect 32968 6866 32996 9318
rect 33060 8974 33088 10066
rect 33336 10062 33364 10406
rect 33784 10260 33836 10266
rect 33784 10202 33836 10208
rect 33324 10056 33376 10062
rect 33230 10024 33286 10033
rect 33324 9998 33376 10004
rect 33230 9959 33232 9968
rect 33284 9959 33286 9968
rect 33232 9930 33284 9936
rect 33796 9722 33824 10202
rect 33784 9716 33836 9722
rect 33784 9658 33836 9664
rect 33324 9376 33376 9382
rect 33324 9318 33376 9324
rect 33140 9172 33192 9178
rect 33140 9114 33192 9120
rect 33048 8968 33100 8974
rect 33048 8910 33100 8916
rect 33060 8634 33088 8910
rect 33048 8628 33100 8634
rect 33048 8570 33100 8576
rect 33152 8362 33180 9114
rect 33336 8974 33364 9318
rect 33796 9178 33824 9658
rect 33784 9172 33836 9178
rect 33784 9114 33836 9120
rect 33324 8968 33376 8974
rect 33324 8910 33376 8916
rect 33140 8356 33192 8362
rect 33140 8298 33192 8304
rect 33336 7857 33364 8910
rect 33600 8288 33652 8294
rect 33600 8230 33652 8236
rect 33968 8288 34020 8294
rect 33968 8230 34020 8236
rect 33508 7948 33560 7954
rect 33508 7890 33560 7896
rect 33322 7848 33378 7857
rect 33322 7783 33378 7792
rect 33520 7546 33548 7890
rect 33508 7540 33560 7546
rect 33508 7482 33560 7488
rect 33048 6996 33100 7002
rect 33048 6938 33100 6944
rect 29000 6860 29052 6866
rect 29000 6802 29052 6808
rect 29644 6860 29696 6866
rect 29644 6802 29696 6808
rect 32956 6860 33008 6866
rect 32956 6802 33008 6808
rect 29012 6458 29040 6802
rect 29644 6656 29696 6662
rect 29644 6598 29696 6604
rect 32864 6656 32916 6662
rect 32864 6598 32916 6604
rect 29000 6452 29052 6458
rect 29000 6394 29052 6400
rect 29012 6254 29040 6394
rect 29274 6352 29330 6361
rect 29274 6287 29330 6296
rect 29288 6254 29316 6287
rect 29000 6248 29052 6254
rect 29000 6190 29052 6196
rect 29276 6248 29328 6254
rect 29276 6190 29328 6196
rect 29460 6112 29512 6118
rect 29460 6054 29512 6060
rect 29274 5672 29330 5681
rect 29274 5607 29330 5616
rect 29000 5568 29052 5574
rect 29000 5510 29052 5516
rect 29012 5166 29040 5510
rect 29288 5166 29316 5607
rect 29472 5273 29500 6054
rect 29656 5846 29684 6598
rect 32876 6361 32904 6598
rect 33060 6458 33088 6938
rect 33520 6798 33548 7482
rect 33612 7002 33640 8230
rect 33980 7750 34008 8230
rect 33968 7744 34020 7750
rect 33968 7686 34020 7692
rect 33980 7206 34008 7686
rect 34256 7410 34284 13495
rect 34440 13326 34468 13806
rect 34428 13320 34480 13326
rect 34428 13262 34480 13268
rect 34440 12986 34468 13262
rect 34428 12980 34480 12986
rect 34428 12922 34480 12928
rect 34532 10713 34560 22335
rect 34624 21434 34652 23310
rect 34716 22234 34744 24908
rect 34796 24890 34848 24896
rect 34980 24676 35032 24682
rect 34980 24618 35032 24624
rect 34992 24410 35020 24618
rect 35360 24410 35388 31826
rect 35452 28801 35480 35566
rect 36188 35290 36216 39335
rect 37554 38312 37610 38321
rect 37554 38247 37610 38256
rect 36176 35284 36228 35290
rect 36176 35226 36228 35232
rect 36176 35148 36228 35154
rect 36176 35090 36228 35096
rect 35532 34944 35584 34950
rect 35532 34886 35584 34892
rect 35544 34542 35572 34886
rect 36188 34542 36216 35090
rect 37568 34746 37596 38247
rect 37556 34740 37608 34746
rect 37556 34682 37608 34688
rect 36268 34672 36320 34678
rect 36266 34640 36268 34649
rect 36320 34640 36322 34649
rect 36266 34575 36322 34584
rect 35532 34536 35584 34542
rect 35532 34478 35584 34484
rect 35900 34536 35952 34542
rect 35900 34478 35952 34484
rect 36176 34536 36228 34542
rect 37924 34536 37976 34542
rect 36176 34478 36228 34484
rect 37554 34504 37610 34513
rect 35912 34202 35940 34478
rect 35900 34196 35952 34202
rect 35900 34138 35952 34144
rect 35990 33688 36046 33697
rect 35990 33623 36046 33632
rect 35808 33380 35860 33386
rect 35808 33322 35860 33328
rect 35820 33114 35848 33322
rect 35808 33108 35860 33114
rect 35808 33050 35860 33056
rect 35806 32600 35862 32609
rect 35806 32535 35862 32544
rect 35622 31376 35678 31385
rect 35622 31311 35678 31320
rect 35438 28792 35494 28801
rect 35494 28750 35572 28778
rect 35636 28762 35664 31311
rect 35820 29866 35848 32535
rect 36004 32026 36032 33623
rect 35992 32020 36044 32026
rect 35992 31962 36044 31968
rect 35820 29850 35940 29866
rect 35820 29844 35952 29850
rect 35820 29838 35900 29844
rect 35900 29786 35952 29792
rect 35808 29708 35860 29714
rect 35808 29650 35860 29656
rect 35820 29186 35848 29650
rect 36084 29504 36136 29510
rect 36084 29446 36136 29452
rect 35820 29158 35940 29186
rect 35808 29028 35860 29034
rect 35808 28970 35860 28976
rect 35438 28727 35494 28736
rect 35440 28620 35492 28626
rect 35440 28562 35492 28568
rect 35452 27878 35480 28562
rect 35440 27872 35492 27878
rect 35440 27814 35492 27820
rect 34980 24404 35032 24410
rect 34980 24346 35032 24352
rect 35348 24404 35400 24410
rect 35348 24346 35400 24352
rect 35360 24290 35388 24346
rect 35268 24262 35388 24290
rect 34940 23964 35236 23984
rect 34996 23962 35020 23964
rect 35076 23962 35100 23964
rect 35156 23962 35180 23964
rect 35018 23910 35020 23962
rect 35082 23910 35094 23962
rect 35156 23910 35158 23962
rect 34996 23908 35020 23910
rect 35076 23908 35100 23910
rect 35156 23908 35180 23910
rect 34940 23888 35236 23908
rect 34796 23588 34848 23594
rect 34796 23530 34848 23536
rect 34808 22982 34836 23530
rect 34796 22976 34848 22982
rect 34796 22918 34848 22924
rect 34704 22228 34756 22234
rect 34704 22170 34756 22176
rect 34808 22114 34836 22918
rect 34940 22876 35236 22896
rect 34996 22874 35020 22876
rect 35076 22874 35100 22876
rect 35156 22874 35180 22876
rect 35018 22822 35020 22874
rect 35082 22822 35094 22874
rect 35156 22822 35158 22874
rect 34996 22820 35020 22822
rect 35076 22820 35100 22822
rect 35156 22820 35180 22822
rect 34940 22800 35236 22820
rect 35164 22568 35216 22574
rect 35164 22510 35216 22516
rect 35176 22438 35204 22510
rect 35164 22432 35216 22438
rect 35164 22374 35216 22380
rect 34808 22086 34838 22114
rect 34810 22030 34838 22086
rect 34796 22024 34848 22030
rect 34796 21966 34848 21972
rect 34808 21894 34836 21966
rect 34796 21888 34848 21894
rect 34796 21830 34848 21836
rect 34940 21788 35236 21808
rect 34996 21786 35020 21788
rect 35076 21786 35100 21788
rect 35156 21786 35180 21788
rect 35018 21734 35020 21786
rect 35082 21734 35094 21786
rect 35156 21734 35158 21786
rect 34996 21732 35020 21734
rect 35076 21732 35100 21734
rect 35156 21732 35180 21734
rect 34940 21712 35236 21732
rect 34888 21480 34940 21486
rect 34624 21406 34836 21434
rect 34888 21422 34940 21428
rect 34612 21140 34664 21146
rect 34612 21082 34664 21088
rect 34624 20602 34652 21082
rect 34612 20596 34664 20602
rect 34612 20538 34664 20544
rect 34624 20330 34652 20538
rect 34612 20324 34664 20330
rect 34612 20266 34664 20272
rect 34612 19848 34664 19854
rect 34664 19796 34744 19802
rect 34612 19790 34744 19796
rect 34624 19774 34744 19790
rect 34612 19712 34664 19718
rect 34612 19654 34664 19660
rect 34624 19378 34652 19654
rect 34612 19372 34664 19378
rect 34612 19314 34664 19320
rect 34716 19242 34744 19774
rect 34704 19236 34756 19242
rect 34704 19178 34756 19184
rect 34716 18970 34744 19178
rect 34704 18964 34756 18970
rect 34704 18906 34756 18912
rect 34808 18850 34836 21406
rect 34900 21146 34928 21422
rect 34888 21140 34940 21146
rect 34888 21082 34940 21088
rect 34940 20700 35236 20720
rect 34996 20698 35020 20700
rect 35076 20698 35100 20700
rect 35156 20698 35180 20700
rect 35018 20646 35020 20698
rect 35082 20646 35094 20698
rect 35156 20646 35158 20698
rect 34996 20644 35020 20646
rect 35076 20644 35100 20646
rect 35156 20644 35180 20646
rect 34940 20624 35236 20644
rect 34940 19612 35236 19632
rect 34996 19610 35020 19612
rect 35076 19610 35100 19612
rect 35156 19610 35180 19612
rect 35018 19558 35020 19610
rect 35082 19558 35094 19610
rect 35156 19558 35158 19610
rect 34996 19556 35020 19558
rect 35076 19556 35100 19558
rect 35156 19556 35180 19558
rect 34940 19536 35236 19556
rect 35164 19372 35216 19378
rect 35164 19314 35216 19320
rect 35176 18970 35204 19314
rect 35164 18964 35216 18970
rect 35164 18906 35216 18912
rect 34716 18822 34836 18850
rect 34612 18352 34664 18358
rect 34612 18294 34664 18300
rect 34624 17202 34652 18294
rect 34612 17196 34664 17202
rect 34612 17138 34664 17144
rect 34612 16652 34664 16658
rect 34612 16594 34664 16600
rect 34624 16250 34652 16594
rect 34612 16244 34664 16250
rect 34612 16186 34664 16192
rect 34624 15706 34652 16186
rect 34612 15700 34664 15706
rect 34612 15642 34664 15648
rect 34612 15564 34664 15570
rect 34612 15506 34664 15512
rect 34624 14822 34652 15506
rect 34612 14816 34664 14822
rect 34612 14758 34664 14764
rect 34624 14482 34652 14758
rect 34612 14476 34664 14482
rect 34612 14418 34664 14424
rect 34624 14074 34652 14418
rect 34612 14068 34664 14074
rect 34612 14010 34664 14016
rect 34624 13530 34652 14010
rect 34612 13524 34664 13530
rect 34612 13466 34664 13472
rect 34610 13424 34666 13433
rect 34610 13359 34666 13368
rect 34624 12764 34652 13359
rect 34716 12866 34744 18822
rect 34940 18524 35236 18544
rect 34996 18522 35020 18524
rect 35076 18522 35100 18524
rect 35156 18522 35180 18524
rect 35018 18470 35020 18522
rect 35082 18470 35094 18522
rect 35156 18470 35158 18522
rect 34996 18468 35020 18470
rect 35076 18468 35100 18470
rect 35156 18468 35180 18470
rect 34940 18448 35236 18468
rect 35072 18148 35124 18154
rect 35072 18090 35124 18096
rect 35084 17882 35112 18090
rect 35072 17876 35124 17882
rect 35072 17818 35124 17824
rect 34940 17436 35236 17456
rect 34996 17434 35020 17436
rect 35076 17434 35100 17436
rect 35156 17434 35180 17436
rect 35018 17382 35020 17434
rect 35082 17382 35094 17434
rect 35156 17382 35158 17434
rect 34996 17380 35020 17382
rect 35076 17380 35100 17382
rect 35156 17380 35180 17382
rect 34940 17360 35236 17380
rect 34978 17232 35034 17241
rect 34978 17167 35034 17176
rect 34992 17134 35020 17167
rect 34980 17128 35032 17134
rect 34980 17070 35032 17076
rect 34940 16348 35236 16368
rect 34996 16346 35020 16348
rect 35076 16346 35100 16348
rect 35156 16346 35180 16348
rect 35018 16294 35020 16346
rect 35082 16294 35094 16346
rect 35156 16294 35158 16346
rect 34996 16292 35020 16294
rect 35076 16292 35100 16294
rect 35156 16292 35180 16294
rect 34940 16272 35236 16292
rect 35268 16130 35296 24262
rect 35348 22976 35400 22982
rect 35348 22918 35400 22924
rect 35360 22574 35388 22918
rect 35348 22568 35400 22574
rect 35348 22510 35400 22516
rect 35452 22114 35480 27814
rect 35544 27418 35572 28750
rect 35624 28756 35676 28762
rect 35624 28698 35676 28704
rect 35820 27962 35848 28970
rect 35912 28914 35940 29158
rect 35912 28886 36032 28914
rect 36004 28422 36032 28886
rect 36096 28762 36124 29446
rect 36084 28756 36136 28762
rect 36084 28698 36136 28704
rect 35992 28416 36044 28422
rect 35992 28358 36044 28364
rect 36004 28121 36032 28358
rect 35990 28112 36046 28121
rect 35990 28047 36046 28056
rect 35820 27934 35940 27962
rect 35808 27872 35860 27878
rect 35808 27814 35860 27820
rect 35716 27464 35768 27470
rect 35544 27390 35664 27418
rect 35716 27406 35768 27412
rect 35532 27328 35584 27334
rect 35532 27270 35584 27276
rect 35544 26926 35572 27270
rect 35532 26920 35584 26926
rect 35532 26862 35584 26868
rect 35544 26586 35572 26862
rect 35636 26858 35664 27390
rect 35624 26852 35676 26858
rect 35624 26794 35676 26800
rect 35622 26752 35678 26761
rect 35622 26687 35678 26696
rect 35532 26580 35584 26586
rect 35532 26522 35584 26528
rect 35636 25673 35664 26687
rect 35622 25664 35678 25673
rect 35622 25599 35678 25608
rect 35624 25288 35676 25294
rect 35624 25230 35676 25236
rect 35636 24018 35664 25230
rect 35728 24682 35756 27406
rect 35820 26897 35848 27814
rect 35912 27130 35940 27934
rect 35900 27124 35952 27130
rect 35900 27066 35952 27072
rect 35806 26888 35862 26897
rect 35806 26823 35862 26832
rect 35808 26784 35860 26790
rect 35808 26726 35860 26732
rect 35716 24676 35768 24682
rect 35716 24618 35768 24624
rect 35820 24290 35848 26726
rect 35912 24818 35940 27066
rect 36084 25968 36136 25974
rect 36084 25910 36136 25916
rect 35900 24812 35952 24818
rect 35900 24754 35952 24760
rect 35716 24268 35768 24274
rect 35820 24262 35940 24290
rect 35716 24210 35768 24216
rect 35544 23990 35664 24018
rect 35544 23526 35572 23990
rect 35624 23724 35676 23730
rect 35624 23666 35676 23672
rect 35532 23520 35584 23526
rect 35532 23462 35584 23468
rect 35544 22234 35572 23462
rect 35636 23322 35664 23666
rect 35728 23662 35756 24210
rect 35808 24200 35860 24206
rect 35808 24142 35860 24148
rect 35820 23866 35848 24142
rect 35808 23860 35860 23866
rect 35808 23802 35860 23808
rect 35912 23746 35940 24262
rect 35820 23718 35940 23746
rect 35716 23656 35768 23662
rect 35716 23598 35768 23604
rect 35820 23338 35848 23718
rect 35624 23316 35676 23322
rect 35624 23258 35676 23264
rect 35728 23310 35848 23338
rect 35636 22574 35664 23258
rect 35624 22568 35676 22574
rect 35624 22510 35676 22516
rect 35728 22409 35756 23310
rect 35808 23180 35860 23186
rect 35808 23122 35860 23128
rect 35820 22438 35848 23122
rect 35808 22432 35860 22438
rect 35714 22400 35770 22409
rect 35808 22374 35860 22380
rect 35714 22335 35770 22344
rect 35532 22228 35584 22234
rect 35532 22170 35584 22176
rect 35716 22228 35768 22234
rect 35716 22170 35768 22176
rect 35452 22086 35572 22114
rect 35544 21842 35572 22086
rect 35728 21978 35756 22170
rect 35820 22098 35848 22374
rect 35808 22092 35860 22098
rect 35808 22034 35860 22040
rect 35900 22024 35952 22030
rect 35728 21972 35900 21978
rect 35728 21966 35952 21972
rect 35728 21950 35940 21966
rect 35360 21814 35572 21842
rect 35360 21570 35388 21814
rect 36096 21672 36124 25910
rect 36188 23798 36216 34478
rect 37924 34478 37976 34484
rect 37554 34439 37610 34448
rect 36268 34128 36320 34134
rect 36268 34070 36320 34076
rect 36280 33658 36308 34070
rect 36268 33652 36320 33658
rect 36268 33594 36320 33600
rect 36268 32972 36320 32978
rect 36268 32914 36320 32920
rect 36280 32570 36308 32914
rect 37568 32570 37596 34439
rect 36268 32564 36320 32570
rect 36268 32506 36320 32512
rect 37556 32564 37608 32570
rect 37556 32506 37608 32512
rect 37372 32360 37424 32366
rect 37372 32302 37424 32308
rect 36820 31748 36872 31754
rect 36820 31690 36872 31696
rect 36268 31680 36320 31686
rect 36268 31622 36320 31628
rect 36280 31482 36308 31622
rect 36832 31482 36860 31690
rect 36268 31476 36320 31482
rect 36268 31418 36320 31424
rect 36820 31476 36872 31482
rect 36820 31418 36872 31424
rect 36268 29572 36320 29578
rect 36268 29514 36320 29520
rect 36280 29306 36308 29514
rect 36268 29300 36320 29306
rect 36268 29242 36320 29248
rect 36636 28620 36688 28626
rect 36636 28562 36688 28568
rect 36648 28014 36676 28562
rect 36636 28008 36688 28014
rect 36634 27976 36636 27985
rect 36688 27976 36690 27985
rect 36634 27911 36690 27920
rect 36268 25288 36320 25294
rect 36266 25256 36268 25265
rect 36320 25256 36322 25265
rect 36266 25191 36322 25200
rect 36268 24200 36320 24206
rect 36268 24142 36320 24148
rect 36176 23792 36228 23798
rect 36176 23734 36228 23740
rect 36004 21644 36124 21672
rect 35360 21542 35480 21570
rect 35348 21412 35400 21418
rect 35348 21354 35400 21360
rect 35360 21146 35388 21354
rect 35348 21140 35400 21146
rect 35348 21082 35400 21088
rect 35360 20466 35388 21082
rect 35348 20460 35400 20466
rect 35348 20402 35400 20408
rect 35360 20058 35388 20402
rect 35348 20052 35400 20058
rect 35348 19994 35400 20000
rect 35348 19712 35400 19718
rect 35348 19654 35400 19660
rect 35360 19174 35388 19654
rect 35348 19168 35400 19174
rect 35348 19110 35400 19116
rect 35348 16992 35400 16998
rect 35348 16934 35400 16940
rect 35360 16794 35388 16934
rect 35348 16788 35400 16794
rect 35348 16730 35400 16736
rect 34808 16102 35296 16130
rect 34808 12968 34836 16102
rect 35348 15428 35400 15434
rect 35348 15370 35400 15376
rect 35256 15360 35308 15366
rect 35256 15302 35308 15308
rect 34940 15260 35236 15280
rect 34996 15258 35020 15260
rect 35076 15258 35100 15260
rect 35156 15258 35180 15260
rect 35018 15206 35020 15258
rect 35082 15206 35094 15258
rect 35156 15206 35158 15258
rect 34996 15204 35020 15206
rect 35076 15204 35100 15206
rect 35156 15204 35180 15206
rect 34940 15184 35236 15204
rect 35268 14958 35296 15302
rect 35256 14952 35308 14958
rect 35256 14894 35308 14900
rect 35256 14816 35308 14822
rect 35360 14770 35388 15370
rect 35308 14764 35388 14770
rect 35256 14758 35388 14764
rect 35268 14742 35388 14758
rect 34940 14172 35236 14192
rect 34996 14170 35020 14172
rect 35076 14170 35100 14172
rect 35156 14170 35180 14172
rect 35018 14118 35020 14170
rect 35082 14118 35094 14170
rect 35156 14118 35158 14170
rect 34996 14116 35020 14118
rect 35076 14116 35100 14118
rect 35156 14116 35180 14118
rect 34940 14096 35236 14116
rect 34940 13084 35236 13104
rect 34996 13082 35020 13084
rect 35076 13082 35100 13084
rect 35156 13082 35180 13084
rect 35018 13030 35020 13082
rect 35082 13030 35094 13082
rect 35156 13030 35158 13082
rect 34996 13028 35020 13030
rect 35076 13028 35100 13030
rect 35156 13028 35180 13030
rect 34940 13008 35236 13028
rect 34808 12940 35204 12968
rect 34716 12838 34836 12866
rect 34624 12736 34744 12764
rect 34518 10704 34574 10713
rect 34518 10639 34574 10648
rect 34716 10305 34744 12736
rect 34702 10296 34758 10305
rect 34702 10231 34758 10240
rect 34808 10146 34836 12838
rect 35176 12186 35204 12940
rect 35268 12442 35296 14742
rect 35348 13456 35400 13462
rect 35348 13398 35400 13404
rect 35360 12782 35388 13398
rect 35348 12776 35400 12782
rect 35348 12718 35400 12724
rect 35360 12442 35388 12718
rect 35256 12436 35308 12442
rect 35256 12378 35308 12384
rect 35348 12436 35400 12442
rect 35348 12378 35400 12384
rect 35176 12158 35296 12186
rect 34940 11996 35236 12016
rect 34996 11994 35020 11996
rect 35076 11994 35100 11996
rect 35156 11994 35180 11996
rect 35018 11942 35020 11994
rect 35082 11942 35094 11994
rect 35156 11942 35158 11994
rect 34996 11940 35020 11942
rect 35076 11940 35100 11942
rect 35156 11940 35180 11942
rect 34940 11920 35236 11940
rect 34940 10908 35236 10928
rect 34996 10906 35020 10908
rect 35076 10906 35100 10908
rect 35156 10906 35180 10908
rect 35018 10854 35020 10906
rect 35082 10854 35094 10906
rect 35156 10854 35158 10906
rect 34996 10852 35020 10854
rect 35076 10852 35100 10854
rect 35156 10852 35180 10854
rect 34940 10832 35236 10852
rect 35164 10464 35216 10470
rect 35164 10406 35216 10412
rect 34612 10124 34664 10130
rect 34612 10066 34664 10072
rect 34716 10118 34836 10146
rect 35176 10130 35204 10406
rect 35164 10124 35216 10130
rect 34520 9512 34572 9518
rect 34520 9454 34572 9460
rect 34428 9444 34480 9450
rect 34428 9386 34480 9392
rect 34336 8356 34388 8362
rect 34336 8298 34388 8304
rect 34348 7834 34376 8298
rect 34440 8090 34468 9386
rect 34428 8084 34480 8090
rect 34428 8026 34480 8032
rect 34532 8022 34560 9454
rect 34624 9382 34652 10066
rect 34612 9376 34664 9382
rect 34612 9318 34664 9324
rect 34612 8968 34664 8974
rect 34612 8910 34664 8916
rect 34520 8016 34572 8022
rect 34520 7958 34572 7964
rect 34348 7806 34560 7834
rect 34244 7404 34296 7410
rect 34244 7346 34296 7352
rect 33968 7200 34020 7206
rect 33968 7142 34020 7148
rect 33600 6996 33652 7002
rect 33600 6938 33652 6944
rect 33600 6860 33652 6866
rect 33600 6802 33652 6808
rect 33508 6792 33560 6798
rect 33508 6734 33560 6740
rect 33520 6458 33548 6734
rect 33612 6458 33640 6802
rect 33048 6452 33100 6458
rect 33048 6394 33100 6400
rect 33508 6452 33560 6458
rect 33508 6394 33560 6400
rect 33600 6452 33652 6458
rect 33600 6394 33652 6400
rect 32862 6352 32918 6361
rect 32862 6287 32918 6296
rect 29736 6180 29788 6186
rect 29736 6122 29788 6128
rect 29644 5840 29696 5846
rect 29644 5782 29696 5788
rect 29458 5264 29514 5273
rect 29458 5199 29514 5208
rect 29000 5160 29052 5166
rect 29000 5102 29052 5108
rect 29276 5160 29328 5166
rect 29276 5102 29328 5108
rect 29276 5024 29328 5030
rect 29276 4966 29328 4972
rect 29460 5024 29512 5030
rect 29460 4966 29512 4972
rect 29288 4622 29316 4966
rect 29368 4684 29420 4690
rect 29368 4626 29420 4632
rect 29276 4616 29328 4622
rect 29276 4558 29328 4564
rect 29288 4146 29316 4558
rect 29276 4140 29328 4146
rect 29276 4082 29328 4088
rect 29380 3738 29408 4626
rect 29472 4049 29500 4966
rect 29644 4140 29696 4146
rect 29644 4082 29696 4088
rect 29458 4040 29514 4049
rect 29458 3975 29514 3984
rect 28632 3732 28684 3738
rect 27620 3188 27672 3194
rect 27620 3130 27672 3136
rect 27988 3188 28040 3194
rect 27988 3130 28040 3136
rect 27250 3088 27306 3097
rect 27250 3023 27306 3032
rect 26608 2984 26660 2990
rect 26608 2926 26660 2932
rect 26884 2984 26936 2990
rect 26884 2926 26936 2932
rect 26620 2854 26648 2926
rect 26608 2848 26660 2854
rect 26608 2790 26660 2796
rect 26620 2650 26648 2790
rect 26240 2644 26292 2650
rect 26240 2586 26292 2592
rect 26608 2644 26660 2650
rect 26608 2586 26660 2592
rect 27264 480 27292 3023
rect 27632 2666 27660 3130
rect 27540 2638 27660 2666
rect 27540 2582 27568 2638
rect 27528 2576 27580 2582
rect 27528 2518 27580 2524
rect 28368 480 28396 3726
rect 28632 3674 28684 3680
rect 28908 3732 28960 3738
rect 28908 3674 28960 3680
rect 29368 3732 29420 3738
rect 29368 3674 29420 3680
rect 28448 3528 28500 3534
rect 28446 3496 28448 3505
rect 28500 3496 28502 3505
rect 28446 3431 28502 3440
rect 28644 3126 28672 3674
rect 29380 3534 29408 3674
rect 29656 3602 29684 4082
rect 29748 3942 29776 6122
rect 30288 6112 30340 6118
rect 30288 6054 30340 6060
rect 30300 5914 30328 6054
rect 30746 5944 30802 5953
rect 30288 5908 30340 5914
rect 30746 5879 30748 5888
rect 30288 5850 30340 5856
rect 30800 5879 30802 5888
rect 30748 5850 30800 5856
rect 30104 5568 30156 5574
rect 30104 5510 30156 5516
rect 29736 3936 29788 3942
rect 29736 3878 29788 3884
rect 29920 3936 29972 3942
rect 29920 3878 29972 3884
rect 29644 3596 29696 3602
rect 29644 3538 29696 3544
rect 28724 3528 28776 3534
rect 28724 3470 28776 3476
rect 29368 3528 29420 3534
rect 29368 3470 29420 3476
rect 28632 3120 28684 3126
rect 28632 3062 28684 3068
rect 28736 2938 28764 3470
rect 28908 3188 28960 3194
rect 28908 3130 28960 3136
rect 28644 2910 28764 2938
rect 28644 2650 28672 2910
rect 28632 2644 28684 2650
rect 28632 2586 28684 2592
rect 28920 2378 28948 3130
rect 29550 2952 29606 2961
rect 29656 2922 29684 3538
rect 29748 3058 29776 3878
rect 29932 3777 29960 3878
rect 29918 3768 29974 3777
rect 29918 3703 29974 3712
rect 30116 3346 30144 5510
rect 30196 5024 30248 5030
rect 30194 4992 30196 5001
rect 30248 4992 30250 5001
rect 30194 4927 30250 4936
rect 30300 4826 30328 5850
rect 31942 5808 31998 5817
rect 30840 5772 30892 5778
rect 31942 5743 31998 5752
rect 30840 5714 30892 5720
rect 30654 5400 30710 5409
rect 30654 5335 30710 5344
rect 30564 5024 30616 5030
rect 30564 4966 30616 4972
rect 30288 4820 30340 4826
rect 30288 4762 30340 4768
rect 30300 4146 30328 4762
rect 30380 4480 30432 4486
rect 30380 4422 30432 4428
rect 30288 4140 30340 4146
rect 30288 4082 30340 4088
rect 30300 3670 30328 4082
rect 30392 4078 30420 4422
rect 30380 4072 30432 4078
rect 30380 4014 30432 4020
rect 30472 3936 30524 3942
rect 30472 3878 30524 3884
rect 30484 3670 30512 3878
rect 30576 3738 30604 4966
rect 30564 3732 30616 3738
rect 30564 3674 30616 3680
rect 30288 3664 30340 3670
rect 30472 3664 30524 3670
rect 30288 3606 30340 3612
rect 30470 3632 30472 3641
rect 30524 3632 30526 3641
rect 30668 3618 30696 5335
rect 30852 5030 30880 5714
rect 31208 5568 31260 5574
rect 31208 5510 31260 5516
rect 31760 5568 31812 5574
rect 31760 5510 31812 5516
rect 31220 5370 31248 5510
rect 31208 5364 31260 5370
rect 31208 5306 31260 5312
rect 30840 5024 30892 5030
rect 30840 4966 30892 4972
rect 30470 3567 30526 3576
rect 30576 3590 30696 3618
rect 30484 3541 30512 3567
rect 30196 3392 30248 3398
rect 30116 3340 30196 3346
rect 30116 3334 30248 3340
rect 30116 3318 30236 3334
rect 30116 3058 30144 3318
rect 29736 3052 29788 3058
rect 29736 2994 29788 3000
rect 30104 3052 30156 3058
rect 30156 3012 30236 3040
rect 30104 2994 30156 3000
rect 29550 2887 29606 2896
rect 29644 2916 29696 2922
rect 29564 2854 29592 2887
rect 29644 2858 29696 2864
rect 29552 2848 29604 2854
rect 29552 2790 29604 2796
rect 29656 2514 29684 2858
rect 30208 2582 30236 3012
rect 30196 2576 30248 2582
rect 30196 2518 30248 2524
rect 29644 2508 29696 2514
rect 29644 2450 29696 2456
rect 28908 2372 28960 2378
rect 28908 2314 28960 2320
rect 29458 2136 29514 2145
rect 29458 2071 29514 2080
rect 29472 480 29500 2071
rect 30576 480 30604 3590
rect 30852 3097 30880 4966
rect 31220 4146 31248 5306
rect 31772 5234 31800 5510
rect 31760 5228 31812 5234
rect 31760 5170 31812 5176
rect 31668 5024 31720 5030
rect 31668 4966 31720 4972
rect 31574 4584 31630 4593
rect 31574 4519 31630 4528
rect 31208 4140 31260 4146
rect 31208 4082 31260 4088
rect 31116 4072 31168 4078
rect 31116 4014 31168 4020
rect 31024 3936 31076 3942
rect 31024 3878 31076 3884
rect 30932 3392 30984 3398
rect 30930 3360 30932 3369
rect 30984 3360 30986 3369
rect 30930 3295 30986 3304
rect 31036 3194 31064 3878
rect 31024 3188 31076 3194
rect 31024 3130 31076 3136
rect 30838 3088 30894 3097
rect 30838 3023 30894 3032
rect 31128 2990 31156 4014
rect 31588 3924 31616 4519
rect 31680 4078 31708 4966
rect 31668 4072 31720 4078
rect 31668 4014 31720 4020
rect 31588 3896 31708 3924
rect 31576 3732 31628 3738
rect 31576 3674 31628 3680
rect 31588 3058 31616 3674
rect 31576 3052 31628 3058
rect 31576 2994 31628 3000
rect 31116 2984 31168 2990
rect 31116 2926 31168 2932
rect 30656 2916 30708 2922
rect 30656 2858 30708 2864
rect 30668 2689 30696 2858
rect 31588 2825 31616 2994
rect 31574 2816 31630 2825
rect 31574 2751 31630 2760
rect 30654 2680 30710 2689
rect 30654 2615 30710 2624
rect 31680 480 31708 3896
rect 31956 3602 31984 5743
rect 32036 5704 32088 5710
rect 32036 5646 32088 5652
rect 32048 5166 32076 5646
rect 32310 5264 32366 5273
rect 32128 5228 32180 5234
rect 32310 5199 32312 5208
rect 32128 5170 32180 5176
rect 32364 5199 32366 5208
rect 32312 5170 32364 5176
rect 32036 5160 32088 5166
rect 32036 5102 32088 5108
rect 32048 4758 32076 5102
rect 32140 4826 32168 5170
rect 32772 5024 32824 5030
rect 32772 4966 32824 4972
rect 32784 4826 32812 4966
rect 32128 4820 32180 4826
rect 32128 4762 32180 4768
rect 32772 4820 32824 4826
rect 32772 4762 32824 4768
rect 32036 4752 32088 4758
rect 32036 4694 32088 4700
rect 32496 4684 32548 4690
rect 32496 4626 32548 4632
rect 33048 4684 33100 4690
rect 33048 4626 33100 4632
rect 32508 4078 32536 4626
rect 32770 4312 32826 4321
rect 32770 4247 32826 4256
rect 32496 4072 32548 4078
rect 32496 4014 32548 4020
rect 32036 3936 32088 3942
rect 32036 3878 32088 3884
rect 32310 3904 32366 3913
rect 32048 3777 32076 3878
rect 32310 3839 32366 3848
rect 32034 3768 32090 3777
rect 32324 3738 32352 3839
rect 32508 3738 32536 4014
rect 32034 3703 32036 3712
rect 32088 3703 32090 3712
rect 32312 3732 32364 3738
rect 32036 3674 32088 3680
rect 32312 3674 32364 3680
rect 32496 3732 32548 3738
rect 32496 3674 32548 3680
rect 31944 3596 31996 3602
rect 31944 3538 31996 3544
rect 31956 3194 31984 3538
rect 31944 3188 31996 3194
rect 31944 3130 31996 3136
rect 32048 3058 32076 3674
rect 32036 3052 32088 3058
rect 32036 2994 32088 3000
rect 32784 480 32812 4247
rect 33060 4146 33088 4626
rect 33980 4622 34008 7142
rect 34256 4826 34284 7346
rect 34532 7206 34560 7806
rect 34520 7200 34572 7206
rect 34520 7142 34572 7148
rect 34624 5273 34652 8910
rect 34716 6361 34744 10118
rect 35164 10066 35216 10072
rect 34796 10056 34848 10062
rect 34796 9998 34848 10004
rect 34808 9450 34836 9998
rect 34940 9820 35236 9840
rect 34996 9818 35020 9820
rect 35076 9818 35100 9820
rect 35156 9818 35180 9820
rect 35018 9766 35020 9818
rect 35082 9766 35094 9818
rect 35156 9766 35158 9818
rect 34996 9764 35020 9766
rect 35076 9764 35100 9766
rect 35156 9764 35180 9766
rect 34940 9744 35236 9764
rect 34888 9512 34940 9518
rect 34888 9454 34940 9460
rect 34796 9444 34848 9450
rect 34796 9386 34848 9392
rect 34900 9382 34928 9454
rect 34888 9376 34940 9382
rect 34808 9324 34888 9330
rect 34808 9318 34940 9324
rect 34808 9302 34928 9318
rect 34808 8838 34836 9302
rect 34796 8832 34848 8838
rect 34796 8774 34848 8780
rect 34808 8362 34836 8774
rect 34940 8732 35236 8752
rect 34996 8730 35020 8732
rect 35076 8730 35100 8732
rect 35156 8730 35180 8732
rect 35018 8678 35020 8730
rect 35082 8678 35094 8730
rect 35156 8678 35158 8730
rect 34996 8676 35020 8678
rect 35076 8676 35100 8678
rect 35156 8676 35180 8678
rect 34940 8656 35236 8676
rect 35164 8424 35216 8430
rect 35164 8366 35216 8372
rect 34796 8356 34848 8362
rect 34796 8298 34848 8304
rect 35176 8090 35204 8366
rect 35268 8265 35296 12158
rect 35360 11898 35388 12378
rect 35348 11892 35400 11898
rect 35348 11834 35400 11840
rect 35346 11792 35402 11801
rect 35346 11727 35402 11736
rect 35254 8256 35310 8265
rect 35254 8191 35310 8200
rect 35164 8084 35216 8090
rect 35164 8026 35216 8032
rect 35256 7948 35308 7954
rect 35256 7890 35308 7896
rect 34796 7812 34848 7818
rect 34796 7754 34848 7760
rect 34808 7002 34836 7754
rect 34940 7644 35236 7664
rect 34996 7642 35020 7644
rect 35076 7642 35100 7644
rect 35156 7642 35180 7644
rect 35018 7590 35020 7642
rect 35082 7590 35094 7642
rect 35156 7590 35158 7642
rect 34996 7588 35020 7590
rect 35076 7588 35100 7590
rect 35156 7588 35180 7590
rect 34940 7568 35236 7588
rect 35164 7404 35216 7410
rect 35164 7346 35216 7352
rect 35072 7200 35124 7206
rect 35070 7168 35072 7177
rect 35124 7168 35126 7177
rect 35070 7103 35126 7112
rect 34796 6996 34848 7002
rect 34796 6938 34848 6944
rect 35176 6934 35204 7346
rect 35268 7342 35296 7890
rect 35256 7336 35308 7342
rect 35256 7278 35308 7284
rect 35164 6928 35216 6934
rect 35164 6870 35216 6876
rect 34940 6556 35236 6576
rect 34996 6554 35020 6556
rect 35076 6554 35100 6556
rect 35156 6554 35180 6556
rect 35018 6502 35020 6554
rect 35082 6502 35094 6554
rect 35156 6502 35158 6554
rect 34996 6500 35020 6502
rect 35076 6500 35100 6502
rect 35156 6500 35180 6502
rect 34940 6480 35236 6500
rect 34702 6352 34758 6361
rect 34702 6287 34758 6296
rect 34940 5468 35236 5488
rect 34996 5466 35020 5468
rect 35076 5466 35100 5468
rect 35156 5466 35180 5468
rect 35018 5414 35020 5466
rect 35082 5414 35094 5466
rect 35156 5414 35158 5466
rect 34996 5412 35020 5414
rect 35076 5412 35100 5414
rect 35156 5412 35180 5414
rect 34940 5392 35236 5412
rect 34610 5264 34666 5273
rect 34610 5199 34666 5208
rect 34520 5024 34572 5030
rect 34520 4966 34572 4972
rect 34244 4820 34296 4826
rect 34244 4762 34296 4768
rect 34244 4684 34296 4690
rect 34244 4626 34296 4632
rect 33968 4616 34020 4622
rect 33968 4558 34020 4564
rect 33048 4140 33100 4146
rect 33048 4082 33100 4088
rect 33980 3942 34008 4558
rect 34256 3942 34284 4626
rect 33600 3936 33652 3942
rect 33600 3878 33652 3884
rect 33968 3936 34020 3942
rect 33968 3878 34020 3884
rect 34244 3936 34296 3942
rect 34244 3878 34296 3884
rect 33140 3664 33192 3670
rect 33138 3632 33140 3641
rect 33192 3632 33194 3641
rect 33138 3567 33194 3576
rect 33612 3398 33640 3878
rect 34060 3596 34112 3602
rect 34060 3538 34112 3544
rect 33600 3392 33652 3398
rect 33600 3334 33652 3340
rect 32954 3088 33010 3097
rect 32954 3023 32956 3032
rect 33008 3023 33010 3032
rect 32956 2994 33008 3000
rect 33612 2854 33640 3334
rect 33600 2848 33652 2854
rect 33600 2790 33652 2796
rect 33612 2514 33640 2790
rect 34072 2650 34100 3538
rect 34242 3360 34298 3369
rect 34242 3295 34298 3304
rect 34256 3194 34284 3295
rect 34532 3194 34560 4966
rect 34624 4826 34652 5199
rect 34612 4820 34664 4826
rect 34612 4762 34664 4768
rect 34940 4380 35236 4400
rect 34996 4378 35020 4380
rect 35076 4378 35100 4380
rect 35156 4378 35180 4380
rect 35018 4326 35020 4378
rect 35082 4326 35094 4378
rect 35156 4326 35158 4378
rect 34996 4324 35020 4326
rect 35076 4324 35100 4326
rect 35156 4324 35180 4326
rect 34940 4304 35236 4324
rect 34612 3936 34664 3942
rect 34612 3878 34664 3884
rect 34624 3738 34652 3878
rect 34612 3732 34664 3738
rect 34612 3674 34664 3680
rect 34940 3292 35236 3312
rect 34996 3290 35020 3292
rect 35076 3290 35100 3292
rect 35156 3290 35180 3292
rect 35018 3238 35020 3290
rect 35082 3238 35094 3290
rect 35156 3238 35158 3290
rect 34996 3236 35020 3238
rect 35076 3236 35100 3238
rect 35156 3236 35180 3238
rect 34940 3216 35236 3236
rect 34244 3188 34296 3194
rect 34244 3130 34296 3136
rect 34520 3188 34572 3194
rect 34520 3130 34572 3136
rect 35162 3088 35218 3097
rect 35162 3023 35218 3032
rect 34888 2848 34940 2854
rect 34794 2816 34850 2825
rect 34888 2790 34940 2796
rect 34794 2751 34850 2760
rect 34808 2650 34836 2751
rect 34060 2644 34112 2650
rect 34060 2586 34112 2592
rect 34796 2644 34848 2650
rect 34796 2586 34848 2592
rect 34808 2514 34836 2586
rect 34900 2553 34928 2790
rect 35176 2650 35204 3023
rect 35164 2644 35216 2650
rect 35164 2586 35216 2592
rect 34886 2544 34942 2553
rect 33600 2508 33652 2514
rect 33600 2450 33652 2456
rect 34796 2508 34848 2514
rect 34886 2479 34942 2488
rect 34796 2450 34848 2456
rect 35176 2446 35204 2586
rect 35164 2440 35216 2446
rect 35164 2382 35216 2388
rect 34940 2204 35236 2224
rect 34996 2202 35020 2204
rect 35076 2202 35100 2204
rect 35156 2202 35180 2204
rect 35018 2150 35020 2202
rect 35082 2150 35094 2202
rect 35156 2150 35158 2202
rect 34996 2148 35020 2150
rect 35076 2148 35100 2150
rect 35156 2148 35180 2150
rect 34940 2128 35236 2148
rect 34978 2000 35034 2009
rect 34978 1935 35034 1944
rect 33874 1864 33930 1873
rect 33874 1799 33930 1808
rect 33888 480 33916 1799
rect 34992 480 35020 1935
rect 35268 649 35296 7278
rect 35360 4049 35388 11727
rect 35452 8838 35480 21542
rect 35624 21480 35676 21486
rect 35624 21422 35676 21428
rect 35532 19916 35584 19922
rect 35532 19858 35584 19864
rect 35544 19378 35572 19858
rect 35532 19372 35584 19378
rect 35532 19314 35584 19320
rect 35636 19281 35664 21422
rect 35806 21312 35862 21321
rect 35806 21247 35862 21256
rect 35820 21146 35848 21247
rect 35808 21140 35860 21146
rect 35808 21082 35860 21088
rect 35716 20936 35768 20942
rect 35716 20878 35768 20884
rect 35820 20890 35848 21082
rect 35728 20534 35756 20878
rect 35820 20862 35940 20890
rect 35912 20602 35940 20862
rect 35900 20596 35952 20602
rect 35900 20538 35952 20544
rect 35716 20528 35768 20534
rect 36004 20482 36032 21644
rect 36188 21486 36216 23734
rect 36280 23526 36308 24142
rect 36268 23520 36320 23526
rect 36268 23462 36320 23468
rect 36280 22778 36308 23462
rect 36728 23316 36780 23322
rect 36728 23258 36780 23264
rect 36268 22772 36320 22778
rect 36268 22714 36320 22720
rect 36740 22234 36768 23258
rect 36728 22228 36780 22234
rect 36728 22170 36780 22176
rect 37384 22114 37412 32302
rect 36268 22092 36320 22098
rect 37384 22086 37504 22114
rect 36268 22034 36320 22040
rect 36280 21690 36308 22034
rect 36268 21684 36320 21690
rect 36268 21626 36320 21632
rect 36176 21480 36228 21486
rect 36176 21422 36228 21428
rect 36280 20942 36308 21626
rect 37372 21344 37424 21350
rect 37370 21312 37372 21321
rect 37424 21312 37426 21321
rect 37370 21247 37426 21256
rect 37186 21176 37242 21185
rect 37186 21111 37242 21120
rect 36268 20936 36320 20942
rect 36268 20878 36320 20884
rect 36084 20800 36136 20806
rect 36084 20742 36136 20748
rect 35716 20470 35768 20476
rect 35820 20454 36032 20482
rect 35714 19952 35770 19961
rect 35714 19887 35770 19896
rect 35622 19272 35678 19281
rect 35622 19207 35678 19216
rect 35728 18850 35756 19887
rect 35544 18822 35756 18850
rect 35544 16182 35572 18822
rect 35716 18760 35768 18766
rect 35716 18702 35768 18708
rect 35728 17882 35756 18702
rect 35820 17898 35848 20454
rect 35992 19168 36044 19174
rect 35992 19110 36044 19116
rect 36004 18426 36032 19110
rect 35992 18420 36044 18426
rect 35992 18362 36044 18368
rect 35716 17876 35768 17882
rect 35820 17870 36032 17898
rect 35716 17818 35768 17824
rect 35806 17776 35862 17785
rect 35806 17711 35862 17720
rect 35624 17196 35676 17202
rect 35624 17138 35676 17144
rect 35636 16794 35664 17138
rect 35624 16788 35676 16794
rect 35624 16730 35676 16736
rect 35820 16658 35848 17711
rect 35808 16652 35860 16658
rect 35808 16594 35860 16600
rect 35624 16584 35676 16590
rect 35624 16526 35676 16532
rect 35636 16250 35664 16526
rect 35820 16266 35848 16594
rect 35820 16250 35940 16266
rect 35624 16244 35676 16250
rect 35820 16244 35952 16250
rect 35820 16238 35900 16244
rect 35624 16186 35676 16192
rect 35900 16186 35952 16192
rect 35532 16176 35584 16182
rect 36004 16130 36032 17870
rect 35532 16118 35584 16124
rect 35820 16102 36032 16130
rect 35624 15496 35676 15502
rect 35624 15438 35676 15444
rect 35532 15020 35584 15026
rect 35532 14962 35584 14968
rect 35544 14618 35572 14962
rect 35636 14822 35664 15438
rect 35624 14816 35676 14822
rect 35624 14758 35676 14764
rect 35532 14612 35584 14618
rect 35532 14554 35584 14560
rect 35530 14240 35586 14249
rect 35530 14175 35586 14184
rect 35544 12753 35572 14175
rect 35636 13802 35664 14758
rect 35624 13796 35676 13802
rect 35624 13738 35676 13744
rect 35636 13530 35664 13738
rect 35624 13524 35676 13530
rect 35624 13466 35676 13472
rect 35820 13433 35848 16102
rect 35992 15360 36044 15366
rect 35992 15302 36044 15308
rect 36004 14385 36032 15302
rect 35990 14376 36046 14385
rect 35990 14311 36046 14320
rect 35806 13424 35862 13433
rect 35806 13359 35862 13368
rect 35806 13152 35862 13161
rect 35806 13087 35862 13096
rect 35530 12744 35586 12753
rect 35530 12679 35586 12688
rect 35716 12708 35768 12714
rect 35716 12650 35768 12656
rect 35622 12472 35678 12481
rect 35622 12407 35678 12416
rect 35532 11008 35584 11014
rect 35532 10950 35584 10956
rect 35544 10606 35572 10950
rect 35532 10600 35584 10606
rect 35532 10542 35584 10548
rect 35544 10266 35572 10542
rect 35532 10260 35584 10266
rect 35532 10202 35584 10208
rect 35440 8832 35492 8838
rect 35440 8774 35492 8780
rect 35440 7744 35492 7750
rect 35440 7686 35492 7692
rect 35452 7002 35480 7686
rect 35440 6996 35492 7002
rect 35440 6938 35492 6944
rect 35452 5914 35480 6938
rect 35544 6798 35572 10202
rect 35636 8537 35664 12407
rect 35728 12238 35756 12650
rect 35716 12232 35768 12238
rect 35820 12209 35848 13087
rect 36004 12238 36032 14311
rect 36096 12481 36124 20742
rect 36280 20602 36308 20878
rect 36268 20596 36320 20602
rect 36268 20538 36320 20544
rect 37200 19310 37228 21111
rect 37476 20874 37504 22086
rect 37464 20868 37516 20874
rect 37464 20810 37516 20816
rect 37936 20505 37964 34478
rect 37922 20496 37978 20505
rect 37922 20431 37978 20440
rect 37188 19304 37240 19310
rect 37188 19246 37240 19252
rect 36268 19168 36320 19174
rect 36266 19136 36268 19145
rect 36820 19168 36872 19174
rect 36320 19136 36322 19145
rect 36820 19110 36872 19116
rect 36266 19071 36322 19080
rect 36832 18873 36860 19110
rect 36818 18864 36874 18873
rect 36818 18799 36874 18808
rect 37094 18864 37150 18873
rect 37094 18799 37150 18808
rect 36820 18692 36872 18698
rect 36820 18634 36872 18640
rect 36832 18426 36860 18634
rect 36820 18420 36872 18426
rect 36820 18362 36872 18368
rect 37108 17338 37136 18799
rect 37096 17332 37148 17338
rect 37096 17274 37148 17280
rect 37108 17134 37136 17274
rect 37096 17128 37148 17134
rect 37096 17070 37148 17076
rect 36452 16992 36504 16998
rect 36452 16934 36504 16940
rect 36176 16448 36228 16454
rect 36176 16390 36228 16396
rect 36188 15366 36216 16390
rect 36176 15360 36228 15366
rect 36176 15302 36228 15308
rect 36464 14618 36492 16934
rect 37094 15464 37150 15473
rect 37094 15399 37150 15408
rect 37108 15162 37136 15399
rect 37096 15156 37148 15162
rect 37096 15098 37148 15104
rect 37108 14958 37136 15098
rect 37096 14952 37148 14958
rect 37096 14894 37148 14900
rect 36636 14816 36688 14822
rect 36636 14758 36688 14764
rect 36452 14612 36504 14618
rect 36452 14554 36504 14560
rect 36648 13841 36676 14758
rect 36634 13832 36690 13841
rect 36634 13767 36690 13776
rect 36820 13388 36872 13394
rect 36820 13330 36872 13336
rect 36832 12986 36860 13330
rect 36820 12980 36872 12986
rect 36820 12922 36872 12928
rect 36082 12472 36138 12481
rect 36082 12407 36138 12416
rect 35992 12232 36044 12238
rect 35716 12174 35768 12180
rect 35806 12200 35862 12209
rect 35728 11762 35756 12174
rect 35992 12174 36044 12180
rect 35806 12135 35862 12144
rect 35806 12064 35862 12073
rect 35806 11999 35862 12008
rect 35716 11756 35768 11762
rect 35716 11698 35768 11704
rect 35820 10248 35848 11999
rect 36004 11898 36032 12174
rect 36820 12096 36872 12102
rect 36820 12038 36872 12044
rect 35992 11892 36044 11898
rect 35992 11834 36044 11840
rect 36832 10810 36860 12038
rect 36820 10804 36872 10810
rect 36820 10746 36872 10752
rect 35728 10220 35848 10248
rect 35728 8974 35756 10220
rect 35808 10124 35860 10130
rect 35808 10066 35860 10072
rect 35716 8968 35768 8974
rect 35716 8910 35768 8916
rect 35716 8832 35768 8838
rect 35716 8774 35768 8780
rect 35622 8528 35678 8537
rect 35622 8463 35678 8472
rect 35622 8256 35678 8265
rect 35622 8191 35678 8200
rect 35636 7449 35664 8191
rect 35622 7440 35678 7449
rect 35622 7375 35678 7384
rect 35624 6860 35676 6866
rect 35624 6802 35676 6808
rect 35532 6792 35584 6798
rect 35532 6734 35584 6740
rect 35544 6390 35572 6734
rect 35636 6458 35664 6802
rect 35624 6452 35676 6458
rect 35624 6394 35676 6400
rect 35532 6384 35584 6390
rect 35532 6326 35584 6332
rect 35440 5908 35492 5914
rect 35440 5850 35492 5856
rect 35728 5137 35756 8774
rect 35820 8634 35848 10066
rect 35990 10024 36046 10033
rect 35990 9959 36046 9968
rect 36004 9178 36032 9959
rect 36268 9376 36320 9382
rect 36268 9318 36320 9324
rect 36820 9376 36872 9382
rect 36820 9318 36872 9324
rect 37096 9376 37148 9382
rect 37096 9318 37148 9324
rect 35992 9172 36044 9178
rect 35992 9114 36044 9120
rect 35808 8628 35860 8634
rect 35808 8570 35860 8576
rect 35820 7818 35848 8570
rect 36004 8090 36032 9114
rect 36280 8974 36308 9318
rect 36268 8968 36320 8974
rect 36268 8910 36320 8916
rect 36280 8430 36308 8910
rect 36832 8634 36860 9318
rect 37108 9042 37136 9318
rect 37096 9036 37148 9042
rect 37096 8978 37148 8984
rect 37108 8634 37136 8978
rect 36820 8628 36872 8634
rect 36820 8570 36872 8576
rect 37096 8628 37148 8634
rect 37096 8570 37148 8576
rect 36268 8424 36320 8430
rect 36268 8366 36320 8372
rect 35992 8084 36044 8090
rect 35992 8026 36044 8032
rect 35990 7984 36046 7993
rect 35990 7919 36046 7928
rect 35808 7812 35860 7818
rect 35808 7754 35860 7760
rect 35808 7404 35860 7410
rect 35808 7346 35860 7352
rect 35820 6662 35848 7346
rect 35808 6656 35860 6662
rect 35808 6598 35860 6604
rect 35900 6656 35952 6662
rect 35900 6598 35952 6604
rect 35912 5522 35940 6598
rect 35820 5494 35940 5522
rect 35714 5128 35770 5137
rect 35714 5063 35770 5072
rect 35346 4040 35402 4049
rect 35346 3975 35402 3984
rect 35440 3596 35492 3602
rect 35440 3538 35492 3544
rect 35348 3392 35400 3398
rect 35348 3334 35400 3340
rect 35360 3058 35388 3334
rect 35452 3058 35480 3538
rect 35348 3052 35400 3058
rect 35348 2994 35400 3000
rect 35440 3052 35492 3058
rect 35440 2994 35492 3000
rect 35360 2650 35388 2994
rect 35348 2644 35400 2650
rect 35348 2586 35400 2592
rect 35820 1737 35848 5494
rect 36004 3913 36032 7919
rect 37278 7848 37334 7857
rect 37278 7783 37334 7792
rect 37292 7546 37320 7783
rect 37280 7540 37332 7546
rect 37280 7482 37332 7488
rect 36176 7336 36228 7342
rect 36176 7278 36228 7284
rect 36188 6662 36216 7278
rect 37278 7168 37334 7177
rect 37278 7103 37334 7112
rect 36176 6656 36228 6662
rect 36176 6598 36228 6604
rect 35990 3904 36046 3913
rect 35990 3839 36046 3848
rect 37186 2952 37242 2961
rect 37292 2922 37320 7103
rect 39394 3904 39450 3913
rect 39394 3839 39450 3848
rect 37186 2887 37242 2896
rect 37280 2916 37332 2922
rect 37002 2680 37058 2689
rect 37002 2615 37004 2624
rect 37056 2615 37058 2624
rect 37004 2586 37056 2592
rect 36082 2544 36138 2553
rect 36082 2479 36138 2488
rect 35806 1728 35862 1737
rect 35806 1663 35862 1672
rect 35254 640 35310 649
rect 35254 575 35310 584
rect 36096 480 36124 2479
rect 37200 480 37228 2887
rect 37280 2858 37332 2864
rect 38292 2916 38344 2922
rect 38292 2858 38344 2864
rect 38304 480 38332 2858
rect 39408 480 39436 3839
rect 570 0 626 480
rect 1674 0 1730 480
rect 2778 0 2834 480
rect 3882 0 3938 480
rect 4986 0 5042 480
rect 6090 0 6146 480
rect 7194 0 7250 480
rect 8298 0 8354 480
rect 9402 0 9458 480
rect 10506 0 10562 480
rect 11610 0 11666 480
rect 12714 0 12770 480
rect 13910 0 13966 480
rect 15014 0 15070 480
rect 16118 0 16174 480
rect 17222 0 17278 480
rect 18326 0 18382 480
rect 19430 0 19486 480
rect 20534 0 20590 480
rect 21638 0 21694 480
rect 22742 0 22798 480
rect 23846 0 23902 480
rect 24950 0 25006 480
rect 26054 0 26110 480
rect 27250 0 27306 480
rect 28354 0 28410 480
rect 29458 0 29514 480
rect 30562 0 30618 480
rect 31666 0 31722 480
rect 32770 0 32826 480
rect 33874 0 33930 480
rect 34978 0 35034 480
rect 36082 0 36138 480
rect 37186 0 37242 480
rect 38290 0 38346 480
rect 39394 0 39450 480
<< via2 >>
rect 36174 39344 36230 39400
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 35622 37032 35678 37088
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 33874 36080 33930 36136
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 27986 33224 28042 33280
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 32034 34620 32036 34640
rect 32036 34620 32088 34640
rect 32088 34620 32090 34640
rect 32034 34584 32090 34620
rect 29826 33088 29882 33144
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 31850 33224 31906 33280
rect 30562 31340 30618 31376
rect 33506 33088 33562 33144
rect 30562 31320 30564 31340
rect 30564 31320 30616 31340
rect 30616 31320 30618 31340
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 34940 33754 34996 33756
rect 35020 33754 35076 33756
rect 35100 33754 35156 33756
rect 35180 33754 35236 33756
rect 34940 33702 34966 33754
rect 34966 33702 34996 33754
rect 35020 33702 35030 33754
rect 35030 33702 35076 33754
rect 35100 33702 35146 33754
rect 35146 33702 35156 33754
rect 35180 33702 35210 33754
rect 35210 33702 35236 33754
rect 34940 33700 34996 33702
rect 35020 33700 35076 33702
rect 35100 33700 35156 33702
rect 35180 33700 35236 33702
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 23294 26288 23350 26344
rect 21822 23976 21878 24032
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 21178 23296 21234 23352
rect 24398 25200 24454 25256
rect 24122 24012 24124 24032
rect 24124 24012 24176 24032
rect 24176 24012 24178 24032
rect 24122 23976 24178 24012
rect 26422 26288 26478 26344
rect 26698 25200 26754 25256
rect 26606 24520 26662 24576
rect 23754 23316 23810 23352
rect 23754 23296 23756 23316
rect 23756 23296 23808 23316
rect 23808 23296 23810 23316
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 21546 23024 21602 23080
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 23846 23060 23848 23080
rect 23848 23060 23900 23080
rect 23900 23060 23902 23080
rect 23846 23024 23902 23060
rect 30654 30232 30710 30288
rect 28722 26732 28724 26752
rect 28724 26732 28776 26752
rect 28776 26732 28778 26752
rect 28722 26696 28778 26732
rect 27158 23296 27214 23352
rect 25870 22636 25926 22672
rect 25870 22616 25872 22636
rect 25872 22616 25924 22636
rect 25924 22616 25926 22636
rect 25778 22208 25834 22264
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 21362 20712 21418 20768
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 3422 20032 3478 20088
rect 23754 20712 23810 20768
rect 22742 20168 22798 20224
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 26054 21936 26110 21992
rect 24122 21292 24124 21312
rect 24124 21292 24176 21312
rect 24176 21292 24178 21312
rect 24122 21256 24178 21292
rect 24674 20168 24730 20224
rect 25042 20204 25044 20224
rect 25044 20204 25096 20224
rect 25096 20204 25098 20224
rect 25042 20168 25098 20204
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 3422 18128 3478 18184
rect 18694 18148 18750 18184
rect 18694 18128 18696 18148
rect 18696 18128 18748 18148
rect 18748 18128 18750 18148
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 5814 15680 5870 15736
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 7838 15816 7894 15872
rect 7746 15680 7802 15736
rect 10138 15972 10194 16008
rect 10138 15952 10140 15972
rect 10140 15952 10192 15972
rect 10192 15952 10194 15972
rect 10046 15816 10102 15872
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 5170 14048 5226 14104
rect 5170 13948 5172 13968
rect 5172 13948 5224 13968
rect 5224 13948 5226 13968
rect 5170 13912 5226 13948
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 7378 14048 7434 14104
rect 7286 13912 7342 13968
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 13542 17076 13544 17096
rect 13544 17076 13596 17096
rect 13596 17076 13598 17096
rect 13542 17040 13598 17076
rect 10782 14864 10838 14920
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 9954 12588 9956 12608
rect 9956 12588 10008 12608
rect 10008 12588 10010 12608
rect 9954 12552 10010 12588
rect 10966 11192 11022 11248
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 2226 6704 2282 6760
rect 2410 5888 2466 5944
rect 3974 6840 4030 6896
rect 2778 6704 2834 6760
rect 3514 6704 3570 6760
rect 7194 8628 7250 8664
rect 7194 8608 7196 8628
rect 7196 8608 7248 8628
rect 7248 8608 7250 8628
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 5170 6704 5226 6760
rect 4434 5888 4490 5944
rect 2410 3440 2466 3496
rect 570 2760 626 2816
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 4342 5092 4398 5128
rect 4342 5072 4344 5092
rect 4344 5072 4396 5092
rect 4396 5072 4398 5092
rect 3974 4664 4030 4720
rect 3882 4528 3938 4584
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 4434 3440 4490 3496
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 4986 4120 5042 4176
rect 4618 3032 4674 3088
rect 4066 2760 4122 2816
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 5630 6160 5686 6216
rect 5446 6060 5448 6080
rect 5448 6060 5500 6080
rect 5500 6060 5502 6080
rect 5446 6024 5502 6060
rect 5446 5228 5502 5264
rect 5446 5208 5448 5228
rect 5448 5208 5500 5228
rect 5500 5208 5502 5228
rect 5998 6704 6054 6760
rect 6826 5888 6882 5944
rect 7562 6024 7618 6080
rect 8390 6196 8392 6216
rect 8392 6196 8444 6216
rect 8444 6196 8446 6216
rect 8390 6160 8446 6196
rect 7286 5616 7342 5672
rect 6826 5344 6882 5400
rect 5630 4664 5686 4720
rect 5998 4548 6054 4584
rect 5998 4528 6000 4548
rect 6000 4528 6052 4548
rect 6052 4528 6054 4548
rect 6182 4276 6238 4312
rect 6182 4256 6184 4276
rect 6184 4256 6236 4276
rect 6236 4256 6238 4276
rect 8022 5072 8078 5128
rect 8114 4800 8170 4856
rect 7102 4120 7158 4176
rect 6826 3884 6828 3904
rect 6828 3884 6880 3904
rect 6880 3884 6882 3904
rect 6826 3848 6882 3884
rect 5538 3440 5594 3496
rect 7010 3440 7066 3496
rect 6090 2760 6146 2816
rect 8574 5344 8630 5400
rect 8482 4684 8538 4720
rect 8482 4664 8484 4684
rect 8484 4664 8536 4684
rect 8536 4664 8538 4684
rect 8482 3848 8538 3904
rect 9126 4428 9128 4448
rect 9128 4428 9180 4448
rect 9180 4428 9182 4448
rect 9126 4392 9182 4428
rect 9034 3032 9090 3088
rect 8942 2932 8944 2952
rect 8944 2932 8996 2952
rect 8996 2932 8998 2952
rect 8942 2896 8998 2932
rect 8666 2760 8722 2816
rect 7102 1808 7158 1864
rect 7194 1400 7250 1456
rect 9218 2388 9220 2408
rect 9220 2388 9272 2408
rect 9272 2388 9274 2408
rect 9218 2352 9274 2388
rect 9678 5888 9734 5944
rect 9494 3984 9550 4040
rect 9678 3732 9734 3768
rect 9678 3712 9680 3732
rect 9680 3712 9732 3732
rect 9732 3712 9734 3732
rect 9862 5636 9918 5672
rect 9862 5616 9864 5636
rect 9864 5616 9916 5636
rect 9916 5616 9918 5636
rect 9770 3168 9826 3224
rect 11150 12552 11206 12608
rect 13818 15952 13874 16008
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 22834 16496 22890 16552
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 12438 14864 12494 14920
rect 10966 8200 11022 8256
rect 10598 6316 10654 6352
rect 10782 6432 10838 6488
rect 10598 6296 10600 6316
rect 10600 6296 10652 6316
rect 10652 6296 10654 6316
rect 10230 3168 10286 3224
rect 10230 2080 10286 2136
rect 10598 5108 10600 5128
rect 10600 5108 10652 5128
rect 10652 5108 10654 5128
rect 10598 5072 10654 5108
rect 10874 5092 10930 5128
rect 10874 5072 10876 5092
rect 10876 5072 10928 5092
rect 10928 5072 10930 5092
rect 10598 3576 10654 3632
rect 11334 10104 11390 10160
rect 14278 12588 14280 12608
rect 14280 12588 14332 12608
rect 14332 12588 14334 12608
rect 14278 12552 14334 12588
rect 13910 12416 13966 12472
rect 15750 12552 15806 12608
rect 13542 11212 13598 11248
rect 13542 11192 13544 11212
rect 13544 11192 13596 11212
rect 13596 11192 13598 11212
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 22926 15136 22982 15192
rect 24398 15308 24400 15328
rect 24400 15308 24452 15328
rect 24452 15308 24454 15328
rect 24398 15272 24454 15308
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 16854 12588 16856 12608
rect 16856 12588 16908 12608
rect 16908 12588 16910 12608
rect 16854 12552 16910 12588
rect 18326 12436 18382 12472
rect 18326 12416 18328 12436
rect 18328 12416 18380 12436
rect 18380 12416 18382 12436
rect 11886 9324 11888 9344
rect 11888 9324 11940 9344
rect 11940 9324 11942 9344
rect 11886 9288 11942 9324
rect 11242 8628 11298 8664
rect 11242 8608 11244 8628
rect 11244 8608 11296 8628
rect 11296 8608 11298 8628
rect 13266 10104 13322 10160
rect 12254 8508 12256 8528
rect 12256 8508 12308 8528
rect 12308 8508 12310 8528
rect 12254 8472 12310 8508
rect 11794 8200 11850 8256
rect 12530 6296 12586 6352
rect 11610 4256 11666 4312
rect 11242 3984 11298 4040
rect 11702 3884 11704 3904
rect 11704 3884 11756 3904
rect 11756 3884 11758 3904
rect 11702 3848 11758 3884
rect 12990 5344 13046 5400
rect 12898 5108 12900 5128
rect 12900 5108 12952 5128
rect 12952 5108 12954 5128
rect 12898 5072 12954 5108
rect 12990 4936 13046 4992
rect 12622 4392 12678 4448
rect 12438 4020 12440 4040
rect 12440 4020 12492 4040
rect 12492 4020 12494 4040
rect 12438 3984 12494 4020
rect 11058 1400 11114 1456
rect 16118 10376 16174 10432
rect 14278 9988 14334 10024
rect 14278 9968 14280 9988
rect 14280 9968 14332 9988
rect 14332 9968 14334 9988
rect 14186 9288 14242 9344
rect 13450 8492 13506 8528
rect 13450 8472 13452 8492
rect 13452 8472 13504 8492
rect 13504 8472 13506 8492
rect 18142 10412 18144 10432
rect 18144 10412 18196 10432
rect 18196 10412 18198 10432
rect 18142 10376 18198 10412
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 21362 12144 21418 12200
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 17590 9968 17646 10024
rect 18050 10004 18052 10024
rect 18052 10004 18104 10024
rect 18104 10004 18106 10024
rect 18050 9968 18106 10004
rect 18694 10104 18750 10160
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 19982 10376 20038 10432
rect 17406 7964 17408 7984
rect 17408 7964 17460 7984
rect 17460 7964 17462 7984
rect 17406 7928 17462 7964
rect 15290 6432 15346 6488
rect 13450 4528 13506 4584
rect 12070 2508 12126 2544
rect 12070 2488 12072 2508
rect 12072 2488 12124 2508
rect 12124 2488 12126 2508
rect 13082 2796 13084 2816
rect 13084 2796 13136 2816
rect 13136 2796 13138 2816
rect 13082 2760 13138 2796
rect 14002 4528 14058 4584
rect 13910 3848 13966 3904
rect 14002 3440 14058 3496
rect 15014 4800 15070 4856
rect 14278 3168 14334 3224
rect 15198 5208 15254 5264
rect 15198 4548 15254 4584
rect 15198 4528 15200 4548
rect 15200 4528 15252 4548
rect 15252 4528 15254 4548
rect 15474 4428 15476 4448
rect 15476 4428 15528 4448
rect 15528 4428 15530 4448
rect 15474 4392 15530 4428
rect 15658 3712 15714 3768
rect 16854 5888 16910 5944
rect 16670 4664 16726 4720
rect 17222 5072 17278 5128
rect 16854 4392 16910 4448
rect 15842 2896 15898 2952
rect 16118 2760 16174 2816
rect 15842 1944 15898 2000
rect 17958 5636 18014 5672
rect 17958 5616 17960 5636
rect 17960 5616 18012 5636
rect 18012 5616 18014 5636
rect 17774 4972 17776 4992
rect 17776 4972 17828 4992
rect 17828 4972 17830 4992
rect 17774 4936 17830 4972
rect 17038 3576 17094 3632
rect 17314 3612 17316 3632
rect 17316 3612 17368 3632
rect 17368 3612 17370 3632
rect 17314 3576 17370 3612
rect 17682 3712 17738 3768
rect 17406 3440 17462 3496
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 20258 10104 20314 10160
rect 18234 7792 18290 7848
rect 18050 4936 18106 4992
rect 17682 3188 17738 3224
rect 17682 3168 17684 3188
rect 17684 3168 17736 3188
rect 17736 3168 17738 3188
rect 17222 2352 17278 2408
rect 18786 7928 18842 7984
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 18878 5772 18934 5808
rect 18878 5752 18880 5772
rect 18880 5752 18932 5772
rect 18932 5752 18934 5772
rect 19338 5888 19394 5944
rect 18418 5208 18474 5264
rect 18878 4664 18934 4720
rect 18602 4392 18658 4448
rect 19338 4936 19394 4992
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 19890 5092 19946 5128
rect 19890 5072 19892 5092
rect 19892 5072 19944 5092
rect 19944 5072 19946 5092
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 19430 3712 19486 3768
rect 20074 3712 20130 3768
rect 19154 3576 19210 3632
rect 25870 12708 25926 12744
rect 25870 12688 25872 12708
rect 25872 12688 25924 12708
rect 25924 12688 25926 12708
rect 25042 12144 25098 12200
rect 24398 11348 24454 11384
rect 24398 11328 24400 11348
rect 24400 11328 24452 11348
rect 24452 11328 24454 11348
rect 25870 10920 25926 10976
rect 26790 21528 26846 21584
rect 26514 21412 26570 21448
rect 26514 21392 26516 21412
rect 26516 21392 26568 21412
rect 26568 21392 26570 21412
rect 27434 21936 27490 21992
rect 33782 31320 33838 31376
rect 34940 32666 34996 32668
rect 35020 32666 35076 32668
rect 35100 32666 35156 32668
rect 35180 32666 35236 32668
rect 34940 32614 34966 32666
rect 34966 32614 34996 32666
rect 35020 32614 35030 32666
rect 35030 32614 35076 32666
rect 35100 32614 35146 32666
rect 35146 32614 35156 32666
rect 35180 32614 35210 32666
rect 35210 32614 35236 32666
rect 34940 32612 34996 32614
rect 35020 32612 35076 32614
rect 35100 32612 35156 32614
rect 35180 32612 35236 32614
rect 34940 31578 34996 31580
rect 35020 31578 35076 31580
rect 35100 31578 35156 31580
rect 35180 31578 35236 31580
rect 34940 31526 34966 31578
rect 34966 31526 34996 31578
rect 35020 31526 35030 31578
rect 35030 31526 35076 31578
rect 35100 31526 35146 31578
rect 35146 31526 35156 31578
rect 35180 31526 35210 31578
rect 35210 31526 35236 31578
rect 34940 31524 34996 31526
rect 35020 31524 35076 31526
rect 35100 31524 35156 31526
rect 35180 31524 35236 31526
rect 34940 30490 34996 30492
rect 35020 30490 35076 30492
rect 35100 30490 35156 30492
rect 35180 30490 35236 30492
rect 34940 30438 34966 30490
rect 34966 30438 34996 30490
rect 35020 30438 35030 30490
rect 35030 30438 35076 30490
rect 35100 30438 35146 30490
rect 35146 30438 35156 30490
rect 35180 30438 35210 30490
rect 35210 30438 35236 30490
rect 34940 30436 34996 30438
rect 35020 30436 35076 30438
rect 35100 30436 35156 30438
rect 35180 30436 35236 30438
rect 34334 29164 34390 29200
rect 34334 29144 34336 29164
rect 34336 29144 34388 29164
rect 34388 29144 34390 29164
rect 32310 28736 32366 28792
rect 34518 28056 34574 28112
rect 29550 25492 29606 25528
rect 29550 25472 29552 25492
rect 29552 25472 29604 25492
rect 29604 25472 29606 25492
rect 31850 25472 31906 25528
rect 31942 25220 31998 25256
rect 31942 25200 31944 25220
rect 31944 25200 31996 25220
rect 31996 25200 31998 25220
rect 29090 21936 29146 21992
rect 29274 21548 29330 21584
rect 29274 21528 29276 21548
rect 29276 21528 29328 21548
rect 29328 21528 29330 21548
rect 28998 21256 29054 21312
rect 28630 20848 28686 20904
rect 29366 20476 29368 20496
rect 29368 20476 29420 20496
rect 29420 20476 29422 20496
rect 29366 20440 29422 20476
rect 27158 17040 27214 17096
rect 28170 17076 28172 17096
rect 28172 17076 28224 17096
rect 28224 17076 28226 17096
rect 28170 17040 28226 17076
rect 26514 16496 26570 16552
rect 26422 15272 26478 15328
rect 26330 15136 26386 15192
rect 30470 21392 30526 21448
rect 32678 26152 32734 26208
rect 32586 25200 32642 25256
rect 33690 25492 33746 25528
rect 33690 25472 33692 25492
rect 33692 25472 33744 25492
rect 33744 25472 33746 25492
rect 32678 23432 32734 23488
rect 32310 20884 32312 20904
rect 32312 20884 32364 20904
rect 32364 20884 32366 20904
rect 32310 20848 32366 20884
rect 34426 23432 34482 23488
rect 34940 29402 34996 29404
rect 35020 29402 35076 29404
rect 35100 29402 35156 29404
rect 35180 29402 35236 29404
rect 34940 29350 34966 29402
rect 34966 29350 34996 29402
rect 35020 29350 35030 29402
rect 35030 29350 35076 29402
rect 35100 29350 35146 29402
rect 35146 29350 35156 29402
rect 35180 29350 35210 29402
rect 35210 29350 35236 29402
rect 34940 29348 34996 29350
rect 35020 29348 35076 29350
rect 35100 29348 35156 29350
rect 35180 29348 35236 29350
rect 34940 28314 34996 28316
rect 35020 28314 35076 28316
rect 35100 28314 35156 28316
rect 35180 28314 35236 28316
rect 34940 28262 34966 28314
rect 34966 28262 34996 28314
rect 35020 28262 35030 28314
rect 35030 28262 35076 28314
rect 35100 28262 35146 28314
rect 35146 28262 35156 28314
rect 35180 28262 35210 28314
rect 35210 28262 35236 28314
rect 34940 28260 34996 28262
rect 35020 28260 35076 28262
rect 35100 28260 35156 28262
rect 35180 28260 35236 28262
rect 34940 27226 34996 27228
rect 35020 27226 35076 27228
rect 35100 27226 35156 27228
rect 35180 27226 35236 27228
rect 34940 27174 34966 27226
rect 34966 27174 34996 27226
rect 35020 27174 35030 27226
rect 35030 27174 35076 27226
rect 35100 27174 35146 27226
rect 35146 27174 35156 27226
rect 35180 27174 35210 27226
rect 35210 27174 35236 27226
rect 34940 27172 34996 27174
rect 35020 27172 35076 27174
rect 35100 27172 35156 27174
rect 35180 27172 35236 27174
rect 34702 26188 34704 26208
rect 34704 26188 34756 26208
rect 34756 26188 34758 26208
rect 34702 26152 34758 26188
rect 34940 26138 34996 26140
rect 35020 26138 35076 26140
rect 35100 26138 35156 26140
rect 35180 26138 35236 26140
rect 34940 26086 34966 26138
rect 34966 26086 34996 26138
rect 35020 26086 35030 26138
rect 35030 26086 35076 26138
rect 35100 26086 35146 26138
rect 35146 26086 35156 26138
rect 35180 26086 35210 26138
rect 35210 26086 35236 26138
rect 34940 26084 34996 26086
rect 35020 26084 35076 26086
rect 35100 26084 35156 26086
rect 35180 26084 35236 26086
rect 34940 25050 34996 25052
rect 35020 25050 35076 25052
rect 35100 25050 35156 25052
rect 35180 25050 35236 25052
rect 34940 24998 34966 25050
rect 34966 24998 34996 25050
rect 35020 24998 35030 25050
rect 35030 24998 35076 25050
rect 35100 24998 35146 25050
rect 35146 24998 35156 25050
rect 35180 24998 35210 25050
rect 35210 24998 35236 25050
rect 34940 24996 34996 24998
rect 35020 24996 35076 24998
rect 35100 24996 35156 24998
rect 35180 24996 35236 24998
rect 34426 22616 34482 22672
rect 28630 15680 28686 15736
rect 27526 14048 27582 14104
rect 28906 14048 28962 14104
rect 26514 11328 26570 11384
rect 26698 11328 26754 11384
rect 27434 13504 27490 13560
rect 28722 12144 28778 12200
rect 27158 10804 27214 10840
rect 27158 10784 27160 10804
rect 27160 10784 27212 10804
rect 27212 10784 27214 10804
rect 29458 11328 29514 11384
rect 28722 10684 28724 10704
rect 28724 10684 28776 10704
rect 28776 10684 28778 10704
rect 28722 10648 28778 10684
rect 29274 10648 29330 10704
rect 26054 10376 26110 10432
rect 21914 9016 21970 9072
rect 21086 7928 21142 7984
rect 20718 7792 20774 7848
rect 20442 7540 20498 7576
rect 20442 7520 20444 7540
rect 20444 7520 20496 7540
rect 20496 7520 20498 7540
rect 22282 7520 22338 7576
rect 20442 6840 20498 6896
rect 21914 6840 21970 6896
rect 23662 7928 23718 7984
rect 22006 5888 22062 5944
rect 20442 5752 20498 5808
rect 20442 4664 20498 4720
rect 19062 3304 19118 3360
rect 18878 3052 18934 3088
rect 18878 3032 18880 3052
rect 18880 3032 18932 3052
rect 18932 3032 18934 3052
rect 19246 3440 19302 3496
rect 20718 5616 20774 5672
rect 22650 6976 22706 7032
rect 22006 5244 22008 5264
rect 22008 5244 22060 5264
rect 22060 5244 22062 5264
rect 22006 5208 22062 5244
rect 25042 6976 25098 7032
rect 24858 6296 24914 6352
rect 24766 6024 24822 6080
rect 23846 5908 23902 5944
rect 23846 5888 23848 5908
rect 23848 5888 23900 5908
rect 23900 5888 23902 5908
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 21822 4936 21878 4992
rect 21270 4428 21272 4448
rect 21272 4428 21324 4448
rect 21324 4428 21326 4448
rect 21270 4392 21326 4428
rect 24122 5228 24178 5264
rect 24122 5208 24124 5228
rect 24124 5208 24176 5228
rect 24176 5208 24178 5228
rect 21638 3712 21694 3768
rect 21362 3596 21418 3632
rect 21362 3576 21364 3596
rect 21364 3576 21416 3596
rect 21416 3576 21418 3596
rect 21454 3476 21456 3496
rect 21456 3476 21508 3496
rect 21508 3476 21510 3496
rect 21454 3440 21510 3476
rect 22650 4120 22706 4176
rect 23110 3884 23112 3904
rect 23112 3884 23164 3904
rect 23164 3884 23166 3904
rect 23110 3848 23166 3884
rect 24214 5072 24270 5128
rect 24030 4972 24032 4992
rect 24032 4972 24084 4992
rect 24084 4972 24086 4992
rect 24030 4936 24086 4972
rect 23662 4800 23718 4856
rect 30654 17040 30710 17096
rect 31574 16496 31630 16552
rect 30194 15680 30250 15736
rect 30562 15700 30618 15736
rect 30562 15680 30564 15700
rect 30564 15680 30616 15700
rect 30616 15680 30618 15700
rect 30746 14884 30802 14920
rect 30746 14864 30748 14884
rect 30748 14864 30800 14884
rect 30800 14864 30802 14884
rect 30286 14612 30342 14648
rect 30286 14592 30288 14612
rect 30288 14592 30340 14612
rect 30340 14592 30342 14612
rect 30378 13776 30434 13832
rect 30102 11348 30158 11384
rect 30102 11328 30104 11348
rect 30104 11328 30156 11348
rect 30156 11328 30158 11348
rect 29734 10920 29790 10976
rect 29642 10784 29698 10840
rect 34518 22344 34574 22400
rect 31850 14592 31906 14648
rect 32310 13504 32366 13560
rect 30010 10648 30066 10704
rect 32310 10648 32366 10704
rect 29550 8472 29606 8528
rect 32402 9036 32458 9072
rect 32402 9016 32404 9036
rect 32404 9016 32456 9036
rect 32456 9016 32458 9036
rect 32862 17176 32918 17232
rect 32954 14864 33010 14920
rect 34058 19080 34114 19136
rect 33690 18808 33746 18864
rect 33506 17176 33562 17232
rect 33690 14356 33692 14376
rect 33692 14356 33744 14376
rect 33744 14356 33746 14376
rect 33690 14320 33746 14356
rect 34242 13504 34298 13560
rect 25962 5616 26018 5672
rect 26514 5752 26570 5808
rect 25778 5208 25834 5264
rect 24858 4936 24914 4992
rect 22190 3440 22246 3496
rect 22742 3304 22798 3360
rect 21822 1808 21878 1864
rect 25594 4156 25596 4176
rect 25596 4156 25648 4176
rect 25648 4156 25650 4176
rect 25594 4120 25650 4156
rect 24950 3848 25006 3904
rect 24582 3440 24638 3496
rect 23846 3032 23902 3088
rect 26974 6060 26976 6080
rect 26976 6060 27028 6080
rect 27028 6060 27030 6080
rect 26974 6024 27030 6060
rect 26698 4936 26754 4992
rect 26882 4800 26938 4856
rect 28538 5888 28594 5944
rect 26698 3984 26754 4040
rect 28354 3884 28356 3904
rect 28356 3884 28408 3904
rect 28408 3884 28410 3904
rect 28354 3848 28410 3884
rect 32678 7828 32680 7848
rect 32680 7828 32732 7848
rect 32732 7828 32734 7848
rect 32678 7792 32734 7828
rect 33230 9988 33286 10024
rect 33230 9968 33232 9988
rect 33232 9968 33284 9988
rect 33284 9968 33286 9988
rect 33322 7792 33378 7848
rect 29274 6296 29330 6352
rect 29274 5616 29330 5672
rect 37554 38256 37610 38312
rect 36266 34620 36268 34640
rect 36268 34620 36320 34640
rect 36320 34620 36322 34640
rect 36266 34584 36322 34620
rect 35990 33632 36046 33688
rect 35806 32544 35862 32600
rect 35622 31320 35678 31376
rect 35438 28736 35494 28792
rect 34940 23962 34996 23964
rect 35020 23962 35076 23964
rect 35100 23962 35156 23964
rect 35180 23962 35236 23964
rect 34940 23910 34966 23962
rect 34966 23910 34996 23962
rect 35020 23910 35030 23962
rect 35030 23910 35076 23962
rect 35100 23910 35146 23962
rect 35146 23910 35156 23962
rect 35180 23910 35210 23962
rect 35210 23910 35236 23962
rect 34940 23908 34996 23910
rect 35020 23908 35076 23910
rect 35100 23908 35156 23910
rect 35180 23908 35236 23910
rect 34940 22874 34996 22876
rect 35020 22874 35076 22876
rect 35100 22874 35156 22876
rect 35180 22874 35236 22876
rect 34940 22822 34966 22874
rect 34966 22822 34996 22874
rect 35020 22822 35030 22874
rect 35030 22822 35076 22874
rect 35100 22822 35146 22874
rect 35146 22822 35156 22874
rect 35180 22822 35210 22874
rect 35210 22822 35236 22874
rect 34940 22820 34996 22822
rect 35020 22820 35076 22822
rect 35100 22820 35156 22822
rect 35180 22820 35236 22822
rect 34940 21786 34996 21788
rect 35020 21786 35076 21788
rect 35100 21786 35156 21788
rect 35180 21786 35236 21788
rect 34940 21734 34966 21786
rect 34966 21734 34996 21786
rect 35020 21734 35030 21786
rect 35030 21734 35076 21786
rect 35100 21734 35146 21786
rect 35146 21734 35156 21786
rect 35180 21734 35210 21786
rect 35210 21734 35236 21786
rect 34940 21732 34996 21734
rect 35020 21732 35076 21734
rect 35100 21732 35156 21734
rect 35180 21732 35236 21734
rect 34940 20698 34996 20700
rect 35020 20698 35076 20700
rect 35100 20698 35156 20700
rect 35180 20698 35236 20700
rect 34940 20646 34966 20698
rect 34966 20646 34996 20698
rect 35020 20646 35030 20698
rect 35030 20646 35076 20698
rect 35100 20646 35146 20698
rect 35146 20646 35156 20698
rect 35180 20646 35210 20698
rect 35210 20646 35236 20698
rect 34940 20644 34996 20646
rect 35020 20644 35076 20646
rect 35100 20644 35156 20646
rect 35180 20644 35236 20646
rect 34940 19610 34996 19612
rect 35020 19610 35076 19612
rect 35100 19610 35156 19612
rect 35180 19610 35236 19612
rect 34940 19558 34966 19610
rect 34966 19558 34996 19610
rect 35020 19558 35030 19610
rect 35030 19558 35076 19610
rect 35100 19558 35146 19610
rect 35146 19558 35156 19610
rect 35180 19558 35210 19610
rect 35210 19558 35236 19610
rect 34940 19556 34996 19558
rect 35020 19556 35076 19558
rect 35100 19556 35156 19558
rect 35180 19556 35236 19558
rect 34610 13368 34666 13424
rect 34940 18522 34996 18524
rect 35020 18522 35076 18524
rect 35100 18522 35156 18524
rect 35180 18522 35236 18524
rect 34940 18470 34966 18522
rect 34966 18470 34996 18522
rect 35020 18470 35030 18522
rect 35030 18470 35076 18522
rect 35100 18470 35146 18522
rect 35146 18470 35156 18522
rect 35180 18470 35210 18522
rect 35210 18470 35236 18522
rect 34940 18468 34996 18470
rect 35020 18468 35076 18470
rect 35100 18468 35156 18470
rect 35180 18468 35236 18470
rect 34940 17434 34996 17436
rect 35020 17434 35076 17436
rect 35100 17434 35156 17436
rect 35180 17434 35236 17436
rect 34940 17382 34966 17434
rect 34966 17382 34996 17434
rect 35020 17382 35030 17434
rect 35030 17382 35076 17434
rect 35100 17382 35146 17434
rect 35146 17382 35156 17434
rect 35180 17382 35210 17434
rect 35210 17382 35236 17434
rect 34940 17380 34996 17382
rect 35020 17380 35076 17382
rect 35100 17380 35156 17382
rect 35180 17380 35236 17382
rect 34978 17176 35034 17232
rect 34940 16346 34996 16348
rect 35020 16346 35076 16348
rect 35100 16346 35156 16348
rect 35180 16346 35236 16348
rect 34940 16294 34966 16346
rect 34966 16294 34996 16346
rect 35020 16294 35030 16346
rect 35030 16294 35076 16346
rect 35100 16294 35146 16346
rect 35146 16294 35156 16346
rect 35180 16294 35210 16346
rect 35210 16294 35236 16346
rect 34940 16292 34996 16294
rect 35020 16292 35076 16294
rect 35100 16292 35156 16294
rect 35180 16292 35236 16294
rect 35990 28056 36046 28112
rect 35622 26696 35678 26752
rect 35622 25608 35678 25664
rect 35806 26832 35862 26888
rect 35714 22344 35770 22400
rect 37554 34448 37610 34504
rect 36634 27956 36636 27976
rect 36636 27956 36688 27976
rect 36688 27956 36690 27976
rect 36634 27920 36690 27956
rect 36266 25236 36268 25256
rect 36268 25236 36320 25256
rect 36320 25236 36322 25256
rect 36266 25200 36322 25236
rect 34940 15258 34996 15260
rect 35020 15258 35076 15260
rect 35100 15258 35156 15260
rect 35180 15258 35236 15260
rect 34940 15206 34966 15258
rect 34966 15206 34996 15258
rect 35020 15206 35030 15258
rect 35030 15206 35076 15258
rect 35100 15206 35146 15258
rect 35146 15206 35156 15258
rect 35180 15206 35210 15258
rect 35210 15206 35236 15258
rect 34940 15204 34996 15206
rect 35020 15204 35076 15206
rect 35100 15204 35156 15206
rect 35180 15204 35236 15206
rect 34940 14170 34996 14172
rect 35020 14170 35076 14172
rect 35100 14170 35156 14172
rect 35180 14170 35236 14172
rect 34940 14118 34966 14170
rect 34966 14118 34996 14170
rect 35020 14118 35030 14170
rect 35030 14118 35076 14170
rect 35100 14118 35146 14170
rect 35146 14118 35156 14170
rect 35180 14118 35210 14170
rect 35210 14118 35236 14170
rect 34940 14116 34996 14118
rect 35020 14116 35076 14118
rect 35100 14116 35156 14118
rect 35180 14116 35236 14118
rect 34940 13082 34996 13084
rect 35020 13082 35076 13084
rect 35100 13082 35156 13084
rect 35180 13082 35236 13084
rect 34940 13030 34966 13082
rect 34966 13030 34996 13082
rect 35020 13030 35030 13082
rect 35030 13030 35076 13082
rect 35100 13030 35146 13082
rect 35146 13030 35156 13082
rect 35180 13030 35210 13082
rect 35210 13030 35236 13082
rect 34940 13028 34996 13030
rect 35020 13028 35076 13030
rect 35100 13028 35156 13030
rect 35180 13028 35236 13030
rect 34518 10648 34574 10704
rect 34702 10240 34758 10296
rect 34940 11994 34996 11996
rect 35020 11994 35076 11996
rect 35100 11994 35156 11996
rect 35180 11994 35236 11996
rect 34940 11942 34966 11994
rect 34966 11942 34996 11994
rect 35020 11942 35030 11994
rect 35030 11942 35076 11994
rect 35100 11942 35146 11994
rect 35146 11942 35156 11994
rect 35180 11942 35210 11994
rect 35210 11942 35236 11994
rect 34940 11940 34996 11942
rect 35020 11940 35076 11942
rect 35100 11940 35156 11942
rect 35180 11940 35236 11942
rect 34940 10906 34996 10908
rect 35020 10906 35076 10908
rect 35100 10906 35156 10908
rect 35180 10906 35236 10908
rect 34940 10854 34966 10906
rect 34966 10854 34996 10906
rect 35020 10854 35030 10906
rect 35030 10854 35076 10906
rect 35100 10854 35146 10906
rect 35146 10854 35156 10906
rect 35180 10854 35210 10906
rect 35210 10854 35236 10906
rect 34940 10852 34996 10854
rect 35020 10852 35076 10854
rect 35100 10852 35156 10854
rect 35180 10852 35236 10854
rect 32862 6296 32918 6352
rect 29458 5208 29514 5264
rect 29458 3984 29514 4040
rect 27250 3032 27306 3088
rect 28446 3476 28448 3496
rect 28448 3476 28500 3496
rect 28500 3476 28502 3496
rect 28446 3440 28502 3476
rect 30746 5908 30802 5944
rect 30746 5888 30748 5908
rect 30748 5888 30800 5908
rect 30800 5888 30802 5908
rect 29550 2896 29606 2952
rect 29918 3712 29974 3768
rect 30194 4972 30196 4992
rect 30196 4972 30248 4992
rect 30248 4972 30250 4992
rect 30194 4936 30250 4972
rect 31942 5752 31998 5808
rect 30654 5344 30710 5400
rect 30470 3612 30472 3632
rect 30472 3612 30524 3632
rect 30524 3612 30526 3632
rect 30470 3576 30526 3612
rect 29458 2080 29514 2136
rect 31574 4528 31630 4584
rect 30930 3340 30932 3360
rect 30932 3340 30984 3360
rect 30984 3340 30986 3360
rect 30930 3304 30986 3340
rect 30838 3032 30894 3088
rect 31574 2760 31630 2816
rect 30654 2624 30710 2680
rect 32310 5228 32366 5264
rect 32310 5208 32312 5228
rect 32312 5208 32364 5228
rect 32364 5208 32366 5228
rect 32770 4256 32826 4312
rect 32310 3848 32366 3904
rect 32034 3732 32090 3768
rect 32034 3712 32036 3732
rect 32036 3712 32088 3732
rect 32088 3712 32090 3732
rect 34940 9818 34996 9820
rect 35020 9818 35076 9820
rect 35100 9818 35156 9820
rect 35180 9818 35236 9820
rect 34940 9766 34966 9818
rect 34966 9766 34996 9818
rect 35020 9766 35030 9818
rect 35030 9766 35076 9818
rect 35100 9766 35146 9818
rect 35146 9766 35156 9818
rect 35180 9766 35210 9818
rect 35210 9766 35236 9818
rect 34940 9764 34996 9766
rect 35020 9764 35076 9766
rect 35100 9764 35156 9766
rect 35180 9764 35236 9766
rect 34940 8730 34996 8732
rect 35020 8730 35076 8732
rect 35100 8730 35156 8732
rect 35180 8730 35236 8732
rect 34940 8678 34966 8730
rect 34966 8678 34996 8730
rect 35020 8678 35030 8730
rect 35030 8678 35076 8730
rect 35100 8678 35146 8730
rect 35146 8678 35156 8730
rect 35180 8678 35210 8730
rect 35210 8678 35236 8730
rect 34940 8676 34996 8678
rect 35020 8676 35076 8678
rect 35100 8676 35156 8678
rect 35180 8676 35236 8678
rect 35346 11736 35402 11792
rect 35254 8200 35310 8256
rect 34940 7642 34996 7644
rect 35020 7642 35076 7644
rect 35100 7642 35156 7644
rect 35180 7642 35236 7644
rect 34940 7590 34966 7642
rect 34966 7590 34996 7642
rect 35020 7590 35030 7642
rect 35030 7590 35076 7642
rect 35100 7590 35146 7642
rect 35146 7590 35156 7642
rect 35180 7590 35210 7642
rect 35210 7590 35236 7642
rect 34940 7588 34996 7590
rect 35020 7588 35076 7590
rect 35100 7588 35156 7590
rect 35180 7588 35236 7590
rect 35070 7148 35072 7168
rect 35072 7148 35124 7168
rect 35124 7148 35126 7168
rect 35070 7112 35126 7148
rect 34940 6554 34996 6556
rect 35020 6554 35076 6556
rect 35100 6554 35156 6556
rect 35180 6554 35236 6556
rect 34940 6502 34966 6554
rect 34966 6502 34996 6554
rect 35020 6502 35030 6554
rect 35030 6502 35076 6554
rect 35100 6502 35146 6554
rect 35146 6502 35156 6554
rect 35180 6502 35210 6554
rect 35210 6502 35236 6554
rect 34940 6500 34996 6502
rect 35020 6500 35076 6502
rect 35100 6500 35156 6502
rect 35180 6500 35236 6502
rect 34702 6296 34758 6352
rect 34940 5466 34996 5468
rect 35020 5466 35076 5468
rect 35100 5466 35156 5468
rect 35180 5466 35236 5468
rect 34940 5414 34966 5466
rect 34966 5414 34996 5466
rect 35020 5414 35030 5466
rect 35030 5414 35076 5466
rect 35100 5414 35146 5466
rect 35146 5414 35156 5466
rect 35180 5414 35210 5466
rect 35210 5414 35236 5466
rect 34940 5412 34996 5414
rect 35020 5412 35076 5414
rect 35100 5412 35156 5414
rect 35180 5412 35236 5414
rect 34610 5208 34666 5264
rect 33138 3612 33140 3632
rect 33140 3612 33192 3632
rect 33192 3612 33194 3632
rect 33138 3576 33194 3612
rect 32954 3052 33010 3088
rect 32954 3032 32956 3052
rect 32956 3032 33008 3052
rect 33008 3032 33010 3052
rect 34242 3304 34298 3360
rect 34940 4378 34996 4380
rect 35020 4378 35076 4380
rect 35100 4378 35156 4380
rect 35180 4378 35236 4380
rect 34940 4326 34966 4378
rect 34966 4326 34996 4378
rect 35020 4326 35030 4378
rect 35030 4326 35076 4378
rect 35100 4326 35146 4378
rect 35146 4326 35156 4378
rect 35180 4326 35210 4378
rect 35210 4326 35236 4378
rect 34940 4324 34996 4326
rect 35020 4324 35076 4326
rect 35100 4324 35156 4326
rect 35180 4324 35236 4326
rect 34940 3290 34996 3292
rect 35020 3290 35076 3292
rect 35100 3290 35156 3292
rect 35180 3290 35236 3292
rect 34940 3238 34966 3290
rect 34966 3238 34996 3290
rect 35020 3238 35030 3290
rect 35030 3238 35076 3290
rect 35100 3238 35146 3290
rect 35146 3238 35156 3290
rect 35180 3238 35210 3290
rect 35210 3238 35236 3290
rect 34940 3236 34996 3238
rect 35020 3236 35076 3238
rect 35100 3236 35156 3238
rect 35180 3236 35236 3238
rect 35162 3032 35218 3088
rect 34794 2760 34850 2816
rect 34886 2488 34942 2544
rect 34940 2202 34996 2204
rect 35020 2202 35076 2204
rect 35100 2202 35156 2204
rect 35180 2202 35236 2204
rect 34940 2150 34966 2202
rect 34966 2150 34996 2202
rect 35020 2150 35030 2202
rect 35030 2150 35076 2202
rect 35100 2150 35146 2202
rect 35146 2150 35156 2202
rect 35180 2150 35210 2202
rect 35210 2150 35236 2202
rect 34940 2148 34996 2150
rect 35020 2148 35076 2150
rect 35100 2148 35156 2150
rect 35180 2148 35236 2150
rect 34978 1944 35034 2000
rect 33874 1808 33930 1864
rect 35806 21256 35862 21312
rect 37370 21292 37372 21312
rect 37372 21292 37424 21312
rect 37424 21292 37426 21312
rect 37370 21256 37426 21292
rect 37186 21120 37242 21176
rect 35714 19896 35770 19952
rect 35622 19216 35678 19272
rect 35806 17720 35862 17776
rect 35530 14184 35586 14240
rect 35990 14320 36046 14376
rect 35806 13368 35862 13424
rect 35806 13096 35862 13152
rect 35530 12688 35586 12744
rect 35622 12416 35678 12472
rect 37922 20440 37978 20496
rect 36266 19116 36268 19136
rect 36268 19116 36320 19136
rect 36320 19116 36322 19136
rect 36266 19080 36322 19116
rect 36818 18808 36874 18864
rect 37094 18808 37150 18864
rect 37094 15408 37150 15464
rect 36634 13776 36690 13832
rect 36082 12416 36138 12472
rect 35806 12144 35862 12200
rect 35806 12008 35862 12064
rect 35622 8472 35678 8528
rect 35622 8200 35678 8256
rect 35622 7384 35678 7440
rect 35990 9968 36046 10024
rect 35990 7928 36046 7984
rect 35714 5072 35770 5128
rect 35346 3984 35402 4040
rect 37278 7792 37334 7848
rect 37278 7112 37334 7168
rect 35990 3848 36046 3904
rect 37186 2896 37242 2952
rect 39394 3848 39450 3904
rect 37002 2644 37058 2680
rect 37002 2624 37004 2644
rect 37004 2624 37056 2644
rect 37056 2624 37058 2644
rect 36082 2488 36138 2544
rect 35806 1672 35862 1728
rect 35254 584 35310 640
<< metal3 >>
rect 36169 39402 36235 39405
rect 39520 39402 40000 39432
rect 36169 39400 40000 39402
rect 36169 39344 36174 39400
rect 36230 39344 40000 39400
rect 36169 39342 40000 39344
rect 36169 39339 36235 39342
rect 39520 39312 40000 39342
rect 37549 38314 37615 38317
rect 39520 38314 40000 38344
rect 37549 38312 40000 38314
rect 37549 38256 37554 38312
rect 37610 38256 40000 38312
rect 37549 38254 40000 38256
rect 37549 38251 37615 38254
rect 39520 38224 40000 38254
rect 19568 37568 19888 37569
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 37503 19888 37504
rect 35617 37090 35683 37093
rect 39520 37090 40000 37120
rect 35617 37088 40000 37090
rect 35617 37032 35622 37088
rect 35678 37032 40000 37088
rect 35617 37030 40000 37032
rect 35617 37027 35683 37030
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 39520 37000 40000 37030
rect 34928 36959 35248 36960
rect 19568 36480 19888 36481
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 33869 36138 33935 36141
rect 33869 36136 35680 36138
rect 33869 36080 33874 36136
rect 33930 36080 35680 36136
rect 33869 36078 35680 36080
rect 33869 36075 33935 36078
rect 35620 36002 35680 36078
rect 39520 36002 40000 36032
rect 35620 35942 40000 36002
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 39520 35912 40000 35942
rect 34928 35871 35248 35872
rect 19568 35392 19888 35393
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 35327 19888 35328
rect 39520 34914 40000 34944
rect 37782 34854 40000 34914
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 34783 35248 34784
rect 32029 34642 32095 34645
rect 36261 34642 36327 34645
rect 32029 34640 36327 34642
rect 32029 34584 32034 34640
rect 32090 34584 36266 34640
rect 36322 34584 36327 34640
rect 32029 34582 36327 34584
rect 32029 34579 32095 34582
rect 36261 34579 36327 34582
rect 37549 34506 37615 34509
rect 37782 34506 37842 34854
rect 39520 34824 40000 34854
rect 37549 34504 37842 34506
rect 37549 34448 37554 34504
rect 37610 34448 37842 34504
rect 37549 34446 37842 34448
rect 37549 34443 37615 34446
rect 19568 34304 19888 34305
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 34928 33760 35248 33761
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 33695 35248 33696
rect 35985 33690 36051 33693
rect 39520 33690 40000 33720
rect 35985 33688 40000 33690
rect 35985 33632 35990 33688
rect 36046 33632 40000 33688
rect 35985 33630 40000 33632
rect 35985 33627 36051 33630
rect 39520 33600 40000 33630
rect 0 33328 480 33448
rect 27981 33282 28047 33285
rect 31845 33282 31911 33285
rect 27981 33280 31911 33282
rect 27981 33224 27986 33280
rect 28042 33224 31850 33280
rect 31906 33224 31911 33280
rect 27981 33222 31911 33224
rect 27981 33219 28047 33222
rect 31845 33219 31911 33222
rect 19568 33216 19888 33217
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 33151 19888 33152
rect 29821 33146 29887 33149
rect 33501 33146 33567 33149
rect 29821 33144 33567 33146
rect 29821 33088 29826 33144
rect 29882 33088 33506 33144
rect 33562 33088 33567 33144
rect 29821 33086 33567 33088
rect 29821 33083 29887 33086
rect 33501 33083 33567 33086
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 34928 32672 35248 32673
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 32607 35248 32608
rect 35801 32602 35867 32605
rect 39520 32602 40000 32632
rect 35801 32600 40000 32602
rect 35801 32544 35806 32600
rect 35862 32544 40000 32600
rect 35801 32542 40000 32544
rect 35801 32539 35867 32542
rect 39520 32512 40000 32542
rect 19568 32128 19888 32129
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 34928 31584 35248 31585
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 31519 35248 31520
rect 30557 31378 30623 31381
rect 33777 31378 33843 31381
rect 30557 31376 33843 31378
rect 30557 31320 30562 31376
rect 30618 31320 33782 31376
rect 33838 31320 33843 31376
rect 30557 31318 33843 31320
rect 30557 31315 30623 31318
rect 33777 31315 33843 31318
rect 35617 31378 35683 31381
rect 39520 31378 40000 31408
rect 35617 31376 40000 31378
rect 35617 31320 35622 31376
rect 35678 31320 40000 31376
rect 35617 31318 40000 31320
rect 35617 31315 35683 31318
rect 39520 31288 40000 31318
rect 19568 31040 19888 31041
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 30975 19888 30976
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 34928 30496 35248 30497
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 30431 35248 30432
rect 30649 30290 30715 30293
rect 39520 30290 40000 30320
rect 30649 30288 40000 30290
rect 30649 30232 30654 30288
rect 30710 30232 40000 30288
rect 30649 30230 40000 30232
rect 30649 30227 30715 30230
rect 39520 30200 40000 30230
rect 19568 29952 19888 29953
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 29887 19888 29888
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 34928 29408 35248 29409
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 29343 35248 29344
rect 34329 29202 34395 29205
rect 39520 29202 40000 29232
rect 34329 29200 40000 29202
rect 34329 29144 34334 29200
rect 34390 29144 40000 29200
rect 34329 29142 40000 29144
rect 34329 29139 34395 29142
rect 39520 29112 40000 29142
rect 19568 28864 19888 28865
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 28799 19888 28800
rect 32305 28794 32371 28797
rect 35433 28794 35499 28797
rect 32305 28792 35499 28794
rect 32305 28736 32310 28792
rect 32366 28736 35438 28792
rect 35494 28736 35499 28792
rect 32305 28734 35499 28736
rect 32305 28731 32371 28734
rect 35433 28731 35499 28734
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 34928 28320 35248 28321
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 28255 35248 28256
rect 34513 28114 34579 28117
rect 35985 28114 36051 28117
rect 34513 28112 36051 28114
rect 34513 28056 34518 28112
rect 34574 28056 35990 28112
rect 36046 28056 36051 28112
rect 34513 28054 36051 28056
rect 34513 28051 34579 28054
rect 35985 28051 36051 28054
rect 36629 27978 36695 27981
rect 39520 27978 40000 28008
rect 36629 27976 40000 27978
rect 36629 27920 36634 27976
rect 36690 27920 40000 27976
rect 36629 27918 40000 27920
rect 36629 27915 36695 27918
rect 39520 27888 40000 27918
rect 19568 27776 19888 27777
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 27711 19888 27712
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 34928 27232 35248 27233
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 27167 35248 27168
rect 35801 26890 35867 26893
rect 39520 26890 40000 26920
rect 35801 26888 40000 26890
rect 35801 26832 35806 26888
rect 35862 26832 40000 26888
rect 35801 26830 40000 26832
rect 35801 26827 35867 26830
rect 39520 26800 40000 26830
rect 28717 26754 28783 26757
rect 35617 26754 35683 26757
rect 28717 26752 35683 26754
rect 28717 26696 28722 26752
rect 28778 26696 35622 26752
rect 35678 26696 35683 26752
rect 28717 26694 35683 26696
rect 28717 26691 28783 26694
rect 35617 26691 35683 26694
rect 19568 26688 19888 26689
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 23289 26346 23355 26349
rect 26417 26346 26483 26349
rect 23289 26344 26483 26346
rect 23289 26288 23294 26344
rect 23350 26288 26422 26344
rect 26478 26288 26483 26344
rect 23289 26286 26483 26288
rect 23289 26283 23355 26286
rect 26417 26283 26483 26286
rect 32673 26210 32739 26213
rect 34697 26210 34763 26213
rect 32673 26208 34763 26210
rect 32673 26152 32678 26208
rect 32734 26152 34702 26208
rect 34758 26152 34763 26208
rect 32673 26150 34763 26152
rect 32673 26147 32739 26150
rect 34697 26147 34763 26150
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 34928 26144 35248 26145
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 26079 35248 26080
rect 35617 25666 35683 25669
rect 39520 25666 40000 25696
rect 35617 25664 40000 25666
rect 35617 25608 35622 25664
rect 35678 25608 40000 25664
rect 35617 25606 40000 25608
rect 35617 25603 35683 25606
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 39520 25576 40000 25606
rect 19568 25535 19888 25536
rect 29545 25530 29611 25533
rect 31845 25530 31911 25533
rect 33685 25530 33751 25533
rect 29545 25528 33751 25530
rect 29545 25472 29550 25528
rect 29606 25472 31850 25528
rect 31906 25472 33690 25528
rect 33746 25472 33751 25528
rect 29545 25470 33751 25472
rect 29545 25467 29611 25470
rect 31845 25467 31911 25470
rect 33685 25467 33751 25470
rect 24393 25258 24459 25261
rect 26693 25258 26759 25261
rect 24393 25256 26759 25258
rect 24393 25200 24398 25256
rect 24454 25200 26698 25256
rect 26754 25200 26759 25256
rect 24393 25198 26759 25200
rect 24393 25195 24459 25198
rect 26693 25195 26759 25198
rect 31937 25258 32003 25261
rect 32581 25258 32647 25261
rect 36261 25258 36327 25261
rect 31937 25256 36327 25258
rect 31937 25200 31942 25256
rect 31998 25200 32586 25256
rect 32642 25200 36266 25256
rect 36322 25200 36327 25256
rect 31937 25198 36327 25200
rect 31937 25195 32003 25198
rect 32581 25195 32647 25198
rect 36261 25195 36327 25198
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 34928 25056 35248 25057
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 24991 35248 24992
rect 26601 24578 26667 24581
rect 39520 24578 40000 24608
rect 26601 24576 40000 24578
rect 26601 24520 26606 24576
rect 26662 24520 40000 24576
rect 26601 24518 40000 24520
rect 26601 24515 26667 24518
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 39520 24488 40000 24518
rect 19568 24447 19888 24448
rect 21817 24034 21883 24037
rect 24117 24034 24183 24037
rect 21817 24032 24183 24034
rect 21817 23976 21822 24032
rect 21878 23976 24122 24032
rect 24178 23976 24183 24032
rect 21817 23974 24183 23976
rect 21817 23971 21883 23974
rect 24117 23971 24183 23974
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 34928 23968 35248 23969
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 23903 35248 23904
rect 32673 23490 32739 23493
rect 27662 23488 32739 23490
rect 27662 23432 32678 23488
rect 32734 23432 32739 23488
rect 27662 23430 32739 23432
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 21173 23354 21239 23357
rect 23749 23354 23815 23357
rect 21173 23352 23815 23354
rect 21173 23296 21178 23352
rect 21234 23296 23754 23352
rect 23810 23296 23815 23352
rect 21173 23294 23815 23296
rect 21173 23291 21239 23294
rect 23749 23291 23815 23294
rect 27153 23354 27219 23357
rect 27662 23354 27722 23430
rect 32673 23427 32739 23430
rect 34421 23490 34487 23493
rect 39520 23490 40000 23520
rect 34421 23488 40000 23490
rect 34421 23432 34426 23488
rect 34482 23432 40000 23488
rect 34421 23430 40000 23432
rect 34421 23427 34487 23430
rect 39520 23400 40000 23430
rect 27153 23352 27722 23354
rect 27153 23296 27158 23352
rect 27214 23296 27722 23352
rect 27153 23294 27722 23296
rect 27153 23291 27219 23294
rect 21541 23082 21607 23085
rect 23841 23082 23907 23085
rect 21541 23080 23907 23082
rect 21541 23024 21546 23080
rect 21602 23024 23846 23080
rect 23902 23024 23907 23080
rect 21541 23022 23907 23024
rect 21541 23019 21607 23022
rect 23841 23019 23907 23022
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 34928 22880 35248 22881
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 22815 35248 22816
rect 25865 22674 25931 22677
rect 34421 22674 34487 22677
rect 25865 22672 34487 22674
rect 25865 22616 25870 22672
rect 25926 22616 34426 22672
rect 34482 22616 34487 22672
rect 25865 22614 34487 22616
rect 25865 22611 25931 22614
rect 34421 22611 34487 22614
rect 34513 22402 34579 22405
rect 35709 22402 35775 22405
rect 34513 22400 35775 22402
rect 34513 22344 34518 22400
rect 34574 22344 35714 22400
rect 35770 22344 35775 22400
rect 34513 22342 35775 22344
rect 34513 22339 34579 22342
rect 35709 22339 35775 22342
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 22271 19888 22272
rect 25773 22266 25839 22269
rect 39520 22266 40000 22296
rect 25773 22264 40000 22266
rect 25773 22208 25778 22264
rect 25834 22208 40000 22264
rect 25773 22206 40000 22208
rect 25773 22203 25839 22206
rect 39520 22176 40000 22206
rect 26049 21994 26115 21997
rect 27429 21994 27495 21997
rect 29085 21994 29151 21997
rect 26049 21992 29151 21994
rect 26049 21936 26054 21992
rect 26110 21936 27434 21992
rect 27490 21936 29090 21992
rect 29146 21936 29151 21992
rect 26049 21934 29151 21936
rect 26049 21931 26115 21934
rect 27429 21931 27495 21934
rect 29085 21931 29151 21934
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 34928 21792 35248 21793
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 21727 35248 21728
rect 26785 21586 26851 21589
rect 29269 21586 29335 21589
rect 26785 21584 29335 21586
rect 26785 21528 26790 21584
rect 26846 21528 29274 21584
rect 29330 21528 29335 21584
rect 26785 21526 29335 21528
rect 26785 21523 26851 21526
rect 29269 21523 29335 21526
rect 26509 21450 26575 21453
rect 30465 21450 30531 21453
rect 26509 21448 30531 21450
rect 26509 21392 26514 21448
rect 26570 21392 30470 21448
rect 30526 21392 30531 21448
rect 26509 21390 30531 21392
rect 26509 21387 26575 21390
rect 30465 21387 30531 21390
rect 24117 21314 24183 21317
rect 28993 21314 29059 21317
rect 24117 21312 29059 21314
rect 24117 21256 24122 21312
rect 24178 21256 28998 21312
rect 29054 21256 29059 21312
rect 24117 21254 29059 21256
rect 24117 21251 24183 21254
rect 28993 21251 29059 21254
rect 35801 21314 35867 21317
rect 37365 21314 37431 21317
rect 35801 21312 37431 21314
rect 35801 21256 35806 21312
rect 35862 21256 37370 21312
rect 37426 21256 37431 21312
rect 35801 21254 37431 21256
rect 35801 21251 35867 21254
rect 37365 21251 37431 21254
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 37181 21178 37247 21181
rect 39520 21178 40000 21208
rect 37181 21176 40000 21178
rect 37181 21120 37186 21176
rect 37242 21120 40000 21176
rect 37181 21118 40000 21120
rect 37181 21115 37247 21118
rect 39520 21088 40000 21118
rect 28625 20906 28691 20909
rect 32305 20906 32371 20909
rect 28625 20904 32371 20906
rect 28625 20848 28630 20904
rect 28686 20848 32310 20904
rect 32366 20848 32371 20904
rect 28625 20846 32371 20848
rect 28625 20843 28691 20846
rect 32305 20843 32371 20846
rect 21357 20770 21423 20773
rect 23749 20770 23815 20773
rect 21357 20768 23815 20770
rect 21357 20712 21362 20768
rect 21418 20712 23754 20768
rect 23810 20712 23815 20768
rect 21357 20710 23815 20712
rect 21357 20707 21423 20710
rect 23749 20707 23815 20710
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 34928 20704 35248 20705
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 20639 35248 20640
rect 29361 20498 29427 20501
rect 35750 20498 35756 20500
rect 29361 20496 35756 20498
rect 29361 20440 29366 20496
rect 29422 20440 35756 20496
rect 29361 20438 35756 20440
rect 29361 20435 29427 20438
rect 35750 20436 35756 20438
rect 35820 20498 35826 20500
rect 37917 20498 37983 20501
rect 35820 20496 37983 20498
rect 35820 20440 37922 20496
rect 37978 20440 37983 20496
rect 35820 20438 37983 20440
rect 35820 20436 35826 20438
rect 37917 20435 37983 20438
rect 22737 20226 22803 20229
rect 24669 20226 24735 20229
rect 25037 20226 25103 20229
rect 22737 20224 25103 20226
rect 22737 20168 22742 20224
rect 22798 20168 24674 20224
rect 24730 20168 25042 20224
rect 25098 20168 25103 20224
rect 22737 20166 25103 20168
rect 22737 20163 22803 20166
rect 24669 20163 24735 20166
rect 25037 20163 25103 20166
rect 19568 20160 19888 20161
rect 0 20090 480 20120
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 3417 20090 3483 20093
rect 0 20088 3483 20090
rect 0 20032 3422 20088
rect 3478 20032 3483 20088
rect 0 20030 3483 20032
rect 0 20000 480 20030
rect 3417 20027 3483 20030
rect 35709 19954 35775 19957
rect 39520 19954 40000 19984
rect 35709 19952 40000 19954
rect 35709 19896 35714 19952
rect 35770 19896 40000 19952
rect 35709 19894 40000 19896
rect 35709 19891 35775 19894
rect 39520 19864 40000 19894
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 34928 19616 35248 19617
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 19551 35248 19552
rect 35617 19276 35683 19277
rect 35566 19274 35572 19276
rect 35526 19214 35572 19274
rect 35636 19272 35683 19276
rect 35678 19216 35683 19272
rect 35566 19212 35572 19214
rect 35636 19212 35683 19216
rect 35617 19211 35683 19212
rect 34053 19138 34119 19141
rect 36261 19138 36327 19141
rect 34053 19136 36327 19138
rect 34053 19080 34058 19136
rect 34114 19080 36266 19136
rect 36322 19080 36327 19136
rect 34053 19078 36327 19080
rect 34053 19075 34119 19078
rect 36261 19075 36327 19078
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 19007 19888 19008
rect 33685 18866 33751 18869
rect 36813 18866 36879 18869
rect 33685 18864 36879 18866
rect 33685 18808 33690 18864
rect 33746 18808 36818 18864
rect 36874 18808 36879 18864
rect 33685 18806 36879 18808
rect 33685 18803 33751 18806
rect 36813 18803 36879 18806
rect 37089 18866 37155 18869
rect 39520 18866 40000 18896
rect 37089 18864 40000 18866
rect 37089 18808 37094 18864
rect 37150 18808 40000 18864
rect 37089 18806 40000 18808
rect 37089 18803 37155 18806
rect 39520 18776 40000 18806
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 34928 18528 35248 18529
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 18463 35248 18464
rect 3417 18186 3483 18189
rect 18689 18186 18755 18189
rect 3417 18184 18755 18186
rect 3417 18128 3422 18184
rect 3478 18128 18694 18184
rect 18750 18128 18755 18184
rect 3417 18126 18755 18128
rect 3417 18123 3483 18126
rect 18689 18123 18755 18126
rect 19568 17984 19888 17985
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 35801 17778 35867 17781
rect 39520 17778 40000 17808
rect 35801 17776 40000 17778
rect 35801 17720 35806 17776
rect 35862 17720 40000 17776
rect 35801 17718 40000 17720
rect 35801 17715 35867 17718
rect 39520 17688 40000 17718
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 34928 17440 35248 17441
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 17375 35248 17376
rect 32857 17234 32923 17237
rect 33501 17234 33567 17237
rect 34973 17234 35039 17237
rect 32857 17232 35039 17234
rect 32857 17176 32862 17232
rect 32918 17176 33506 17232
rect 33562 17176 34978 17232
rect 35034 17176 35039 17232
rect 32857 17174 35039 17176
rect 32857 17171 32923 17174
rect 33501 17171 33567 17174
rect 34973 17171 35039 17174
rect 13537 17098 13603 17101
rect 27153 17098 27219 17101
rect 13537 17096 27219 17098
rect 13537 17040 13542 17096
rect 13598 17040 27158 17096
rect 27214 17040 27219 17096
rect 13537 17038 27219 17040
rect 13537 17035 13603 17038
rect 27153 17035 27219 17038
rect 28165 17098 28231 17101
rect 30649 17098 30715 17101
rect 28165 17096 30715 17098
rect 28165 17040 28170 17096
rect 28226 17040 30654 17096
rect 30710 17040 30715 17096
rect 28165 17038 30715 17040
rect 28165 17035 28231 17038
rect 30649 17035 30715 17038
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 16831 19888 16832
rect 22829 16554 22895 16557
rect 26509 16554 26575 16557
rect 22829 16552 26575 16554
rect 22829 16496 22834 16552
rect 22890 16496 26514 16552
rect 26570 16496 26575 16552
rect 22829 16494 26575 16496
rect 22829 16491 22895 16494
rect 26509 16491 26575 16494
rect 31569 16554 31635 16557
rect 39520 16554 40000 16584
rect 31569 16552 40000 16554
rect 31569 16496 31574 16552
rect 31630 16496 40000 16552
rect 31569 16494 40000 16496
rect 31569 16491 31635 16494
rect 39520 16464 40000 16494
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 34928 16352 35248 16353
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 16287 35248 16288
rect 10133 16010 10199 16013
rect 13813 16010 13879 16013
rect 10133 16008 13879 16010
rect 10133 15952 10138 16008
rect 10194 15952 13818 16008
rect 13874 15952 13879 16008
rect 10133 15950 13879 15952
rect 10133 15947 10199 15950
rect 13813 15947 13879 15950
rect 7833 15874 7899 15877
rect 10041 15874 10107 15877
rect 7833 15872 10107 15874
rect 7833 15816 7838 15872
rect 7894 15816 10046 15872
rect 10102 15816 10107 15872
rect 7833 15814 10107 15816
rect 7833 15811 7899 15814
rect 10041 15811 10107 15814
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 5809 15738 5875 15741
rect 7741 15738 7807 15741
rect 5809 15736 7807 15738
rect 5809 15680 5814 15736
rect 5870 15680 7746 15736
rect 7802 15680 7807 15736
rect 5809 15678 7807 15680
rect 5809 15675 5875 15678
rect 7741 15675 7807 15678
rect 28625 15738 28691 15741
rect 30189 15738 30255 15741
rect 30557 15738 30623 15741
rect 28625 15736 30623 15738
rect 28625 15680 28630 15736
rect 28686 15680 30194 15736
rect 30250 15680 30562 15736
rect 30618 15680 30623 15736
rect 28625 15678 30623 15680
rect 28625 15675 28691 15678
rect 30189 15675 30255 15678
rect 30557 15675 30623 15678
rect 37089 15466 37155 15469
rect 39520 15466 40000 15496
rect 37089 15464 40000 15466
rect 37089 15408 37094 15464
rect 37150 15408 40000 15464
rect 37089 15406 40000 15408
rect 37089 15403 37155 15406
rect 39520 15376 40000 15406
rect 24393 15330 24459 15333
rect 26417 15330 26483 15333
rect 24393 15328 26483 15330
rect 24393 15272 24398 15328
rect 24454 15272 26422 15328
rect 26478 15272 26483 15328
rect 24393 15270 26483 15272
rect 24393 15267 24459 15270
rect 26417 15267 26483 15270
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 34928 15264 35248 15265
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 15199 35248 15200
rect 22921 15194 22987 15197
rect 26325 15194 26391 15197
rect 22921 15192 26391 15194
rect 22921 15136 22926 15192
rect 22982 15136 26330 15192
rect 26386 15136 26391 15192
rect 22921 15134 26391 15136
rect 22921 15131 22987 15134
rect 26325 15131 26391 15134
rect 10777 14922 10843 14925
rect 12433 14922 12499 14925
rect 10777 14920 12499 14922
rect 10777 14864 10782 14920
rect 10838 14864 12438 14920
rect 12494 14864 12499 14920
rect 10777 14862 12499 14864
rect 10777 14859 10843 14862
rect 12433 14859 12499 14862
rect 30741 14922 30807 14925
rect 32949 14922 33015 14925
rect 30741 14920 33015 14922
rect 30741 14864 30746 14920
rect 30802 14864 32954 14920
rect 33010 14864 33015 14920
rect 30741 14862 33015 14864
rect 30741 14859 30807 14862
rect 32949 14859 33015 14862
rect 19568 14720 19888 14721
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 30281 14650 30347 14653
rect 31845 14650 31911 14653
rect 30281 14648 31911 14650
rect 30281 14592 30286 14648
rect 30342 14592 31850 14648
rect 31906 14592 31911 14648
rect 30281 14590 31911 14592
rect 30281 14587 30347 14590
rect 31845 14587 31911 14590
rect 33685 14378 33751 14381
rect 35985 14378 36051 14381
rect 33685 14376 36051 14378
rect 33685 14320 33690 14376
rect 33746 14320 35990 14376
rect 36046 14320 36051 14376
rect 33685 14318 36051 14320
rect 33685 14315 33751 14318
rect 35985 14315 36051 14318
rect 35525 14242 35591 14245
rect 39520 14242 40000 14272
rect 35525 14240 40000 14242
rect 35525 14184 35530 14240
rect 35586 14184 40000 14240
rect 35525 14182 40000 14184
rect 35525 14179 35591 14182
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 34928 14176 35248 14177
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 39520 14152 40000 14182
rect 34928 14111 35248 14112
rect 5165 14106 5231 14109
rect 7373 14106 7439 14109
rect 5165 14104 7439 14106
rect 5165 14048 5170 14104
rect 5226 14048 7378 14104
rect 7434 14048 7439 14104
rect 5165 14046 7439 14048
rect 5165 14043 5231 14046
rect 7373 14043 7439 14046
rect 27521 14106 27587 14109
rect 28901 14106 28967 14109
rect 27521 14104 28967 14106
rect 27521 14048 27526 14104
rect 27582 14048 28906 14104
rect 28962 14048 28967 14104
rect 27521 14046 28967 14048
rect 27521 14043 27587 14046
rect 28901 14043 28967 14046
rect 5165 13970 5231 13973
rect 7281 13970 7347 13973
rect 5165 13968 7347 13970
rect 5165 13912 5170 13968
rect 5226 13912 7286 13968
rect 7342 13912 7347 13968
rect 5165 13910 7347 13912
rect 5165 13907 5231 13910
rect 7281 13907 7347 13910
rect 30373 13834 30439 13837
rect 36629 13834 36695 13837
rect 30373 13832 36695 13834
rect 30373 13776 30378 13832
rect 30434 13776 36634 13832
rect 36690 13776 36695 13832
rect 30373 13774 36695 13776
rect 30373 13771 30439 13774
rect 36629 13771 36695 13774
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 13567 19888 13568
rect 27429 13562 27495 13565
rect 32305 13562 32371 13565
rect 34237 13562 34303 13565
rect 27429 13560 34303 13562
rect 27429 13504 27434 13560
rect 27490 13504 32310 13560
rect 32366 13504 34242 13560
rect 34298 13504 34303 13560
rect 27429 13502 34303 13504
rect 27429 13499 27495 13502
rect 32305 13499 32371 13502
rect 34237 13499 34303 13502
rect 34605 13426 34671 13429
rect 35801 13426 35867 13429
rect 34605 13424 35867 13426
rect 34605 13368 34610 13424
rect 34666 13368 35806 13424
rect 35862 13368 35867 13424
rect 34605 13366 35867 13368
rect 34605 13363 34671 13366
rect 35801 13363 35867 13366
rect 35801 13154 35867 13157
rect 39520 13154 40000 13184
rect 35801 13152 40000 13154
rect 35801 13096 35806 13152
rect 35862 13096 40000 13152
rect 35801 13094 40000 13096
rect 35801 13091 35867 13094
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 34928 13088 35248 13089
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 39520 13064 40000 13094
rect 34928 13023 35248 13024
rect 25865 12746 25931 12749
rect 35525 12746 35591 12749
rect 25865 12744 35591 12746
rect 25865 12688 25870 12744
rect 25926 12688 35530 12744
rect 35586 12688 35591 12744
rect 25865 12686 35591 12688
rect 25865 12683 25931 12686
rect 35525 12683 35591 12686
rect 9949 12610 10015 12613
rect 11145 12610 11211 12613
rect 9949 12608 11211 12610
rect 9949 12552 9954 12608
rect 10010 12552 11150 12608
rect 11206 12552 11211 12608
rect 9949 12550 11211 12552
rect 9949 12547 10015 12550
rect 11145 12547 11211 12550
rect 14273 12610 14339 12613
rect 15745 12610 15811 12613
rect 16849 12610 16915 12613
rect 14273 12608 16915 12610
rect 14273 12552 14278 12608
rect 14334 12552 15750 12608
rect 15806 12552 16854 12608
rect 16910 12552 16915 12608
rect 14273 12550 16915 12552
rect 14273 12547 14339 12550
rect 15745 12547 15811 12550
rect 16849 12547 16915 12550
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 13905 12474 13971 12477
rect 18321 12474 18387 12477
rect 13905 12472 18387 12474
rect 13905 12416 13910 12472
rect 13966 12416 18326 12472
rect 18382 12416 18387 12472
rect 13905 12414 18387 12416
rect 13905 12411 13971 12414
rect 18321 12411 18387 12414
rect 35617 12474 35683 12477
rect 36077 12474 36143 12477
rect 35617 12472 36143 12474
rect 35617 12416 35622 12472
rect 35678 12416 36082 12472
rect 36138 12416 36143 12472
rect 35617 12414 36143 12416
rect 35617 12411 35683 12414
rect 36077 12411 36143 12414
rect 21357 12202 21423 12205
rect 25037 12202 25103 12205
rect 21357 12200 25103 12202
rect 21357 12144 21362 12200
rect 21418 12144 25042 12200
rect 25098 12144 25103 12200
rect 21357 12142 25103 12144
rect 21357 12139 21423 12142
rect 25037 12139 25103 12142
rect 28717 12202 28783 12205
rect 35801 12202 35867 12205
rect 28717 12200 35867 12202
rect 28717 12144 28722 12200
rect 28778 12144 35806 12200
rect 35862 12144 35867 12200
rect 28717 12142 35867 12144
rect 28717 12139 28783 12142
rect 35801 12139 35867 12142
rect 35801 12066 35867 12069
rect 39520 12066 40000 12096
rect 35801 12064 40000 12066
rect 35801 12008 35806 12064
rect 35862 12008 40000 12064
rect 35801 12006 40000 12008
rect 35801 12003 35867 12006
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 34928 12000 35248 12001
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 39520 11976 40000 12006
rect 34928 11935 35248 11936
rect 35341 11794 35407 11797
rect 35566 11794 35572 11796
rect 35341 11792 35572 11794
rect 35341 11736 35346 11792
rect 35402 11736 35572 11792
rect 35341 11734 35572 11736
rect 35341 11731 35407 11734
rect 35566 11732 35572 11734
rect 35636 11732 35642 11796
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 11391 19888 11392
rect 24393 11386 24459 11389
rect 26509 11386 26575 11389
rect 24393 11384 26575 11386
rect 24393 11328 24398 11384
rect 24454 11328 26514 11384
rect 26570 11328 26575 11384
rect 24393 11326 26575 11328
rect 24393 11323 24459 11326
rect 26509 11323 26575 11326
rect 26693 11386 26759 11389
rect 29453 11386 29519 11389
rect 30097 11386 30163 11389
rect 26693 11384 30163 11386
rect 26693 11328 26698 11384
rect 26754 11328 29458 11384
rect 29514 11328 30102 11384
rect 30158 11328 30163 11384
rect 26693 11326 30163 11328
rect 26693 11323 26759 11326
rect 29453 11323 29519 11326
rect 30097 11323 30163 11326
rect 10961 11250 11027 11253
rect 13537 11250 13603 11253
rect 10961 11248 13603 11250
rect 10961 11192 10966 11248
rect 11022 11192 13542 11248
rect 13598 11192 13603 11248
rect 10961 11190 13603 11192
rect 10961 11187 11027 11190
rect 13537 11187 13603 11190
rect 25865 10978 25931 10981
rect 29729 10978 29795 10981
rect 25865 10976 29795 10978
rect 25865 10920 25870 10976
rect 25926 10920 29734 10976
rect 29790 10920 29795 10976
rect 25865 10918 29795 10920
rect 25865 10915 25931 10918
rect 29729 10915 29795 10918
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 34928 10912 35248 10913
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 10847 35248 10848
rect 27153 10842 27219 10845
rect 29637 10842 29703 10845
rect 39520 10842 40000 10872
rect 27153 10840 29703 10842
rect 27153 10784 27158 10840
rect 27214 10784 29642 10840
rect 29698 10784 29703 10840
rect 27153 10782 29703 10784
rect 27153 10779 27219 10782
rect 29637 10779 29703 10782
rect 35390 10782 40000 10842
rect 28717 10706 28783 10709
rect 29269 10706 29335 10709
rect 30005 10706 30071 10709
rect 32305 10706 32371 10709
rect 28717 10704 32371 10706
rect 28717 10648 28722 10704
rect 28778 10648 29274 10704
rect 29330 10648 30010 10704
rect 30066 10648 32310 10704
rect 32366 10648 32371 10704
rect 28717 10646 32371 10648
rect 28717 10643 28783 10646
rect 29269 10643 29335 10646
rect 30005 10643 30071 10646
rect 32305 10643 32371 10646
rect 34513 10706 34579 10709
rect 35390 10706 35450 10782
rect 39520 10752 40000 10782
rect 34513 10704 35450 10706
rect 34513 10648 34518 10704
rect 34574 10648 35450 10704
rect 34513 10646 35450 10648
rect 34513 10643 34579 10646
rect 16113 10434 16179 10437
rect 18137 10434 18203 10437
rect 16113 10432 18203 10434
rect 16113 10376 16118 10432
rect 16174 10376 18142 10432
rect 18198 10376 18203 10432
rect 16113 10374 18203 10376
rect 16113 10371 16179 10374
rect 18137 10371 18203 10374
rect 19977 10434 20043 10437
rect 26049 10434 26115 10437
rect 19977 10432 26115 10434
rect 19977 10376 19982 10432
rect 20038 10376 26054 10432
rect 26110 10376 26115 10432
rect 19977 10374 26115 10376
rect 19977 10371 20043 10374
rect 26049 10371 26115 10374
rect 19568 10368 19888 10369
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 34697 10298 34763 10301
rect 34697 10296 36186 10298
rect 34697 10240 34702 10296
rect 34758 10240 36186 10296
rect 34697 10238 36186 10240
rect 34697 10235 34763 10238
rect 11329 10162 11395 10165
rect 13261 10162 13327 10165
rect 11329 10160 13327 10162
rect 11329 10104 11334 10160
rect 11390 10104 13266 10160
rect 13322 10104 13327 10160
rect 11329 10102 13327 10104
rect 11329 10099 11395 10102
rect 13261 10099 13327 10102
rect 18689 10162 18755 10165
rect 20253 10162 20319 10165
rect 18689 10160 20319 10162
rect 18689 10104 18694 10160
rect 18750 10104 20258 10160
rect 20314 10104 20319 10160
rect 18689 10102 20319 10104
rect 18689 10099 18755 10102
rect 20253 10099 20319 10102
rect 14273 10026 14339 10029
rect 17585 10026 17651 10029
rect 18045 10026 18111 10029
rect 14273 10024 18111 10026
rect 14273 9968 14278 10024
rect 14334 9968 17590 10024
rect 17646 9968 18050 10024
rect 18106 9968 18111 10024
rect 14273 9966 18111 9968
rect 14273 9963 14339 9966
rect 17585 9963 17651 9966
rect 18045 9963 18111 9966
rect 33225 10026 33291 10029
rect 35985 10026 36051 10029
rect 33225 10024 36051 10026
rect 33225 9968 33230 10024
rect 33286 9968 35990 10024
rect 36046 9968 36051 10024
rect 33225 9966 36051 9968
rect 33225 9963 33291 9966
rect 35985 9963 36051 9966
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 34928 9824 35248 9825
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 9759 35248 9760
rect 36126 9754 36186 10238
rect 39520 9754 40000 9784
rect 36126 9694 40000 9754
rect 39520 9664 40000 9694
rect 11881 9346 11947 9349
rect 14181 9346 14247 9349
rect 11881 9344 14247 9346
rect 11881 9288 11886 9344
rect 11942 9288 14186 9344
rect 14242 9288 14247 9344
rect 11881 9286 14247 9288
rect 11881 9283 11947 9286
rect 14181 9283 14247 9286
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 21909 9074 21975 9077
rect 32397 9074 32463 9077
rect 21909 9072 32463 9074
rect 21909 9016 21914 9072
rect 21970 9016 32402 9072
rect 32458 9016 32463 9072
rect 21909 9014 32463 9016
rect 21909 9011 21975 9014
rect 32397 9011 32463 9014
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 34928 8736 35248 8737
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 8671 35248 8672
rect 7189 8666 7255 8669
rect 11237 8666 11303 8669
rect 7189 8664 11303 8666
rect 7189 8608 7194 8664
rect 7250 8608 11242 8664
rect 11298 8608 11303 8664
rect 7189 8606 11303 8608
rect 7189 8603 7255 8606
rect 11237 8603 11303 8606
rect 12249 8530 12315 8533
rect 13445 8530 13511 8533
rect 29545 8530 29611 8533
rect 12249 8528 29611 8530
rect 12249 8472 12254 8528
rect 12310 8472 13450 8528
rect 13506 8472 29550 8528
rect 29606 8472 29611 8528
rect 12249 8470 29611 8472
rect 12249 8467 12315 8470
rect 13445 8467 13511 8470
rect 29545 8467 29611 8470
rect 35617 8530 35683 8533
rect 39520 8530 40000 8560
rect 35617 8528 40000 8530
rect 35617 8472 35622 8528
rect 35678 8472 40000 8528
rect 35617 8470 40000 8472
rect 35617 8467 35683 8470
rect 39520 8440 40000 8470
rect 10961 8258 11027 8261
rect 11789 8258 11855 8261
rect 10961 8256 11855 8258
rect 10961 8200 10966 8256
rect 11022 8200 11794 8256
rect 11850 8200 11855 8256
rect 10961 8198 11855 8200
rect 10961 8195 11027 8198
rect 11789 8195 11855 8198
rect 35249 8258 35315 8261
rect 35617 8258 35683 8261
rect 35249 8256 35683 8258
rect 35249 8200 35254 8256
rect 35310 8200 35622 8256
rect 35678 8200 35683 8256
rect 35249 8198 35683 8200
rect 35249 8195 35315 8198
rect 35617 8195 35683 8198
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 17401 7986 17467 7989
rect 18781 7986 18847 7989
rect 21081 7986 21147 7989
rect 17401 7984 21147 7986
rect 17401 7928 17406 7984
rect 17462 7928 18786 7984
rect 18842 7928 21086 7984
rect 21142 7928 21147 7984
rect 17401 7926 21147 7928
rect 17401 7923 17467 7926
rect 18781 7923 18847 7926
rect 21081 7923 21147 7926
rect 23657 7986 23723 7989
rect 35985 7986 36051 7989
rect 23657 7984 36051 7986
rect 23657 7928 23662 7984
rect 23718 7928 35990 7984
rect 36046 7928 36051 7984
rect 23657 7926 36051 7928
rect 23657 7923 23723 7926
rect 35985 7923 36051 7926
rect 18229 7850 18295 7853
rect 20713 7850 20779 7853
rect 18229 7848 20779 7850
rect 18229 7792 18234 7848
rect 18290 7792 20718 7848
rect 20774 7792 20779 7848
rect 18229 7790 20779 7792
rect 18229 7787 18295 7790
rect 20713 7787 20779 7790
rect 32673 7850 32739 7853
rect 33317 7850 33383 7853
rect 37273 7850 37339 7853
rect 32673 7848 37339 7850
rect 32673 7792 32678 7848
rect 32734 7792 33322 7848
rect 33378 7792 37278 7848
rect 37334 7792 37339 7848
rect 32673 7790 37339 7792
rect 32673 7787 32739 7790
rect 33317 7787 33383 7790
rect 37273 7787 37339 7790
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 34928 7648 35248 7649
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 7583 35248 7584
rect 20437 7578 20503 7581
rect 22277 7578 22343 7581
rect 20437 7576 22343 7578
rect 20437 7520 20442 7576
rect 20498 7520 22282 7576
rect 22338 7520 22343 7576
rect 20437 7518 22343 7520
rect 20437 7515 20503 7518
rect 22277 7515 22343 7518
rect 35617 7442 35683 7445
rect 39520 7442 40000 7472
rect 35617 7440 40000 7442
rect 35617 7384 35622 7440
rect 35678 7384 40000 7440
rect 35617 7382 40000 7384
rect 35617 7379 35683 7382
rect 39520 7352 40000 7382
rect 35065 7170 35131 7173
rect 37273 7170 37339 7173
rect 35065 7168 37339 7170
rect 35065 7112 35070 7168
rect 35126 7112 37278 7168
rect 37334 7112 37339 7168
rect 35065 7110 37339 7112
rect 35065 7107 35131 7110
rect 37273 7107 37339 7110
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 22645 7034 22711 7037
rect 25037 7034 25103 7037
rect 22645 7032 25103 7034
rect 22645 6976 22650 7032
rect 22706 6976 25042 7032
rect 25098 6976 25103 7032
rect 22645 6974 25103 6976
rect 22645 6971 22711 6974
rect 25037 6971 25103 6974
rect 3969 6898 4035 6901
rect 3374 6896 4035 6898
rect 3374 6840 3974 6896
rect 4030 6840 4035 6896
rect 3374 6838 4035 6840
rect 0 6762 480 6792
rect 2221 6762 2287 6765
rect 2773 6762 2839 6765
rect 3374 6762 3434 6838
rect 3969 6835 4035 6838
rect 20437 6898 20503 6901
rect 21909 6898 21975 6901
rect 20437 6896 21975 6898
rect 20437 6840 20442 6896
rect 20498 6840 21914 6896
rect 21970 6840 21975 6896
rect 20437 6838 21975 6840
rect 20437 6835 20503 6838
rect 21909 6835 21975 6838
rect 0 6760 3434 6762
rect 0 6704 2226 6760
rect 2282 6704 2778 6760
rect 2834 6704 3434 6760
rect 0 6702 3434 6704
rect 3509 6762 3575 6765
rect 5165 6762 5231 6765
rect 5993 6762 6059 6765
rect 3509 6760 6059 6762
rect 3509 6704 3514 6760
rect 3570 6704 5170 6760
rect 5226 6704 5998 6760
rect 6054 6704 6059 6760
rect 3509 6702 6059 6704
rect 0 6672 480 6702
rect 2221 6699 2287 6702
rect 2773 6699 2839 6702
rect 3509 6699 3575 6702
rect 5165 6699 5231 6702
rect 5993 6699 6059 6702
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 34928 6560 35248 6561
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 6495 35248 6496
rect 10777 6490 10843 6493
rect 15285 6490 15351 6493
rect 10777 6488 15351 6490
rect 10777 6432 10782 6488
rect 10838 6432 15290 6488
rect 15346 6432 15351 6488
rect 10777 6430 15351 6432
rect 10777 6427 10843 6430
rect 15285 6427 15351 6430
rect 10593 6354 10659 6357
rect 12525 6354 12591 6357
rect 10593 6352 12591 6354
rect 10593 6296 10598 6352
rect 10654 6296 12530 6352
rect 12586 6296 12591 6352
rect 10593 6294 12591 6296
rect 10593 6291 10659 6294
rect 12525 6291 12591 6294
rect 24853 6354 24919 6357
rect 29269 6354 29335 6357
rect 24853 6352 29335 6354
rect 24853 6296 24858 6352
rect 24914 6296 29274 6352
rect 29330 6296 29335 6352
rect 24853 6294 29335 6296
rect 24853 6291 24919 6294
rect 29269 6291 29335 6294
rect 32857 6354 32923 6357
rect 34697 6354 34763 6357
rect 39520 6354 40000 6384
rect 32857 6352 40000 6354
rect 32857 6296 32862 6352
rect 32918 6296 34702 6352
rect 34758 6296 40000 6352
rect 32857 6294 40000 6296
rect 32857 6291 32923 6294
rect 34697 6291 34763 6294
rect 39520 6264 40000 6294
rect 5625 6218 5691 6221
rect 8385 6218 8451 6221
rect 5625 6216 8451 6218
rect 5625 6160 5630 6216
rect 5686 6160 8390 6216
rect 8446 6160 8451 6216
rect 5625 6158 8451 6160
rect 5625 6155 5691 6158
rect 8385 6155 8451 6158
rect 5441 6082 5507 6085
rect 7557 6082 7623 6085
rect 5441 6080 7623 6082
rect 5441 6024 5446 6080
rect 5502 6024 7562 6080
rect 7618 6024 7623 6080
rect 5441 6022 7623 6024
rect 5441 6019 5507 6022
rect 7557 6019 7623 6022
rect 24761 6082 24827 6085
rect 26969 6082 27035 6085
rect 24761 6080 27035 6082
rect 24761 6024 24766 6080
rect 24822 6024 26974 6080
rect 27030 6024 27035 6080
rect 24761 6022 27035 6024
rect 24761 6019 24827 6022
rect 26969 6019 27035 6022
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 2405 5946 2471 5949
rect 4429 5946 4495 5949
rect 2405 5944 4495 5946
rect 2405 5888 2410 5944
rect 2466 5888 4434 5944
rect 4490 5888 4495 5944
rect 2405 5886 4495 5888
rect 2405 5883 2471 5886
rect 4429 5883 4495 5886
rect 6821 5946 6887 5949
rect 9673 5946 9739 5949
rect 6821 5944 9739 5946
rect 6821 5888 6826 5944
rect 6882 5888 9678 5944
rect 9734 5888 9739 5944
rect 6821 5886 9739 5888
rect 6821 5883 6887 5886
rect 9673 5883 9739 5886
rect 16849 5946 16915 5949
rect 19333 5946 19399 5949
rect 16849 5944 19399 5946
rect 16849 5888 16854 5944
rect 16910 5888 19338 5944
rect 19394 5888 19399 5944
rect 16849 5886 19399 5888
rect 16849 5883 16915 5886
rect 19333 5883 19399 5886
rect 22001 5946 22067 5949
rect 23841 5946 23907 5949
rect 22001 5944 23907 5946
rect 22001 5888 22006 5944
rect 22062 5888 23846 5944
rect 23902 5888 23907 5944
rect 22001 5886 23907 5888
rect 22001 5883 22067 5886
rect 23841 5883 23907 5886
rect 28533 5946 28599 5949
rect 30741 5946 30807 5949
rect 28533 5944 30807 5946
rect 28533 5888 28538 5944
rect 28594 5888 30746 5944
rect 30802 5888 30807 5944
rect 28533 5886 30807 5888
rect 28533 5883 28599 5886
rect 30741 5883 30807 5886
rect 18873 5810 18939 5813
rect 20437 5810 20503 5813
rect 18873 5808 20503 5810
rect 18873 5752 18878 5808
rect 18934 5752 20442 5808
rect 20498 5752 20503 5808
rect 18873 5750 20503 5752
rect 18873 5747 18939 5750
rect 20437 5747 20503 5750
rect 26509 5810 26575 5813
rect 31937 5810 32003 5813
rect 26509 5808 32003 5810
rect 26509 5752 26514 5808
rect 26570 5752 31942 5808
rect 31998 5752 32003 5808
rect 26509 5750 32003 5752
rect 26509 5747 26575 5750
rect 31937 5747 32003 5750
rect 7281 5674 7347 5677
rect 9857 5674 9923 5677
rect 7281 5672 9923 5674
rect 7281 5616 7286 5672
rect 7342 5616 9862 5672
rect 9918 5616 9923 5672
rect 7281 5614 9923 5616
rect 7281 5611 7347 5614
rect 9857 5611 9923 5614
rect 17953 5674 18019 5677
rect 20713 5674 20779 5677
rect 17953 5672 20779 5674
rect 17953 5616 17958 5672
rect 18014 5616 20718 5672
rect 20774 5616 20779 5672
rect 17953 5614 20779 5616
rect 17953 5611 18019 5614
rect 20713 5611 20779 5614
rect 25957 5674 26023 5677
rect 29269 5674 29335 5677
rect 25957 5672 29335 5674
rect 25957 5616 25962 5672
rect 26018 5616 29274 5672
rect 29330 5616 29335 5672
rect 25957 5614 29335 5616
rect 25957 5611 26023 5614
rect 29269 5611 29335 5614
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 34928 5472 35248 5473
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 5407 35248 5408
rect 6821 5402 6887 5405
rect 8569 5402 8635 5405
rect 6821 5400 8635 5402
rect 6821 5344 6826 5400
rect 6882 5344 8574 5400
rect 8630 5344 8635 5400
rect 6821 5342 8635 5344
rect 6821 5339 6887 5342
rect 8569 5339 8635 5342
rect 12985 5402 13051 5405
rect 30649 5402 30715 5405
rect 12985 5400 30715 5402
rect 12985 5344 12990 5400
rect 13046 5344 30654 5400
rect 30710 5344 30715 5400
rect 12985 5342 30715 5344
rect 12985 5339 13051 5342
rect 30649 5339 30715 5342
rect 5441 5266 5507 5269
rect 15193 5266 15259 5269
rect 5441 5264 15259 5266
rect 5441 5208 5446 5264
rect 5502 5208 15198 5264
rect 15254 5208 15259 5264
rect 5441 5206 15259 5208
rect 5441 5203 5507 5206
rect 15193 5203 15259 5206
rect 18413 5266 18479 5269
rect 22001 5266 22067 5269
rect 24117 5266 24183 5269
rect 18413 5264 21834 5266
rect 18413 5208 18418 5264
rect 18474 5208 21834 5264
rect 18413 5206 21834 5208
rect 18413 5203 18479 5206
rect 4337 5130 4403 5133
rect 8017 5130 8083 5133
rect 10593 5130 10659 5133
rect 4337 5128 7850 5130
rect 4337 5072 4342 5128
rect 4398 5072 7850 5128
rect 4337 5070 7850 5072
rect 4337 5067 4403 5070
rect 7790 4994 7850 5070
rect 8017 5128 10659 5130
rect 8017 5072 8022 5128
rect 8078 5072 10598 5128
rect 10654 5072 10659 5128
rect 8017 5070 10659 5072
rect 8017 5067 8083 5070
rect 10593 5067 10659 5070
rect 10869 5130 10935 5133
rect 12893 5130 12959 5133
rect 10869 5128 12959 5130
rect 10869 5072 10874 5128
rect 10930 5072 12898 5128
rect 12954 5072 12959 5128
rect 10869 5070 12959 5072
rect 10869 5067 10935 5070
rect 12893 5067 12959 5070
rect 17217 5130 17283 5133
rect 19885 5130 19951 5133
rect 17217 5128 19951 5130
rect 17217 5072 17222 5128
rect 17278 5072 19890 5128
rect 19946 5072 19951 5128
rect 17217 5070 19951 5072
rect 21774 5130 21834 5206
rect 22001 5264 24183 5266
rect 22001 5208 22006 5264
rect 22062 5208 24122 5264
rect 24178 5208 24183 5264
rect 22001 5206 24183 5208
rect 22001 5203 22067 5206
rect 24117 5203 24183 5206
rect 25773 5266 25839 5269
rect 29453 5266 29519 5269
rect 25773 5264 29519 5266
rect 25773 5208 25778 5264
rect 25834 5208 29458 5264
rect 29514 5208 29519 5264
rect 25773 5206 29519 5208
rect 25773 5203 25839 5206
rect 29453 5203 29519 5206
rect 32305 5266 32371 5269
rect 34605 5266 34671 5269
rect 32305 5264 34671 5266
rect 32305 5208 32310 5264
rect 32366 5208 34610 5264
rect 34666 5208 34671 5264
rect 32305 5206 34671 5208
rect 32305 5203 32371 5206
rect 34605 5203 34671 5206
rect 24209 5130 24275 5133
rect 21774 5128 24275 5130
rect 21774 5072 24214 5128
rect 24270 5072 24275 5128
rect 21774 5070 24275 5072
rect 17217 5067 17283 5070
rect 19885 5067 19951 5070
rect 24209 5067 24275 5070
rect 35709 5130 35775 5133
rect 39520 5130 40000 5160
rect 35709 5128 40000 5130
rect 35709 5072 35714 5128
rect 35770 5072 40000 5128
rect 35709 5070 40000 5072
rect 35709 5067 35775 5070
rect 39520 5040 40000 5070
rect 12985 4994 13051 4997
rect 7790 4992 13051 4994
rect 7790 4936 12990 4992
rect 13046 4936 13051 4992
rect 7790 4934 13051 4936
rect 12985 4931 13051 4934
rect 17769 4994 17835 4997
rect 18045 4994 18111 4997
rect 19333 4994 19399 4997
rect 17769 4992 19399 4994
rect 17769 4936 17774 4992
rect 17830 4936 18050 4992
rect 18106 4936 19338 4992
rect 19394 4936 19399 4992
rect 17769 4934 19399 4936
rect 17769 4931 17835 4934
rect 18045 4931 18111 4934
rect 19333 4931 19399 4934
rect 21817 4994 21883 4997
rect 24025 4994 24091 4997
rect 24853 4994 24919 4997
rect 21817 4992 24919 4994
rect 21817 4936 21822 4992
rect 21878 4936 24030 4992
rect 24086 4936 24858 4992
rect 24914 4936 24919 4992
rect 21817 4934 24919 4936
rect 21817 4931 21883 4934
rect 24025 4931 24091 4934
rect 24853 4931 24919 4934
rect 26693 4994 26759 4997
rect 30189 4994 30255 4997
rect 26693 4992 30255 4994
rect 26693 4936 26698 4992
rect 26754 4936 30194 4992
rect 30250 4936 30255 4992
rect 26693 4934 30255 4936
rect 26693 4931 26759 4934
rect 30189 4931 30255 4934
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 8109 4858 8175 4861
rect 15009 4858 15075 4861
rect 8109 4856 15075 4858
rect 8109 4800 8114 4856
rect 8170 4800 15014 4856
rect 15070 4800 15075 4856
rect 8109 4798 15075 4800
rect 8109 4795 8175 4798
rect 15009 4795 15075 4798
rect 23657 4858 23723 4861
rect 26877 4858 26943 4861
rect 23657 4856 26943 4858
rect 23657 4800 23662 4856
rect 23718 4800 26882 4856
rect 26938 4800 26943 4856
rect 23657 4798 26943 4800
rect 23657 4795 23723 4798
rect 26877 4795 26943 4798
rect 3969 4722 4035 4725
rect 5625 4722 5691 4725
rect 3969 4720 5691 4722
rect 3969 4664 3974 4720
rect 4030 4664 5630 4720
rect 5686 4664 5691 4720
rect 3969 4662 5691 4664
rect 3969 4659 4035 4662
rect 5625 4659 5691 4662
rect 8477 4722 8543 4725
rect 16665 4722 16731 4725
rect 8477 4720 16731 4722
rect 8477 4664 8482 4720
rect 8538 4664 16670 4720
rect 16726 4664 16731 4720
rect 8477 4662 16731 4664
rect 8477 4659 8543 4662
rect 16665 4659 16731 4662
rect 18873 4722 18939 4725
rect 20437 4722 20503 4725
rect 18873 4720 20503 4722
rect 18873 4664 18878 4720
rect 18934 4664 20442 4720
rect 20498 4664 20503 4720
rect 18873 4662 20503 4664
rect 18873 4659 18939 4662
rect 20437 4659 20503 4662
rect 3877 4586 3943 4589
rect 5993 4586 6059 4589
rect 3877 4584 6059 4586
rect 3877 4528 3882 4584
rect 3938 4528 5998 4584
rect 6054 4528 6059 4584
rect 3877 4526 6059 4528
rect 3877 4523 3943 4526
rect 5993 4523 6059 4526
rect 13445 4586 13511 4589
rect 13997 4586 14063 4589
rect 13445 4584 14063 4586
rect 13445 4528 13450 4584
rect 13506 4528 14002 4584
rect 14058 4528 14063 4584
rect 13445 4526 14063 4528
rect 13445 4523 13511 4526
rect 13997 4523 14063 4526
rect 15193 4586 15259 4589
rect 31569 4586 31635 4589
rect 15193 4584 31635 4586
rect 15193 4528 15198 4584
rect 15254 4528 31574 4584
rect 31630 4528 31635 4584
rect 15193 4526 31635 4528
rect 15193 4523 15259 4526
rect 31569 4523 31635 4526
rect 9121 4450 9187 4453
rect 12617 4450 12683 4453
rect 9121 4448 12683 4450
rect 9121 4392 9126 4448
rect 9182 4392 12622 4448
rect 12678 4392 12683 4448
rect 9121 4390 12683 4392
rect 9121 4387 9187 4390
rect 12617 4387 12683 4390
rect 15469 4450 15535 4453
rect 16849 4450 16915 4453
rect 15469 4448 16915 4450
rect 15469 4392 15474 4448
rect 15530 4392 16854 4448
rect 16910 4392 16915 4448
rect 15469 4390 16915 4392
rect 15469 4387 15535 4390
rect 16849 4387 16915 4390
rect 18597 4450 18663 4453
rect 21265 4450 21331 4453
rect 18597 4448 21331 4450
rect 18597 4392 18602 4448
rect 18658 4392 21270 4448
rect 21326 4392 21331 4448
rect 18597 4390 21331 4392
rect 18597 4387 18663 4390
rect 21265 4387 21331 4390
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 34928 4384 35248 4385
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 4319 35248 4320
rect 6177 4314 6243 4317
rect 11605 4314 11671 4317
rect 32765 4314 32831 4317
rect 6177 4312 32831 4314
rect 6177 4256 6182 4312
rect 6238 4256 11610 4312
rect 11666 4256 32770 4312
rect 32826 4256 32831 4312
rect 6177 4254 32831 4256
rect 6177 4251 6243 4254
rect 11605 4251 11671 4254
rect 32765 4251 32831 4254
rect 4981 4178 5047 4181
rect 7097 4178 7163 4181
rect 4981 4176 7163 4178
rect 4981 4120 4986 4176
rect 5042 4120 7102 4176
rect 7158 4120 7163 4176
rect 4981 4118 7163 4120
rect 4981 4115 5047 4118
rect 7097 4115 7163 4118
rect 22645 4178 22711 4181
rect 25589 4178 25655 4181
rect 22645 4176 25655 4178
rect 22645 4120 22650 4176
rect 22706 4120 25594 4176
rect 25650 4120 25655 4176
rect 22645 4118 25655 4120
rect 22645 4115 22711 4118
rect 25589 4115 25655 4118
rect 9489 4042 9555 4045
rect 11237 4042 11303 4045
rect 12433 4042 12499 4045
rect 9489 4040 11303 4042
rect 9489 3984 9494 4040
rect 9550 3984 11242 4040
rect 11298 3984 11303 4040
rect 9489 3982 11303 3984
rect 9489 3979 9555 3982
rect 11237 3979 11303 3982
rect 11470 4040 12499 4042
rect 11470 3984 12438 4040
rect 12494 3984 12499 4040
rect 11470 3982 12499 3984
rect 6821 3906 6887 3909
rect 8477 3906 8543 3909
rect 11470 3906 11530 3982
rect 12433 3979 12499 3982
rect 26693 4042 26759 4045
rect 29453 4042 29519 4045
rect 26693 4040 29519 4042
rect 26693 3984 26698 4040
rect 26754 3984 29458 4040
rect 29514 3984 29519 4040
rect 26693 3982 29519 3984
rect 26693 3979 26759 3982
rect 29453 3979 29519 3982
rect 35341 4042 35407 4045
rect 39520 4042 40000 4072
rect 35341 4040 40000 4042
rect 35341 3984 35346 4040
rect 35402 3984 40000 4040
rect 35341 3982 40000 3984
rect 35341 3979 35407 3982
rect 39520 3952 40000 3982
rect 6821 3904 11530 3906
rect 6821 3848 6826 3904
rect 6882 3848 8482 3904
rect 8538 3848 11530 3904
rect 6821 3846 11530 3848
rect 11697 3906 11763 3909
rect 13905 3906 13971 3909
rect 11697 3904 13971 3906
rect 11697 3848 11702 3904
rect 11758 3848 13910 3904
rect 13966 3848 13971 3904
rect 11697 3846 13971 3848
rect 6821 3843 6887 3846
rect 8477 3843 8543 3846
rect 11697 3843 11763 3846
rect 13905 3843 13971 3846
rect 23105 3906 23171 3909
rect 24945 3906 25011 3909
rect 23105 3904 25011 3906
rect 23105 3848 23110 3904
rect 23166 3848 24950 3904
rect 25006 3848 25011 3904
rect 23105 3846 25011 3848
rect 23105 3843 23171 3846
rect 24945 3843 25011 3846
rect 28349 3906 28415 3909
rect 32305 3906 32371 3909
rect 28349 3904 32371 3906
rect 28349 3848 28354 3904
rect 28410 3848 32310 3904
rect 32366 3848 32371 3904
rect 28349 3846 32371 3848
rect 28349 3843 28415 3846
rect 32305 3843 32371 3846
rect 35985 3906 36051 3909
rect 39389 3906 39455 3909
rect 35985 3904 39455 3906
rect 35985 3848 35990 3904
rect 36046 3848 39394 3904
rect 39450 3848 39455 3904
rect 35985 3846 39455 3848
rect 35985 3843 36051 3846
rect 39389 3843 39455 3846
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 9673 3770 9739 3773
rect 15653 3770 15719 3773
rect 9673 3768 15719 3770
rect 9673 3712 9678 3768
rect 9734 3712 15658 3768
rect 15714 3712 15719 3768
rect 9673 3710 15719 3712
rect 9673 3707 9739 3710
rect 15653 3707 15719 3710
rect 17677 3770 17743 3773
rect 19425 3770 19491 3773
rect 17677 3768 19491 3770
rect 17677 3712 17682 3768
rect 17738 3712 19430 3768
rect 19486 3712 19491 3768
rect 17677 3710 19491 3712
rect 17677 3707 17743 3710
rect 19425 3707 19491 3710
rect 20069 3770 20135 3773
rect 21633 3770 21699 3773
rect 20069 3768 21699 3770
rect 20069 3712 20074 3768
rect 20130 3712 21638 3768
rect 21694 3712 21699 3768
rect 20069 3710 21699 3712
rect 20069 3707 20135 3710
rect 21633 3707 21699 3710
rect 29913 3770 29979 3773
rect 32029 3770 32095 3773
rect 29913 3768 32095 3770
rect 29913 3712 29918 3768
rect 29974 3712 32034 3768
rect 32090 3712 32095 3768
rect 29913 3710 32095 3712
rect 29913 3707 29979 3710
rect 32029 3707 32095 3710
rect 10593 3634 10659 3637
rect 17033 3634 17099 3637
rect 10593 3632 17099 3634
rect 10593 3576 10598 3632
rect 10654 3576 17038 3632
rect 17094 3576 17099 3632
rect 10593 3574 17099 3576
rect 10593 3571 10659 3574
rect 17033 3571 17099 3574
rect 17309 3634 17375 3637
rect 19149 3634 19215 3637
rect 17309 3632 19215 3634
rect 17309 3576 17314 3632
rect 17370 3576 19154 3632
rect 19210 3576 19215 3632
rect 17309 3574 19215 3576
rect 17309 3571 17375 3574
rect 19149 3571 19215 3574
rect 21357 3634 21423 3637
rect 30465 3634 30531 3637
rect 33133 3634 33199 3637
rect 21357 3632 30531 3634
rect 21357 3576 21362 3632
rect 21418 3576 30470 3632
rect 30526 3576 30531 3632
rect 21357 3574 30531 3576
rect 21357 3571 21423 3574
rect 30465 3571 30531 3574
rect 30606 3632 33199 3634
rect 30606 3576 33138 3632
rect 33194 3576 33199 3632
rect 30606 3574 33199 3576
rect 2405 3498 2471 3501
rect 4429 3498 4495 3501
rect 2405 3496 4495 3498
rect 2405 3440 2410 3496
rect 2466 3440 4434 3496
rect 4490 3440 4495 3496
rect 2405 3438 4495 3440
rect 2405 3435 2471 3438
rect 4429 3435 4495 3438
rect 5533 3498 5599 3501
rect 7005 3498 7071 3501
rect 5533 3496 7071 3498
rect 5533 3440 5538 3496
rect 5594 3440 7010 3496
rect 7066 3440 7071 3496
rect 5533 3438 7071 3440
rect 5533 3435 5599 3438
rect 7005 3435 7071 3438
rect 13997 3498 14063 3501
rect 17401 3498 17467 3501
rect 13997 3496 17467 3498
rect 13997 3440 14002 3496
rect 14058 3440 17406 3496
rect 17462 3440 17467 3496
rect 13997 3438 17467 3440
rect 13997 3435 14063 3438
rect 17401 3435 17467 3438
rect 19241 3498 19307 3501
rect 21449 3498 21515 3501
rect 19241 3496 21515 3498
rect 19241 3440 19246 3496
rect 19302 3440 21454 3496
rect 21510 3440 21515 3496
rect 19241 3438 21515 3440
rect 19241 3435 19307 3438
rect 21449 3435 21515 3438
rect 22185 3498 22251 3501
rect 24577 3498 24643 3501
rect 22185 3496 24643 3498
rect 22185 3440 22190 3496
rect 22246 3440 24582 3496
rect 24638 3440 24643 3496
rect 22185 3438 24643 3440
rect 22185 3435 22251 3438
rect 24577 3435 24643 3438
rect 28441 3498 28507 3501
rect 30606 3498 30666 3574
rect 33133 3571 33199 3574
rect 28441 3496 30666 3498
rect 28441 3440 28446 3496
rect 28502 3440 30666 3496
rect 28441 3438 30666 3440
rect 28441 3435 28507 3438
rect 19057 3362 19123 3365
rect 22737 3362 22803 3365
rect 19057 3360 22803 3362
rect 19057 3304 19062 3360
rect 19118 3304 22742 3360
rect 22798 3304 22803 3360
rect 19057 3302 22803 3304
rect 19057 3299 19123 3302
rect 22737 3299 22803 3302
rect 30925 3362 30991 3365
rect 34237 3362 34303 3365
rect 30925 3360 34303 3362
rect 30925 3304 30930 3360
rect 30986 3304 34242 3360
rect 34298 3304 34303 3360
rect 30925 3302 34303 3304
rect 30925 3299 30991 3302
rect 34237 3299 34303 3302
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 34928 3296 35248 3297
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 3231 35248 3232
rect 9765 3226 9831 3229
rect 10225 3226 10291 3229
rect 8894 3224 10291 3226
rect 8894 3168 9770 3224
rect 9826 3168 10230 3224
rect 10286 3168 10291 3224
rect 8894 3166 10291 3168
rect 4613 3090 4679 3093
rect 8894 3090 8954 3166
rect 9765 3163 9831 3166
rect 10225 3163 10291 3166
rect 14273 3226 14339 3229
rect 17677 3226 17743 3229
rect 14273 3224 17743 3226
rect 14273 3168 14278 3224
rect 14334 3168 17682 3224
rect 17738 3168 17743 3224
rect 14273 3166 17743 3168
rect 14273 3163 14339 3166
rect 17677 3163 17743 3166
rect 4613 3088 8954 3090
rect 4613 3032 4618 3088
rect 4674 3032 8954 3088
rect 4613 3030 8954 3032
rect 9029 3090 9095 3093
rect 18873 3090 18939 3093
rect 23841 3090 23907 3093
rect 9029 3088 16130 3090
rect 9029 3032 9034 3088
rect 9090 3032 16130 3088
rect 9029 3030 16130 3032
rect 4613 3027 4679 3030
rect 9029 3027 9095 3030
rect 8937 2954 9003 2957
rect 15837 2954 15903 2957
rect 8937 2952 15903 2954
rect 8937 2896 8942 2952
rect 8998 2896 15842 2952
rect 15898 2896 15903 2952
rect 8937 2894 15903 2896
rect 16070 2954 16130 3030
rect 18873 3088 23907 3090
rect 18873 3032 18878 3088
rect 18934 3032 23846 3088
rect 23902 3032 23907 3088
rect 18873 3030 23907 3032
rect 18873 3027 18939 3030
rect 23841 3027 23907 3030
rect 27245 3090 27311 3093
rect 30833 3090 30899 3093
rect 32949 3090 33015 3093
rect 35157 3090 35223 3093
rect 27245 3088 35223 3090
rect 27245 3032 27250 3088
rect 27306 3032 30838 3088
rect 30894 3032 32954 3088
rect 33010 3032 35162 3088
rect 35218 3032 35223 3088
rect 27245 3030 35223 3032
rect 27245 3027 27311 3030
rect 30833 3027 30899 3030
rect 32949 3027 33015 3030
rect 35157 3027 35223 3030
rect 29545 2954 29611 2957
rect 37181 2954 37247 2957
rect 16070 2952 37247 2954
rect 16070 2896 29550 2952
rect 29606 2896 37186 2952
rect 37242 2896 37247 2952
rect 16070 2894 37247 2896
rect 8937 2891 9003 2894
rect 15837 2891 15903 2894
rect 29545 2891 29611 2894
rect 37181 2891 37247 2894
rect 565 2818 631 2821
rect 4061 2818 4127 2821
rect 565 2816 4127 2818
rect 565 2760 570 2816
rect 626 2760 4066 2816
rect 4122 2760 4127 2816
rect 565 2758 4127 2760
rect 565 2755 631 2758
rect 4061 2755 4127 2758
rect 6085 2818 6151 2821
rect 8661 2818 8727 2821
rect 6085 2816 8727 2818
rect 6085 2760 6090 2816
rect 6146 2760 8666 2816
rect 8722 2760 8727 2816
rect 6085 2758 8727 2760
rect 6085 2755 6151 2758
rect 8661 2755 8727 2758
rect 13077 2818 13143 2821
rect 16113 2818 16179 2821
rect 13077 2816 16179 2818
rect 13077 2760 13082 2816
rect 13138 2760 16118 2816
rect 16174 2760 16179 2816
rect 13077 2758 16179 2760
rect 13077 2755 13143 2758
rect 16113 2755 16179 2758
rect 31569 2818 31635 2821
rect 34789 2818 34855 2821
rect 31569 2816 34855 2818
rect 31569 2760 31574 2816
rect 31630 2760 34794 2816
rect 34850 2760 34855 2816
rect 31569 2758 34855 2760
rect 31569 2755 31635 2758
rect 34789 2755 34855 2758
rect 35750 2756 35756 2820
rect 35820 2818 35826 2820
rect 39520 2818 40000 2848
rect 35820 2758 40000 2818
rect 35820 2756 35826 2758
rect 19568 2752 19888 2753
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 39520 2728 40000 2758
rect 19568 2687 19888 2688
rect 30649 2682 30715 2685
rect 36997 2682 37063 2685
rect 30649 2680 37063 2682
rect 30649 2624 30654 2680
rect 30710 2624 37002 2680
rect 37058 2624 37063 2680
rect 30649 2622 37063 2624
rect 30649 2619 30715 2622
rect 36997 2619 37063 2622
rect 12065 2546 12131 2549
rect 34881 2546 34947 2549
rect 36077 2546 36143 2549
rect 12065 2544 36143 2546
rect 12065 2488 12070 2544
rect 12126 2488 34886 2544
rect 34942 2488 36082 2544
rect 36138 2488 36143 2544
rect 12065 2486 36143 2488
rect 12065 2483 12131 2486
rect 34881 2483 34947 2486
rect 36077 2483 36143 2486
rect 9213 2410 9279 2413
rect 17217 2410 17283 2413
rect 9213 2408 17283 2410
rect 9213 2352 9218 2408
rect 9274 2352 17222 2408
rect 17278 2352 17283 2408
rect 9213 2350 17283 2352
rect 9213 2347 9279 2350
rect 17217 2347 17283 2350
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 34928 2208 35248 2209
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2143 35248 2144
rect 10225 2138 10291 2141
rect 29453 2138 29519 2141
rect 10225 2136 29519 2138
rect 10225 2080 10230 2136
rect 10286 2080 29458 2136
rect 29514 2080 29519 2136
rect 10225 2078 29519 2080
rect 10225 2075 10291 2078
rect 29453 2075 29519 2078
rect 15837 2002 15903 2005
rect 34973 2002 35039 2005
rect 15837 2000 35039 2002
rect 15837 1944 15842 2000
rect 15898 1944 34978 2000
rect 35034 1944 35039 2000
rect 15837 1942 35039 1944
rect 15837 1939 15903 1942
rect 34973 1939 35039 1942
rect 7097 1866 7163 1869
rect 21817 1866 21883 1869
rect 33869 1866 33935 1869
rect 7097 1864 33935 1866
rect 7097 1808 7102 1864
rect 7158 1808 21822 1864
rect 21878 1808 33874 1864
rect 33930 1808 33935 1864
rect 7097 1806 33935 1808
rect 7097 1803 7163 1806
rect 21817 1803 21883 1806
rect 33869 1803 33935 1806
rect 35801 1730 35867 1733
rect 39520 1730 40000 1760
rect 35801 1728 40000 1730
rect 35801 1672 35806 1728
rect 35862 1672 40000 1728
rect 35801 1670 40000 1672
rect 35801 1667 35867 1670
rect 39520 1640 40000 1670
rect 7189 1458 7255 1461
rect 11053 1458 11119 1461
rect 7189 1456 11119 1458
rect 7189 1400 7194 1456
rect 7250 1400 11058 1456
rect 11114 1400 11119 1456
rect 7189 1398 11119 1400
rect 7189 1395 7255 1398
rect 11053 1395 11119 1398
rect 35249 642 35315 645
rect 39520 642 40000 672
rect 35249 640 40000 642
rect 35249 584 35254 640
rect 35310 584 40000 640
rect 35249 582 40000 584
rect 35249 579 35315 582
rect 39520 552 40000 582
<< via3 >>
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 34936 33756 35000 33760
rect 34936 33700 34940 33756
rect 34940 33700 34996 33756
rect 34996 33700 35000 33756
rect 34936 33696 35000 33700
rect 35016 33756 35080 33760
rect 35016 33700 35020 33756
rect 35020 33700 35076 33756
rect 35076 33700 35080 33756
rect 35016 33696 35080 33700
rect 35096 33756 35160 33760
rect 35096 33700 35100 33756
rect 35100 33700 35156 33756
rect 35156 33700 35160 33756
rect 35096 33696 35160 33700
rect 35176 33756 35240 33760
rect 35176 33700 35180 33756
rect 35180 33700 35236 33756
rect 35236 33700 35240 33756
rect 35176 33696 35240 33700
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 34936 32668 35000 32672
rect 34936 32612 34940 32668
rect 34940 32612 34996 32668
rect 34996 32612 35000 32668
rect 34936 32608 35000 32612
rect 35016 32668 35080 32672
rect 35016 32612 35020 32668
rect 35020 32612 35076 32668
rect 35076 32612 35080 32668
rect 35016 32608 35080 32612
rect 35096 32668 35160 32672
rect 35096 32612 35100 32668
rect 35100 32612 35156 32668
rect 35156 32612 35160 32668
rect 35096 32608 35160 32612
rect 35176 32668 35240 32672
rect 35176 32612 35180 32668
rect 35180 32612 35236 32668
rect 35236 32612 35240 32668
rect 35176 32608 35240 32612
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 34936 31580 35000 31584
rect 34936 31524 34940 31580
rect 34940 31524 34996 31580
rect 34996 31524 35000 31580
rect 34936 31520 35000 31524
rect 35016 31580 35080 31584
rect 35016 31524 35020 31580
rect 35020 31524 35076 31580
rect 35076 31524 35080 31580
rect 35016 31520 35080 31524
rect 35096 31580 35160 31584
rect 35096 31524 35100 31580
rect 35100 31524 35156 31580
rect 35156 31524 35160 31580
rect 35096 31520 35160 31524
rect 35176 31580 35240 31584
rect 35176 31524 35180 31580
rect 35180 31524 35236 31580
rect 35236 31524 35240 31580
rect 35176 31520 35240 31524
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 34936 30492 35000 30496
rect 34936 30436 34940 30492
rect 34940 30436 34996 30492
rect 34996 30436 35000 30492
rect 34936 30432 35000 30436
rect 35016 30492 35080 30496
rect 35016 30436 35020 30492
rect 35020 30436 35076 30492
rect 35076 30436 35080 30492
rect 35016 30432 35080 30436
rect 35096 30492 35160 30496
rect 35096 30436 35100 30492
rect 35100 30436 35156 30492
rect 35156 30436 35160 30492
rect 35096 30432 35160 30436
rect 35176 30492 35240 30496
rect 35176 30436 35180 30492
rect 35180 30436 35236 30492
rect 35236 30436 35240 30492
rect 35176 30432 35240 30436
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 34936 29404 35000 29408
rect 34936 29348 34940 29404
rect 34940 29348 34996 29404
rect 34996 29348 35000 29404
rect 34936 29344 35000 29348
rect 35016 29404 35080 29408
rect 35016 29348 35020 29404
rect 35020 29348 35076 29404
rect 35076 29348 35080 29404
rect 35016 29344 35080 29348
rect 35096 29404 35160 29408
rect 35096 29348 35100 29404
rect 35100 29348 35156 29404
rect 35156 29348 35160 29404
rect 35096 29344 35160 29348
rect 35176 29404 35240 29408
rect 35176 29348 35180 29404
rect 35180 29348 35236 29404
rect 35236 29348 35240 29404
rect 35176 29344 35240 29348
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 34936 28316 35000 28320
rect 34936 28260 34940 28316
rect 34940 28260 34996 28316
rect 34996 28260 35000 28316
rect 34936 28256 35000 28260
rect 35016 28316 35080 28320
rect 35016 28260 35020 28316
rect 35020 28260 35076 28316
rect 35076 28260 35080 28316
rect 35016 28256 35080 28260
rect 35096 28316 35160 28320
rect 35096 28260 35100 28316
rect 35100 28260 35156 28316
rect 35156 28260 35160 28316
rect 35096 28256 35160 28260
rect 35176 28316 35240 28320
rect 35176 28260 35180 28316
rect 35180 28260 35236 28316
rect 35236 28260 35240 28316
rect 35176 28256 35240 28260
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 34936 27228 35000 27232
rect 34936 27172 34940 27228
rect 34940 27172 34996 27228
rect 34996 27172 35000 27228
rect 34936 27168 35000 27172
rect 35016 27228 35080 27232
rect 35016 27172 35020 27228
rect 35020 27172 35076 27228
rect 35076 27172 35080 27228
rect 35016 27168 35080 27172
rect 35096 27228 35160 27232
rect 35096 27172 35100 27228
rect 35100 27172 35156 27228
rect 35156 27172 35160 27228
rect 35096 27168 35160 27172
rect 35176 27228 35240 27232
rect 35176 27172 35180 27228
rect 35180 27172 35236 27228
rect 35236 27172 35240 27228
rect 35176 27168 35240 27172
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 34936 26140 35000 26144
rect 34936 26084 34940 26140
rect 34940 26084 34996 26140
rect 34996 26084 35000 26140
rect 34936 26080 35000 26084
rect 35016 26140 35080 26144
rect 35016 26084 35020 26140
rect 35020 26084 35076 26140
rect 35076 26084 35080 26140
rect 35016 26080 35080 26084
rect 35096 26140 35160 26144
rect 35096 26084 35100 26140
rect 35100 26084 35156 26140
rect 35156 26084 35160 26140
rect 35096 26080 35160 26084
rect 35176 26140 35240 26144
rect 35176 26084 35180 26140
rect 35180 26084 35236 26140
rect 35236 26084 35240 26140
rect 35176 26080 35240 26084
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 34936 25052 35000 25056
rect 34936 24996 34940 25052
rect 34940 24996 34996 25052
rect 34996 24996 35000 25052
rect 34936 24992 35000 24996
rect 35016 25052 35080 25056
rect 35016 24996 35020 25052
rect 35020 24996 35076 25052
rect 35076 24996 35080 25052
rect 35016 24992 35080 24996
rect 35096 25052 35160 25056
rect 35096 24996 35100 25052
rect 35100 24996 35156 25052
rect 35156 24996 35160 25052
rect 35096 24992 35160 24996
rect 35176 25052 35240 25056
rect 35176 24996 35180 25052
rect 35180 24996 35236 25052
rect 35236 24996 35240 25052
rect 35176 24992 35240 24996
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 34936 23964 35000 23968
rect 34936 23908 34940 23964
rect 34940 23908 34996 23964
rect 34996 23908 35000 23964
rect 34936 23904 35000 23908
rect 35016 23964 35080 23968
rect 35016 23908 35020 23964
rect 35020 23908 35076 23964
rect 35076 23908 35080 23964
rect 35016 23904 35080 23908
rect 35096 23964 35160 23968
rect 35096 23908 35100 23964
rect 35100 23908 35156 23964
rect 35156 23908 35160 23964
rect 35096 23904 35160 23908
rect 35176 23964 35240 23968
rect 35176 23908 35180 23964
rect 35180 23908 35236 23964
rect 35236 23908 35240 23964
rect 35176 23904 35240 23908
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 34936 22876 35000 22880
rect 34936 22820 34940 22876
rect 34940 22820 34996 22876
rect 34996 22820 35000 22876
rect 34936 22816 35000 22820
rect 35016 22876 35080 22880
rect 35016 22820 35020 22876
rect 35020 22820 35076 22876
rect 35076 22820 35080 22876
rect 35016 22816 35080 22820
rect 35096 22876 35160 22880
rect 35096 22820 35100 22876
rect 35100 22820 35156 22876
rect 35156 22820 35160 22876
rect 35096 22816 35160 22820
rect 35176 22876 35240 22880
rect 35176 22820 35180 22876
rect 35180 22820 35236 22876
rect 35236 22820 35240 22876
rect 35176 22816 35240 22820
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 34936 21788 35000 21792
rect 34936 21732 34940 21788
rect 34940 21732 34996 21788
rect 34996 21732 35000 21788
rect 34936 21728 35000 21732
rect 35016 21788 35080 21792
rect 35016 21732 35020 21788
rect 35020 21732 35076 21788
rect 35076 21732 35080 21788
rect 35016 21728 35080 21732
rect 35096 21788 35160 21792
rect 35096 21732 35100 21788
rect 35100 21732 35156 21788
rect 35156 21732 35160 21788
rect 35096 21728 35160 21732
rect 35176 21788 35240 21792
rect 35176 21732 35180 21788
rect 35180 21732 35236 21788
rect 35236 21732 35240 21788
rect 35176 21728 35240 21732
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 34936 20700 35000 20704
rect 34936 20644 34940 20700
rect 34940 20644 34996 20700
rect 34996 20644 35000 20700
rect 34936 20640 35000 20644
rect 35016 20700 35080 20704
rect 35016 20644 35020 20700
rect 35020 20644 35076 20700
rect 35076 20644 35080 20700
rect 35016 20640 35080 20644
rect 35096 20700 35160 20704
rect 35096 20644 35100 20700
rect 35100 20644 35156 20700
rect 35156 20644 35160 20700
rect 35096 20640 35160 20644
rect 35176 20700 35240 20704
rect 35176 20644 35180 20700
rect 35180 20644 35236 20700
rect 35236 20644 35240 20700
rect 35176 20640 35240 20644
rect 35756 20436 35820 20500
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 34936 19612 35000 19616
rect 34936 19556 34940 19612
rect 34940 19556 34996 19612
rect 34996 19556 35000 19612
rect 34936 19552 35000 19556
rect 35016 19612 35080 19616
rect 35016 19556 35020 19612
rect 35020 19556 35076 19612
rect 35076 19556 35080 19612
rect 35016 19552 35080 19556
rect 35096 19612 35160 19616
rect 35096 19556 35100 19612
rect 35100 19556 35156 19612
rect 35156 19556 35160 19612
rect 35096 19552 35160 19556
rect 35176 19612 35240 19616
rect 35176 19556 35180 19612
rect 35180 19556 35236 19612
rect 35236 19556 35240 19612
rect 35176 19552 35240 19556
rect 35572 19272 35636 19276
rect 35572 19216 35622 19272
rect 35622 19216 35636 19272
rect 35572 19212 35636 19216
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 34936 18524 35000 18528
rect 34936 18468 34940 18524
rect 34940 18468 34996 18524
rect 34996 18468 35000 18524
rect 34936 18464 35000 18468
rect 35016 18524 35080 18528
rect 35016 18468 35020 18524
rect 35020 18468 35076 18524
rect 35076 18468 35080 18524
rect 35016 18464 35080 18468
rect 35096 18524 35160 18528
rect 35096 18468 35100 18524
rect 35100 18468 35156 18524
rect 35156 18468 35160 18524
rect 35096 18464 35160 18468
rect 35176 18524 35240 18528
rect 35176 18468 35180 18524
rect 35180 18468 35236 18524
rect 35236 18468 35240 18524
rect 35176 18464 35240 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 34936 17436 35000 17440
rect 34936 17380 34940 17436
rect 34940 17380 34996 17436
rect 34996 17380 35000 17436
rect 34936 17376 35000 17380
rect 35016 17436 35080 17440
rect 35016 17380 35020 17436
rect 35020 17380 35076 17436
rect 35076 17380 35080 17436
rect 35016 17376 35080 17380
rect 35096 17436 35160 17440
rect 35096 17380 35100 17436
rect 35100 17380 35156 17436
rect 35156 17380 35160 17436
rect 35096 17376 35160 17380
rect 35176 17436 35240 17440
rect 35176 17380 35180 17436
rect 35180 17380 35236 17436
rect 35236 17380 35240 17436
rect 35176 17376 35240 17380
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 34936 16348 35000 16352
rect 34936 16292 34940 16348
rect 34940 16292 34996 16348
rect 34996 16292 35000 16348
rect 34936 16288 35000 16292
rect 35016 16348 35080 16352
rect 35016 16292 35020 16348
rect 35020 16292 35076 16348
rect 35076 16292 35080 16348
rect 35016 16288 35080 16292
rect 35096 16348 35160 16352
rect 35096 16292 35100 16348
rect 35100 16292 35156 16348
rect 35156 16292 35160 16348
rect 35096 16288 35160 16292
rect 35176 16348 35240 16352
rect 35176 16292 35180 16348
rect 35180 16292 35236 16348
rect 35236 16292 35240 16348
rect 35176 16288 35240 16292
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 34936 15260 35000 15264
rect 34936 15204 34940 15260
rect 34940 15204 34996 15260
rect 34996 15204 35000 15260
rect 34936 15200 35000 15204
rect 35016 15260 35080 15264
rect 35016 15204 35020 15260
rect 35020 15204 35076 15260
rect 35076 15204 35080 15260
rect 35016 15200 35080 15204
rect 35096 15260 35160 15264
rect 35096 15204 35100 15260
rect 35100 15204 35156 15260
rect 35156 15204 35160 15260
rect 35096 15200 35160 15204
rect 35176 15260 35240 15264
rect 35176 15204 35180 15260
rect 35180 15204 35236 15260
rect 35236 15204 35240 15260
rect 35176 15200 35240 15204
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 34936 14172 35000 14176
rect 34936 14116 34940 14172
rect 34940 14116 34996 14172
rect 34996 14116 35000 14172
rect 34936 14112 35000 14116
rect 35016 14172 35080 14176
rect 35016 14116 35020 14172
rect 35020 14116 35076 14172
rect 35076 14116 35080 14172
rect 35016 14112 35080 14116
rect 35096 14172 35160 14176
rect 35096 14116 35100 14172
rect 35100 14116 35156 14172
rect 35156 14116 35160 14172
rect 35096 14112 35160 14116
rect 35176 14172 35240 14176
rect 35176 14116 35180 14172
rect 35180 14116 35236 14172
rect 35236 14116 35240 14172
rect 35176 14112 35240 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 34936 13084 35000 13088
rect 34936 13028 34940 13084
rect 34940 13028 34996 13084
rect 34996 13028 35000 13084
rect 34936 13024 35000 13028
rect 35016 13084 35080 13088
rect 35016 13028 35020 13084
rect 35020 13028 35076 13084
rect 35076 13028 35080 13084
rect 35016 13024 35080 13028
rect 35096 13084 35160 13088
rect 35096 13028 35100 13084
rect 35100 13028 35156 13084
rect 35156 13028 35160 13084
rect 35096 13024 35160 13028
rect 35176 13084 35240 13088
rect 35176 13028 35180 13084
rect 35180 13028 35236 13084
rect 35236 13028 35240 13084
rect 35176 13024 35240 13028
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 34936 11996 35000 12000
rect 34936 11940 34940 11996
rect 34940 11940 34996 11996
rect 34996 11940 35000 11996
rect 34936 11936 35000 11940
rect 35016 11996 35080 12000
rect 35016 11940 35020 11996
rect 35020 11940 35076 11996
rect 35076 11940 35080 11996
rect 35016 11936 35080 11940
rect 35096 11996 35160 12000
rect 35096 11940 35100 11996
rect 35100 11940 35156 11996
rect 35156 11940 35160 11996
rect 35096 11936 35160 11940
rect 35176 11996 35240 12000
rect 35176 11940 35180 11996
rect 35180 11940 35236 11996
rect 35236 11940 35240 11996
rect 35176 11936 35240 11940
rect 35572 11732 35636 11796
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 34936 10908 35000 10912
rect 34936 10852 34940 10908
rect 34940 10852 34996 10908
rect 34996 10852 35000 10908
rect 34936 10848 35000 10852
rect 35016 10908 35080 10912
rect 35016 10852 35020 10908
rect 35020 10852 35076 10908
rect 35076 10852 35080 10908
rect 35016 10848 35080 10852
rect 35096 10908 35160 10912
rect 35096 10852 35100 10908
rect 35100 10852 35156 10908
rect 35156 10852 35160 10908
rect 35096 10848 35160 10852
rect 35176 10908 35240 10912
rect 35176 10852 35180 10908
rect 35180 10852 35236 10908
rect 35236 10852 35240 10908
rect 35176 10848 35240 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 34936 9820 35000 9824
rect 34936 9764 34940 9820
rect 34940 9764 34996 9820
rect 34996 9764 35000 9820
rect 34936 9760 35000 9764
rect 35016 9820 35080 9824
rect 35016 9764 35020 9820
rect 35020 9764 35076 9820
rect 35076 9764 35080 9820
rect 35016 9760 35080 9764
rect 35096 9820 35160 9824
rect 35096 9764 35100 9820
rect 35100 9764 35156 9820
rect 35156 9764 35160 9820
rect 35096 9760 35160 9764
rect 35176 9820 35240 9824
rect 35176 9764 35180 9820
rect 35180 9764 35236 9820
rect 35236 9764 35240 9820
rect 35176 9760 35240 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 34936 8732 35000 8736
rect 34936 8676 34940 8732
rect 34940 8676 34996 8732
rect 34996 8676 35000 8732
rect 34936 8672 35000 8676
rect 35016 8732 35080 8736
rect 35016 8676 35020 8732
rect 35020 8676 35076 8732
rect 35076 8676 35080 8732
rect 35016 8672 35080 8676
rect 35096 8732 35160 8736
rect 35096 8676 35100 8732
rect 35100 8676 35156 8732
rect 35156 8676 35160 8732
rect 35096 8672 35160 8676
rect 35176 8732 35240 8736
rect 35176 8676 35180 8732
rect 35180 8676 35236 8732
rect 35236 8676 35240 8732
rect 35176 8672 35240 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 34936 7644 35000 7648
rect 34936 7588 34940 7644
rect 34940 7588 34996 7644
rect 34996 7588 35000 7644
rect 34936 7584 35000 7588
rect 35016 7644 35080 7648
rect 35016 7588 35020 7644
rect 35020 7588 35076 7644
rect 35076 7588 35080 7644
rect 35016 7584 35080 7588
rect 35096 7644 35160 7648
rect 35096 7588 35100 7644
rect 35100 7588 35156 7644
rect 35156 7588 35160 7644
rect 35096 7584 35160 7588
rect 35176 7644 35240 7648
rect 35176 7588 35180 7644
rect 35180 7588 35236 7644
rect 35236 7588 35240 7644
rect 35176 7584 35240 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 34936 6556 35000 6560
rect 34936 6500 34940 6556
rect 34940 6500 34996 6556
rect 34996 6500 35000 6556
rect 34936 6496 35000 6500
rect 35016 6556 35080 6560
rect 35016 6500 35020 6556
rect 35020 6500 35076 6556
rect 35076 6500 35080 6556
rect 35016 6496 35080 6500
rect 35096 6556 35160 6560
rect 35096 6500 35100 6556
rect 35100 6500 35156 6556
rect 35156 6500 35160 6556
rect 35096 6496 35160 6500
rect 35176 6556 35240 6560
rect 35176 6500 35180 6556
rect 35180 6500 35236 6556
rect 35236 6500 35240 6556
rect 35176 6496 35240 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 34936 5468 35000 5472
rect 34936 5412 34940 5468
rect 34940 5412 34996 5468
rect 34996 5412 35000 5468
rect 34936 5408 35000 5412
rect 35016 5468 35080 5472
rect 35016 5412 35020 5468
rect 35020 5412 35076 5468
rect 35076 5412 35080 5468
rect 35016 5408 35080 5412
rect 35096 5468 35160 5472
rect 35096 5412 35100 5468
rect 35100 5412 35156 5468
rect 35156 5412 35160 5468
rect 35096 5408 35160 5412
rect 35176 5468 35240 5472
rect 35176 5412 35180 5468
rect 35180 5412 35236 5468
rect 35236 5412 35240 5468
rect 35176 5408 35240 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 34936 4380 35000 4384
rect 34936 4324 34940 4380
rect 34940 4324 34996 4380
rect 34996 4324 35000 4380
rect 34936 4320 35000 4324
rect 35016 4380 35080 4384
rect 35016 4324 35020 4380
rect 35020 4324 35076 4380
rect 35076 4324 35080 4380
rect 35016 4320 35080 4324
rect 35096 4380 35160 4384
rect 35096 4324 35100 4380
rect 35100 4324 35156 4380
rect 35156 4324 35160 4380
rect 35096 4320 35160 4324
rect 35176 4380 35240 4384
rect 35176 4324 35180 4380
rect 35180 4324 35236 4380
rect 35236 4324 35240 4380
rect 35176 4320 35240 4324
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 34936 3292 35000 3296
rect 34936 3236 34940 3292
rect 34940 3236 34996 3292
rect 34996 3236 35000 3292
rect 34936 3232 35000 3236
rect 35016 3292 35080 3296
rect 35016 3236 35020 3292
rect 35020 3236 35076 3292
rect 35076 3236 35080 3292
rect 35016 3232 35080 3236
rect 35096 3292 35160 3296
rect 35096 3236 35100 3292
rect 35100 3236 35156 3292
rect 35156 3236 35160 3292
rect 35096 3232 35160 3236
rect 35176 3292 35240 3296
rect 35176 3236 35180 3292
rect 35180 3236 35236 3292
rect 35236 3236 35240 3292
rect 35176 3232 35240 3236
rect 35756 2756 35820 2820
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 34936 2204 35000 2208
rect 34936 2148 34940 2204
rect 34940 2148 34996 2204
rect 34996 2148 35000 2204
rect 34936 2144 35000 2148
rect 35016 2204 35080 2208
rect 35016 2148 35020 2204
rect 35020 2148 35076 2204
rect 35076 2148 35080 2204
rect 35016 2144 35080 2148
rect 35096 2204 35160 2208
rect 35096 2148 35100 2204
rect 35100 2148 35156 2204
rect 35156 2148 35160 2204
rect 35096 2144 35160 2148
rect 35176 2204 35240 2208
rect 35176 2148 35180 2204
rect 35180 2148 35236 2204
rect 35236 2148 35240 2204
rect 35176 2144 35240 2148
<< metal4 >>
rect 4208 37024 4528 37584
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2128 4528 2144
rect 19568 37568 19888 37584
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 36480 19888 37504
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 35392 19888 36416
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 34304 19888 35328
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 33216 19888 34240
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 31040 19888 32064
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 28864 19888 29888
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 27776 19888 28800
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 26688 19888 27712
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 25600 19888 26624
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 24512 19888 25536
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20160 19888 21184
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2128 19888 2688
rect 34928 37024 35248 37584
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 35936 35248 36960
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 34848 35248 35872
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 33760 35248 34784
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 32672 35248 33696
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 31584 35248 32608
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 30496 35248 31520
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 29408 35248 30432
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 28320 35248 29344
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 27232 35248 28256
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 26144 35248 27168
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 25056 35248 26080
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 23968 35248 24992
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 22880 35248 23904
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 21792 35248 22816
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 20704 35248 21728
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 19616 35248 20640
rect 35755 20500 35821 20501
rect 35755 20436 35756 20500
rect 35820 20436 35821 20500
rect 35755 20435 35821 20436
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 18528 35248 19552
rect 35571 19276 35637 19277
rect 35571 19212 35572 19276
rect 35636 19212 35637 19276
rect 35571 19211 35637 19212
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 17440 35248 18464
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 16352 35248 17376
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 15264 35248 16288
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 14176 35248 15200
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 13088 35248 14112
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 12000 35248 13024
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 10912 35248 11936
rect 35574 11797 35634 19211
rect 35571 11796 35637 11797
rect 35571 11732 35572 11796
rect 35636 11732 35637 11796
rect 35571 11731 35637 11732
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 9824 35248 10848
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 8736 35248 9760
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 7648 35248 8672
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 6560 35248 7584
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 5472 35248 6496
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 4384 35248 5408
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 3296 35248 4320
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 2208 35248 3232
rect 35758 2821 35818 20435
rect 35755 2820 35821 2821
rect 35755 2756 35756 2820
rect 35820 2756 35821 2820
rect 35755 2755 35821 2756
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2128 35248 2144
use scs8hd_fill_2  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_9
timestamp 1586364061
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2116 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
timestamp 1586364061
transform 1 0 1748 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
timestamp 1586364061
transform 1 0 1564 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_13 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2300 0 -1 2720
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_1_30
timestamp 1586364061
transform 1 0 3864 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_26
timestamp 1586364061
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
timestamp 1586364061
transform 1 0 3680 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
timestamp 1586364061
transform 1 0 4048 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_130 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1586364061
transform 1 0 5980 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_51
timestamp 1586364061
transform 1 0 5796 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
timestamp 1586364061
transform 1 0 6348 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_55
timestamp 1586364061
transform 1 0 6164 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_59
timestamp 1586364061
transform 1 0 6532 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
timestamp 1586364061
transform 1 0 6900 0 1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_82
timestamp 1586364061
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_76
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
timestamp 1586364061
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__69__A
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 222 592
use scs8hd_or2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 498 592
use scs8hd_fill_1  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9844 0 -1 2720
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9384 0 1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_0_104
timestamp 1586364061
transform 1 0 10672 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_109
timestamp 1586364061
transform 1 0 11132 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_108
timestamp 1586364061
transform 1 0 11040 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_113
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11316 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _70_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_117
timestamp 1586364061
transform 1 0 11868 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__70__A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_131
timestamp 1586364061
transform 1 0 13156 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_127
timestamp 1586364061
transform 1 0 12788 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13340 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 12972 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 13708 0 1 2720
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12880 0 -1 2720
box -38 -48 1786 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13892 0 1 2720
box -38 -48 2246 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16284 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 16652 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_163
timestamp 1586364061
transform 1 0 16100 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_167
timestamp 1586364061
transform 1 0 16468 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 17388 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_175
timestamp 1586364061
transform 1 0 17204 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_179
timestamp 1586364061
transform 1 0 17572 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_183
timestamp 1586364061
transform 1 0 17940 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 18216 0 1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_194
timestamp 1586364061
transform 1 0 18952 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_190
timestamp 1586364061
transform 1 0 18584 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 18768 0 1 2720
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19320 0 1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18584 0 -1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_0_209
timestamp 1586364061
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_221
timestamp 1586364061
transform 1 0 21436 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_217
timestamp 1586364061
transform 1 0 21068 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 21252 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21620 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_1_234
timestamp 1586364061
transform 1 0 22632 0 1 2720
box -38 -48 406 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21804 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 23092 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_237
timestamp 1586364061
transform 1 0 22908 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_241
timestamp 1586364061
transform 1 0 23276 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_245
timestamp 1586364061
transform 1 0 23644 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
timestamp 1586364061
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
timestamp 1586364061
transform 1 0 24288 0 -1 2720
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 26036 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 25668 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_271
timestamp 1586364061
transform 1 0 26036 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_264
timestamp 1586364061
transform 1 0 25392 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_273
timestamp 1586364061
transform 1 0 26220 0 1 2720
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 26588 0 1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 27140 0 -1 2720
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
timestamp 1586364061
transform 1 0 26404 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 26588 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 28520 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_275
timestamp 1586364061
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_280
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_296
timestamp 1586364061
transform 1 0 28336 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 28980 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 29072 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_302
timestamp 1586364061
transform 1 0 28888 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_300
timestamp 1586364061
transform 1 0 28704 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 29440 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_306
timestamp 1586364061
transform 1 0 29256 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_306
timestamp 1586364061
transform 1 0 29256 0 1 2720
box -38 -48 314 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 29532 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_322
timestamp 1586364061
transform 1 0 30728 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_318
timestamp 1586364061
transform 1 0 30360 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_311
timestamp 1586364061
transform 1 0 29716 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 30544 0 1 2720
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 29992 0 -1 2720
box -38 -48 1786 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 31096 0 1 2720
box -38 -48 2246 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 32752 0 -1 2720
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 30912 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 32292 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 31924 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_333
timestamp 1586364061
transform 1 0 31740 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_337
timestamp 1586364061
transform 1 0 32108 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_342
timestamp 1586364061
transform 1 0 32568 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_354
timestamp 1586364061
transform 1 0 33672 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_350
timestamp 1586364061
transform 1 0 33304 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 33856 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 33488 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_362
timestamp 1586364061
transform 1 0 34408 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_358
timestamp 1586364061
transform 1 0 34040 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_363
timestamp 1586364061
transform 1 0 34500 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 34224 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 34776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 34592 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 34868 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_0_368
timestamp 1586364061
transform 1 0 34960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 35144 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_376
timestamp 1586364061
transform 1 0 35696 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_382
timestamp 1586364061
transform 1 0 36248 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 36432 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 35880 0 1 2720
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 35420 0 -1 2720
box -38 -48 866 592
use scs8hd_decap_8  FILLER_0_393 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 37260 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_386
timestamp 1586364061
transform 1 0 36616 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 36800 0 -1 2720
box -38 -48 222 592
use scs8hd_conb_1  _48_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 36984 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_392 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 37168 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_380
timestamp 1586364061
transform 1 0 36064 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_401
timestamp 1586364061
transform 1 0 37996 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_404
timestamp 1586364061
transform 1 0 38272 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_1_404
timestamp 1586364061
transform 1 0 38272 0 1 2720
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
timestamp 1586364061
transform 1 0 1472 0 -1 3808
box -38 -48 1786 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use scs8hd_fill_2  FILLER_2_41
timestamp 1586364061
transform 1 0 4876 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
timestamp 1586364061
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_49
timestamp 1586364061
transform 1 0 5612 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_45
timestamp 1586364061
transform 1 0 5244 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 5428 0 -1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
timestamp 1586364061
transform 1 0 5980 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
timestamp 1586364061
transform 1 0 5796 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
timestamp 1586364061
transform 1 0 7912 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_72
timestamp 1586364061
transform 1 0 7728 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_76
timestamp 1586364061
transform 1 0 8096 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1586364061
transform 1 0 8280 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _69_
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_conb_1  _41_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_96
timestamp 1586364061
transform 1 0 9936 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10120 0 -1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_100
timestamp 1586364061
transform 1 0 10304 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_123
timestamp 1586364061
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13156 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 14168 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 14536 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_127
timestamp 1586364061
transform 1 0 12788 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_140
timestamp 1586364061
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_144
timestamp 1586364061
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_148
timestamp 1586364061
transform 1 0 14720 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_158
timestamp 1586364061
transform 1 0 15640 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_152
timestamp 1586364061
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14904 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 15456 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15824 0 -1 3808
box -38 -48 866 592
use scs8hd_fill_2  FILLER_2_173
timestamp 1586364061
transform 1 0 17020 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_169
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 222 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 17388 0 -1 3808
box -38 -48 2246 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17204 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 19780 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 20148 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_201
timestamp 1586364061
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_205
timestamp 1586364061
transform 1 0 19964 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_209
timestamp 1586364061
transform 1 0 20332 0 -1 3808
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
timestamp 1586364061
transform 1 0 23276 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21896 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 22264 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 22632 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_224
timestamp 1586364061
transform 1 0 21712 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_228
timestamp 1586364061
transform 1 0 22080 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_232
timestamp 1586364061
transform 1 0 22448 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_236
timestamp 1586364061
transform 1 0 22816 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
timestamp 1586364061
transform 1 0 25208 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
timestamp 1586364061
transform 1 0 25576 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 26128 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_260
timestamp 1586364061
transform 1 0 25024 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_264
timestamp 1586364061
transform 1 0 25392 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_268
timestamp 1586364061
transform 1 0 25760 0 -1 3808
box -38 -48 406 592
use scs8hd_or2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 498 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 27968 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 27784 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
timestamp 1586364061
transform 1 0 27140 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_274
timestamp 1586364061
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_281
timestamp 1586364061
transform 1 0 26956 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_285
timestamp 1586364061
transform 1 0 27324 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_289
timestamp 1586364061
transform 1 0 27692 0 -1 3808
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 29532 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 29256 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_301
timestamp 1586364061
transform 1 0 28796 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_305
timestamp 1586364061
transform 1 0 29164 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_308
timestamp 1586364061
transform 1 0 29440 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_332
timestamp 1586364061
transform 1 0 31648 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_328
timestamp 1586364061
transform 1 0 31280 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 31464 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 31832 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 32108 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_341
timestamp 1586364061
transform 1 0 32476 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_345
timestamp 1586364061
transform 1 0 32844 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 33028 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 32660 0 -1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 33212 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 35144 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_368
timestamp 1586364061
transform 1 0 34960 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_372
timestamp 1586364061
transform 1 0 35328 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 35512 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_376
timestamp 1586364061
transform 1 0 35696 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_388
timestamp 1586364061
transform 1 0 36800 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_396
timestamp 1586364061
transform 1 0 37536 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_398
timestamp 1586364061
transform 1 0 37720 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_406
timestamp 1586364061
transform 1 0 38456 0 -1 3808
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1786 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
timestamp 1586364061
transform 1 0 3312 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_22
timestamp 1586364061
transform 1 0 3128 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _64_
timestamp 1586364061
transform 1 0 3864 0 1 3808
box -38 -48 406 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1586364061
transform 1 0 5060 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__64__A
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1586364061
transform 1 0 3680 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_26
timestamp 1586364061
transform 1 0 3496 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_34
timestamp 1586364061
transform 1 0 4232 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_38
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_42
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__67__A
timestamp 1586364061
transform 1 0 6072 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__68__A
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_52
timestamp 1586364061
transform 1 0 5888 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_56
timestamp 1586364061
transform 1 0 6256 0 1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_3_71
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_77
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_104
timestamp 1586364061
transform 1 0 10672 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_100
timestamp 1586364061
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10488 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10856 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 11040 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_112
timestamp 1586364061
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_116
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_120
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 12972 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_127
timestamp 1586364061
transform 1 0 12788 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_131
timestamp 1586364061
transform 1 0 13156 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_157
timestamp 1586364061
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_161
timestamp 1586364061
transform 1 0 15916 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_175
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18216 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 18400 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_192
timestamp 1586364061
transform 1 0 18768 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 18952 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 19320 0 1 3808
box -38 -48 222 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 19504 0 1 3808
box -38 -48 2246 592
use scs8hd_fill_2  FILLER_3_228
timestamp 1586364061
transform 1 0 22080 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_224
timestamp 1586364061
transform 1 0 21712 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1586364061
transform 1 0 22264 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1586364061
transform 1 0 21896 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_240
timestamp 1586364061
transform 1 0 23184 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_236
timestamp 1586364061
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1786 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1586364061
transform 1 0 26128 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 25944 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 25576 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_264
timestamp 1586364061
transform 1 0 25392 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_268
timestamp 1586364061
transform 1 0 25760 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 27692 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 27416 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 28244 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_281
timestamp 1586364061
transform 1 0 26956 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_285
timestamp 1586364061
transform 1 0 27324 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_288
timestamp 1586364061
transform 1 0 27600 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_293
timestamp 1586364061
transform 1 0 28060 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_297
timestamp 1586364061
transform 1 0 28428 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 29440 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 28980 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 30452 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 28612 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_301
timestamp 1586364061
transform 1 0 28796 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_306
timestamp 1586364061
transform 1 0 29256 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_317
timestamp 1586364061
transform 1 0 30268 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_321
timestamp 1586364061
transform 1 0 30636 0 1 3808
box -38 -48 222 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 31004 0 1 3808
box -38 -48 2246 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 30820 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 33948 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 33396 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 34316 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_349
timestamp 1586364061
transform 1 0 33212 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_353
timestamp 1586364061
transform 1 0 33580 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_359
timestamp 1586364061
transform 1 0 34132 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_363
timestamp 1586364061
transform 1 0 34500 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_367
timestamp 1586364061
transform 1 0 34868 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_379
timestamp 1586364061
transform 1 0 35972 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_391
timestamp 1586364061
transform 1 0 37076 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_3_403
timestamp 1586364061
transform 1 0 38180 0 1 3808
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1786 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
timestamp 1586364061
transform 1 0 3312 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_22
timestamp 1586364061
transform 1 0 3128 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1586364061
transform 1 0 4232 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 5244 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 5612 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_26
timestamp 1586364061
transform 1 0 3496 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_43
timestamp 1586364061
transform 1 0 5060 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_47
timestamp 1586364061
transform 1 0 5428 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_2  _67_
timestamp 1586364061
transform 1 0 5796 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_59
timestamp 1586364061
transform 1 0 6532 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_55
timestamp 1586364061
transform 1 0 6164 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 6348 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 6716 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_2  _68_
timestamp 1586364061
transform 1 0 6900 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_67
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 7452 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_71
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 866 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11960 0 -1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 11776 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11408 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_110
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_114
timestamp 1586364061
transform 1 0 11592 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13892 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14260 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_137
timestamp 1586364061
transform 1 0 13708 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16744 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_163
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_168
timestamp 1586364061
transform 1 0 16560 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_172
timestamp 1586364061
transform 1 0 16928 0 -1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 17296 0 -1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 17112 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_195
timestamp 1586364061
transform 1 0 19044 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_199
timestamp 1586364061
transform 1 0 19412 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 19504 0 -1 4896
box -38 -48 222 592
use scs8hd_conb_1  _46_
timestamp 1586364061
transform 1 0 19780 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_210
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_4  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_221
timestamp 1586364061
transform 1 0 21436 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1586364061
transform 1 0 21252 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1586364061
transform 1 0 21620 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1586364061
transform 1 0 21804 0 -1 4896
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
timestamp 1586364061
transform 1 0 23368 0 -1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
timestamp 1586364061
transform 1 0 23184 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
timestamp 1586364061
transform 1 0 22816 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_234
timestamp 1586364061
transform 1 0 22632 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_238
timestamp 1586364061
transform 1 0 23000 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 25668 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 26128 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_261
timestamp 1586364061
transform 1 0 25116 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_265
timestamp 1586364061
transform 1 0 25484 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_269
timestamp 1586364061
transform 1 0 25852 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_280
timestamp 1586364061
transform 1 0 26864 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_274
timestamp 1586364061
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 27048 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 26680 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_284
timestamp 1586364061
transform 1 0 27232 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 27416 0 -1 4896
box -38 -48 866 592
use scs8hd_fill_2  FILLER_4_295
timestamp 1586364061
transform 1 0 28244 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 28428 0 -1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 29256 0 -1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 28796 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_299
timestamp 1586364061
transform 1 0 28612 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_303
timestamp 1586364061
transform 1 0 28980 0 -1 4896
box -38 -48 314 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 32108 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 31648 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 31188 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_325
timestamp 1586364061
transform 1 0 31004 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_329
timestamp 1586364061
transform 1 0 31372 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_334
timestamp 1586364061
transform 1 0 31832 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_346
timestamp 1586364061
transform 1 0 32936 0 -1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 33948 0 -1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 33120 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 33488 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_350
timestamp 1586364061
transform 1 0 33304 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_354
timestamp 1586364061
transform 1 0 33672 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_376
timestamp 1586364061
transform 1 0 35696 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_4_388
timestamp 1586364061
transform 1 0 36800 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_396
timestamp 1586364061
transform 1 0 37536 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_398
timestamp 1586364061
transform 1 0 37720 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_406
timestamp 1586364061
transform 1 0 38456 0 -1 4896
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1586364061
transform 1 0 2116 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
timestamp 1586364061
transform 1 0 1564 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
timestamp 1586364061
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
timestamp 1586364061
transform 1 0 3128 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_20
timestamp 1586364061
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_24
timestamp 1586364061
transform 1 0 3312 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 3496 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _65_
timestamp 1586364061
transform 1 0 3680 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_32
timestamp 1586364061
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__65__A
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_36
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_44
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _66_
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_48
timestamp 1586364061
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__66__A
timestamp 1586364061
transform 1 0 5336 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 5704 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_52
timestamp 1586364061
transform 1 0 5888 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_71
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_78
timestamp 1586364061
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_75
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 8096 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _71_
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_83
timestamp 1586364061
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_87
timestamp 1586364061
transform 1 0 9108 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 9292 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__71__A
timestamp 1586364061
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 9476 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_95
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_99
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_107
timestamp 1586364061
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_111
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_115
timestamp 1586364061
transform 1 0 11684 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 13156 0 1 4896
box -38 -48 2246 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 12972 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12604 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_127
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 15548 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 15916 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_155
timestamp 1586364061
transform 1 0 15364 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_163
timestamp 1586364061
transform 1 0 16100 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_175
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 18216 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_194
timestamp 1586364061
transform 1 0 18952 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_190
timestamp 1586364061
transform 1 0 18584 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 18768 0 1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 19320 0 1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 21252 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 21620 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_217
timestamp 1586364061
transform 1 0 21068 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_221
timestamp 1586364061
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1586364061
transform 1 0 21988 0 1 4896
box -38 -48 866 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_225
timestamp 1586364061
transform 1 0 21804 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_236
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_240
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1586364061
transform 1 0 25208 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 25024 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_254
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_258
timestamp 1586364061
transform 1 0 24840 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_271
timestamp 1586364061
transform 1 0 26036 0 1 4896
box -38 -48 406 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1586364061
transform 1 0 27324 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
timestamp 1586364061
transform 1 0 28336 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1586364061
transform 1 0 27140 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1586364061
transform 1 0 26772 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 26404 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_277
timestamp 1586364061
transform 1 0 26588 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_281
timestamp 1586364061
transform 1 0 26956 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_294
timestamp 1586364061
transform 1 0 28152 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_298
timestamp 1586364061
transform 1 0 28520 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_302
timestamp 1586364061
transform 1 0 28888 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
timestamp 1586364061
transform 1 0 28704 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
timestamp 1586364061
transform 1 0 29256 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_310
timestamp 1586364061
transform 1 0 29624 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
timestamp 1586364061
transform 1 0 29808 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_314
timestamp 1586364061
transform 1 0 29992 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 30176 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_322
timestamp 1586364061
transform 1 0 30728 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 30360 0 1 4896
box -38 -48 406 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 31648 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__72__A
timestamp 1586364061
transform 1 0 30912 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 31464 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 32660 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_326
timestamp 1586364061
transform 1 0 31096 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_341
timestamp 1586364061
transform 1 0 32476 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_345
timestamp 1586364061
transform 1 0 32844 0 1 4896
box -38 -48 406 592
use scs8hd_conb_1  _49_
timestamp 1586364061
transform 1 0 33212 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_352
timestamp 1586364061
transform 1 0 33488 0 1 4896
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_5_364
timestamp 1586364061
transform 1 0 34592 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_367
timestamp 1586364061
transform 1 0 34868 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_379
timestamp 1586364061
transform 1 0 35972 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_391
timestamp 1586364061
transform 1 0 37076 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_5_403
timestamp 1586364061
transform 1 0 38180 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_9
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_22
timestamp 1586364061
transform 1 0 3128 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 3312 0 -1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
timestamp 1586364061
transform 1 0 2300 0 1 5984
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_7_32
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_30
timestamp 1586364061
transform 1 0 3864 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_26
timestamp 1586364061
transform 1 0 3496 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1586364061
transform 1 0 3680 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_1  FILLER_7_44
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_40
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_36
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 5060 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_49
timestamp 1586364061
transform 1 0 5612 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_49
timestamp 1586364061
transform 1 0 5612 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_45
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 5428 0 -1 5984
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
timestamp 1586364061
transform 1 0 5244 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_55
timestamp 1586364061
transform 1 0 6164 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 5980 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6348 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1586364061
transform 1 0 6532 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_72
timestamp 1586364061
transform 1 0 7728 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 7912 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 7544 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_83
timestamp 1586364061
transform 1 0 8740 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_75
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 8096 0 -1 5984
box -38 -48 406 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
timestamp 1586364061
transform 1 0 8372 0 1 5984
box -38 -48 406 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9568 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_87
timestamp 1586364061
transform 1 0 9108 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_90
timestamp 1586364061
transform 1 0 9384 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10212 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_97
timestamp 1586364061
transform 1 0 10028 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_94
timestamp 1586364061
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 866 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_107
timestamp 1586364061
transform 1 0 10948 0 1 5984
box -38 -48 406 592
use scs8hd_decap_6  FILLER_6_108 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11040 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_6_101
timestamp 1586364061
transform 1 0 10396 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 10580 0 -1 5984
box -38 -48 222 592
use scs8hd_conb_1  _40_
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_111
timestamp 1586364061
transform 1 0 11316 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11592 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 11776 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_136
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_132
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_125
timestamp 1586364061
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 13156 0 -1 5984
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13340 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_6_146
timestamp 1586364061
transform 1 0 14536 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_142
timestamp 1586364061
transform 1 0 14168 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14720 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 1786 592
use scs8hd_decap_3  FILLER_6_150
timestamp 1586364061
transform 1 0 14904 0 -1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_3  FILLER_7_167
timestamp 1586364061
transform 1 0 16468 0 1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_168
timestamp 1586364061
transform 1 0 16560 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_172
timestamp 1586364061
transform 1 0 16928 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16744 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use scs8hd_conb_1  _44_
timestamp 1586364061
transform 1 0 16928 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_177
timestamp 1586364061
transform 1 0 17388 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17204 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17572 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 17756 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_1  FILLER_6_198
timestamp 1586364061
transform 1 0 19320 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_194
timestamp 1586364061
transform 1 0 18952 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18768 0 -1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_7_207
timestamp 1586364061
transform 1 0 20148 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_203
timestamp 1586364061
transform 1 0 19780 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_206
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 19872 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 19964 0 1 5984
box -38 -48 222 592
use scs8hd_conb_1  _45_
timestamp 1586364061
transform 1 0 19412 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_223
timestamp 1586364061
transform 1 0 21620 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_219
timestamp 1586364061
transform 1 0 21252 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_215
timestamp 1586364061
transform 1 0 20884 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 21068 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 21436 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 21804 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1586364061
transform 1 0 21988 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_236
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_238
timestamp 1586364061
transform 1 0 23000 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_234
timestamp 1586364061
transform 1 0 22632 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 23184 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1586364061
transform 1 0 22816 0 -1 5984
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1586364061
transform 1 0 23368 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_258
timestamp 1586364061
transform 1 0 24840 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_254
timestamp 1586364061
transform 1 0 24472 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_255
timestamp 1586364061
transform 1 0 24564 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 24748 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 24380 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 24656 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_266
timestamp 1586364061
transform 1 0 25576 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_262
timestamp 1586364061
transform 1 0 25208 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_267
timestamp 1586364061
transform 1 0 25668 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_259
timestamp 1586364061
transform 1 0 24932 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 25116 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 25760 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 25392 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 25024 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_6_272
timestamp 1586364061
transform 1 0 26128 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 25944 0 -1 5984
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1586364061
transform 1 0 25944 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_283
timestamp 1586364061
transform 1 0 27140 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_279
timestamp 1586364061
transform 1 0 26772 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_285
timestamp 1586364061
transform 1 0 27324 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
timestamp 1586364061
transform 1 0 26956 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 27324 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_296
timestamp 1586364061
transform 1 0 28336 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_289
timestamp 1586364061
transform 1 0 27692 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1586364061
transform 1 0 27876 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 27508 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
timestamp 1586364061
transform 1 0 28520 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1586364061
transform 1 0 27508 0 1 5984
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
timestamp 1586364061
transform 1 0 28060 0 -1 5984
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_7_310
timestamp 1586364061
transform 1 0 29624 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_304
timestamp 1586364061
transform 1 0 29072 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_300
timestamp 1586364061
transform 1 0 28704 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
timestamp 1586364061
transform 1 0 28888 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
timestamp 1586364061
transform 1 0 29256 0 1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
timestamp 1586364061
transform 1 0 29808 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 29992 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_312
timestamp 1586364061
transform 1 0 29808 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_314
timestamp 1586364061
transform 1 0 29992 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  _72_
timestamp 1586364061
transform 1 0 30544 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 30360 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 30176 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 30544 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_316
timestamp 1586364061
transform 1 0 30176 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_318
timestamp 1586364061
transform 1 0 30360 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_322
timestamp 1586364061
transform 1 0 30728 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_334
timestamp 1586364061
transform 1 0 31832 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_334
timestamp 1586364061
transform 1 0 31832 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_328
timestamp 1586364061
transform 1 0 31280 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_324
timestamp 1586364061
transform 1 0 30912 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 31648 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 31096 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_347
timestamp 1586364061
transform 1 0 33028 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_342
timestamp 1586364061
transform 1 0 32568 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 32844 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use scs8hd_conb_1  _50_
timestamp 1586364061
transform 1 0 32108 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_340
timestamp 1586364061
transform 1 0 32384 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_355
timestamp 1586364061
transform 1 0 33764 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_351
timestamp 1586364061
transform 1 0 33396 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 33580 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 33212 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_367
timestamp 1586364061
transform 1 0 34868 0 1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_7_363
timestamp 1586364061
transform 1 0 34500 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_370
timestamp 1586364061
transform 1 0 35144 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_6_364
timestamp 1586364061
transform 1 0 34592 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 35236 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 35236 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_352
timestamp 1586364061
transform 1 0 33488 0 -1 5984
box -38 -48 1142 592
use scs8hd_conb_1  _54_
timestamp 1586364061
transform 1 0 35420 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 35880 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_373
timestamp 1586364061
transform 1 0 35420 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_385
timestamp 1586364061
transform 1 0 36524 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_376
timestamp 1586364061
transform 1 0 35696 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_380
timestamp 1586364061
transform 1 0 36064 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_392
timestamp 1586364061
transform 1 0 37168 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_6_398
timestamp 1586364061
transform 1 0 37720 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_406
timestamp 1586364061
transform 1 0 38456 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_404
timestamp 1586364061
transform 1 0 38272 0 1 5984
box -38 -48 314 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_7
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_10
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 6532 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
timestamp 1586364061
transform 1 0 5980 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 6348 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_51
timestamp 1586364061
transform 1 0 5796 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_55
timestamp 1586364061
transform 1 0 6164 0 -1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10028 0 -1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_78
timestamp 1586364061
transform 1 0 8280 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_82
timestamp 1586364061
transform 1 0 8648 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_90
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 406 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12512 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 12328 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11960 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_116
timestamp 1586364061
transform 1 0 11776 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_120
timestamp 1586364061
transform 1 0 12144 0 -1 7072
box -38 -48 222 592
use scs8hd_conb_1  _42_
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 13524 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13892 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_133
timestamp 1586364061
transform 1 0 13340 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_137
timestamp 1586364061
transform 1 0 13708 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_144
timestamp 1586364061
transform 1 0 14352 0 -1 7072
box -38 -48 774 592
use scs8hd_conb_1  _37_
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use scs8hd_conb_1  _43_
timestamp 1586364061
transform 1 0 16652 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_152
timestamp 1586364061
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_157
timestamp 1586364061
transform 1 0 15548 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_8_172
timestamp 1586364061
transform 1 0 16928 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 19228 0 -1 7072
box -38 -48 406 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 17664 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18676 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17112 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_176
timestamp 1586364061
transform 1 0 17296 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_189
timestamp 1586364061
transform 1 0 18492 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_193
timestamp 1586364061
transform 1 0 18860 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_201
timestamp 1586364061
transform 1 0 19596 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_8_213
timestamp 1586364061
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_223
timestamp 1586364061
transform 1 0 21620 0 -1 7072
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 22080 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 21896 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_247
timestamp 1586364061
transform 1 0 23828 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1586364061
transform 1 0 24840 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 24012 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 26220 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 24380 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 25852 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_255
timestamp 1586364061
transform 1 0 24564 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_267
timestamp 1586364061
transform 1 0 25668 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_271
timestamp 1586364061
transform 1 0 26036 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
timestamp 1586364061
transform 1 0 28244 0 -1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
timestamp 1586364061
transform 1 0 27048 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 27508 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_280
timestamp 1586364061
transform 1 0 26864 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_284
timestamp 1586364061
transform 1 0 27232 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_6  FILLER_8_289
timestamp 1586364061
transform 1 0 27692 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_8_314
timestamp 1586364061
transform 1 0 29992 0 -1 7072
box -38 -48 1142 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 32844 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 32660 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_326
timestamp 1586364061
transform 1 0 31096 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_334
timestamp 1586364061
transform 1 0 31832 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_337
timestamp 1586364061
transform 1 0 32108 0 -1 7072
box -38 -48 590 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 35236 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 35052 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 34684 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_354
timestamp 1586364061
transform 1 0 33672 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_362
timestamp 1586364061
transform 1 0 34408 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_367
timestamp 1586364061
transform 1 0 34868 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 36248 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 36616 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_380
timestamp 1586364061
transform 1 0 36064 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_384
timestamp 1586364061
transform 1 0 36432 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_388
timestamp 1586364061
transform 1 0 36800 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_396
timestamp 1586364061
transform 1 0 37536 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_398
timestamp 1586364061
transform 1 0 37720 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_406
timestamp 1586364061
transform 1 0 38456 0 -1 7072
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
timestamp 1586364061
transform 1 0 2944 0 1 7072
box -38 -48 1786 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
timestamp 1586364061
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 2392 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_9_11
timestamp 1586364061
transform 1 0 2116 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_16
timestamp 1586364061
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
timestamp 1586364061
transform 1 0 5612 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
timestamp 1586364061
transform 1 0 5336 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_44
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_48
timestamp 1586364061
transform 1 0 5520 0 1 7072
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_81
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_85
timestamp 1586364061
transform 1 0 8924 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_90
timestamp 1586364061
transform 1 0 9384 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_113
timestamp 1586364061
transform 1 0 11500 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_117
timestamp 1586364061
transform 1 0 11868 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 12880 0 1 7072
box -38 -48 2246 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 12696 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 16652 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_152
timestamp 1586364061
transform 1 0 15088 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_156
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_160
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_9_168
timestamp 1586364061
transform 1 0 16560 0 1 7072
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_203
timestamp 1586364061
transform 1 0 19780 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
timestamp 1586364061
transform 1 0 19964 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_207
timestamp 1586364061
transform 1 0 20148 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
timestamp 1586364061
transform 1 0 20332 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 20516 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_219
timestamp 1586364061
transform 1 0 21252 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_215
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_223
timestamp 1586364061
transform 1 0 21620 0 1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 21436 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 22264 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_229
timestamp 1586364061
transform 1 0 22172 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_236
timestamp 1586364061
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_240
timestamp 1586364061
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 26128 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 25760 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_264
timestamp 1586364061
transform 1 0 25392 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_270
timestamp 1586364061
transform 1 0 25944 0 1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
timestamp 1586364061
transform 1 0 26680 0 1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
timestamp 1586364061
transform 1 0 26496 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_274
timestamp 1586364061
transform 1 0 26312 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_297
timestamp 1586364061
transform 1 0 28428 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _47_
timestamp 1586364061
transform 1 0 29256 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
timestamp 1586364061
transform 1 0 28612 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
timestamp 1586364061
transform 1 0 28980 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_301
timestamp 1586364061
transform 1 0 28796 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_309
timestamp 1586364061
transform 1 0 29532 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_321
timestamp 1586364061
transform 1 0 30636 0 1 7072
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 32108 0 1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 31924 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 31556 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_329
timestamp 1586364061
transform 1 0 31372 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_333
timestamp 1586364061
transform 1 0 31740 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 35236 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 34040 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 34592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_356
timestamp 1586364061
transform 1 0 33856 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_360
timestamp 1586364061
transform 1 0 34224 0 1 7072
box -38 -48 406 592
use scs8hd_decap_4  FILLER_9_367
timestamp 1586364061
transform 1 0 34868 0 1 7072
box -38 -48 406 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 35420 0 1 7072
box -38 -48 2246 592
use scs8hd_decap_8  FILLER_9_397
timestamp 1586364061
transform 1 0 37628 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_405
timestamp 1586364061
transform 1 0 38364 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
timestamp 1586364061
transform 1 0 2944 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_19
timestamp 1586364061
transform 1 0 2852 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_22
timestamp 1586364061
transform 1 0 3128 0 -1 8160
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
timestamp 1586364061
transform 1 0 4968 0 -1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_30
timestamp 1586364061
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_36
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 590 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6900 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_61
timestamp 1586364061
transform 1 0 6716 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_65
timestamp 1586364061
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9844 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_78
timestamp 1586364061
transform 1 0 8280 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_82
timestamp 1586364061
transform 1 0 8648 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_90
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_97
timestamp 1586364061
transform 1 0 10028 0 -1 8160
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 10304 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_121
timestamp 1586364061
transform 1 0 12236 0 -1 8160
box -38 -48 406 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 12696 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13984 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 14352 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_125
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_128
timestamp 1586364061
transform 1 0 12880 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_138
timestamp 1586364061
transform 1 0 13800 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_142
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_146
timestamp 1586364061
transform 1 0 14536 0 -1 8160
box -38 -48 590 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_152
timestamp 1586364061
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_173
timestamp 1586364061
transform 1 0 17020 0 -1 8160
box -38 -48 314 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 17848 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 19044 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17664 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 17296 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_178
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_191
timestamp 1586364061
transform 1 0 18676 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_3  FILLER_10_197
timestamp 1586364061
transform 1 0 19228 0 -1 8160
box -38 -48 314 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use scs8hd_or2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
timestamp 1586364061
transform 1 0 19504 0 -1 8160
box -38 -48 498 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_205
timestamp 1586364061
transform 1 0 19964 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_213
timestamp 1586364061
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_219
timestamp 1586364061
transform 1 0 21252 0 -1 8160
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 23368 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 23184 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_231
timestamp 1586364061
transform 1 0 22356 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 25300 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
timestamp 1586364061
transform 1 0 26220 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 25668 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_261
timestamp 1586364061
transform 1 0 25116 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_265
timestamp 1586364061
transform 1 0 25484 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_269
timestamp 1586364061
transform 1 0 25852 0 -1 8160
box -38 -48 406 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1586364061
transform 1 0 26588 0 -1 8160
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
timestamp 1586364061
transform 1 0 28244 0 -1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_286
timestamp 1586364061
transform 1 0 27416 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_294
timestamp 1586364061
transform 1 0 28152 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 30452 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_314
timestamp 1586364061
transform 1 0 29992 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_318
timestamp 1586364061
transform 1 0 30360 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_321
timestamp 1586364061
transform 1 0 30636 0 -1 8160
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 32936 0 -1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 32568 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 31096 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_325
timestamp 1586364061
transform 1 0 31004 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_328
timestamp 1586364061
transform 1 0 31280 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_4  FILLER_10_337
timestamp 1586364061
transform 1 0 32108 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_341
timestamp 1586364061
transform 1 0 32476 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_344
timestamp 1586364061
transform 1 0 32752 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 35236 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 34868 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_365
timestamp 1586364061
transform 1 0 34684 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_369
timestamp 1586364061
transform 1 0 35052 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 35420 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 36432 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_382
timestamp 1586364061
transform 1 0 36248 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_386
timestamp 1586364061
transform 1 0 36616 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_10_394
timestamp 1586364061
transform 1 0 37352 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_398
timestamp 1586364061
transform 1 0 37720 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_406
timestamp 1586364061
transform 1 0 38456 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_11_23
timestamp 1586364061
transform 1 0 3220 0 1 8160
box -38 -48 314 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1586364061
transform 1 0 4048 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 3496 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_28
timestamp 1586364061
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_41
timestamp 1586364061
transform 1 0 4876 0 1 8160
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_81
timestamp 1586364061
transform 1 0 8556 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 12696 0 1 8160
box -38 -48 2246 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 16744 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16284 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_150
timestamp 1586364061
transform 1 0 14904 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_156
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_163
timestamp 1586364061
transform 1 0 16100 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_167
timestamp 1586364061
transform 1 0 16468 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_178
timestamp 1586364061
transform 1 0 17480 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_174
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 18216 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 17296 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_192
timestamp 1586364061
transform 1 0 18768 0 1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_188
timestamp 1586364061
transform 1 0 18400 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
timestamp 1586364061
transform 1 0 20976 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_214
timestamp 1586364061
transform 1 0 20792 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_218
timestamp 1586364061
transform 1 0 21160 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_222
timestamp 1586364061
transform 1 0 21528 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_11_234
timestamp 1586364061
transform 1 0 22632 0 1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_11_242
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
timestamp 1586364061
transform 1 0 24196 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
timestamp 1586364061
transform 1 0 26128 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
timestamp 1586364061
transform 1 0 24012 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_270
timestamp 1586364061
transform 1 0 25944 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
timestamp 1586364061
transform 1 0 26680 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
timestamp 1586364061
transform 1 0 26496 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_274
timestamp 1586364061
transform 1 0 26312 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_297
timestamp 1586364061
transform 1 0 28428 0 1 8160
box -38 -48 774 592
use scs8hd_conb_1  _51_
timestamp 1586364061
transform 1 0 30084 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 30544 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 29900 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_306
timestamp 1586364061
transform 1 0 29256 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_312
timestamp 1586364061
transform 1 0 29808 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_318
timestamp 1586364061
transform 1 0 30360 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_322
timestamp 1586364061
transform 1 0 30728 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 31096 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 33028 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 30912 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_345
timestamp 1586364061
transform 1 0 32844 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_356
timestamp 1586364061
transform 1 0 33856 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_349
timestamp 1586364061
transform 1 0 33212 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 34224 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 33396 0 1 8160
box -38 -48 222 592
use scs8hd_conb_1  _52_
timestamp 1586364061
transform 1 0 33580 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_367
timestamp 1586364061
transform 1 0 34868 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_362
timestamp 1586364061
transform 1 0 34408 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 34592 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 35052 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 36984 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_388
timestamp 1586364061
transform 1 0 36800 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_392
timestamp 1586364061
transform 1 0 37168 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_404
timestamp 1586364061
transform 1 0 38272 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6900 0 -1 9248
box -38 -48 1786 592
use scs8hd_decap_6  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_62
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 130 592
use scs8hd_conb_1  _39_
timestamp 1586364061
transform 1 0 9936 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_82
timestamp 1586364061
transform 1 0 8648 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_90
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_12_99
timestamp 1586364061
transform 1 0 10212 0 -1 9248
box -38 -48 590 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11684 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11500 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11132 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_107
timestamp 1586364061
transform 1 0 10948 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_111
timestamp 1586364061
transform 1 0 11316 0 -1 9248
box -38 -48 222 592
use scs8hd_conb_1  _38_
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_134
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_138
timestamp 1586364061
transform 1 0 13800 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15916 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 15456 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16928 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_158
timestamp 1586364061
transform 1 0 15640 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_170
timestamp 1586364061
transform 1 0 16744 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
timestamp 1586364061
transform 1 0 19228 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 17572 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_174
timestamp 1586364061
transform 1 0 17112 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_181
timestamp 1586364061
transform 1 0 17756 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_195
timestamp 1586364061
transform 1 0 19044 0 -1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
timestamp 1586364061
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1586364061
transform 1 0 19872 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_199
timestamp 1586364061
transform 1 0 19412 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_203
timestamp 1586364061
transform 1 0 19780 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_206
timestamp 1586364061
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_210
timestamp 1586364061
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_234
timestamp 1586364061
transform 1 0 22632 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_12_246
timestamp 1586364061
transform 1 0 23736 0 -1 9248
box -38 -48 406 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1586364061
transform 1 0 24840 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
timestamp 1586364061
transform 1 0 26220 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 24656 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_250
timestamp 1586364061
transform 1 0 24104 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_253
timestamp 1586364061
transform 1 0 24380 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_12_267
timestamp 1586364061
transform 1 0 25668 0 -1 9248
box -38 -48 590 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_295
timestamp 1586364061
transform 1 0 28244 0 -1 9248
box -38 -48 1142 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 30452 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 29992 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 29624 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_307
timestamp 1586364061
transform 1 0 29348 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_312
timestamp 1586364061
transform 1 0 29808 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_316
timestamp 1586364061
transform 1 0 30176 0 -1 9248
box -38 -48 314 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 32568 0 -1 9248
box -38 -48 2246 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 32384 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_328
timestamp 1586364061
transform 1 0 31280 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_12_337
timestamp 1586364061
transform 1 0 32108 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 35144 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_366
timestamp 1586364061
transform 1 0 34776 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_372
timestamp 1586364061
transform 1 0 35328 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 35512 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_383
timestamp 1586364061
transform 1 0 36340 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_12_395
timestamp 1586364061
transform 1 0 37444 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_398
timestamp 1586364061
transform 1 0 37720 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_406
timestamp 1586364061
transform 1 0 38456 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1586364061
transform 1 0 6440 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_64
timestamp 1586364061
transform 1 0 6992 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_60
timestamp 1586364061
transform 1 0 6624 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_69
timestamp 1586364061
transform 1 0 7452 0 1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_13_66
timestamp 1586364061
transform 1 0 7176 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 7268 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1586364061
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 866 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 7728 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_81
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_76
timestamp 1586364061
transform 1 0 8096 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_80
timestamp 1586364061
transform 1 0 8464 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_76
timestamp 1586364061
transform 1 0 8096 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1586364061
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1586364061
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 8280 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_91
timestamp 1586364061
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_85
timestamp 1586364061
transform 1 0 8924 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_92
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_84
timestamp 1586364061
transform 1 0 8832 0 1 9248
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_97
timestamp 1586364061
transform 1 0 10028 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_97
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 406 592
use scs8hd_conb_1  _36_
timestamp 1586364061
transform 1 0 9752 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_106
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_103
timestamp 1586364061
transform 1 0 10580 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_101
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_110
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 11408 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_121
timestamp 1586364061
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_133
timestamp 1586364061
transform 1 0 13340 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13156 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_140
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_136
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_148
timestamp 1586364061
transform 1 0 14720 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_144
timestamp 1586364061
transform 1 0 14352 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 14536 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_158
timestamp 1586364061
transform 1 0 15640 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_152
timestamp 1586364061
transform 1 0 15088 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14904 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 15824 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 15456 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_171
timestamp 1586364061
transform 1 0 16836 0 -1 10336
box -38 -48 774 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16008 0 -1 10336
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_13_181
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1586364061
transform 1 0 17572 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_1  FILLER_14_192
timestamp 1586364061
transform 1 0 18768 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_188
timestamp 1586364061
transform 1 0 18400 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_3  FILLER_13_188
timestamp 1586364061
transform 1 0 18400 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 18860 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 18676 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 18216 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 866 592
use scs8hd_fill_1  FILLER_14_195
timestamp 1586364061
transform 1 0 19044 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
timestamp 1586364061
transform 1 0 19136 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_14_208
timestamp 1586364061
transform 1 0 20240 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_204
timestamp 1586364061
transform 1 0 19872 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_200
timestamp 1586364061
transform 1 0 19504 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_202
timestamp 1586364061
transform 1 0 19688 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1586364061
transform 1 0 20056 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
timestamp 1586364061
transform 1 0 19872 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1586364061
transform 1 0 20056 0 1 9248
box -38 -48 866 592
use scs8hd_fill_1  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
timestamp 1586364061
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
timestamp 1586364061
transform 1 0 20884 0 1 9248
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
timestamp 1586364061
transform 1 0 20976 0 -1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_234
timestamp 1586364061
transform 1 0 22632 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_242
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_235
timestamp 1586364061
transform 1 0 22724 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_247
timestamp 1586364061
transform 1 0 23828 0 -1 10336
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
timestamp 1586364061
transform 1 0 25300 0 1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
timestamp 1586364061
transform 1 0 25116 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 406 592
use scs8hd_decap_4  FILLER_14_259
timestamp 1586364061
transform 1 0 24932 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_265
timestamp 1586364061
transform 1 0 25484 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_273
timestamp 1586364061
transform 1 0 26220 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_282
timestamp 1586364061
transform 1 0 27048 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_294
timestamp 1586364061
transform 1 0 28152 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_288
timestamp 1586364061
transform 1 0 27600 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 28888 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 28888 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_300
timestamp 1586364061
transform 1 0 28704 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_304
timestamp 1586364061
transform 1 0 29072 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_306
timestamp 1586364061
transform 1 0 29256 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_306
timestamp 1586364061
transform 1 0 29256 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 29440 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_310
timestamp 1586364061
transform 1 0 29624 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_310
timestamp 1586364061
transform 1 0 29624 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_313
timestamp 1586364061
transform 1 0 29900 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 29716 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 29808 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 30084 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 29992 0 -1 10336
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 30268 0 1 9248
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_14_327
timestamp 1586364061
transform 1 0 31188 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_323
timestamp 1586364061
transform 1 0 30820 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 31004 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_337
timestamp 1586364061
transform 1 0 32108 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_14_335
timestamp 1586364061
transform 1 0 31924 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_340
timestamp 1586364061
transform 1 0 32384 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_336
timestamp 1586364061
transform 1 0 32016 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 32200 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 32568 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_346
timestamp 1586364061
transform 1 0 32936 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_343
timestamp 1586364061
transform 1 0 32660 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 32752 0 -1 10336
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 32752 0 1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_358
timestamp 1586364061
transform 1 0 34040 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_357
timestamp 1586364061
transform 1 0 33948 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_353
timestamp 1586364061
transform 1 0 33580 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 34132 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 33764 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 33212 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_1  FILLER_14_369
timestamp 1586364061
transform 1 0 35052 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_366
timestamp 1586364061
transform 1 0 34776 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_361
timestamp 1586364061
transform 1 0 34316 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 34868 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 34592 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 35144 0 -1 10336
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 34868 0 1 9248
box -38 -48 1786 592
use scs8hd_conb_1  _53_
timestamp 1586364061
transform 1 0 37352 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 36800 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_386
timestamp 1586364061
transform 1 0 36616 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_390
timestamp 1586364061
transform 1 0 36984 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_13_397
timestamp 1586364061
transform 1 0 37628 0 1 9248
box -38 -48 774 592
use scs8hd_decap_8  FILLER_14_389
timestamp 1586364061
transform 1 0 36892 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_405
timestamp 1586364061
transform 1 0 38364 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_398
timestamp 1586364061
transform 1 0 37720 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_406
timestamp 1586364061
transform 1 0 38456 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_75
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_88
timestamp 1586364061
transform 1 0 9200 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_108
timestamp 1586364061
transform 1 0 11040 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use scs8hd_or2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 498 592
use scs8hd_decap_4  FILLER_15_116
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_112
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_137
timestamp 1586364061
transform 1 0 13708 0 1 10336
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_15_149
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 14904 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_152
timestamp 1586364061
transform 1 0 15088 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 866 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 18584 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
timestamp 1586364061
transform 1 0 18952 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_15_188
timestamp 1586364061
transform 1 0 18400 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_192
timestamp 1586364061
transform 1 0 18768 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 130 592
use scs8hd_clkbuf_16  clkbuf_1_0__f_clk tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20792 0 1 10336
box -38 -48 1878 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
timestamp 1586364061
transform 1 0 20608 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_206
timestamp 1586364061
transform 1 0 20056 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_210
timestamp 1586364061
transform 1 0 20424 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_15_234
timestamp 1586364061
transform 1 0 22632 0 1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_15_242
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 774 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
timestamp 1586364061
transform 1 0 25668 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1586364061
transform 1 0 24380 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
timestamp 1586364061
transform 1 0 26220 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1586364061
transform 1 0 25116 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_255
timestamp 1586364061
transform 1 0 24564 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_259
timestamp 1586364061
transform 1 0 24932 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_263
timestamp 1586364061
transform 1 0 25300 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_271
timestamp 1586364061
transform 1 0 26036 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_275
timestamp 1586364061
transform 1 0 26404 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
timestamp 1586364061
transform 1 0 26772 0 1 10336
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
timestamp 1586364061
transform 1 0 26956 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_285
timestamp 1586364061
transform 1 0 27324 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
timestamp 1586364061
transform 1 0 27508 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_289
timestamp 1586364061
transform 1 0 27692 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
timestamp 1586364061
transform 1 0 27876 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_297
timestamp 1586364061
transform 1 0 28428 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_293
timestamp 1586364061
transform 1 0 28060 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 28244 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 29808 0 1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 29624 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
timestamp 1586364061
transform 1 0 28980 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 28612 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_301
timestamp 1586364061
transform 1 0 28796 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_306
timestamp 1586364061
transform 1 0 29256 0 1 10336
box -38 -48 406 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 32292 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 32844 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 32108 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_331
timestamp 1586364061
transform 1 0 31556 0 1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_15_343
timestamp 1586364061
transform 1 0 32660 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_347
timestamp 1586364061
transform 1 0 33028 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 35236 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 33212 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_351
timestamp 1586364061
transform 1 0 33396 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_15_363
timestamp 1586364061
transform 1 0 34500 0 1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_15_367
timestamp 1586364061
transform 1 0 34868 0 1 10336
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 35420 0 1 10336
box -38 -48 1786 592
use scs8hd_decap_12  FILLER_15_392
timestamp 1586364061
transform 1 0 37168 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_404
timestamp 1586364061
transform 1 0 38272 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
timestamp 1586364061
transform 1 0 7084 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_64
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 9936 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
timestamp 1586364061
transform 1 0 9292 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_88
timestamp 1586364061
transform 1 0 9200 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_91
timestamp 1586364061
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 11040 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_100
timestamp 1586364061
transform 1 0 10304 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_104
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 406 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 13524 0 -1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_127
timestamp 1586364061
transform 1 0 12788 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_131
timestamp 1586364061
transform 1 0 13156 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_139
timestamp 1586364061
transform 1 0 13892 0 -1 11424
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 15456 0 -1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_151
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 19228 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
timestamp 1586364061
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 18400 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_175
timestamp 1586364061
transform 1 0 17204 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_183
timestamp 1586364061
transform 1 0 17940 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_186
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_190
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_195
timestamp 1586364061
transform 1 0 19044 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1586364061
transform 1 0 20332 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 19596 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 19964 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_199
timestamp 1586364061
transform 1 0 19412 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_203
timestamp 1586364061
transform 1 0 19780 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_207
timestamp 1586364061
transform 1 0 20148 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_211
timestamp 1586364061
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
timestamp 1586364061
transform 1 0 23920 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
timestamp 1586364061
transform 1 0 23552 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_234
timestamp 1586364061
transform 1 0 22632 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_242
timestamp 1586364061
transform 1 0 23368 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_246
timestamp 1586364061
transform 1 0 23736 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1586364061
transform 1 0 24380 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
timestamp 1586364061
transform 1 0 25668 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_250
timestamp 1586364061
transform 1 0 24104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_16_262
timestamp 1586364061
transform 1 0 25208 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_266
timestamp 1586364061
transform 1 0 25576 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_269
timestamp 1586364061
transform 1 0 25852 0 -1 11424
box -38 -48 590 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
timestamp 1586364061
transform 1 0 27140 0 -1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
timestamp 1586364061
transform 1 0 26680 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_280
timestamp 1586364061
transform 1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1586364061
transform 1 0 29624 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
timestamp 1586364061
transform 1 0 29256 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_302
timestamp 1586364061
transform 1 0 28888 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_308
timestamp 1586364061
transform 1 0 29440 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_319
timestamp 1586364061
transform 1 0 30452 0 -1 11424
box -38 -48 1142 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 32108 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_331
timestamp 1586364061
transform 1 0 31556 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_335
timestamp 1586364061
transform 1 0 31924 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_341
timestamp 1586364061
transform 1 0 32476 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_353
timestamp 1586364061
transform 1 0 33580 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_365
timestamp 1586364061
transform 1 0 34684 0 -1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 35420 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_375
timestamp 1586364061
transform 1 0 35604 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_387
timestamp 1586364061
transform 1 0 36708 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_395
timestamp 1586364061
transform 1 0 37444 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_398
timestamp 1586364061
transform 1 0 37720 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_406
timestamp 1586364061
transform 1 0 38456 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
timestamp 1586364061
transform 1 0 9292 0 1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
timestamp 1586364061
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 8740 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_81
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_85
timestamp 1586364061
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_108
timestamp 1586364061
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_112
timestamp 1586364061
transform 1 0 11408 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
timestamp 1586364061
transform 1 0 14720 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_142
timestamp 1586364061
transform 1 0 14168 0 1 11424
box -38 -48 590 592
use scs8hd_conb_1  _35_
timestamp 1586364061
transform 1 0 14904 0 1 11424
box -38 -48 314 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1586364061
transform 1 0 15916 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
timestamp 1586364061
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_153
timestamp 1586364061
transform 1 0 15180 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_157
timestamp 1586364061
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_170
timestamp 1586364061
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 18584 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 17296 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_174
timestamp 1586364061
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_178
timestamp 1586364061
transform 1 0 17480 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_188
timestamp 1586364061
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_192
timestamp 1586364061
transform 1 0 18768 0 1 11424
box -38 -48 774 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1586364061
transform 1 0 20332 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1586364061
transform 1 0 20148 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1586364061
transform 1 0 19780 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_clkbuf_1_0__f_clk_A
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_200
timestamp 1586364061
transform 1 0 19504 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_205
timestamp 1586364061
transform 1 0 19964 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_218
timestamp 1586364061
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_222
timestamp 1586364061
transform 1 0 21528 0 1 11424
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
timestamp 1586364061
transform 1 0 23920 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
timestamp 1586364061
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_234
timestamp 1586364061
transform 1 0 22632 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_240
timestamp 1586364061
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
timestamp 1586364061
transform 1 0 25668 0 1 11424
box -38 -48 1786 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 28060 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
timestamp 1586364061
transform 1 0 27600 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_286
timestamp 1586364061
transform 1 0 27416 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_290
timestamp 1586364061
transform 1 0 27784 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_297
timestamp 1586364061
transform 1 0 28428 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
timestamp 1586364061
transform 1 0 29256 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
timestamp 1586364061
transform 1 0 28980 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 28612 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_301
timestamp 1586364061
transform 1 0 28796 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_325
timestamp 1586364061
transform 1 0 31004 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_337
timestamp 1586364061
transform 1 0 32108 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 35236 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_349
timestamp 1586364061
transform 1 0 33212 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_17_361
timestamp 1586364061
transform 1 0 34316 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_365
timestamp 1586364061
transform 1 0 34684 0 1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_17_367
timestamp 1586364061
transform 1 0 34868 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 35604 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 35972 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_373
timestamp 1586364061
transform 1 0 35420 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_377
timestamp 1586364061
transform 1 0 35788 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_381
timestamp 1586364061
transform 1 0 36156 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_393
timestamp 1586364061
transform 1 0 37260 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_405
timestamp 1586364061
transform 1 0 38364 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
timestamp 1586364061
transform 1 0 6624 0 -1 12512
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 406 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_79
timestamp 1586364061
transform 1 0 8372 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_91
timestamp 1586364061
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11316 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11684 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_106
timestamp 1586364061
transform 1 0 10856 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_110
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_113
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 13892 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_136
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
timestamp 1586364061
transform 1 0 15364 0 -1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1586364061
transform 1 0 17848 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 18860 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_174
timestamp 1586364061
transform 1 0 17112 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_191
timestamp 1586364061
transform 1 0 18676 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_195
timestamp 1586364061
transform 1 0 19044 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_207
timestamp 1586364061
transform 1 0 20148 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_203
timestamp 1586364061
transform 1 0 19780 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_199
timestamp 1586364061
transform 1 0 19412 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1586364061
transform 1 0 19964 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 19596 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
timestamp 1586364061
transform 1 0 20516 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_213
timestamp 1586364061
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
timestamp 1586364061
transform 1 0 21068 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_219
timestamp 1586364061
transform 1 0 21252 0 -1 12512
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
timestamp 1586364061
transform 1 0 23736 0 -1 12512
box -38 -48 1786 592
use scs8hd_decap_12  FILLER_18_231
timestamp 1586364061
transform 1 0 22356 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_18_243
timestamp 1586364061
transform 1 0 23460 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
timestamp 1586364061
transform 1 0 25668 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1586364061
transform 1 0 26220 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_265
timestamp 1586364061
transform 1 0 25484 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_269
timestamp 1586364061
transform 1 0 25852 0 -1 12512
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1586364061
transform 1 0 28428 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_295
timestamp 1586364061
transform 1 0 28244 0 -1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
timestamp 1586364061
transform 1 0 28980 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
timestamp 1586364061
transform 1 0 28796 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_299
timestamp 1586364061
transform 1 0 28612 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_322
timestamp 1586364061
transform 1 0 30728 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
timestamp 1586364061
transform 1 0 32660 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
timestamp 1586364061
transform 1 0 33028 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
timestamp 1586364061
transform 1 0 32292 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_334
timestamp 1586364061
transform 1 0 31832 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_337
timestamp 1586364061
transform 1 0 32108 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_341
timestamp 1586364061
transform 1 0 32476 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_345
timestamp 1586364061
transform 1 0 32844 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1586364061
transform 1 0 35236 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_12  FILLER_18_349
timestamp 1586364061
transform 1 0 33212 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_361
timestamp 1586364061
transform 1 0 34316 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_369
timestamp 1586364061
transform 1 0 35052 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 36248 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_380
timestamp 1586364061
transform 1 0 36064 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_384
timestamp 1586364061
transform 1 0 36432 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_396
timestamp 1586364061
transform 1 0 37536 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_398
timestamp 1586364061
transform 1 0 37720 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_406
timestamp 1586364061
transform 1 0 38456 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_19_47
timestamp 1586364061
transform 1 0 5428 0 1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_46
timestamp 1586364061
transform 1 0 5336 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_19_56
timestamp 1586364061
transform 1 0 6256 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_52
timestamp 1586364061
transform 1 0 5888 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
timestamp 1586364061
transform 1 0 6072 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
timestamp 1586364061
transform 1 0 5704 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_73
timestamp 1586364061
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_69
timestamp 1586364061
transform 1 0 7452 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
timestamp 1586364061
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
timestamp 1586364061
transform 1 0 5704 0 -1 13600
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_20_81
timestamp 1586364061
transform 1 0 8556 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_81
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
timestamp 1586364061
transform 1 0 8188 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_20_89
timestamp 1586364061
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_85
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
timestamp 1586364061
transform 1 0 9108 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
timestamp 1586364061
transform 1 0 9292 0 1 12512
box -38 -48 406 592
use scs8hd_decap_4  FILLER_20_99
timestamp 1586364061
transform 1 0 10212 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_97
timestamp 1586364061
transform 1 0 10028 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_93
timestamp 1586364061
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 9844 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_6  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 10580 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 11316 0 -1 13600
box -38 -48 866 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_120
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_116
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_112
timestamp 1586364061
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_120
timestamp 1586364061
transform 1 0 12144 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_132
timestamp 1586364061
transform 1 0 13248 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_6  FILLER_19_131
timestamp 1586364061
transform 1 0 13156 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_127
timestamp 1586364061
transform 1 0 12788 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 12972 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_138
timestamp 1586364061
transform 1 0 13800 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_19_148
timestamp 1586364061
transform 1 0 14720 0 1 12512
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 13892 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 13708 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1586364061
transform 1 0 13892 0 1 12512
box -38 -48 866 592
use scs8hd_decap_12  FILLER_20_141
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_158
timestamp 1586364061
transform 1 0 15640 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_168
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_164
timestamp 1586364061
transform 1 0 16192 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 16008 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
timestamp 1586364061
transform 1 0 16652 0 -1 13600
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_192
timestamp 1586364061
transform 1 0 18768 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_188
timestamp 1586364061
transform 1 0 18400 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_190
timestamp 1586364061
transform 1 0 18584 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 18400 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1586364061
transform 1 0 18768 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_196
timestamp 1586364061
transform 1 0 19136 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 18952 0 -1 13600
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1586364061
transform 1 0 18952 0 1 12512
box -38 -48 866 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1586364061
transform 1 0 19228 0 -1 13600
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
timestamp 1586364061
transform 1 0 20516 0 1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
timestamp 1586364061
transform 1 0 20332 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
timestamp 1586364061
transform 1 0 19964 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_203
timestamp 1586364061
transform 1 0 19780 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_207
timestamp 1586364061
transform 1 0 20148 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
timestamp 1586364061
transform 1 0 23460 0 -1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
timestamp 1586364061
transform 1 0 23828 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_230
timestamp 1586364061
transform 1 0 22264 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_19_242
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_234
timestamp 1586364061
transform 1 0 22632 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_242
timestamp 1586364061
transform 1 0 23368 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_259
timestamp 1586364061
transform 1 0 24932 0 1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_19_253
timestamp 1586364061
transform 1 0 24380 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_249
timestamp 1586364061
transform 1 0 24012 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_clkbuf_1_1__f_clk_A
timestamp 1586364061
transform 1 0 25024 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
timestamp 1586364061
transform 1 0 24196 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 25392 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 25392 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_262
timestamp 1586364061
transform 1 0 25208 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_262
timestamp 1586364061
transform 1 0 25208 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 25760 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 25760 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_266
timestamp 1586364061
transform 1 0 25576 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_266
timestamp 1586364061
transform 1 0 25576 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_270
timestamp 1586364061
transform 1 0 25944 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 26036 0 -1 13600
box -38 -48 406 592
use scs8hd_clkbuf_16  clkbuf_1_1__f_clk
timestamp 1586364061
transform 1 0 25944 0 1 12512
box -38 -48 1878 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1586364061
transform 1 0 26588 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_3  FILLER_20_286
timestamp 1586364061
transform 1 0 27416 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_290
timestamp 1586364061
transform 1 0 27784 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1586364061
transform 1 0 27968 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1586364061
transform 1 0 27692 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_298
timestamp 1586364061
transform 1 0 28520 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_298
timestamp 1586364061
transform 1 0 28520 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_294
timestamp 1586364061
transform 1 0 28152 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1586364061
transform 1 0 28336 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_308
timestamp 1586364061
transform 1 0 29440 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_302
timestamp 1586364061
transform 1 0 28888 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_19_302
timestamp 1586364061
transform 1 0 28888 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1586364061
transform 1 0 28704 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 29624 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 29256 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1586364061
transform 1 0 28704 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1586364061
transform 1 0 29256 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_317
timestamp 1586364061
transform 1 0 30268 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_312
timestamp 1586364061
transform 1 0 29808 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_319
timestamp 1586364061
transform 1 0 30452 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_315
timestamp 1586364061
transform 1 0 30084 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 30452 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 30268 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
timestamp 1586364061
transform 1 0 30636 0 1 12512
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 29900 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_321
timestamp 1586364061
transform 1 0 30636 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_20_333
timestamp 1586364061
transform 1 0 31740 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_19_332
timestamp 1586364061
transform 1 0 31648 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_328
timestamp 1586364061
transform 1 0 31280 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
timestamp 1586364061
transform 1 0 31464 0 1 12512
box -38 -48 222 592
use scs8hd_or2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
timestamp 1586364061
transform 1 0 30820 0 1 12512
box -38 -48 498 592
use scs8hd_fill_2  FILLER_20_341
timestamp 1586364061
transform 1 0 32476 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_337
timestamp 1586364061
transform 1 0 32108 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
timestamp 1586364061
transform 1 0 32292 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
timestamp 1586364061
transform 1 0 32016 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 32016 0 -1 13600
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
timestamp 1586364061
transform 1 0 32200 0 1 12512
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
timestamp 1586364061
transform 1 0 32660 0 -1 13600
box -38 -48 1786 592
use scs8hd_decap_3  FILLER_19_357
timestamp 1586364061
transform 1 0 33948 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 34224 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_362
timestamp 1586364061
transform 1 0 34408 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_362
timestamp 1586364061
transform 1 0 34408 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 34592 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
timestamp 1586364061
transform 1 0 34592 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_367
timestamp 1586364061
transform 1 0 34868 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_366
timestamp 1586364061
transform 1 0 34776 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 35144 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 34960 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_372
timestamp 1586364061
transform 1 0 35328 0 1 12512
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 35144 0 -1 13600
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 35420 0 1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 37628 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_392
timestamp 1586364061
transform 1 0 37168 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_20_389
timestamp 1586364061
transform 1 0 36892 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_404
timestamp 1586364061
transform 1 0 38272 0 1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_398
timestamp 1586364061
transform 1 0 37720 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_406
timestamp 1586364061
transform 1 0 38456 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  FILLER_21_35
timestamp 1586364061
transform 1 0 4324 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_40
timestamp 1586364061
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1586364061
transform 1 0 6900 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_72
timestamp 1586364061
transform 1 0 7728 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_84
timestamp 1586364061
transform 1 0 8832 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_80
timestamp 1586364061
transform 1 0 8464 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_76
timestamp 1586364061
transform 1 0 8096 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
timestamp 1586364061
transform 1 0 8648 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 8280 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_93
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_89
timestamp 1586364061
transform 1 0 9292 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 9108 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 11040 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_106
timestamp 1586364061
transform 1 0 10856 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 774 592
use scs8hd_decap_12  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_21_147
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 590 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
timestamp 1586364061
transform 1 0 15456 0 1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
timestamp 1586364061
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_153
timestamp 1586364061
transform 1 0 15180 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1586364061
transform 1 0 18124 0 1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_21_198
timestamp 1586364061
transform 1 0 19320 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_194
timestamp 1586364061
transform 1 0 18952 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
timestamp 1586364061
transform 1 0 19688 0 1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
timestamp 1586364061
transform 1 0 19504 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_221
timestamp 1586364061
transform 1 0 21436 0 1 13600
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
timestamp 1586364061
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_233
timestamp 1586364061
transform 1 0 22540 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_237
timestamp 1586364061
transform 1 0 22908 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_240
timestamp 1586364061
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1586364061
transform 1 0 25392 0 1 13600
box -38 -48 866 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1586364061
transform 1 0 26220 0 1 13600
box -38 -48 866 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1586364061
transform 1 0 27048 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 28060 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 28428 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_291
timestamp 1586364061
transform 1 0 27876 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_295
timestamp 1586364061
transform 1 0 28244 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_306
timestamp 1586364061
transform 1 0 29256 0 1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_21_303
timestamp 1586364061
transform 1 0 28980 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_299
timestamp 1586364061
transform 1 0 28612 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 28796 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 29164 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_314
timestamp 1586364061
transform 1 0 29992 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 29808 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_322
timestamp 1586364061
transform 1 0 30728 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_318
timestamp 1586364061
transform 1 0 30360 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 30544 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 30176 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
timestamp 1586364061
transform 1 0 32292 0 1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
timestamp 1586364061
transform 1 0 32108 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 31740 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_330
timestamp 1586364061
transform 1 0 31464 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_335
timestamp 1586364061
transform 1 0 31924 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 35328 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 34776 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
timestamp 1586364061
transform 1 0 34500 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 35144 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_358
timestamp 1586364061
transform 1 0 34040 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_362
timestamp 1586364061
transform 1 0 34408 0 1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_21_365
timestamp 1586364061
transform 1 0 34684 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_21_367
timestamp 1586364061
transform 1 0 34868 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_391
timestamp 1586364061
transform 1 0 37076 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 38824 0 1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_21_403
timestamp 1586364061
transform 1 0 38180 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_22_46
timestamp 1586364061
transform 1 0 5336 0 -1 14688
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
timestamp 1586364061
transform 1 0 5796 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
timestamp 1586364061
transform 1 0 7728 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_50
timestamp 1586364061
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_70
timestamp 1586364061
transform 1 0 7544 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_74
timestamp 1586364061
transform 1 0 7912 0 -1 14688
box -38 -48 590 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 10028 0 -1 14688
box -38 -48 406 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 9844 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 11132 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10580 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_101
timestamp 1586364061
transform 1 0 10396 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_105
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_113
timestamp 1586364061
transform 1 0 11500 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_125
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_137
timestamp 1586364061
transform 1 0 13708 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_22_149
timestamp 1586364061
transform 1 0 14812 0 -1 14688
box -38 -48 406 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
timestamp 1586364061
transform 1 0 15456 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 16192 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_158
timestamp 1586364061
transform 1 0 15640 0 -1 14688
box -38 -48 590 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
timestamp 1586364061
transform 1 0 17940 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 17756 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_175
timestamp 1586364061
transform 1 0 17204 0 -1 14688
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_202
timestamp 1586364061
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
timestamp 1586364061
transform 1 0 23644 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 22816 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_235
timestamp 1586364061
transform 1 0 22724 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_22_238
timestamp 1586364061
transform 1 0 23000 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_244
timestamp 1586364061
transform 1 0 23552 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_247
timestamp 1586364061
transform 1 0 23828 0 -1 14688
box -38 -48 314 592
use scs8hd_clkbuf_16  clkbuf_0_clk
timestamp 1586364061
transform 1 0 24104 0 -1 14688
box -38 -48 1878 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 26220 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_270
timestamp 1586364061
transform 1 0 25944 0 -1 14688
box -38 -48 314 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1586364061
transform 1 0 26680 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 27692 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 28060 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 28428 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_287
timestamp 1586364061
transform 1 0 27508 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_291
timestamp 1586364061
transform 1 0 27876 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_295
timestamp 1586364061
transform 1 0 28244 0 -1 14688
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1586364061
transform 1 0 29808 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_12  FILLER_22_299
timestamp 1586364061
transform 1 0 28612 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_22_311
timestamp 1586364061
transform 1 0 29716 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_321
timestamp 1586364061
transform 1 0 30636 0 -1 14688
box -38 -48 1142 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1586364061
transform 1 0 32936 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 32016 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 32752 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 32384 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 31832 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_333
timestamp 1586364061
transform 1 0 31740 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_337
timestamp 1586364061
transform 1 0 32108 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_342
timestamp 1586364061
transform 1 0 32568 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
timestamp 1586364061
transform 1 0 34500 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
timestamp 1586364061
transform 1 0 34040 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_355
timestamp 1586364061
transform 1 0 33764 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_360
timestamp 1586364061
transform 1 0 34224 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 37628 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 36432 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_382
timestamp 1586364061
transform 1 0 36248 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_386
timestamp 1586364061
transform 1 0 36616 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  FILLER_22_394
timestamp 1586364061
transform 1 0 37352 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 38824 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_398
timestamp 1586364061
transform 1 0 37720 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_406
timestamp 1586364061
transform 1 0 38456 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_286
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 9292 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 8924 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_81
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_87
timestamp 1586364061
transform 1 0 9108 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_91
timestamp 1586364061
transform 1 0 9476 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_95
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_287
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 11316 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 11684 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_108
timestamp 1586364061
transform 1 0 11040 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_113
timestamp 1586364061
transform 1 0 11500 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_117
timestamp 1586364061
transform 1 0 11868 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_121
timestamp 1586364061
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_147
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_159
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_171
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_288
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
timestamp 1586364061
transform 1 0 18952 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_192
timestamp 1586364061
transform 1 0 18768 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_215
timestamp 1586364061
transform 1 0 20884 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_23_227
timestamp 1586364061
transform 1 0 21988 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_231
timestamp 1586364061
transform 1 0 22356 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_238
timestamp 1586364061
transform 1 0 23000 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_234
timestamp 1586364061
transform 1 0 22632 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_289
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 23920 0 1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
timestamp 1586364061
transform 1 0 24472 0 1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
timestamp 1586364061
transform 1 0 24288 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_250
timestamp 1586364061
transform 1 0 24104 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_273
timestamp 1586364061
transform 1 0 26220 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_278
timestamp 1586364061
transform 1 0 26680 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 26496 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_285
timestamp 1586364061
transform 1 0 27324 0 1 14688
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
timestamp 1586364061
transform 1 0 26956 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_293
timestamp 1586364061
transform 1 0 28060 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_289
timestamp 1586364061
transform 1 0 27692 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
timestamp 1586364061
transform 1 0 27876 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 27508 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_297
timestamp 1586364061
transform 1 0 28428 0 1 14688
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 28244 0 1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
timestamp 1586364061
transform 1 0 30452 0 1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_290
timestamp 1586364061
transform 1 0 29164 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
timestamp 1586364061
transform 1 0 29440 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
timestamp 1586364061
transform 1 0 30268 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
timestamp 1586364061
transform 1 0 29900 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
timestamp 1586364061
transform 1 0 28980 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_306
timestamp 1586364061
transform 1 0 29256 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_310
timestamp 1586364061
transform 1 0 29624 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_315
timestamp 1586364061
transform 1 0 30084 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1586364061
transform 1 0 32936 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 32476 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_338
timestamp 1586364061
transform 1 0 32200 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_343
timestamp 1586364061
transform 1 0 32660 0 1 14688
box -38 -48 314 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1586364061
transform 1 0 34868 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_291
timestamp 1586364061
transform 1 0 34776 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 34592 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 33948 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_355
timestamp 1586364061
transform 1 0 33764 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_359
timestamp 1586364061
transform 1 0 34132 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_363
timestamp 1586364061
transform 1 0 34500 0 1 14688
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 36432 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 36984 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 35880 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 36248 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_376
timestamp 1586364061
transform 1 0 35696 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_380
timestamp 1586364061
transform 1 0 36064 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_388
timestamp 1586364061
transform 1 0 36800 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_392
timestamp 1586364061
transform 1 0 37168 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 38824 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_404
timestamp 1586364061
transform 1 0 38272 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_292
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_46
timestamp 1586364061
transform 1 0 5336 0 -1 15776
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
timestamp 1586364061
transform 1 0 6348 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
timestamp 1586364061
transform 1 0 6164 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_54
timestamp 1586364061
transform 1 0 6072 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_76
timestamp 1586364061
transform 1 0 8096 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 8648 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 8280 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_88
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_293
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 11316 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11132 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_108
timestamp 1586364061
transform 1 0 11040 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
timestamp 1586364061
transform 1 0 13248 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_130
timestamp 1586364061
transform 1 0 13064 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_134
timestamp 1586364061
transform 1 0 13432 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_24_146
timestamp 1586364061
transform 1 0 14536 0 -1 15776
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_294
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_152
timestamp 1586364061
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_166
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
timestamp 1586364061
transform 1 0 19136 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_178
timestamp 1586364061
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_24_190
timestamp 1586364061
transform 1 0 18584 0 -1 15776
box -38 -48 590 592
use scs8hd_decap_12  FILLER_24_198
timestamp 1586364061
transform 1 0 19320 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_295
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_210
timestamp 1586364061
transform 1 0 20424 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1586364061
transform 1 0 22816 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 22356 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
timestamp 1586364061
transform 1 0 23828 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_229
timestamp 1586364061
transform 1 0 22172 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_233
timestamp 1586364061
transform 1 0 22540 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_245
timestamp 1586364061
transform 1 0 23644 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1586364061
transform 1 0 24380 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 25392 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 26220 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_249
timestamp 1586364061
transform 1 0 24012 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_262
timestamp 1586364061
transform 1 0 25208 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_266
timestamp 1586364061
transform 1 0 25576 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_272
timestamp 1586364061
transform 1 0 26128 0 -1 15776
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_296
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 27508 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_285
timestamp 1586364061
transform 1 0 27324 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_289
timestamp 1586364061
transform 1 0 27692 0 -1 15776
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
timestamp 1586364061
transform 1 0 29164 0 -1 15776
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_24_301
timestamp 1586364061
transform 1 0 28796 0 -1 15776
box -38 -48 406 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1586364061
transform 1 0 32476 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_297
timestamp 1586364061
transform 1 0 32016 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 32292 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1586364061
transform 1 0 31832 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_324
timestamp 1586364061
transform 1 0 30912 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_332
timestamp 1586364061
transform 1 0 31648 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_337
timestamp 1586364061
transform 1 0 32108 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_354
timestamp 1586364061
transform 1 0 33672 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_350
timestamp 1586364061
transform 1 0 33304 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 33856 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 33488 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_366
timestamp 1586364061
transform 1 0 34776 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_362
timestamp 1586364061
transform 1 0 34408 0 -1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 34868 0 -1 15776
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
timestamp 1586364061
transform 1 0 34040 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_369
timestamp 1586364061
transform 1 0 35052 0 -1 15776
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1586364061
transform 1 0 35144 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_298
timestamp 1586364061
transform 1 0 37628 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 36156 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_379
timestamp 1586364061
transform 1 0 35972 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_383
timestamp 1586364061
transform 1 0 36340 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_24_395
timestamp 1586364061
transform 1 0 37444 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 38824 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_398
timestamp 1586364061
transform 1 0 37720 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_24_406
timestamp 1586364061
transform 1 0 38456 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
timestamp 1586364061
transform 1 0 7176 0 1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_299
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
timestamp 1586364061
transform 1 0 6992 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
timestamp 1586364061
transform 1 0 9752 0 1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
timestamp 1586364061
transform 1 0 9568 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
timestamp 1586364061
transform 1 0 9200 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_85
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_90
timestamp 1586364061
transform 1 0 9384 0 1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_300
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_113
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_117
timestamp 1586364061
transform 1 0 11868 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_142
timestamp 1586364061
transform 1 0 14168 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_154
timestamp 1586364061
transform 1 0 15272 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_166
timestamp 1586364061
transform 1 0 16376 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_301
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_25_178
timestamp 1586364061
transform 1 0 17480 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_182
timestamp 1586364061
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_25_222
timestamp 1586364061
transform 1 0 21528 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_226
timestamp 1586364061
transform 1 0 21896 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 21712 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1586364061
transform 1 0 21988 0 1 15776
box -38 -48 866 592
use scs8hd_fill_2  FILLER_25_240
timestamp 1586364061
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_236
timestamp 1586364061
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 23920 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_302
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
timestamp 1586364061
transform 1 0 24472 0 1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
timestamp 1586364061
transform 1 0 24288 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_250
timestamp 1586364061
transform 1 0 24104 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_273
timestamp 1586364061
transform 1 0 26220 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1586364061
transform 1 0 26956 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
timestamp 1586364061
transform 1 0 28336 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 26772 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 26404 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_277
timestamp 1586364061
transform 1 0 26588 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_290
timestamp 1586364061
transform 1 0 27784 0 1 15776
box -38 -48 590 592
use scs8hd_fill_2  FILLER_25_298
timestamp 1586364061
transform 1 0 28520 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1586364061
transform 1 0 30084 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_303
timestamp 1586364061
transform 1 0 29164 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
timestamp 1586364061
transform 1 0 28704 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 29900 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 29532 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_302
timestamp 1586364061
transform 1 0 28888 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_25_306
timestamp 1586364061
transform 1 0 29256 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_311
timestamp 1586364061
transform 1 0 29716 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_324
timestamp 1586364061
transform 1 0 30912 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
timestamp 1586364061
transform 1 0 31096 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_332
timestamp 1586364061
transform 1 0 31648 0 1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_25_328
timestamp 1586364061
transform 1 0 31280 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_335
timestamp 1586364061
transform 1 0 31924 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1586364061
transform 1 0 31740 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1586364061
transform 1 0 32108 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_339
timestamp 1586364061
transform 1 0 32292 0 1 15776
box -38 -48 314 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 32568 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_346
timestamp 1586364061
transform 1 0 32936 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_350
timestamp 1586364061
transform 1 0 33304 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 33488 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 33120 0 1 15776
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 33672 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_362
timestamp 1586364061
transform 1 0 34408 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_358
timestamp 1586364061
transform 1 0 34040 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 34224 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_367
timestamp 1586364061
transform 1 0 34868 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 34592 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_304
timestamp 1586364061
transform 1 0 34776 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 35236 0 1 15776
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 35420 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 35972 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_377
timestamp 1586364061
transform 1 0 35788 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_381
timestamp 1586364061
transform 1 0 36156 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_393
timestamp 1586364061
transform 1 0 37260 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 38824 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_405
timestamp 1586364061
transform 1 0 38364 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_305
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use scs8hd_decap_8  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_312
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_70
timestamp 1586364061
transform 1 0 7544 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_64
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 7636 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
timestamp 1586364061
transform 1 0 7176 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
timestamp 1586364061
transform 1 0 7728 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1586364061
transform 1 0 7820 0 -1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 1786 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_306
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_82
timestamp 1586364061
transform 1 0 8648 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_8  FILLER_27_93
timestamp 1586364061
transform 1 0 9660 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_101
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_107
timestamp 1586364061
transform 1 0 10948 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_313
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 11316 0 -1 16864
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13248 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_130
timestamp 1586364061
transform 1 0 13064 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_134
timestamp 1586364061
transform 1 0 13432 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_26_146
timestamp 1586364061
transform 1 0 14536 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_136
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_148
timestamp 1586364061
transform 1 0 14720 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_307
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_152
timestamp 1586364061
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_166
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_160
timestamp 1586364061
transform 1 0 15824 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_172
timestamp 1586364061
transform 1 0 16928 0 1 16864
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_314
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_178
timestamp 1586364061
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_27_180
timestamp 1586364061
transform 1 0 17664 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_209
timestamp 1586364061
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_204
timestamp 1586364061
transform 1 0 19872 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 20148 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 20516 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_223
timestamp 1586364061
transform 1 0 21620 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 21436 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_308
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 20700 0 1 16864
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_27_232
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 22632 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_240
timestamp 1586364061
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_236
timestamp 1586364061
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_247
timestamp 1586364061
transform 1 0 23828 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_243
timestamp 1586364061
transform 1 0 23460 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
timestamp 1586364061
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
timestamp 1586364061
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
timestamp 1586364061
transform 1 0 23920 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_315
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 21712 0 -1 16864
box -38 -48 1786 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
timestamp 1586364061
transform 1 0 25208 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_250
timestamp 1586364061
transform 1 0 24104 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_260
timestamp 1586364061
transform 1 0 25024 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_264
timestamp 1586364061
transform 1 0 25392 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_26_272
timestamp 1586364061
transform 1 0 26128 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_264
timestamp 1586364061
transform 1 0 25392 0 1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_284
timestamp 1586364061
transform 1 0 27232 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_276
timestamp 1586364061
transform 1 0 26496 0 1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_26_284
timestamp 1586364061
transform 1 0 27232 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_280
timestamp 1586364061
transform 1 0 26864 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1586364061
transform 1 0 27048 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 27048 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_309
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_297
timestamp 1586364061
transform 1 0 28428 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_288
timestamp 1586364061
transform 1 0 27600 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1586364061
transform 1 0 27416 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
timestamp 1586364061
transform 1 0 28152 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 27416 0 -1 16864
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1586364061
transform 1 0 27600 0 1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
timestamp 1586364061
transform 1 0 28336 0 -1 16864
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
timestamp 1586364061
transform 1 0 29256 0 1 16864
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_316
timestamp 1586364061
transform 1 0 29164 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
timestamp 1586364061
transform 1 0 28980 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
timestamp 1586364061
transform 1 0 28612 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 30268 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_315
timestamp 1586364061
transform 1 0 30084 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_319
timestamp 1586364061
transform 1 0 30452 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_301
timestamp 1586364061
transform 1 0 28796 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_329
timestamp 1586364061
transform 1 0 31372 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_325
timestamp 1586364061
transform 1 0 31004 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_332
timestamp 1586364061
transform 1 0 31648 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_328
timestamp 1586364061
transform 1 0 31280 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_323
timestamp 1586364061
transform 1 0 30820 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 31556 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
timestamp 1586364061
transform 1 0 31188 0 1 16864
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
timestamp 1586364061
transform 1 0 30912 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_27_342
timestamp 1586364061
transform 1 0 32568 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_335
timestamp 1586364061
transform 1 0 31924 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 31740 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_310
timestamp 1586364061
transform 1 0 32016 0 -1 16864
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1586364061
transform 1 0 31740 0 1 16864
box -38 -48 866 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1586364061
transform 1 0 32108 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_4  FILLER_27_347
timestamp 1586364061
transform 1 0 33028 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_346
timestamp 1586364061
transform 1 0 32936 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 32844 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_351
timestamp 1586364061
transform 1 0 33396 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_356
timestamp 1586364061
transform 1 0 33856 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_350
timestamp 1586364061
transform 1 0 33304 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 33672 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 33120 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 33488 0 1 16864
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 33672 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_364
timestamp 1586364061
transform 1 0 34592 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_358
timestamp 1586364061
transform 1 0 34040 0 1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 34040 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 34408 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_317
timestamp 1586364061
transform 1 0 34776 0 1 16864
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1586364061
transform 1 0 34868 0 1 16864
box -38 -48 866 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1586364061
transform 1 0 34224 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_26_369
timestamp 1586364061
transform 1 0 35052 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 35236 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_380
timestamp 1586364061
transform 1 0 36064 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_376
timestamp 1586364061
transform 1 0 35696 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_373
timestamp 1586364061
transform 1 0 35420 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 35604 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 35880 0 1 16864
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 36432 0 1 16864
box -38 -48 406 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 35788 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_388
timestamp 1586364061
transform 1 0 36800 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_393
timestamp 1586364061
transform 1 0 37260 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 36984 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_311
timestamp 1586364061
transform 1 0 37628 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_392
timestamp 1586364061
transform 1 0 37168 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_381
timestamp 1586364061
transform 1 0 36156 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 38824 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 38824 0 1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_26_398
timestamp 1586364061
transform 1 0 37720 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_26_406
timestamp 1586364061
transform 1 0 38456 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_27_404
timestamp 1586364061
transform 1 0 38272 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_318
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
timestamp 1586364061
transform 1 0 7912 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_319
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_76
timestamp 1586364061
transform 1 0 8096 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_28_88
timestamp 1586364061
transform 1 0 9200 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11316 0 -1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_107
timestamp 1586364061
transform 1 0 10948 0 -1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 13248 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_130
timestamp 1586364061
transform 1 0 13064 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_134
timestamp 1586364061
transform 1 0 13432 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_28_146
timestamp 1586364061
transform 1 0 14536 0 -1 17952
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_320
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_152
timestamp 1586364061
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18860 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_178
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_28_190
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_195
timestamp 1586364061
transform 1 0 19044 0 -1 17952
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 21436 0 -1 17952
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_321
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_28_207
timestamp 1586364061
transform 1 0 20148 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_213
timestamp 1586364061
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 590 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
timestamp 1586364061
transform 1 0 23920 0 -1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
timestamp 1586364061
transform 1 0 23644 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_240
timestamp 1586364061
transform 1 0 23184 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_244
timestamp 1586364061
transform 1 0 23552 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_247
timestamp 1586364061
transform 1 0 23828 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_267
timestamp 1586364061
transform 1 0 25668 0 -1 17952
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
timestamp 1586364061
transform 1 0 28152 0 -1 17952
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_322
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1586364061
transform 1 0 27600 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_28_290
timestamp 1586364061
transform 1 0 27784 0 -1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
timestamp 1586364061
transform 1 0 30084 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_313
timestamp 1586364061
transform 1 0 29900 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_317
timestamp 1586364061
transform 1 0 30268 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_332
timestamp 1586364061
transform 1 0 31648 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_328
timestamp 1586364061
transform 1 0 31280 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_323
timestamp 1586364061
transform 1 0 30820 0 -1 17952
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
timestamp 1586364061
transform 1 0 30912 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_6  FILLER_28_337
timestamp 1586364061
transform 1 0 32108 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_335
timestamp 1586364061
transform 1 0 31924 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 31740 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_323
timestamp 1586364061
transform 1 0 32016 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 32660 0 -1 17952
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1586364061
transform 1 0 32844 0 -1 17952
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 34408 0 -1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 33856 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 34224 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_354
timestamp 1586364061
transform 1 0 33672 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_358
timestamp 1586364061
transform 1 0 34040 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_324
timestamp 1586364061
transform 1 0 37628 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_381
timestamp 1586364061
transform 1 0 36156 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_28_393
timestamp 1586364061
transform 1 0 37260 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 38824 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_398
timestamp 1586364061
transform 1 0 37720 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_28_406
timestamp 1586364061
transform 1 0 38456 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_325
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_98
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_326
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_147
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18860 0 1 17952
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_327
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18676 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_29_190
timestamp 1586364061
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_212
timestamp 1586364061
transform 1 0 20608 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_328
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_224
timestamp 1586364061
transform 1 0 21712 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_236
timestamp 1586364061
transform 1 0 22816 0 1 17952
box -38 -48 774 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 25760 0 1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 25576 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_29_265
timestamp 1586364061
transform 1 0 25484 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1586364061
transform 1 0 28428 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
timestamp 1586364061
transform 1 0 28060 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_287
timestamp 1586364061
transform 1 0 27508 0 1 17952
box -38 -48 590 592
use scs8hd_fill_2  FILLER_29_295
timestamp 1586364061
transform 1 0 28244 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1586364061
transform 1 0 29256 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_329
timestamp 1586364061
transform 1 0 29164 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
timestamp 1586364061
transform 1 0 30728 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
timestamp 1586364061
transform 1 0 28796 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1586364061
transform 1 0 30268 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_299
timestamp 1586364061
transform 1 0 28612 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_303
timestamp 1586364061
transform 1 0 28980 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_315
timestamp 1586364061
transform 1 0 30084 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_319
timestamp 1586364061
transform 1 0 30452 0 1 17952
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
timestamp 1586364061
transform 1 0 30912 0 1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
timestamp 1586364061
transform 1 0 32844 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_343
timestamp 1586364061
transform 1 0 32660 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_347
timestamp 1586364061
transform 1 0 33028 0 1 17952
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 33672 0 1 17952
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 34868 0 1 17952
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_330
timestamp 1586364061
transform 1 0 34776 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 34592 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
timestamp 1586364061
transform 1 0 33212 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 34224 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_351
timestamp 1586364061
transform 1 0 33396 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_358
timestamp 1586364061
transform 1 0 34040 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_362
timestamp 1586364061
transform 1 0 34408 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 36800 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_386
timestamp 1586364061
transform 1 0 36616 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_390
timestamp 1586364061
transform 1 0 36984 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 38824 0 1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_29_402
timestamp 1586364061
transform 1 0 38088 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_406
timestamp 1586364061
transform 1 0 38456 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_331
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_332
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_333
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_334
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 25760 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_267
timestamp 1586364061
transform 1 0 25668 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_270
timestamp 1586364061
transform 1 0 25944 0 -1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_335
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_274
timestamp 1586364061
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_30_288
timestamp 1586364061
transform 1 0 27600 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_30_296
timestamp 1586364061
transform 1 0 28336 0 -1 19040
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
timestamp 1586364061
transform 1 0 28796 0 -1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1586364061
transform 1 0 28612 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_320
timestamp 1586364061
transform 1 0 30544 0 -1 19040
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
timestamp 1586364061
transform 1 0 32660 0 -1 19040
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_336
timestamp 1586364061
transform 1 0 32016 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
timestamp 1586364061
transform 1 0 30912 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_326
timestamp 1586364061
transform 1 0 31096 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_334
timestamp 1586364061
transform 1 0 31832 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_337
timestamp 1586364061
transform 1 0 32108 0 -1 19040
box -38 -48 590 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 35144 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 34868 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_362
timestamp 1586364061
transform 1 0 34408 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_366
timestamp 1586364061
transform 1 0 34776 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_369
timestamp 1586364061
transform 1 0 35052 0 -1 19040
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_337
timestamp 1586364061
transform 1 0 37628 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 36156 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_379
timestamp 1586364061
transform 1 0 35972 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_383
timestamp 1586364061
transform 1 0 36340 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_30_395
timestamp 1586364061
transform 1 0 37444 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 38824 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_398
timestamp 1586364061
transform 1 0 37720 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_406
timestamp 1586364061
transform 1 0 38456 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_338
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_339
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_171
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_340
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_341
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 22816 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_234
timestamp 1586364061
transform 1 0 22632 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_238
timestamp 1586364061
transform 1 0 23000 0 1 19040
box -38 -48 590 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_281
timestamp 1586364061
transform 1 0 26956 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_293
timestamp 1586364061
transform 1 0 28060 0 1 19040
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
timestamp 1586364061
transform 1 0 29716 0 1 19040
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_342
timestamp 1586364061
transform 1 0 29164 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
timestamp 1586364061
transform 1 0 29532 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_306
timestamp 1586364061
transform 1 0 29256 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 32476 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_330
timestamp 1586364061
transform 1 0 31464 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_31_338
timestamp 1586364061
transform 1 0 32200 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_343
timestamp 1586364061
transform 1 0 32660 0 1 19040
box -38 -48 774 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 33672 0 1 19040
box -38 -48 406 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 34868 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_343
timestamp 1586364061
transform 1 0 34776 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 34592 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 34224 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 33488 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_351
timestamp 1586364061
transform 1 0 33396 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_358
timestamp 1586364061
transform 1 0 34040 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_362
timestamp 1586364061
transform 1 0 34408 0 1 19040
box -38 -48 222 592
use scs8hd_or2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
timestamp 1586364061
transform 1 0 36432 0 1 19040
box -38 -48 498 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
timestamp 1586364061
transform 1 0 37076 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 35880 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
timestamp 1586364061
transform 1 0 36248 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_376
timestamp 1586364061
transform 1 0 35696 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_380
timestamp 1586364061
transform 1 0 36064 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_389
timestamp 1586364061
transform 1 0 36892 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_393
timestamp 1586364061
transform 1 0 37260 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 38824 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_405
timestamp 1586364061
transform 1 0 38364 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_344
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_345
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_129
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_141
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_346
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_347
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 22448 0 -1 20128
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_231
timestamp 1586364061
transform 1 0 22356 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 24380 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 26128 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_255
timestamp 1586364061
transform 1 0 24564 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_32_267
timestamp 1586364061
transform 1 0 25668 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_271
timestamp 1586364061
transform 1 0 26036 0 -1 20128
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_348
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 26680 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 28336 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 27048 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_274
timestamp 1586364061
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_280
timestamp 1586364061
transform 1 0 26864 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_284
timestamp 1586364061
transform 1 0 27232 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_32_298
timestamp 1586364061
transform 1 0 28520 0 -1 20128
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
timestamp 1586364061
transform 1 0 29716 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 29348 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_306
timestamp 1586364061
transform 1 0 29256 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_309
timestamp 1586364061
transform 1 0 29532 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_313
timestamp 1586364061
transform 1 0 29900 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_349
timestamp 1586364061
transform 1 0 32016 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 32568 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 32936 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_325
timestamp 1586364061
transform 1 0 31004 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_3  FILLER_32_333
timestamp 1586364061
transform 1 0 31740 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_32_337
timestamp 1586364061
transform 1 0 32108 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_341
timestamp 1586364061
transform 1 0 32476 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_344
timestamp 1586364061
transform 1 0 32752 0 -1 20128
box -38 -48 222 592
use scs8hd_conb_1  _55_
timestamp 1586364061
transform 1 0 33672 0 -1 20128
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 34684 0 -1 20128
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 34500 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 33304 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_348
timestamp 1586364061
transform 1 0 33120 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_352
timestamp 1586364061
transform 1 0 33488 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_357
timestamp 1586364061
transform 1 0 33948 0 -1 20128
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_350
timestamp 1586364061
transform 1 0 37628 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_384
timestamp 1586364061
transform 1 0 36432 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_32_396
timestamp 1586364061
transform 1 0 37536 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 38824 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_398
timestamp 1586364061
transform 1 0 37720 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_406
timestamp 1586364061
transform 1 0 38456 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_357
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_351
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_358
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_352
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_359
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_159
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_353
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_34_210
timestamp 1586364061
transform 1 0 20424 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_6  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_217
timestamp 1586364061
transform 1 0 21068 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_214
timestamp 1586364061
transform 1 0 20792 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
timestamp 1586364061
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
timestamp 1586364061
transform 1 0 21252 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
timestamp 1586364061
transform 1 0 20884 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_360
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_221
timestamp 1586364061
transform 1 0 21436 0 1 20128
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1786 592
use scs8hd_decap_6  FILLER_34_234
timestamp 1586364061
transform 1 0 22632 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_33_233
timestamp 1586364061
transform 1 0 22540 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 22632 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_240
timestamp 1586364061
transform 1 0 23184 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_236
timestamp 1586364061
transform 1 0 22816 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 23184 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23000 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_354
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 23368 0 -1 21216
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 26128 0 1 20128
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 25944 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 26220 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 25576 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 25852 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_264
timestamp 1586364061
transform 1 0 25392 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_268
timestamp 1586364061
transform 1 0 25760 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_261
timestamp 1586364061
transform 1 0 25116 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_271
timestamp 1586364061
transform 1 0 26036 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_285
timestamp 1586364061
transform 1 0 27324 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_361
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_1  FILLER_34_295
timestamp 1586364061
transform 1 0 28244 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_34_289
timestamp 1586364061
transform 1 0 27692 0 -1 21216
box -38 -48 590 592
use scs8hd_decap_4  FILLER_33_298
timestamp 1586364061
transform 1 0 28520 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_295
timestamp 1586364061
transform 1 0 28244 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_291
timestamp 1586364061
transform 1 0 27876 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 27508 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 28336 0 1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 28336 0 -1 21216
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_33_306
timestamp 1586364061
transform 1 0 29256 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_302
timestamp 1586364061
transform 1 0 28888 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 28980 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_355
timestamp 1586364061
transform 1 0 29164 0 1 20128
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 29348 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_315
timestamp 1586364061
transform 1 0 30084 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_316
timestamp 1586364061
transform 1 0 30176 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 30268 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_319
timestamp 1586364061
transform 1 0 30452 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_320
timestamp 1586364061
transform 1 0 30544 0 1 20128
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 30360 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 30636 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_326
timestamp 1586364061
transform 1 0 31096 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_334
timestamp 1586364061
transform 1 0 31832 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_328
timestamp 1586364061
transform 1 0 31280 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 31832 0 -1 21216
box -38 -48 222 592
use scs8hd_conb_1  _58_
timestamp 1586364061
transform 1 0 31556 0 1 20128
box -38 -48 314 592
use scs8hd_conb_1  _33_
timestamp 1586364061
transform 1 0 30820 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_337
timestamp 1586364061
transform 1 0 32108 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_338
timestamp 1586364061
transform 1 0 32200 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 32292 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 32016 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 32384 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_362
timestamp 1586364061
transform 1 0 32016 0 -1 21216
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 32568 0 1 20128
box -38 -48 866 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 32476 0 -1 21216
box -38 -48 2246 592
use scs8hd_decap_4  FILLER_33_355
timestamp 1586364061
transform 1 0 33764 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_351
timestamp 1586364061
transform 1 0 33396 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 33580 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_365
timestamp 1586364061
transform 1 0 34684 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_362
timestamp 1586364061
transform 1 0 34408 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_359
timestamp 1586364061
transform 1 0 34132 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 34224 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 34592 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 34868 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_356
timestamp 1586364061
transform 1 0 34776 0 1 20128
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 34868 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_369
timestamp 1586364061
transform 1 0 35052 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 35236 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_384
timestamp 1586364061
transform 1 0 36432 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_380
timestamp 1586364061
transform 1 0 36064 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_376
timestamp 1586364061
transform 1 0 35696 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 36248 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 35880 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 35420 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_3  FILLER_34_394
timestamp 1586364061
transform 1 0 37352 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 36616 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_363
timestamp 1586364061
transform 1 0 37628 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_382
timestamp 1586364061
transform 1 0 36248 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_388
timestamp 1586364061
transform 1 0 36800 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 38824 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 38824 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_6  FILLER_33_400
timestamp 1586364061
transform 1 0 37904 0 1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_33_406
timestamp 1586364061
transform 1 0 38456 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_34_398
timestamp 1586364061
transform 1 0 37720 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_406
timestamp 1586364061
transform 1 0 38456 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_364
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_365
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_147
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_159
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_171
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_366
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
timestamp 1586364061
transform 1 0 20976 0 1 21216
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
timestamp 1586364061
transform 1 0 20792 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
timestamp 1586364061
transform 1 0 20424 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
timestamp 1586364061
transform 1 0 20056 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_204
timestamp 1586364061
transform 1 0 19872 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_212
timestamp 1586364061
transform 1 0 20608 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_367
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 23000 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_235
timestamp 1586364061
transform 1 0 22724 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_240
timestamp 1586364061
transform 1 0 23184 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_258
timestamp 1586364061
transform 1 0 24840 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_254
timestamp 1586364061
transform 1 0 24472 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 25024 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 24656 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_265
timestamp 1586364061
transform 1 0 25484 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 25668 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 26036 0 1 21216
box -38 -48 222 592
use scs8hd_conb_1  _34_
timestamp 1586364061
transform 1 0 25208 0 1 21216
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 26220 0 1 21216
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 28152 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_292
timestamp 1586364061
transform 1 0 27968 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_296
timestamp 1586364061
transform 1 0 28336 0 1 21216
box -38 -48 314 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 29256 0 1 21216
box -38 -48 2246 592
use scs8hd_tapvpwrvgnd_1  PHY_368
timestamp 1586364061
transform 1 0 29164 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 28980 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 28612 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_301
timestamp 1586364061
transform 1 0 28796 0 1 21216
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 32200 0 1 21216
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 32016 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 31648 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_330
timestamp 1586364061
transform 1 0 31464 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_334
timestamp 1586364061
transform 1 0 31832 0 1 21216
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 34868 0 1 21216
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_369
timestamp 1586364061
transform 1 0 34776 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 34316 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_357
timestamp 1586364061
transform 1 0 33948 0 1 21216
box -38 -48 406 592
use scs8hd_decap_3  FILLER_35_363
timestamp 1586364061
transform 1 0 34500 0 1 21216
box -38 -48 314 592
use scs8hd_conb_1  _56_
timestamp 1586364061
transform 1 0 37352 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 36800 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_386
timestamp 1586364061
transform 1 0 36616 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_390
timestamp 1586364061
transform 1 0 36984 0 1 21216
box -38 -48 406 592
use scs8hd_decap_8  FILLER_35_397
timestamp 1586364061
transform 1 0 37628 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 38824 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_405
timestamp 1586364061
transform 1 0 38364 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_370
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_371
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_372
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_373
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1586364061
transform 1 0 23368 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 23184 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_234
timestamp 1586364061
transform 1 0 22632 0 -1 22304
box -38 -48 590 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 24932 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 24380 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 26220 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_255
timestamp 1586364061
transform 1 0 24564 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_36_261
timestamp 1586364061
transform 1 0 25116 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_267
timestamp 1586364061
transform 1 0 25668 0 -1 22304
box -38 -48 590 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 26772 0 -1 22304
box -38 -48 2246 592
use scs8hd_tapvpwrvgnd_1  PHY_374
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 314 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 29716 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 29532 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 29164 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 30728 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_303
timestamp 1586364061
transform 1 0 28980 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_307
timestamp 1586364061
transform 1 0 29348 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_320
timestamp 1586364061
transform 1 0 30544 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 32108 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_375
timestamp 1586364061
transform 1 0 32016 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 31832 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_324
timestamp 1586364061
transform 1 0 30912 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_36_332
timestamp 1586364061
transform 1 0 31648 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_346
timestamp 1586364061
transform 1 0 32936 0 -1 22304
box -38 -48 406 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 34316 0 -1 22304
box -38 -48 2246 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 34132 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 33764 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 33396 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_350
timestamp 1586364061
transform 1 0 33304 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_353
timestamp 1586364061
transform 1 0 33580 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_357
timestamp 1586364061
transform 1 0 33948 0 -1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_376
timestamp 1586364061
transform 1 0 37628 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 36708 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_385
timestamp 1586364061
transform 1 0 36524 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_389
timestamp 1586364061
transform 1 0 36892 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 38824 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_398
timestamp 1586364061
transform 1 0 37720 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_1  FILLER_36_406
timestamp 1586364061
transform 1 0 38456 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_377
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_378
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_147
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_159
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_171
timestamp 1586364061
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_379
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 774 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1586364061
transform 1 0 21528 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
timestamp 1586364061
transform 1 0 20884 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
timestamp 1586364061
transform 1 0 20516 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 20148 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_204
timestamp 1586364061
transform 1 0 19872 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_209
timestamp 1586364061
transform 1 0 20332 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_213
timestamp 1586364061
transform 1 0 20700 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_217
timestamp 1586364061
transform 1 0 21068 0 1 22304
box -38 -48 314 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_380
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 22540 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 23000 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_231
timestamp 1586364061
transform 1 0 22356 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_235
timestamp 1586364061
transform 1 0 22724 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_240
timestamp 1586364061
transform 1 0 23184 0 1 22304
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 25208 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 25760 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 24656 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 25024 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_254
timestamp 1586364061
transform 1 0 24472 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_258
timestamp 1586364061
transform 1 0 24840 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_266
timestamp 1586364061
transform 1 0 25576 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_270
timestamp 1586364061
transform 1 0 25944 0 1 22304
box -38 -48 406 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 26864 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 26680 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 27876 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 28244 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 26312 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_276
timestamp 1586364061
transform 1 0 26496 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_289
timestamp 1586364061
transform 1 0 27692 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_293
timestamp 1586364061
transform 1 0 28060 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_297
timestamp 1586364061
transform 1 0 28428 0 1 22304
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 29256 0 1 22304
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_381
timestamp 1586364061
transform 1 0 29164 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 28980 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 28612 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_301
timestamp 1586364061
transform 1 0 28796 0 1 22304
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 32200 0 1 22304
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 32016 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 31648 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_325
timestamp 1586364061
transform 1 0 31004 0 1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_37_331
timestamp 1586364061
transform 1 0 31556 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_334
timestamp 1586364061
transform 1 0 31832 0 1 22304
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 35328 0 1 22304
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_382
timestamp 1586364061
transform 1 0 34776 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 35144 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 34592 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 34224 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_357
timestamp 1586364061
transform 1 0 33948 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_362
timestamp 1586364061
transform 1 0 34408 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_367
timestamp 1586364061
transform 1 0 34868 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_391
timestamp 1586364061
transform 1 0 37076 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 38824 0 1 22304
box -38 -48 314 592
use scs8hd_decap_4  FILLER_37_403
timestamp 1586364061
transform 1 0 38180 0 1 22304
box -38 -48 406 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_383
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_384
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_141
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_385
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_166
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_178
timestamp 1586364061
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_386
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 20608 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_202
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_38_210
timestamp 1586364061
transform 1 0 20424 0 -1 23392
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1586364061
transform 1 0 23368 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 22816 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 23184 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_234
timestamp 1586364061
transform 1 0 22632 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_238
timestamp 1586364061
transform 1 0 23000 0 -1 23392
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 24932 0 -1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 24380 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 24748 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_255
timestamp 1586364061
transform 1 0 24564 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 27876 0 -1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_387
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 27600 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 26864 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 28428 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_6  FILLER_38_282
timestamp 1586364061
transform 1 0 27048 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_38_290
timestamp 1586364061
transform 1 0 27784 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_295
timestamp 1586364061
transform 1 0 28244 0 -1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 28980 0 -1 23392
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 28796 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_299
timestamp 1586364061
transform 1 0 28612 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_322
timestamp 1586364061
transform 1 0 30728 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_388
timestamp 1586364061
transform 1 0 32016 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_334
timestamp 1586364061
transform 1 0 31832 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_337
timestamp 1586364061
transform 1 0 32108 0 -1 23392
box -38 -48 1142 592
use scs8hd_conb_1  _57_
timestamp 1586364061
transform 1 0 34132 0 -1 23392
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 35144 0 -1 23392
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 34868 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_349
timestamp 1586364061
transform 1 0 33212 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_38_357
timestamp 1586364061
transform 1 0 33948 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_362
timestamp 1586364061
transform 1 0 34408 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_366
timestamp 1586364061
transform 1 0 34776 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_369
timestamp 1586364061
transform 1 0 35052 0 -1 23392
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_389
timestamp 1586364061
transform 1 0 37628 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_389
timestamp 1586364061
transform 1 0 36892 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 38824 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_398
timestamp 1586364061
transform 1 0 37720 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_38_406
timestamp 1586364061
transform 1 0 38456 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_396
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_27
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_39
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_390
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_51
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_397
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_391
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_147
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_398
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_159
timestamp 1586364061
transform 1 0 15732 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_171
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_392
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_196
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_206
timestamp 1586364061
transform 1 0 20056 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 19872 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
timestamp 1586364061
transform 1 0 20516 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 20608 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_210
timestamp 1586364061
transform 1 0 20424 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_210
timestamp 1586364061
transform 1 0 20424 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_213
timestamp 1586364061
transform 1 0 20700 0 -1 24480
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_399
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 20976 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_214
timestamp 1586364061
transform 1 0 20792 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 314 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1586364061
transform 1 0 21160 0 1 23392
box -38 -48 866 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1586364061
transform 1 0 21160 0 -1 24480
box -38 -48 866 592
use scs8hd_decap_8  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_4  FILLER_39_231
timestamp 1586364061
transform 1 0 22356 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_227
timestamp 1586364061
transform 1 0 21988 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 22172 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_241
timestamp 1586364061
transform 1 0 23276 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_237
timestamp 1586364061
transform 1 0 22908 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 23092 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 22724 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1586364061
transform 1 0 22724 0 -1 24480
box -38 -48 866 592
use scs8hd_decap_6  FILLER_40_244
timestamp 1586364061
transform 1 0 23552 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 23828 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_393
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_249
timestamp 1586364061
transform 1 0 24012 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1586364061
transform 1 0 24104 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 24196 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 866 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1586364061
transform 1 0 24288 0 -1 24480
box -38 -48 866 592
use scs8hd_decap_8  FILLER_40_265
timestamp 1586364061
transform 1 0 25484 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_40_261
timestamp 1586364061
transform 1 0 25116 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_266
timestamp 1586364061
transform 1 0 25576 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_262
timestamp 1586364061
transform 1 0 25208 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 25760 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 25392 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_273
timestamp 1586364061
transform 1 0 26220 0 -1 24480
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 25944 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_400
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 26496 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 26680 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_274
timestamp 1586364061
transform 1 0 26312 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_278
timestamp 1586364061
transform 1 0 26680 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 26956 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_280
timestamp 1586364061
transform 1 0 26864 0 -1 24480
box -38 -48 406 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 27324 0 -1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 27324 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_283
timestamp 1586364061
transform 1 0 27140 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_284
timestamp 1586364061
transform 1 0 27232 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_293
timestamp 1586364061
transform 1 0 28060 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_289
timestamp 1586364061
transform 1 0 27692 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_297
timestamp 1586364061
transform 1 0 28428 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_287
timestamp 1586364061
transform 1 0 27508 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 27876 0 -1 24480
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 27600 0 1 23392
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 28428 0 -1 24480
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_39_301
timestamp 1586364061
transform 1 0 28796 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 28980 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 28612 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_394
timestamp 1586364061
transform 1 0 29164 0 1 23392
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 29256 0 1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_316
timestamp 1586364061
transform 1 0 30176 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_319
timestamp 1586364061
transform 1 0 30452 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_315
timestamp 1586364061
transform 1 0 30084 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 30636 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 30268 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 30360 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_320
timestamp 1586364061
transform 1 0 30544 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_40_332
timestamp 1586364061
transform 1 0 31648 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 31832 0 -1 24480
box -38 -48 222 592
use scs8hd_conb_1  _32_
timestamp 1586364061
transform 1 0 30820 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_345
timestamp 1586364061
transform 1 0 32844 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_40_337
timestamp 1586364061
transform 1 0 32108 0 -1 24480
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 33028 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 32660 0 -1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_401
timestamp 1586364061
transform 1 0 32016 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_338
timestamp 1586364061
transform 1 0 32200 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_326
timestamp 1586364061
transform 1 0 31096 0 1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_357
timestamp 1586364061
transform 1 0 33948 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_353
timestamp 1586364061
transform 1 0 33580 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_349
timestamp 1586364061
transform 1 0 33212 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_350
timestamp 1586364061
transform 1 0 33304 0 1 23392
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 33396 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 34408 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 34224 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 34040 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_358
timestamp 1586364061
transform 1 0 34040 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_362
timestamp 1586364061
transform 1 0 34408 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_360
timestamp 1586364061
transform 1 0 34224 0 -1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_395
timestamp 1586364061
transform 1 0 34776 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 34868 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 34592 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_364
timestamp 1586364061
transform 1 0 34592 0 -1 24480
box -38 -48 314 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 34868 0 1 23392
box -38 -48 866 592
use scs8hd_decap_3  FILLER_40_369
timestamp 1586364061
transform 1 0 35052 0 -1 24480
box -38 -48 314 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 35328 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_39_384
timestamp 1586364061
transform 1 0 36432 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_380
timestamp 1586364061
transform 1 0 36064 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_376
timestamp 1586364061
transform 1 0 35696 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 36248 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 35880 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_393
timestamp 1586364061
transform 1 0 37260 0 -1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 36616 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_402
timestamp 1586364061
transform 1 0 37628 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_381
timestamp 1586364061
transform 1 0 36156 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_388
timestamp 1586364061
transform 1 0 36800 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 38824 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 38824 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_6  FILLER_39_400
timestamp 1586364061
transform 1 0 37904 0 1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_39_406
timestamp 1586364061
transform 1 0 38456 0 1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_40_398
timestamp 1586364061
transform 1 0 37720 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_1  FILLER_40_406
timestamp 1586364061
transform 1 0 38456 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_403
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_404
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_405
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
timestamp 1586364061
transform 1 0 20516 0 1 24480
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
timestamp 1586364061
transform 1 0 20332 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
timestamp 1586364061
transform 1 0 19964 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_204
timestamp 1586364061
transform 1 0 19872 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_207
timestamp 1586364061
transform 1 0 20148 0 1 24480
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_406
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
timestamp 1586364061
transform 1 0 23368 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_230
timestamp 1586364061
transform 1 0 22264 0 1 24480
box -38 -48 1142 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1586364061
transform 1 0 25024 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1586364061
transform 1 0 24196 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1586364061
transform 1 0 24564 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 26036 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_249
timestamp 1586364061
transform 1 0 24012 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_253
timestamp 1586364061
transform 1 0 24380 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_273
timestamp 1586364061
transform 1 0 26220 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1586364061
transform 1 0 26588 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 26404 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 27600 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 27968 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 28336 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_286
timestamp 1586364061
transform 1 0 27416 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_290
timestamp 1586364061
transform 1 0 27784 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_294
timestamp 1586364061
transform 1 0 28152 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_298
timestamp 1586364061
transform 1 0 28520 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_302
timestamp 1586364061
transform 1 0 28888 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 28704 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_306
timestamp 1586364061
transform 1 0 29256 0 1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_407
timestamp 1586364061
transform 1 0 29164 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_311
timestamp 1586364061
transform 1 0 29716 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 29532 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_315
timestamp 1586364061
transform 1 0 30084 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 29900 0 1 24480
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 30176 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_320
timestamp 1586364061
transform 1 0 30544 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 30728 0 1 24480
box -38 -48 222 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 31832 0 1 24480
box -38 -48 2246 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 31648 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 31280 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_324
timestamp 1586364061
transform 1 0 30912 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_330
timestamp 1586364061
transform 1 0 31464 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 34868 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_408
timestamp 1586364061
transform 1 0 34776 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 34408 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_358
timestamp 1586364061
transform 1 0 34040 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_364
timestamp 1586364061
transform 1 0 34592 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 35880 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 36248 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_376
timestamp 1586364061
transform 1 0 35696 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_380
timestamp 1586364061
transform 1 0 36064 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_384
timestamp 1586364061
transform 1 0 36432 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_396
timestamp 1586364061
transform 1 0 37536 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 38824 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_41_404
timestamp 1586364061
transform 1 0 38272 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_409
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_68
timestamp 1586364061
transform 1 0 7360 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_410
timestamp 1586364061
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_80
timestamp 1586364061
transform 1 0 8464 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_93
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_105
timestamp 1586364061
transform 1 0 10764 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_117
timestamp 1586364061
transform 1 0 11868 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_129
timestamp 1586364061
transform 1 0 12972 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_141
timestamp 1586364061
transform 1 0 14076 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_411
timestamp 1586364061
transform 1 0 15180 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_154
timestamp 1586364061
transform 1 0 15272 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_166
timestamp 1586364061
transform 1 0 16376 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_178
timestamp 1586364061
transform 1 0 17480 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_190
timestamp 1586364061
transform 1 0 18584 0 -1 25568
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
timestamp 1586364061
transform 1 0 20884 0 -1 25568
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_412
timestamp 1586364061
transform 1 0 20792 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_202
timestamp 1586364061
transform 1 0 19688 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_1  FILLER_42_210
timestamp 1586364061
transform 1 0 20424 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_1  FILLER_42_213
timestamp 1586364061
transform 1 0 20700 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
timestamp 1586364061
transform 1 0 23552 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_234
timestamp 1586364061
transform 1 0 22632 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_246
timestamp 1586364061
transform 1 0 23736 0 -1 25568
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1586364061
transform 1 0 24104 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1586364061
transform 1 0 25484 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_259
timestamp 1586364061
transform 1 0 24932 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_263
timestamp 1586364061
transform 1 0 25300 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_42_267
timestamp 1586364061
transform 1 0 25668 0 -1 25568
box -38 -48 590 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1586364061
transform 1 0 27876 0 -1 25568
box -38 -48 866 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 26772 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_413
timestamp 1586364061
transform 1 0 26404 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
timestamp 1586364061
transform 1 0 27324 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_276
timestamp 1586364061
transform 1 0 26496 0 -1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_42_283
timestamp 1586364061
transform 1 0 27140 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_287
timestamp 1586364061
transform 1 0 27508 0 -1 25568
box -38 -48 406 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 29532 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 29256 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_42_300
timestamp 1586364061
transform 1 0 28704 0 -1 25568
box -38 -48 590 592
use scs8hd_fill_1  FILLER_42_308
timestamp 1586364061
transform 1 0 29440 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_318
timestamp 1586364061
transform 1 0 30360 0 -1 25568
box -38 -48 1142 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 32660 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_414
timestamp 1586364061
transform 1 0 32016 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 31832 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 32384 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_330
timestamp 1586364061
transform 1 0 31464 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_3  FILLER_42_337
timestamp 1586364061
transform 1 0 32108 0 -1 25568
box -38 -48 314 592
use scs8hd_fill_1  FILLER_42_342
timestamp 1586364061
transform 1 0 32568 0 -1 25568
box -38 -48 130 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 34408 0 -1 25568
box -38 -48 2246 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 33672 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 34224 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_352
timestamp 1586364061
transform 1 0 33488 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_356
timestamp 1586364061
transform 1 0 33856 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_415
timestamp 1586364061
transform 1 0 37628 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_386
timestamp 1586364061
transform 1 0 36616 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_3  FILLER_42_394
timestamp 1586364061
transform 1 0 37352 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 38824 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_8  FILLER_42_398
timestamp 1586364061
transform 1 0 37720 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_1  FILLER_42_406
timestamp 1586364061
transform 1 0 38456 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_3  PHY_86
timestamp 1586364061
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_43_3
timestamp 1586364061
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_15
timestamp 1586364061
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_27
timestamp 1586364061
transform 1 0 3588 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_39
timestamp 1586364061
transform 1 0 4692 0 1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_416
timestamp 1586364061
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_43_51
timestamp 1586364061
transform 1 0 5796 0 1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_43_59
timestamp 1586364061
transform 1 0 6532 0 1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_43_62
timestamp 1586364061
transform 1 0 6808 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_74
timestamp 1586364061
transform 1 0 7912 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_86
timestamp 1586364061
transform 1 0 9016 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_98
timestamp 1586364061
transform 1 0 10120 0 1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_417
timestamp 1586364061
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_43_110
timestamp 1586364061
transform 1 0 11224 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_123
timestamp 1586364061
transform 1 0 12420 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_135
timestamp 1586364061
transform 1 0 13524 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_147
timestamp 1586364061
transform 1 0 14628 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_159
timestamp 1586364061
transform 1 0 15732 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_171
timestamp 1586364061
transform 1 0 16836 0 1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_418
timestamp 1586364061
transform 1 0 17940 0 1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_43_184
timestamp 1586364061
transform 1 0 18032 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_196
timestamp 1586364061
transform 1 0 19136 0 1 25568
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
timestamp 1586364061
transform 1 0 20884 0 1 25568
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
timestamp 1586364061
transform 1 0 20700 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
timestamp 1586364061
transform 1 0 20332 0 1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_43_208
timestamp 1586364061
transform 1 0 20240 0 1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_43_211
timestamp 1586364061
transform 1 0 20516 0 1 25568
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
timestamp 1586364061
transform 1 0 23920 0 1 25568
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_419
timestamp 1586364061
transform 1 0 23552 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
timestamp 1586364061
transform 1 0 23368 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
timestamp 1586364061
transform 1 0 22816 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_234
timestamp 1586364061
transform 1 0 22632 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_238
timestamp 1586364061
transform 1 0 23000 0 1 25568
box -38 -48 406 592
use scs8hd_decap_3  FILLER_43_245
timestamp 1586364061
transform 1 0 23644 0 1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
timestamp 1586364061
transform 1 0 26220 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
timestamp 1586364061
transform 1 0 25852 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_267
timestamp 1586364061
transform 1 0 25668 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_271
timestamp 1586364061
transform 1 0 26036 0 1 25568
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
timestamp 1586364061
transform 1 0 26404 0 1 25568
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_43_294
timestamp 1586364061
transform 1 0 28152 0 1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_43_298
timestamp 1586364061
transform 1 0 28520 0 1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_43_310
timestamp 1586364061
transform 1 0 29624 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_301
timestamp 1586364061
transform 1 0 28796 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 28612 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 28980 0 1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_420
timestamp 1586364061
transform 1 0 29164 0 1 25568
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 29256 0 1 25568
box -38 -48 406 592
use scs8hd_fill_2  FILLER_43_314
timestamp 1586364061
transform 1 0 29992 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 29808 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 30176 0 1 25568
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 30360 0 1 25568
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 32384 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 33028 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_43_337
timestamp 1586364061
transform 1 0 32108 0 1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_43_342
timestamp 1586364061
transform 1 0 32568 0 1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_43_346
timestamp 1586364061
transform 1 0 32936 0 1 25568
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 34868 0 1 25568
box -38 -48 866 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 33212 0 1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_421
timestamp 1586364061
transform 1 0 34776 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 34592 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 34224 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_358
timestamp 1586364061
transform 1 0 34040 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_362
timestamp 1586364061
transform 1 0 34408 0 1 25568
box -38 -48 222 592
use scs8hd_conb_1  _61_
timestamp 1586364061
transform 1 0 36432 0 1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 35880 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 36248 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_376
timestamp 1586364061
transform 1 0 35696 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_380
timestamp 1586364061
transform 1 0 36064 0 1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_43_387
timestamp 1586364061
transform 1 0 36708 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_87
timestamp 1586364061
transform -1 0 38824 0 1 25568
box -38 -48 314 592
use scs8hd_decap_8  FILLER_43_399
timestamp 1586364061
transform 1 0 37812 0 1 25568
box -38 -48 774 592
use scs8hd_decap_3  PHY_88
timestamp 1586364061
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_44_3
timestamp 1586364061
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_15
timestamp 1586364061
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_422
timestamp 1586364061
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_4  FILLER_44_27
timestamp 1586364061
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use scs8hd_decap_12  FILLER_44_32
timestamp 1586364061
transform 1 0 4048 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_44
timestamp 1586364061
transform 1 0 5152 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_56
timestamp 1586364061
transform 1 0 6256 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_68
timestamp 1586364061
transform 1 0 7360 0 -1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_423
timestamp 1586364061
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_44_80
timestamp 1586364061
transform 1 0 8464 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_93
timestamp 1586364061
transform 1 0 9660 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_105
timestamp 1586364061
transform 1 0 10764 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_117
timestamp 1586364061
transform 1 0 11868 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_129
timestamp 1586364061
transform 1 0 12972 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_141
timestamp 1586364061
transform 1 0 14076 0 -1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_424
timestamp 1586364061
transform 1 0 15180 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_44_154
timestamp 1586364061
transform 1 0 15272 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_166
timestamp 1586364061
transform 1 0 16376 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_178
timestamp 1586364061
transform 1 0 17480 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_190
timestamp 1586364061
transform 1 0 18584 0 -1 26656
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
timestamp 1586364061
transform 1 0 21436 0 -1 26656
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_425
timestamp 1586364061
transform 1 0 20792 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
timestamp 1586364061
transform 1 0 21068 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_44_202
timestamp 1586364061
transform 1 0 19688 0 -1 26656
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_44_215
timestamp 1586364061
transform 1 0 20884 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_219
timestamp 1586364061
transform 1 0 21252 0 -1 26656
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
timestamp 1586364061
transform 1 0 23920 0 -1 26656
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
timestamp 1586364061
transform 1 0 23736 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_6  FILLER_44_240
timestamp 1586364061
transform 1 0 23184 0 -1 26656
box -38 -48 590 592
use scs8hd_decap_8  FILLER_44_267
timestamp 1586364061
transform 1 0 25668 0 -1 26656
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
timestamp 1586364061
transform 1 0 26496 0 -1 26656
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_426
timestamp 1586364061
transform 1 0 26404 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 28520 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_44_295
timestamp 1586364061
transform 1 0 28244 0 -1 26656
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 28980 0 -1 26656
box -38 -48 1786 592
use scs8hd_decap_3  FILLER_44_300
timestamp 1586364061
transform 1 0 28704 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_8  FILLER_44_322
timestamp 1586364061
transform 1 0 30728 0 -1 26656
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 32384 0 -1 26656
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_427
timestamp 1586364061
transform 1 0 32016 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 31832 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 31464 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_332
timestamp 1586364061
transform 1 0 31648 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_44_337
timestamp 1586364061
transform 1 0 32108 0 -1 26656
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 34868 0 -1 26656
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 34316 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 34684 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_359
timestamp 1586364061
transform 1 0 34132 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_363
timestamp 1586364061
transform 1 0 34500 0 -1 26656
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_428
timestamp 1586364061
transform 1 0 37628 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_8  FILLER_44_386
timestamp 1586364061
transform 1 0 36616 0 -1 26656
box -38 -48 774 592
use scs8hd_decap_3  FILLER_44_394
timestamp 1586364061
transform 1 0 37352 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_3  PHY_89
timestamp 1586364061
transform -1 0 38824 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_8  FILLER_44_398
timestamp 1586364061
transform 1 0 37720 0 -1 26656
box -38 -48 774 592
use scs8hd_fill_1  FILLER_44_406
timestamp 1586364061
transform 1 0 38456 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_3  PHY_90
timestamp 1586364061
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_45_3
timestamp 1586364061
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_15
timestamp 1586364061
transform 1 0 2484 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_27
timestamp 1586364061
transform 1 0 3588 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_39
timestamp 1586364061
transform 1 0 4692 0 1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_429
timestamp 1586364061
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use scs8hd_decap_8  FILLER_45_51
timestamp 1586364061
transform 1 0 5796 0 1 26656
box -38 -48 774 592
use scs8hd_fill_2  FILLER_45_59
timestamp 1586364061
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_45_62
timestamp 1586364061
transform 1 0 6808 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_74
timestamp 1586364061
transform 1 0 7912 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_86
timestamp 1586364061
transform 1 0 9016 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_98
timestamp 1586364061
transform 1 0 10120 0 1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_430
timestamp 1586364061
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_45_110
timestamp 1586364061
transform 1 0 11224 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_123
timestamp 1586364061
transform 1 0 12420 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_135
timestamp 1586364061
transform 1 0 13524 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_147
timestamp 1586364061
transform 1 0 14628 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_159
timestamp 1586364061
transform 1 0 15732 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_171
timestamp 1586364061
transform 1 0 16836 0 1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_431
timestamp 1586364061
transform 1 0 17940 0 1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_45_184
timestamp 1586364061
transform 1 0 18032 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_196
timestamp 1586364061
transform 1 0 19136 0 1 26656
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1586364061
transform 1 0 21620 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1586364061
transform 1 0 21252 0 1 26656
box -38 -48 222 592
use scs8hd_decap_8  FILLER_45_208
timestamp 1586364061
transform 1 0 20240 0 1 26656
box -38 -48 774 592
use scs8hd_decap_3  FILLER_45_216
timestamp 1586364061
transform 1 0 20976 0 1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_45_221
timestamp 1586364061
transform 1 0 21436 0 1 26656
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1586364061
transform 1 0 21804 0 1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_432
timestamp 1586364061
transform 1 0 23552 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
timestamp 1586364061
transform 1 0 23092 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_234
timestamp 1586364061
transform 1 0 22632 0 1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_45_238
timestamp 1586364061
transform 1 0 23000 0 1 26656
box -38 -48 130 592
use scs8hd_decap_3  FILLER_45_241
timestamp 1586364061
transform 1 0 23276 0 1 26656
box -38 -48 314 592
use scs8hd_decap_4  FILLER_45_245
timestamp 1586364061
transform 1 0 23644 0 1 26656
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
timestamp 1586364061
transform 1 0 24656 0 1 26656
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
timestamp 1586364061
transform 1 0 24472 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
timestamp 1586364061
transform 1 0 24104 0 1 26656
box -38 -48 222 592
use scs8hd_fill_1  FILLER_45_249
timestamp 1586364061
transform 1 0 24012 0 1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_45_252
timestamp 1586364061
transform 1 0 24288 0 1 26656
box -38 -48 222 592
use scs8hd_or2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
timestamp 1586364061
transform 1 0 27968 0 1 26656
box -38 -48 498 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
timestamp 1586364061
transform 1 0 27784 0 1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_45_275
timestamp 1586364061
transform 1 0 26404 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_45_287
timestamp 1586364061
transform 1 0 27508 0 1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_45_297
timestamp 1586364061
transform 1 0 28428 0 1 26656
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 29256 0 1 26656
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_433
timestamp 1586364061
transform 1 0 29164 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 28980 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
timestamp 1586364061
transform 1 0 28612 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_301
timestamp 1586364061
transform 1 0 28796 0 1 26656
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 31740 0 1 26656
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 31556 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 31188 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_325
timestamp 1586364061
transform 1 0 31004 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_329
timestamp 1586364061
transform 1 0 31372 0 1 26656
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 34960 0 1 26656
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_434
timestamp 1586364061
transform 1 0 34776 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 34592 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 33856 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 34224 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_352
timestamp 1586364061
transform 1 0 33488 0 1 26656
box -38 -48 406 592
use scs8hd_fill_2  FILLER_45_358
timestamp 1586364061
transform 1 0 34040 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_362
timestamp 1586364061
transform 1 0 34408 0 1 26656
box -38 -48 222 592
use scs8hd_fill_1  FILLER_45_367
timestamp 1586364061
transform 1 0 34868 0 1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_45_387
timestamp 1586364061
transform 1 0 36708 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_3  PHY_91
timestamp 1586364061
transform -1 0 38824 0 1 26656
box -38 -48 314 592
use scs8hd_decap_8  FILLER_45_399
timestamp 1586364061
transform 1 0 37812 0 1 26656
box -38 -48 774 592
use scs8hd_decap_3  PHY_92
timestamp 1586364061
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_94
timestamp 1586364061
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use scs8hd_decap_12  FILLER_46_3
timestamp 1586364061
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_15
timestamp 1586364061
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_3
timestamp 1586364061
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_15
timestamp 1586364061
transform 1 0 2484 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_435
timestamp 1586364061
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_46_27
timestamp 1586364061
transform 1 0 3588 0 -1 27744
box -38 -48 406 592
use scs8hd_decap_12  FILLER_46_32
timestamp 1586364061
transform 1 0 4048 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_44
timestamp 1586364061
transform 1 0 5152 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_27
timestamp 1586364061
transform 1 0 3588 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_39
timestamp 1586364061
transform 1 0 4692 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_442
timestamp 1586364061
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_56
timestamp 1586364061
transform 1 0 6256 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_68
timestamp 1586364061
transform 1 0 7360 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_47_51
timestamp 1586364061
transform 1 0 5796 0 1 27744
box -38 -48 774 592
use scs8hd_fill_2  FILLER_47_59
timestamp 1586364061
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_47_62
timestamp 1586364061
transform 1 0 6808 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_74
timestamp 1586364061
transform 1 0 7912 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_436
timestamp 1586364061
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_80
timestamp 1586364061
transform 1 0 8464 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_93
timestamp 1586364061
transform 1 0 9660 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_86
timestamp 1586364061
transform 1 0 9016 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_98
timestamp 1586364061
transform 1 0 10120 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_443
timestamp 1586364061
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_105
timestamp 1586364061
transform 1 0 10764 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_117
timestamp 1586364061
transform 1 0 11868 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_110
timestamp 1586364061
transform 1 0 11224 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_123
timestamp 1586364061
transform 1 0 12420 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_129
timestamp 1586364061
transform 1 0 12972 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_141
timestamp 1586364061
transform 1 0 14076 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_135
timestamp 1586364061
transform 1 0 13524 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_147
timestamp 1586364061
transform 1 0 14628 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_437
timestamp 1586364061
transform 1 0 15180 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_154
timestamp 1586364061
transform 1 0 15272 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_166
timestamp 1586364061
transform 1 0 16376 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_159
timestamp 1586364061
transform 1 0 15732 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_171
timestamp 1586364061
transform 1 0 16836 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_444
timestamp 1586364061
transform 1 0 17940 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_178
timestamp 1586364061
transform 1 0 17480 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_190
timestamp 1586364061
transform 1 0 18584 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_184
timestamp 1586364061
transform 1 0 18032 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_196
timestamp 1586364061
transform 1 0 19136 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_438
timestamp 1586364061
transform 1 0 20792 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_202
timestamp 1586364061
transform 1 0 19688 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_46_215
timestamp 1586364061
transform 1 0 20884 0 -1 27744
box -38 -48 774 592
use scs8hd_fill_2  FILLER_46_223
timestamp 1586364061
transform 1 0 21620 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_47_208
timestamp 1586364061
transform 1 0 20240 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_220
timestamp 1586364061
transform 1 0 21344 0 1 27744
box -38 -48 1142 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
timestamp 1586364061
transform 1 0 23092 0 -1 27744
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_445
timestamp 1586364061
transform 1 0 23552 0 1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1586364061
transform 1 0 21804 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_46_227
timestamp 1586364061
transform 1 0 21988 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_46_243
timestamp 1586364061
transform 1 0 23460 0 -1 27744
box -38 -48 774 592
use scs8hd_decap_12  FILLER_47_232
timestamp 1586364061
transform 1 0 22448 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_245
timestamp 1586364061
transform 1 0 23644 0 1 27744
box -38 -48 1142 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
timestamp 1586364061
transform 1 0 24380 0 -1 27744
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
timestamp 1586364061
transform 1 0 24932 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_251
timestamp 1586364061
transform 1 0 24196 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_257
timestamp 1586364061
transform 1 0 24748 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_46_261
timestamp 1586364061
transform 1 0 25116 0 -1 27744
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_46_273
timestamp 1586364061
transform 1 0 26220 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_47_257
timestamp 1586364061
transform 1 0 24748 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_269
timestamp 1586364061
transform 1 0 25852 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_47_281
timestamp 1586364061
transform 1 0 26956 0 1 27744
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_439
timestamp 1586364061
transform 1 0 26404 0 -1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_297
timestamp 1586364061
transform 1 0 28428 0 1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_47_289
timestamp 1586364061
transform 1 0 27692 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_46_294
timestamp 1586364061
transform 1 0 28152 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_46_288
timestamp 1586364061
transform 1 0 27600 0 -1 27744
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 27968 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 28336 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 27968 0 1 27744
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 28520 0 -1 27744
box -38 -48 866 592
use scs8hd_conb_1  _63_
timestamp 1586364061
transform 1 0 28152 0 1 27744
box -38 -48 314 592
use scs8hd_decap_12  FILLER_46_276
timestamp 1586364061
transform 1 0 26496 0 -1 27744
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_47_301
timestamp 1586364061
transform 1 0 28796 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_307
timestamp 1586364061
transform 1 0 29348 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 28980 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 28612 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 29532 0 -1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_446
timestamp 1586364061
transform 1 0 29164 0 1 27744
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 29256 0 1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_319
timestamp 1586364061
transform 1 0 30452 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_315
timestamp 1586364061
transform 1 0 30084 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_311
timestamp 1586364061
transform 1 0 29716 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 29900 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 30636 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 30268 0 1 27744
box -38 -48 222 592
use scs8hd_conb_1  _59_
timestamp 1586364061
transform 1 0 30084 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_12  FILLER_46_318
timestamp 1586364061
transform 1 0 30360 0 -1 27744
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_47_331
timestamp 1586364061
transform 1 0 31556 0 1 27744
box -38 -48 222 592
use scs8hd_decap_6  FILLER_47_323
timestamp 1586364061
transform 1 0 30820 0 1 27744
box -38 -48 590 592
use scs8hd_decap_4  FILLER_46_330
timestamp 1586364061
transform 1 0 31464 0 -1 27744
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 31372 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_335
timestamp 1586364061
transform 1 0 31924 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 31832 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 31740 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 32108 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_440
timestamp 1586364061
transform 1 0 32016 0 -1 27744
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 32292 0 1 27744
box -38 -48 866 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 32108 0 -1 27744
box -38 -48 866 592
use scs8hd_decap_8  FILLER_46_346
timestamp 1586364061
transform 1 0 32936 0 -1 27744
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 33856 0 -1 27744
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_447
timestamp 1586364061
transform 1 0 34776 0 1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__73__A
timestamp 1586364061
transform 1 0 35236 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_354
timestamp 1586364061
transform 1 0 33672 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_47_348
timestamp 1586364061
transform 1 0 33120 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_47_360
timestamp 1586364061
transform 1 0 34224 0 1 27744
box -38 -48 590 592
use scs8hd_decap_4  FILLER_47_367
timestamp 1586364061
transform 1 0 34868 0 1 27744
box -38 -48 406 592
use scs8hd_decap_4  FILLER_47_381
timestamp 1586364061
transform 1 0 36156 0 1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_47_377
timestamp 1586364061
transform 1 0 35788 0 1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_46_379
timestamp 1586364061
transform 1 0 35972 0 -1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_46_375
timestamp 1586364061
transform 1 0 35604 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 35788 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 35972 0 1 27744
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 35420 0 1 27744
box -38 -48 406 592
use scs8hd_conb_1  _62_
timestamp 1586364061
transform 1 0 36340 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  FILLER_46_394
timestamp 1586364061
transform 1 0 37352 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_8  FILLER_46_386
timestamp 1586364061
transform 1 0 36616 0 -1 27744
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 36524 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_441
timestamp 1586364061
transform 1 0 37628 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_47_387
timestamp 1586364061
transform 1 0 36708 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_3  PHY_93
timestamp 1586364061
transform -1 0 38824 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_95
timestamp 1586364061
transform -1 0 38824 0 1 27744
box -38 -48 314 592
use scs8hd_decap_8  FILLER_46_398
timestamp 1586364061
transform 1 0 37720 0 -1 27744
box -38 -48 774 592
use scs8hd_fill_1  FILLER_46_406
timestamp 1586364061
transform 1 0 38456 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_8  FILLER_47_399
timestamp 1586364061
transform 1 0 37812 0 1 27744
box -38 -48 774 592
use scs8hd_decap_3  PHY_96
timestamp 1586364061
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_48_3
timestamp 1586364061
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_15
timestamp 1586364061
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_448
timestamp 1586364061
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_4  FILLER_48_27
timestamp 1586364061
transform 1 0 3588 0 -1 28832
box -38 -48 406 592
use scs8hd_decap_12  FILLER_48_32
timestamp 1586364061
transform 1 0 4048 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_44
timestamp 1586364061
transform 1 0 5152 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_56
timestamp 1586364061
transform 1 0 6256 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_68
timestamp 1586364061
transform 1 0 7360 0 -1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_449
timestamp 1586364061
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_48_80
timestamp 1586364061
transform 1 0 8464 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_93
timestamp 1586364061
transform 1 0 9660 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_105
timestamp 1586364061
transform 1 0 10764 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_117
timestamp 1586364061
transform 1 0 11868 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_129
timestamp 1586364061
transform 1 0 12972 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_141
timestamp 1586364061
transform 1 0 14076 0 -1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_450
timestamp 1586364061
transform 1 0 15180 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_48_154
timestamp 1586364061
transform 1 0 15272 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_166
timestamp 1586364061
transform 1 0 16376 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_178
timestamp 1586364061
transform 1 0 17480 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_190
timestamp 1586364061
transform 1 0 18584 0 -1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_451
timestamp 1586364061
transform 1 0 20792 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_48_202
timestamp 1586364061
transform 1 0 19688 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_215
timestamp 1586364061
transform 1 0 20884 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_227
timestamp 1586364061
transform 1 0 21988 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_239
timestamp 1586364061
transform 1 0 23092 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_251
timestamp 1586364061
transform 1 0 24196 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_263
timestamp 1586364061
transform 1 0 25300 0 -1 28832
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 27968 0 -1 28832
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_452
timestamp 1586364061
transform 1 0 26404 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 27600 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_48_276
timestamp 1586364061
transform 1 0 26496 0 -1 28832
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_48_290
timestamp 1586364061
transform 1 0 27784 0 -1 28832
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 30452 0 -1 28832
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 29992 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_48_311
timestamp 1586364061
transform 1 0 29716 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_3  FILLER_48_316
timestamp 1586364061
transform 1 0 30176 0 -1 28832
box -38 -48 314 592
use scs8hd_conb_1  _60_
timestamp 1586364061
transform 1 0 32384 0 -1 28832
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_453
timestamp 1586364061
transform 1 0 32016 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_48_323
timestamp 1586364061
transform 1 0 30820 0 -1 28832
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_48_335
timestamp 1586364061
transform 1 0 31924 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_3  FILLER_48_337
timestamp 1586364061
transform 1 0 32108 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_48_343
timestamp 1586364061
transform 1 0 32660 0 -1 28832
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 34868 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 34224 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_355
timestamp 1586364061
transform 1 0 33764 0 -1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_48_359
timestamp 1586364061
transform 1 0 34132 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_4  FILLER_48_362
timestamp 1586364061
transform 1 0 34408 0 -1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_48_366
timestamp 1586364061
transform 1 0 34776 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_4  FILLER_48_369
timestamp 1586364061
transform 1 0 35052 0 -1 28832
box -38 -48 406 592
use scs8hd_buf_2  _73_
timestamp 1586364061
transform 1 0 35420 0 -1 28832
box -38 -48 406 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 36524 0 -1 28832
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_454
timestamp 1586364061
transform 1 0 37628 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__74__A
timestamp 1586364061
transform 1 0 35972 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_377
timestamp 1586364061
transform 1 0 35788 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_381
timestamp 1586364061
transform 1 0 36156 0 -1 28832
box -38 -48 406 592
use scs8hd_decap_8  FILLER_48_389
timestamp 1586364061
transform 1 0 36892 0 -1 28832
box -38 -48 774 592
use scs8hd_decap_3  PHY_97
timestamp 1586364061
transform -1 0 38824 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_8  FILLER_48_398
timestamp 1586364061
transform 1 0 37720 0 -1 28832
box -38 -48 774 592
use scs8hd_fill_1  FILLER_48_406
timestamp 1586364061
transform 1 0 38456 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_3  PHY_98
timestamp 1586364061
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_49_3
timestamp 1586364061
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_15
timestamp 1586364061
transform 1 0 2484 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_27
timestamp 1586364061
transform 1 0 3588 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_39
timestamp 1586364061
transform 1 0 4692 0 1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_455
timestamp 1586364061
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use scs8hd_decap_8  FILLER_49_51
timestamp 1586364061
transform 1 0 5796 0 1 28832
box -38 -48 774 592
use scs8hd_fill_2  FILLER_49_59
timestamp 1586364061
transform 1 0 6532 0 1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_49_62
timestamp 1586364061
transform 1 0 6808 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_74
timestamp 1586364061
transform 1 0 7912 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_86
timestamp 1586364061
transform 1 0 9016 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_98
timestamp 1586364061
transform 1 0 10120 0 1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_456
timestamp 1586364061
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_49_110
timestamp 1586364061
transform 1 0 11224 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_123
timestamp 1586364061
transform 1 0 12420 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_135
timestamp 1586364061
transform 1 0 13524 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_147
timestamp 1586364061
transform 1 0 14628 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_159
timestamp 1586364061
transform 1 0 15732 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_171
timestamp 1586364061
transform 1 0 16836 0 1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_457
timestamp 1586364061
transform 1 0 17940 0 1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_49_184
timestamp 1586364061
transform 1 0 18032 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_196
timestamp 1586364061
transform 1 0 19136 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_208
timestamp 1586364061
transform 1 0 20240 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_220
timestamp 1586364061
transform 1 0 21344 0 1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_458
timestamp 1586364061
transform 1 0 23552 0 1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_49_232
timestamp 1586364061
transform 1 0 22448 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_245
timestamp 1586364061
transform 1 0 23644 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_257
timestamp 1586364061
transform 1 0 24748 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_269
timestamp 1586364061
transform 1 0 25852 0 1 28832
box -38 -48 1142 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 27600 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 27416 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_281
timestamp 1586364061
transform 1 0 26956 0 1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_49_285
timestamp 1586364061
transform 1 0 27324 0 1 28832
box -38 -48 130 592
use scs8hd_fill_2  FILLER_49_297
timestamp 1586364061
transform 1 0 28428 0 1 28832
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1586364061
transform 1 0 29992 0 1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_459
timestamp 1586364061
transform 1 0 29164 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 28612 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 29808 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 29440 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 28980 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_301
timestamp 1586364061
transform 1 0 28796 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_306
timestamp 1586364061
transform 1 0 29256 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_310
timestamp 1586364061
transform 1 0 29624 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
timestamp 1586364061
transform 1 0 31004 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
timestamp 1586364061
transform 1 0 31372 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 32108 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_323
timestamp 1586364061
transform 1 0 30820 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_327
timestamp 1586364061
transform 1 0 31188 0 1 28832
box -38 -48 222 592
use scs8hd_decap_6  FILLER_49_331
timestamp 1586364061
transform 1 0 31556 0 1 28832
box -38 -48 590 592
use scs8hd_decap_12  FILLER_49_339
timestamp 1586364061
transform 1 0 32292 0 1 28832
box -38 -48 1142 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 33672 0 1 28832
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 34868 0 1 28832
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_460
timestamp 1586364061
transform 1 0 34776 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 34592 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 34224 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 33488 0 1 28832
box -38 -48 222 592
use scs8hd_fill_1  FILLER_49_351
timestamp 1586364061
transform 1 0 33396 0 1 28832
box -38 -48 130 592
use scs8hd_fill_2  FILLER_49_358
timestamp 1586364061
transform 1 0 34040 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_362
timestamp 1586364061
transform 1 0 34408 0 1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_49_386
timestamp 1586364061
transform 1 0 36616 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_3  PHY_99
timestamp 1586364061
transform -1 0 38824 0 1 28832
box -38 -48 314 592
use scs8hd_decap_8  FILLER_49_398
timestamp 1586364061
transform 1 0 37720 0 1 28832
box -38 -48 774 592
use scs8hd_fill_1  FILLER_49_406
timestamp 1586364061
transform 1 0 38456 0 1 28832
box -38 -48 130 592
use scs8hd_decap_3  PHY_100
timestamp 1586364061
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_50_3
timestamp 1586364061
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_15
timestamp 1586364061
transform 1 0 2484 0 -1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_461
timestamp 1586364061
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_4  FILLER_50_27
timestamp 1586364061
transform 1 0 3588 0 -1 29920
box -38 -48 406 592
use scs8hd_decap_12  FILLER_50_32
timestamp 1586364061
transform 1 0 4048 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_44
timestamp 1586364061
transform 1 0 5152 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_56
timestamp 1586364061
transform 1 0 6256 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_68
timestamp 1586364061
transform 1 0 7360 0 -1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_462
timestamp 1586364061
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_50_80
timestamp 1586364061
transform 1 0 8464 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_93
timestamp 1586364061
transform 1 0 9660 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_105
timestamp 1586364061
transform 1 0 10764 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_117
timestamp 1586364061
transform 1 0 11868 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_129
timestamp 1586364061
transform 1 0 12972 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_141
timestamp 1586364061
transform 1 0 14076 0 -1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_463
timestamp 1586364061
transform 1 0 15180 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_50_154
timestamp 1586364061
transform 1 0 15272 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_166
timestamp 1586364061
transform 1 0 16376 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_178
timestamp 1586364061
transform 1 0 17480 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_190
timestamp 1586364061
transform 1 0 18584 0 -1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_464
timestamp 1586364061
transform 1 0 20792 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_50_202
timestamp 1586364061
transform 1 0 19688 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_215
timestamp 1586364061
transform 1 0 20884 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_227
timestamp 1586364061
transform 1 0 21988 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_239
timestamp 1586364061
transform 1 0 23092 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_251
timestamp 1586364061
transform 1 0 24196 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_263
timestamp 1586364061
transform 1 0 25300 0 -1 29920
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 28152 0 -1 29920
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_465
timestamp 1586364061
transform 1 0 26404 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 27600 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_50_276
timestamp 1586364061
transform 1 0 26496 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_50_290
timestamp 1586364061
transform 1 0 27784 0 -1 29920
box -38 -48 406 592
use scs8hd_or2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
timestamp 1586364061
transform 1 0 30636 0 -1 29920
box -38 -48 498 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
timestamp 1586364061
transform 1 0 30084 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_313
timestamp 1586364061
transform 1 0 29900 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_50_317
timestamp 1586364061
transform 1 0 30268 0 -1 29920
box -38 -48 406 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 32108 0 -1 29920
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_466
timestamp 1586364061
transform 1 0 32016 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_8  FILLER_50_326
timestamp 1586364061
transform 1 0 31096 0 -1 29920
box -38 -48 774 592
use scs8hd_fill_2  FILLER_50_334
timestamp 1586364061
transform 1 0 31832 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_8  FILLER_50_341
timestamp 1586364061
transform 1 0 32476 0 -1 29920
box -38 -48 774 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1586364061
transform 1 0 34224 0 -1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 35236 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 33212 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 34040 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 33580 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_351
timestamp 1586364061
transform 1 0 33396 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_3  FILLER_50_355
timestamp 1586364061
transform 1 0 33764 0 -1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_50_369
timestamp 1586364061
transform 1 0 35052 0 -1 29920
box -38 -48 222 592
use scs8hd_buf_2  _74_
timestamp 1586364061
transform 1 0 35788 0 -1 29920
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_467
timestamp 1586364061
transform 1 0 37628 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 35604 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_373
timestamp 1586364061
transform 1 0 35420 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_50_381
timestamp 1586364061
transform 1 0 36156 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_50_393
timestamp 1586364061
transform 1 0 37260 0 -1 29920
box -38 -48 406 592
use scs8hd_decap_3  PHY_101
timestamp 1586364061
transform -1 0 38824 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_8  FILLER_50_398
timestamp 1586364061
transform 1 0 37720 0 -1 29920
box -38 -48 774 592
use scs8hd_fill_1  FILLER_50_406
timestamp 1586364061
transform 1 0 38456 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_3  PHY_102
timestamp 1586364061
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_51_3
timestamp 1586364061
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_15
timestamp 1586364061
transform 1 0 2484 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_27
timestamp 1586364061
transform 1 0 3588 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_39
timestamp 1586364061
transform 1 0 4692 0 1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_468
timestamp 1586364061
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use scs8hd_decap_8  FILLER_51_51
timestamp 1586364061
transform 1 0 5796 0 1 29920
box -38 -48 774 592
use scs8hd_fill_2  FILLER_51_59
timestamp 1586364061
transform 1 0 6532 0 1 29920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_51_62
timestamp 1586364061
transform 1 0 6808 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_74
timestamp 1586364061
transform 1 0 7912 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_86
timestamp 1586364061
transform 1 0 9016 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_98
timestamp 1586364061
transform 1 0 10120 0 1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_469
timestamp 1586364061
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_51_110
timestamp 1586364061
transform 1 0 11224 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_123
timestamp 1586364061
transform 1 0 12420 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_135
timestamp 1586364061
transform 1 0 13524 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_147
timestamp 1586364061
transform 1 0 14628 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_159
timestamp 1586364061
transform 1 0 15732 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_171
timestamp 1586364061
transform 1 0 16836 0 1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_470
timestamp 1586364061
transform 1 0 17940 0 1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_51_184
timestamp 1586364061
transform 1 0 18032 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_196
timestamp 1586364061
transform 1 0 19136 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_208
timestamp 1586364061
transform 1 0 20240 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_220
timestamp 1586364061
transform 1 0 21344 0 1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_471
timestamp 1586364061
transform 1 0 23552 0 1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_51_232
timestamp 1586364061
transform 1 0 22448 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_245
timestamp 1586364061
transform 1 0 23644 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_257
timestamp 1586364061
transform 1 0 24748 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_269
timestamp 1586364061
transform 1 0 25852 0 1 29920
box -38 -48 1142 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 28060 0 1 29920
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 27876 0 1 29920
box -38 -48 222 592
use scs8hd_decap_8  FILLER_51_281
timestamp 1586364061
transform 1 0 26956 0 1 29920
box -38 -48 774 592
use scs8hd_fill_2  FILLER_51_289
timestamp 1586364061
transform 1 0 27692 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_297
timestamp 1586364061
transform 1 0 28428 0 1 29920
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 29348 0 1 29920
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_472
timestamp 1586364061
transform 1 0 29164 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 28980 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
timestamp 1586364061
transform 1 0 28612 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_301
timestamp 1586364061
transform 1 0 28796 0 1 29920
box -38 -48 222 592
use scs8hd_fill_1  FILLER_51_306
timestamp 1586364061
transform 1 0 29256 0 1 29920
box -38 -48 130 592
use scs8hd_decap_4  FILLER_51_326
timestamp 1586364061
transform 1 0 31096 0 1 29920
box -38 -48 406 592
use scs8hd_fill_1  FILLER_51_330
timestamp 1586364061
transform 1 0 31464 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 31556 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_333
timestamp 1586364061
transform 1 0 31740 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 31924 0 1 29920
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 32108 0 1 29920
box -38 -48 406 592
use scs8hd_fill_2  FILLER_51_341
timestamp 1586364061
transform 1 0 32476 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_345
timestamp 1586364061
transform 1 0 32844 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 33028 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 32660 0 1 29920
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1586364061
transform 1 0 33212 0 1 29920
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 34868 0 1 29920
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_473
timestamp 1586364061
transform 1 0 34776 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 34408 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_358
timestamp 1586364061
transform 1 0 34040 0 1 29920
box -38 -48 406 592
use scs8hd_fill_2  FILLER_51_364
timestamp 1586364061
transform 1 0 34592 0 1 29920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_51_386
timestamp 1586364061
transform 1 0 36616 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_3  PHY_103
timestamp 1586364061
transform -1 0 38824 0 1 29920
box -38 -48 314 592
use scs8hd_decap_8  FILLER_51_398
timestamp 1586364061
transform 1 0 37720 0 1 29920
box -38 -48 774 592
use scs8hd_fill_1  FILLER_51_406
timestamp 1586364061
transform 1 0 38456 0 1 29920
box -38 -48 130 592
use scs8hd_decap_3  PHY_104
timestamp 1586364061
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_106
timestamp 1586364061
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use scs8hd_decap_12  FILLER_52_3
timestamp 1586364061
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_15
timestamp 1586364061
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_3
timestamp 1586364061
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_15
timestamp 1586364061
transform 1 0 2484 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_474
timestamp 1586364061
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_52_27
timestamp 1586364061
transform 1 0 3588 0 -1 31008
box -38 -48 406 592
use scs8hd_decap_12  FILLER_52_32
timestamp 1586364061
transform 1 0 4048 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_44
timestamp 1586364061
transform 1 0 5152 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_27
timestamp 1586364061
transform 1 0 3588 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_39
timestamp 1586364061
transform 1 0 4692 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_481
timestamp 1586364061
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_56
timestamp 1586364061
transform 1 0 6256 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_68
timestamp 1586364061
transform 1 0 7360 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_53_51
timestamp 1586364061
transform 1 0 5796 0 1 31008
box -38 -48 774 592
use scs8hd_fill_2  FILLER_53_59
timestamp 1586364061
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_53_62
timestamp 1586364061
transform 1 0 6808 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_74
timestamp 1586364061
transform 1 0 7912 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_475
timestamp 1586364061
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_80
timestamp 1586364061
transform 1 0 8464 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_93
timestamp 1586364061
transform 1 0 9660 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_86
timestamp 1586364061
transform 1 0 9016 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_98
timestamp 1586364061
transform 1 0 10120 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_482
timestamp 1586364061
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_105
timestamp 1586364061
transform 1 0 10764 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_117
timestamp 1586364061
transform 1 0 11868 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_110
timestamp 1586364061
transform 1 0 11224 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_123
timestamp 1586364061
transform 1 0 12420 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_129
timestamp 1586364061
transform 1 0 12972 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_141
timestamp 1586364061
transform 1 0 14076 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_135
timestamp 1586364061
transform 1 0 13524 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_147
timestamp 1586364061
transform 1 0 14628 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_476
timestamp 1586364061
transform 1 0 15180 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_154
timestamp 1586364061
transform 1 0 15272 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_166
timestamp 1586364061
transform 1 0 16376 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_159
timestamp 1586364061
transform 1 0 15732 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_171
timestamp 1586364061
transform 1 0 16836 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_483
timestamp 1586364061
transform 1 0 17940 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_178
timestamp 1586364061
transform 1 0 17480 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_190
timestamp 1586364061
transform 1 0 18584 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_184
timestamp 1586364061
transform 1 0 18032 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_196
timestamp 1586364061
transform 1 0 19136 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_477
timestamp 1586364061
transform 1 0 20792 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_202
timestamp 1586364061
transform 1 0 19688 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_215
timestamp 1586364061
transform 1 0 20884 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_208
timestamp 1586364061
transform 1 0 20240 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_220
timestamp 1586364061
transform 1 0 21344 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_484
timestamp 1586364061
transform 1 0 23552 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_227
timestamp 1586364061
transform 1 0 21988 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_239
timestamp 1586364061
transform 1 0 23092 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_232
timestamp 1586364061
transform 1 0 22448 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_245
timestamp 1586364061
transform 1 0 23644 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_251
timestamp 1586364061
transform 1 0 24196 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_263
timestamp 1586364061
transform 1 0 25300 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_257
timestamp 1586364061
transform 1 0 24748 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_269
timestamp 1586364061
transform 1 0 25852 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_478
timestamp 1586364061
transform 1 0 26404 0 -1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 28520 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 28152 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_276
timestamp 1586364061
transform 1 0 26496 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_288
timestamp 1586364061
transform 1 0 27600 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_281
timestamp 1586364061
transform 1 0 26956 0 1 31008
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_53_293
timestamp 1586364061
transform 1 0 28060 0 1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_53_296
timestamp 1586364061
transform 1 0 28336 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
timestamp 1586364061
transform 1 0 28888 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_300
timestamp 1586364061
transform 1 0 28704 0 1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_53_304
timestamp 1586364061
transform 1 0 29072 0 1 31008
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_485
timestamp 1586364061
transform 1 0 29164 0 1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 29348 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1586364061
transform 1 0 29440 0 1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_52_306
timestamp 1586364061
transform 1 0 29256 0 -1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_53_306
timestamp 1586364061
transform 1 0 29256 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_310
timestamp 1586364061
transform 1 0 29624 0 1 31008
box -38 -48 222 592
use scs8hd_decap_6  FILLER_52_300
timestamp 1586364061
transform 1 0 28704 0 -1 31008
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1586364061
transform 1 0 29808 0 1 31008
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1586364061
transform 1 0 29992 0 1 31008
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
timestamp 1586364061
transform 1 0 29532 0 -1 31008
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_53_327
timestamp 1586364061
transform 1 0 31188 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_323
timestamp 1586364061
transform 1 0 30820 0 1 31008
box -38 -48 222 592
use scs8hd_decap_3  FILLER_52_328
timestamp 1586364061
transform 1 0 31280 0 -1 31008
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 31004 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 31556 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 31372 0 1 31008
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1586364061
transform 1 0 31556 0 1 31008
box -38 -48 866 592
use scs8hd_decap_4  FILLER_53_340
timestamp 1586364061
transform 1 0 32384 0 1 31008
box -38 -48 406 592
use scs8hd_fill_1  FILLER_52_337
timestamp 1586364061
transform 1 0 32108 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_3  FILLER_52_333
timestamp 1586364061
transform 1 0 31740 0 -1 31008
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_479
timestamp 1586364061
transform 1 0 32016 0 -1 31008
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1586364061
transform 1 0 32200 0 -1 31008
box -38 -48 866 592
use scs8hd_decap_4  FILLER_53_347
timestamp 1586364061
transform 1 0 33028 0 1 31008
box -38 -48 406 592
use scs8hd_fill_1  FILLER_53_344
timestamp 1586364061
transform 1 0 32752 0 1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_52_347
timestamp 1586364061
transform 1 0 33028 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
timestamp 1586364061
transform 1 0 32844 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 33488 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 33212 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_53_351
timestamp 1586364061
transform 1 0 33396 0 1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 34224 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 34224 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 33856 0 1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_52_359
timestamp 1586364061
transform 1 0 34132 0 -1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_53_354
timestamp 1586364061
transform 1 0 33672 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_358
timestamp 1586364061
transform 1 0 34040 0 1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_52_351
timestamp 1586364061
transform 1 0 33396 0 -1 31008
box -38 -48 774 592
use scs8hd_fill_2  FILLER_53_362
timestamp 1586364061
transform 1 0 34408 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 34592 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_486
timestamp 1586364061
transform 1 0 34776 0 1 31008
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 34868 0 1 31008
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 34408 0 -1 31008
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_480
timestamp 1586364061
transform 1 0 37628 0 -1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__75__A
timestamp 1586364061
transform 1 0 36800 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_381
timestamp 1586364061
transform 1 0 36156 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_52_393
timestamp 1586364061
transform 1 0 37260 0 -1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_386
timestamp 1586364061
transform 1 0 36616 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_53_390
timestamp 1586364061
transform 1 0 36984 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_3  PHY_105
timestamp 1586364061
transform -1 0 38824 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_107
timestamp 1586364061
transform -1 0 38824 0 1 31008
box -38 -48 314 592
use scs8hd_decap_8  FILLER_52_398
timestamp 1586364061
transform 1 0 37720 0 -1 31008
box -38 -48 774 592
use scs8hd_fill_1  FILLER_52_406
timestamp 1586364061
transform 1 0 38456 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_53_402
timestamp 1586364061
transform 1 0 38088 0 1 31008
box -38 -48 406 592
use scs8hd_fill_1  FILLER_53_406
timestamp 1586364061
transform 1 0 38456 0 1 31008
box -38 -48 130 592
use scs8hd_decap_3  PHY_108
timestamp 1586364061
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_54_3
timestamp 1586364061
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_15
timestamp 1586364061
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_487
timestamp 1586364061
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_4  FILLER_54_27
timestamp 1586364061
transform 1 0 3588 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_12  FILLER_54_32
timestamp 1586364061
transform 1 0 4048 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_44
timestamp 1586364061
transform 1 0 5152 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_56
timestamp 1586364061
transform 1 0 6256 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_68
timestamp 1586364061
transform 1 0 7360 0 -1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_488
timestamp 1586364061
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_54_80
timestamp 1586364061
transform 1 0 8464 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_93
timestamp 1586364061
transform 1 0 9660 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_105
timestamp 1586364061
transform 1 0 10764 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_117
timestamp 1586364061
transform 1 0 11868 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_129
timestamp 1586364061
transform 1 0 12972 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_141
timestamp 1586364061
transform 1 0 14076 0 -1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_489
timestamp 1586364061
transform 1 0 15180 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_54_154
timestamp 1586364061
transform 1 0 15272 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_166
timestamp 1586364061
transform 1 0 16376 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_178
timestamp 1586364061
transform 1 0 17480 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_190
timestamp 1586364061
transform 1 0 18584 0 -1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_490
timestamp 1586364061
transform 1 0 20792 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_54_202
timestamp 1586364061
transform 1 0 19688 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_215
timestamp 1586364061
transform 1 0 20884 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_227
timestamp 1586364061
transform 1 0 21988 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_239
timestamp 1586364061
transform 1 0 23092 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_251
timestamp 1586364061
transform 1 0 24196 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_263
timestamp 1586364061
transform 1 0 25300 0 -1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_491
timestamp 1586364061
transform 1 0 26404 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_54_276
timestamp 1586364061
transform 1 0 26496 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_288
timestamp 1586364061
transform 1 0 27600 0 -1 32096
box -38 -48 1142 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1586364061
transform 1 0 29992 0 -1 32096
box -38 -48 866 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
timestamp 1586364061
transform 1 0 28888 0 -1 32096
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
timestamp 1586364061
transform 1 0 29532 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_300
timestamp 1586364061
transform 1 0 28704 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_54_306
timestamp 1586364061
transform 1 0 29256 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_3  FILLER_54_311
timestamp 1586364061
transform 1 0 29716 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_4  FILLER_54_327
timestamp 1586364061
transform 1 0 31188 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_2  FILLER_54_323
timestamp 1586364061
transform 1 0 30820 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1586364061
transform 1 0 31004 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 31556 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_337
timestamp 1586364061
transform 1 0 32108 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_54_333
timestamp 1586364061
transform 1 0 31740 0 -1 32096
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_492
timestamp 1586364061
transform 1 0 32016 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_4  FILLER_54_341
timestamp 1586364061
transform 1 0 32476 0 -1 32096
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1586364061
transform 1 0 32292 0 -1 32096
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
timestamp 1586364061
transform 1 0 32844 0 -1 32096
box -38 -48 406 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1586364061
transform 1 0 34224 0 -1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
timestamp 1586364061
transform 1 0 35236 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 34040 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 33396 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_349
timestamp 1586364061
transform 1 0 33212 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_353
timestamp 1586364061
transform 1 0 33580 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_1  FILLER_54_357
timestamp 1586364061
transform 1 0 33948 0 -1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_54_369
timestamp 1586364061
transform 1 0 35052 0 -1 32096
box -38 -48 222 592
use scs8hd_buf_2  _75_
timestamp 1586364061
transform 1 0 35788 0 -1 32096
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_493
timestamp 1586364061
transform 1 0 37628 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_4  FILLER_54_373
timestamp 1586364061
transform 1 0 35420 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_12  FILLER_54_381
timestamp 1586364061
transform 1 0 36156 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_54_393
timestamp 1586364061
transform 1 0 37260 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_3  PHY_109
timestamp 1586364061
transform -1 0 38824 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_8  FILLER_54_398
timestamp 1586364061
transform 1 0 37720 0 -1 32096
box -38 -48 774 592
use scs8hd_fill_1  FILLER_54_406
timestamp 1586364061
transform 1 0 38456 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_3  PHY_110
timestamp 1586364061
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_55_3
timestamp 1586364061
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_15
timestamp 1586364061
transform 1 0 2484 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_27
timestamp 1586364061
transform 1 0 3588 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_39
timestamp 1586364061
transform 1 0 4692 0 1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_494
timestamp 1586364061
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use scs8hd_decap_8  FILLER_55_51
timestamp 1586364061
transform 1 0 5796 0 1 32096
box -38 -48 774 592
use scs8hd_fill_2  FILLER_55_59
timestamp 1586364061
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_55_62
timestamp 1586364061
transform 1 0 6808 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_74
timestamp 1586364061
transform 1 0 7912 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_86
timestamp 1586364061
transform 1 0 9016 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_98
timestamp 1586364061
transform 1 0 10120 0 1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_495
timestamp 1586364061
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_55_110
timestamp 1586364061
transform 1 0 11224 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_123
timestamp 1586364061
transform 1 0 12420 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_135
timestamp 1586364061
transform 1 0 13524 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_147
timestamp 1586364061
transform 1 0 14628 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_159
timestamp 1586364061
transform 1 0 15732 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_171
timestamp 1586364061
transform 1 0 16836 0 1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_496
timestamp 1586364061
transform 1 0 17940 0 1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_55_184
timestamp 1586364061
transform 1 0 18032 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_196
timestamp 1586364061
transform 1 0 19136 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_208
timestamp 1586364061
transform 1 0 20240 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_220
timestamp 1586364061
transform 1 0 21344 0 1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_497
timestamp 1586364061
transform 1 0 23552 0 1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_55_232
timestamp 1586364061
transform 1 0 22448 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_245
timestamp 1586364061
transform 1 0 23644 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_257
timestamp 1586364061
transform 1 0 24748 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_269
timestamp 1586364061
transform 1 0 25852 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_281
timestamp 1586364061
transform 1 0 26956 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_55_293
timestamp 1586364061
transform 1 0 28060 0 1 32096
box -38 -48 590 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
timestamp 1586364061
transform 1 0 29624 0 1 32096
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_498
timestamp 1586364061
transform 1 0 29164 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
timestamp 1586364061
transform 1 0 29440 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
timestamp 1586364061
transform 1 0 28980 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
timestamp 1586364061
transform 1 0 28612 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_301
timestamp 1586364061
transform 1 0 28796 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_306
timestamp 1586364061
transform 1 0 29256 0 1 32096
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
timestamp 1586364061
transform 1 0 32108 0 1 32096
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1586364061
transform 1 0 32660 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1586364061
transform 1 0 31924 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
timestamp 1586364061
transform 1 0 31556 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 33028 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_329
timestamp 1586364061
transform 1 0 31372 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_333
timestamp 1586364061
transform 1 0 31740 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_341
timestamp 1586364061
transform 1 0 32476 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_345
timestamp 1586364061
transform 1 0 32844 0 1 32096
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1586364061
transform 1 0 33212 0 1 32096
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
timestamp 1586364061
transform 1 0 34868 0 1 32096
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_499
timestamp 1586364061
transform 1 0 34776 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
timestamp 1586364061
transform 1 0 34592 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
timestamp 1586364061
transform 1 0 34224 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_358
timestamp 1586364061
transform 1 0 34040 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_362
timestamp 1586364061
transform 1 0 34408 0 1 32096
box -38 -48 222 592
use scs8hd_buf_2  _76_
timestamp 1586364061
transform 1 0 37352 0 1 32096
box -38 -48 406 592
use scs8hd_decap_8  FILLER_55_386
timestamp 1586364061
transform 1 0 36616 0 1 32096
box -38 -48 774 592
use scs8hd_decap_3  PHY_111
timestamp 1586364061
transform -1 0 38824 0 1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__76__A
timestamp 1586364061
transform 1 0 37904 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_398
timestamp 1586364061
transform 1 0 37720 0 1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_55_402
timestamp 1586364061
transform 1 0 38088 0 1 32096
box -38 -48 406 592
use scs8hd_fill_1  FILLER_55_406
timestamp 1586364061
transform 1 0 38456 0 1 32096
box -38 -48 130 592
use scs8hd_decap_3  PHY_112
timestamp 1586364061
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_56_3
timestamp 1586364061
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_15
timestamp 1586364061
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_500
timestamp 1586364061
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_4  FILLER_56_27
timestamp 1586364061
transform 1 0 3588 0 -1 33184
box -38 -48 406 592
use scs8hd_decap_12  FILLER_56_32
timestamp 1586364061
transform 1 0 4048 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_44
timestamp 1586364061
transform 1 0 5152 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_56
timestamp 1586364061
transform 1 0 6256 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_68
timestamp 1586364061
transform 1 0 7360 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_501
timestamp 1586364061
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_56_80
timestamp 1586364061
transform 1 0 8464 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_93
timestamp 1586364061
transform 1 0 9660 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_105
timestamp 1586364061
transform 1 0 10764 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_117
timestamp 1586364061
transform 1 0 11868 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_129
timestamp 1586364061
transform 1 0 12972 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_141
timestamp 1586364061
transform 1 0 14076 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_502
timestamp 1586364061
transform 1 0 15180 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_56_154
timestamp 1586364061
transform 1 0 15272 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_166
timestamp 1586364061
transform 1 0 16376 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_178
timestamp 1586364061
transform 1 0 17480 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_190
timestamp 1586364061
transform 1 0 18584 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_503
timestamp 1586364061
transform 1 0 20792 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_56_202
timestamp 1586364061
transform 1 0 19688 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_215
timestamp 1586364061
transform 1 0 20884 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_227
timestamp 1586364061
transform 1 0 21988 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_239
timestamp 1586364061
transform 1 0 23092 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_251
timestamp 1586364061
transform 1 0 24196 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_263
timestamp 1586364061
transform 1 0 25300 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_504
timestamp 1586364061
transform 1 0 26404 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1586364061
transform 1 0 27968 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_12  FILLER_56_276
timestamp 1586364061
transform 1 0 26496 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_56_288
timestamp 1586364061
transform 1 0 27600 0 -1 33184
box -38 -48 406 592
use scs8hd_decap_12  FILLER_56_294
timestamp 1586364061
transform 1 0 28152 0 -1 33184
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
timestamp 1586364061
transform 1 0 29532 0 -1 33184
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
timestamp 1586364061
transform 1 0 29348 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_1  FILLER_56_306
timestamp 1586364061
transform 1 0 29256 0 -1 33184
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1586364061
transform 1 0 32108 0 -1 33184
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_505
timestamp 1586364061
transform 1 0 32016 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 31832 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_6  FILLER_56_328
timestamp 1586364061
transform 1 0 31280 0 -1 33184
box -38 -48 590 592
use scs8hd_decap_3  FILLER_56_346
timestamp 1586364061
transform 1 0 32936 0 -1 33184
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
timestamp 1586364061
transform 1 0 34684 0 -1 33184
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
timestamp 1586364061
transform 1 0 34500 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
timestamp 1586364061
transform 1 0 34132 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 33212 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_8  FILLER_56_351
timestamp 1586364061
transform 1 0 33396 0 -1 33184
box -38 -48 774 592
use scs8hd_fill_2  FILLER_56_361
timestamp 1586364061
transform 1 0 34316 0 -1 33184
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_506
timestamp 1586364061
transform 1 0 37628 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_56_384
timestamp 1586364061
transform 1 0 36432 0 -1 33184
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_56_396
timestamp 1586364061
transform 1 0 37536 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_3  PHY_113
timestamp 1586364061
transform -1 0 38824 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_8  FILLER_56_398
timestamp 1586364061
transform 1 0 37720 0 -1 33184
box -38 -48 774 592
use scs8hd_fill_1  FILLER_56_406
timestamp 1586364061
transform 1 0 38456 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_3  PHY_114
timestamp 1586364061
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_57_3
timestamp 1586364061
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_15
timestamp 1586364061
transform 1 0 2484 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_27
timestamp 1586364061
transform 1 0 3588 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_39
timestamp 1586364061
transform 1 0 4692 0 1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_507
timestamp 1586364061
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use scs8hd_decap_8  FILLER_57_51
timestamp 1586364061
transform 1 0 5796 0 1 33184
box -38 -48 774 592
use scs8hd_fill_2  FILLER_57_59
timestamp 1586364061
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use scs8hd_decap_12  FILLER_57_62
timestamp 1586364061
transform 1 0 6808 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_74
timestamp 1586364061
transform 1 0 7912 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_86
timestamp 1586364061
transform 1 0 9016 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_98
timestamp 1586364061
transform 1 0 10120 0 1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_508
timestamp 1586364061
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_57_110
timestamp 1586364061
transform 1 0 11224 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_123
timestamp 1586364061
transform 1 0 12420 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_135
timestamp 1586364061
transform 1 0 13524 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_147
timestamp 1586364061
transform 1 0 14628 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_159
timestamp 1586364061
transform 1 0 15732 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_171
timestamp 1586364061
transform 1 0 16836 0 1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_509
timestamp 1586364061
transform 1 0 17940 0 1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_57_184
timestamp 1586364061
transform 1 0 18032 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_196
timestamp 1586364061
transform 1 0 19136 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_208
timestamp 1586364061
transform 1 0 20240 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_220
timestamp 1586364061
transform 1 0 21344 0 1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_510
timestamp 1586364061
transform 1 0 23552 0 1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_57_232
timestamp 1586364061
transform 1 0 22448 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_245
timestamp 1586364061
transform 1 0 23644 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_257
timestamp 1586364061
transform 1 0 24748 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_269
timestamp 1586364061
transform 1 0 25852 0 1 33184
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1586364061
transform 1 0 27968 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1586364061
transform 1 0 27600 0 1 33184
box -38 -48 222 592
use scs8hd_decap_6  FILLER_57_281
timestamp 1586364061
transform 1 0 26956 0 1 33184
box -38 -48 590 592
use scs8hd_fill_1  FILLER_57_287
timestamp 1586364061
transform 1 0 27508 0 1 33184
box -38 -48 130 592
use scs8hd_fill_2  FILLER_57_290
timestamp 1586364061
transform 1 0 27784 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_294
timestamp 1586364061
transform 1 0 28152 0 1 33184
box -38 -48 406 592
use scs8hd_fill_1  FILLER_57_298
timestamp 1586364061
transform 1 0 28520 0 1 33184
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
timestamp 1586364061
transform 1 0 29624 0 1 33184
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_511
timestamp 1586364061
transform 1 0 29164 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
timestamp 1586364061
transform 1 0 29440 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
timestamp 1586364061
transform 1 0 28980 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
timestamp 1586364061
transform 1 0 28612 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_301
timestamp 1586364061
transform 1 0 28796 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_306
timestamp 1586364061
transform 1 0 29256 0 1 33184
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1586364061
transform 1 0 32108 0 1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
timestamp 1586364061
transform 1 0 31924 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
timestamp 1586364061
transform 1 0 31556 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_329
timestamp 1586364061
transform 1 0 31372 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_333
timestamp 1586364061
transform 1 0 31740 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_346
timestamp 1586364061
transform 1 0 32936 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_358
timestamp 1586364061
transform 1 0 34040 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_350
timestamp 1586364061
transform 1 0 33304 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 33120 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__77__A
timestamp 1586364061
transform 1 0 33488 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
timestamp 1586364061
transform 1 0 34224 0 1 33184
box -38 -48 222 592
use scs8hd_buf_2  _77_
timestamp 1586364061
transform 1 0 33672 0 1 33184
box -38 -48 406 592
use scs8hd_fill_2  FILLER_57_362
timestamp 1586364061
transform 1 0 34408 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
timestamp 1586364061
transform 1 0 34592 0 1 33184
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_512
timestamp 1586364061
transform 1 0 34776 0 1 33184
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
timestamp 1586364061
transform 1 0 34868 0 1 33184
box -38 -48 1786 592
use scs8hd_decap_12  FILLER_57_386
timestamp 1586364061
transform 1 0 36616 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_3  PHY_115
timestamp 1586364061
transform -1 0 38824 0 1 33184
box -38 -48 314 592
use scs8hd_decap_8  FILLER_57_398
timestamp 1586364061
transform 1 0 37720 0 1 33184
box -38 -48 774 592
use scs8hd_fill_1  FILLER_57_406
timestamp 1586364061
transform 1 0 38456 0 1 33184
box -38 -48 130 592
use scs8hd_decap_3  PHY_116
timestamp 1586364061
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_58_3
timestamp 1586364061
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_15
timestamp 1586364061
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_513
timestamp 1586364061
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_4  FILLER_58_27
timestamp 1586364061
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_12  FILLER_58_32
timestamp 1586364061
transform 1 0 4048 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_44
timestamp 1586364061
transform 1 0 5152 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_56
timestamp 1586364061
transform 1 0 6256 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_68
timestamp 1586364061
transform 1 0 7360 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_514
timestamp 1586364061
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_58_80
timestamp 1586364061
transform 1 0 8464 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_93
timestamp 1586364061
transform 1 0 9660 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_105
timestamp 1586364061
transform 1 0 10764 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_117
timestamp 1586364061
transform 1 0 11868 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_129
timestamp 1586364061
transform 1 0 12972 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_141
timestamp 1586364061
transform 1 0 14076 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_515
timestamp 1586364061
transform 1 0 15180 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_58_154
timestamp 1586364061
transform 1 0 15272 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_166
timestamp 1586364061
transform 1 0 16376 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_178
timestamp 1586364061
transform 1 0 17480 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_190
timestamp 1586364061
transform 1 0 18584 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_516
timestamp 1586364061
transform 1 0 20792 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_58_202
timestamp 1586364061
transform 1 0 19688 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_215
timestamp 1586364061
transform 1 0 20884 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_227
timestamp 1586364061
transform 1 0 21988 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_239
timestamp 1586364061
transform 1 0 23092 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_251
timestamp 1586364061
transform 1 0 24196 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_263
timestamp 1586364061
transform 1 0 25300 0 -1 34272
box -38 -48 1142 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1586364061
transform 1 0 27968 0 -1 34272
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_517
timestamp 1586364061
transform 1 0 26404 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_58_276
timestamp 1586364061
transform 1 0 26496 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_58_288
timestamp 1586364061
transform 1 0 27600 0 -1 34272
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
timestamp 1586364061
transform 1 0 29532 0 -1 34272
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_58_301
timestamp 1586364061
transform 1 0 28796 0 -1 34272
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
timestamp 1586364061
transform 1 0 32108 0 -1 34272
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_518
timestamp 1586364061
transform 1 0 32016 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 31832 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_6  FILLER_58_328
timestamp 1586364061
transform 1 0 31280 0 -1 34272
box -38 -48 590 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
timestamp 1586364061
transform 1 0 34684 0 -1 34272
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
timestamp 1586364061
transform 1 0 34500 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 34132 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_58_356
timestamp 1586364061
transform 1 0 33856 0 -1 34272
box -38 -48 314 592
use scs8hd_fill_2  FILLER_58_361
timestamp 1586364061
transform 1 0 34316 0 -1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_519
timestamp 1586364061
transform 1 0 37628 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_58_384
timestamp 1586364061
transform 1 0 36432 0 -1 34272
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_58_396
timestamp 1586364061
transform 1 0 37536 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_3  PHY_117
timestamp 1586364061
transform -1 0 38824 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_8  FILLER_58_398
timestamp 1586364061
transform 1 0 37720 0 -1 34272
box -38 -48 774 592
use scs8hd_fill_1  FILLER_58_406
timestamp 1586364061
transform 1 0 38456 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_3  PHY_118
timestamp 1586364061
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_120
timestamp 1586364061
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_59_3
timestamp 1586364061
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_15
timestamp 1586364061
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_3
timestamp 1586364061
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_15
timestamp 1586364061
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_526
timestamp 1586364061
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_27
timestamp 1586364061
transform 1 0 3588 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_39
timestamp 1586364061
transform 1 0 4692 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_60_27
timestamp 1586364061
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use scs8hd_decap_12  FILLER_60_32
timestamp 1586364061
transform 1 0 4048 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_44
timestamp 1586364061
transform 1 0 5152 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_520
timestamp 1586364061
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use scs8hd_decap_8  FILLER_59_51
timestamp 1586364061
transform 1 0 5796 0 1 34272
box -38 -48 774 592
use scs8hd_fill_2  FILLER_59_59
timestamp 1586364061
transform 1 0 6532 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_59_62
timestamp 1586364061
transform 1 0 6808 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_74
timestamp 1586364061
transform 1 0 7912 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_56
timestamp 1586364061
transform 1 0 6256 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_68
timestamp 1586364061
transform 1 0 7360 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_527
timestamp 1586364061
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_86
timestamp 1586364061
transform 1 0 9016 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_98
timestamp 1586364061
transform 1 0 10120 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_80
timestamp 1586364061
transform 1 0 8464 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_93
timestamp 1586364061
transform 1 0 9660 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_521
timestamp 1586364061
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_110
timestamp 1586364061
transform 1 0 11224 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_123
timestamp 1586364061
transform 1 0 12420 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_105
timestamp 1586364061
transform 1 0 10764 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_117
timestamp 1586364061
transform 1 0 11868 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_135
timestamp 1586364061
transform 1 0 13524 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_147
timestamp 1586364061
transform 1 0 14628 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_129
timestamp 1586364061
transform 1 0 12972 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_141
timestamp 1586364061
transform 1 0 14076 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_528
timestamp 1586364061
transform 1 0 15180 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_159
timestamp 1586364061
transform 1 0 15732 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_171
timestamp 1586364061
transform 1 0 16836 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_154
timestamp 1586364061
transform 1 0 15272 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_166
timestamp 1586364061
transform 1 0 16376 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_522
timestamp 1586364061
transform 1 0 17940 0 1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_184
timestamp 1586364061
transform 1 0 18032 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_196
timestamp 1586364061
transform 1 0 19136 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_178
timestamp 1586364061
transform 1 0 17480 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_190
timestamp 1586364061
transform 1 0 18584 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_529
timestamp 1586364061
transform 1 0 20792 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_208
timestamp 1586364061
transform 1 0 20240 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_220
timestamp 1586364061
transform 1 0 21344 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_202
timestamp 1586364061
transform 1 0 19688 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_215
timestamp 1586364061
transform 1 0 20884 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_523
timestamp 1586364061
transform 1 0 23552 0 1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_232
timestamp 1586364061
transform 1 0 22448 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_245
timestamp 1586364061
transform 1 0 23644 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_227
timestamp 1586364061
transform 1 0 21988 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_239
timestamp 1586364061
transform 1 0 23092 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_257
timestamp 1586364061
transform 1 0 24748 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_269
timestamp 1586364061
transform 1 0 25852 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_251
timestamp 1586364061
transform 1 0 24196 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_263
timestamp 1586364061
transform 1 0 25300 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_530
timestamp 1586364061
transform 1 0 26404 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_281
timestamp 1586364061
transform 1 0 26956 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_59_293
timestamp 1586364061
transform 1 0 28060 0 1 34272
box -38 -48 774 592
use scs8hd_decap_12  FILLER_60_276
timestamp 1586364061
transform 1 0 26496 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_288
timestamp 1586364061
transform 1 0 27600 0 -1 35360
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_59_310
timestamp 1586364061
transform 1 0 29624 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_306
timestamp 1586364061
transform 1 0 29256 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_301
timestamp 1586364061
transform 1 0 28796 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 28980 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
timestamp 1586364061
transform 1 0 29440 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_524
timestamp 1586364061
transform 1 0 29164 0 1 34272
box -38 -48 130 592
use scs8hd_fill_1  FILLER_60_318
timestamp 1586364061
transform 1 0 30360 0 -1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_60_314
timestamp 1586364061
transform 1 0 29992 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 29808 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
timestamp 1586364061
transform 1 0 30176 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
timestamp 1586364061
transform 1 0 29808 0 1 34272
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1586364061
transform 1 0 30452 0 -1 35360
box -38 -48 866 592
use scs8hd_decap_12  FILLER_60_300
timestamp 1586364061
transform 1 0 28704 0 -1 35360
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
timestamp 1586364061
transform 1 0 29992 0 1 34272
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_531
timestamp 1586364061
transform 1 0 32016 0 -1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 33028 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 31924 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 32660 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_333
timestamp 1586364061
transform 1 0 31740 0 1 34272
box -38 -48 222 592
use scs8hd_decap_6  FILLER_59_337
timestamp 1586364061
transform 1 0 32108 0 1 34272
box -38 -48 590 592
use scs8hd_fill_2  FILLER_59_345
timestamp 1586364061
transform 1 0 32844 0 1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_60_328
timestamp 1586364061
transform 1 0 31280 0 -1 35360
box -38 -48 774 592
use scs8hd_decap_12  FILLER_60_337
timestamp 1586364061
transform 1 0 32108 0 -1 35360
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_60_359
timestamp 1586364061
transform 1 0 34132 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_8  FILLER_60_351
timestamp 1586364061
transform 1 0 33396 0 -1 35360
box -38 -48 774 592
use scs8hd_fill_2  FILLER_59_358
timestamp 1586364061
transform 1 0 34040 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 33212 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 34224 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 34224 0 1 34272
box -38 -48 222 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1586364061
transform 1 0 33212 0 1 34272
box -38 -48 866 592
use scs8hd_fill_2  FILLER_60_371
timestamp 1586364061
transform 1 0 35236 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_362
timestamp 1586364061
transform 1 0 34408 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
timestamp 1586364061
transform 1 0 34592 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_525
timestamp 1586364061
transform 1 0 34776 0 1 34272
box -38 -48 130 592
use scs8hd_mux2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1586364061
transform 1 0 34408 0 -1 35360
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
timestamp 1586364061
transform 1 0 34868 0 1 34272
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_60_375
timestamp 1586364061
transform 1 0 35604 0 -1 35360
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
timestamp 1586364061
transform 1 0 35420 0 -1 35360
box -38 -48 222 592
use scs8hd_buf_2  _80_
timestamp 1586364061
transform 1 0 35972 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_60_395
timestamp 1586364061
transform 1 0 37444 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_59_390
timestamp 1586364061
transform 1 0 36984 0 1 34272
box -38 -48 406 592
use scs8hd_fill_2  FILLER_59_386
timestamp 1586364061
transform 1 0 36616 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__80__A
timestamp 1586364061
transform 1 0 36800 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_532
timestamp 1586364061
transform 1 0 37628 0 -1 35360
box -38 -48 130 592
use scs8hd_buf_2  _79_
timestamp 1586364061
transform 1 0 37352 0 1 34272
box -38 -48 406 592
use scs8hd_decap_12  FILLER_60_383
timestamp 1586364061
transform 1 0 36340 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_3  PHY_119
timestamp 1586364061
transform -1 0 38824 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_121
timestamp 1586364061
transform -1 0 38824 0 -1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__79__A
timestamp 1586364061
transform 1 0 37904 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_398
timestamp 1586364061
transform 1 0 37720 0 1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_59_402
timestamp 1586364061
transform 1 0 38088 0 1 34272
box -38 -48 406 592
use scs8hd_fill_1  FILLER_59_406
timestamp 1586364061
transform 1 0 38456 0 1 34272
box -38 -48 130 592
use scs8hd_decap_8  FILLER_60_398
timestamp 1586364061
transform 1 0 37720 0 -1 35360
box -38 -48 774 592
use scs8hd_fill_1  FILLER_60_406
timestamp 1586364061
transform 1 0 38456 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_3  PHY_122
timestamp 1586364061
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_61_3
timestamp 1586364061
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_15
timestamp 1586364061
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_27
timestamp 1586364061
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_39
timestamp 1586364061
transform 1 0 4692 0 1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_533
timestamp 1586364061
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use scs8hd_decap_8  FILLER_61_51
timestamp 1586364061
transform 1 0 5796 0 1 35360
box -38 -48 774 592
use scs8hd_fill_2  FILLER_61_59
timestamp 1586364061
transform 1 0 6532 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_62
timestamp 1586364061
transform 1 0 6808 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_74
timestamp 1586364061
transform 1 0 7912 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_86
timestamp 1586364061
transform 1 0 9016 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_98
timestamp 1586364061
transform 1 0 10120 0 1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_534
timestamp 1586364061
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_61_110
timestamp 1586364061
transform 1 0 11224 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_123
timestamp 1586364061
transform 1 0 12420 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_135
timestamp 1586364061
transform 1 0 13524 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_147
timestamp 1586364061
transform 1 0 14628 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_159
timestamp 1586364061
transform 1 0 15732 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_171
timestamp 1586364061
transform 1 0 16836 0 1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_535
timestamp 1586364061
transform 1 0 17940 0 1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_61_184
timestamp 1586364061
transform 1 0 18032 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_196
timestamp 1586364061
transform 1 0 19136 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_208
timestamp 1586364061
transform 1 0 20240 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_220
timestamp 1586364061
transform 1 0 21344 0 1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_536
timestamp 1586364061
transform 1 0 23552 0 1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_61_232
timestamp 1586364061
transform 1 0 22448 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_245
timestamp 1586364061
transform 1 0 23644 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_257
timestamp 1586364061
transform 1 0 24748 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_269
timestamp 1586364061
transform 1 0 25852 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_281
timestamp 1586364061
transform 1 0 26956 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_293
timestamp 1586364061
transform 1 0 28060 0 1 35360
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
timestamp 1586364061
transform 1 0 30176 0 1 35360
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_537
timestamp 1586364061
transform 1 0 29164 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
timestamp 1586364061
transform 1 0 29992 0 1 35360
box -38 -48 222 592
use scs8hd_decap_8  FILLER_61_306
timestamp 1586364061
transform 1 0 29256 0 1 35360
box -38 -48 774 592
use scs8hd_decap_12  FILLER_61_335
timestamp 1586364061
transform 1 0 31924 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_347
timestamp 1586364061
transform 1 0 33028 0 1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_538
timestamp 1586364061
transform 1 0 34776 0 1 35360
box -38 -48 130 592
use scs8hd_decap_6  FILLER_61_359
timestamp 1586364061
transform 1 0 34132 0 1 35360
box -38 -48 590 592
use scs8hd_fill_1  FILLER_61_365
timestamp 1586364061
transform 1 0 34684 0 1 35360
box -38 -48 130 592
use scs8hd_decap_6  FILLER_61_367
timestamp 1586364061
transform 1 0 34868 0 1 35360
box -38 -48 590 592
use scs8hd_buf_2  _78_
timestamp 1586364061
transform 1 0 35420 0 1 35360
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__78__A
timestamp 1586364061
transform 1 0 35972 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_377
timestamp 1586364061
transform 1 0 35788 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_381
timestamp 1586364061
transform 1 0 36156 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_393
timestamp 1586364061
transform 1 0 37260 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_3  PHY_123
timestamp 1586364061
transform -1 0 38824 0 1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_61_405
timestamp 1586364061
transform 1 0 38364 0 1 35360
box -38 -48 222 592
use scs8hd_decap_3  PHY_124
timestamp 1586364061
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_62_3
timestamp 1586364061
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_15
timestamp 1586364061
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_539
timestamp 1586364061
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_4  FILLER_62_27
timestamp 1586364061
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use scs8hd_decap_12  FILLER_62_32
timestamp 1586364061
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_44
timestamp 1586364061
transform 1 0 5152 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_56
timestamp 1586364061
transform 1 0 6256 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_68
timestamp 1586364061
transform 1 0 7360 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_540
timestamp 1586364061
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_80
timestamp 1586364061
transform 1 0 8464 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_93
timestamp 1586364061
transform 1 0 9660 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_105
timestamp 1586364061
transform 1 0 10764 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_117
timestamp 1586364061
transform 1 0 11868 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_129
timestamp 1586364061
transform 1 0 12972 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_141
timestamp 1586364061
transform 1 0 14076 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_541
timestamp 1586364061
transform 1 0 15180 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_154
timestamp 1586364061
transform 1 0 15272 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_166
timestamp 1586364061
transform 1 0 16376 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_178
timestamp 1586364061
transform 1 0 17480 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_190
timestamp 1586364061
transform 1 0 18584 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_542
timestamp 1586364061
transform 1 0 20792 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_202
timestamp 1586364061
transform 1 0 19688 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_215
timestamp 1586364061
transform 1 0 20884 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_227
timestamp 1586364061
transform 1 0 21988 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_239
timestamp 1586364061
transform 1 0 23092 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_251
timestamp 1586364061
transform 1 0 24196 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_263
timestamp 1586364061
transform 1 0 25300 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_543
timestamp 1586364061
transform 1 0 26404 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_276
timestamp 1586364061
transform 1 0 26496 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_288
timestamp 1586364061
transform 1 0 27600 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_300
timestamp 1586364061
transform 1 0 28704 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_312
timestamp 1586364061
transform 1 0 29808 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_544
timestamp 1586364061
transform 1 0 32016 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_324
timestamp 1586364061
transform 1 0 30912 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_337
timestamp 1586364061
transform 1 0 32108 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_349
timestamp 1586364061
transform 1 0 33212 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_361
timestamp 1586364061
transform 1 0 34316 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_545
timestamp 1586364061
transform 1 0 37628 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_373
timestamp 1586364061
transform 1 0 35420 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_385
timestamp 1586364061
transform 1 0 36524 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_3  PHY_125
timestamp 1586364061
transform -1 0 38824 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_8  FILLER_62_398
timestamp 1586364061
transform 1 0 37720 0 -1 36448
box -38 -48 774 592
use scs8hd_fill_1  FILLER_62_406
timestamp 1586364061
transform 1 0 38456 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_3  PHY_126
timestamp 1586364061
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_3
timestamp 1586364061
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_15
timestamp 1586364061
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_27
timestamp 1586364061
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_39
timestamp 1586364061
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_546
timestamp 1586364061
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use scs8hd_decap_8  FILLER_63_51
timestamp 1586364061
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use scs8hd_fill_2  FILLER_63_59
timestamp 1586364061
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_63_62
timestamp 1586364061
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_74
timestamp 1586364061
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_86
timestamp 1586364061
transform 1 0 9016 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_98
timestamp 1586364061
transform 1 0 10120 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_547
timestamp 1586364061
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_110
timestamp 1586364061
transform 1 0 11224 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_123
timestamp 1586364061
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_135
timestamp 1586364061
transform 1 0 13524 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_147
timestamp 1586364061
transform 1 0 14628 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_159
timestamp 1586364061
transform 1 0 15732 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_171
timestamp 1586364061
transform 1 0 16836 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_548
timestamp 1586364061
transform 1 0 17940 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_184
timestamp 1586364061
transform 1 0 18032 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_196
timestamp 1586364061
transform 1 0 19136 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_208
timestamp 1586364061
transform 1 0 20240 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_220
timestamp 1586364061
transform 1 0 21344 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_549
timestamp 1586364061
transform 1 0 23552 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_232
timestamp 1586364061
transform 1 0 22448 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_245
timestamp 1586364061
transform 1 0 23644 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_257
timestamp 1586364061
transform 1 0 24748 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_269
timestamp 1586364061
transform 1 0 25852 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_281
timestamp 1586364061
transform 1 0 26956 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_293
timestamp 1586364061
transform 1 0 28060 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_550
timestamp 1586364061
transform 1 0 29164 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_306
timestamp 1586364061
transform 1 0 29256 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_318
timestamp 1586364061
transform 1 0 30360 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_330
timestamp 1586364061
transform 1 0 31464 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_342
timestamp 1586364061
transform 1 0 32568 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_551
timestamp 1586364061
transform 1 0 34776 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_354
timestamp 1586364061
transform 1 0 33672 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_367
timestamp 1586364061
transform 1 0 34868 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_379
timestamp 1586364061
transform 1 0 35972 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_391
timestamp 1586364061
transform 1 0 37076 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_3  PHY_127
timestamp 1586364061
transform -1 0 38824 0 1 36448
box -38 -48 314 592
use scs8hd_decap_4  FILLER_63_403
timestamp 1586364061
transform 1 0 38180 0 1 36448
box -38 -48 406 592
use scs8hd_decap_3  PHY_128
timestamp 1586364061
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_64_3
timestamp 1586364061
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_15
timestamp 1586364061
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_552
timestamp 1586364061
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_4  FILLER_64_27
timestamp 1586364061
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use scs8hd_decap_12  FILLER_64_32
timestamp 1586364061
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_44
timestamp 1586364061
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_553
timestamp 1586364061
transform 1 0 6808 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_56
timestamp 1586364061
transform 1 0 6256 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_63
timestamp 1586364061
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_554
timestamp 1586364061
transform 1 0 9660 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_75
timestamp 1586364061
transform 1 0 8004 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_64_87
timestamp 1586364061
transform 1 0 9108 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_94
timestamp 1586364061
transform 1 0 9752 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_555
timestamp 1586364061
transform 1 0 12512 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_106
timestamp 1586364061
transform 1 0 10856 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_64_118
timestamp 1586364061
transform 1 0 11960 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_125
timestamp 1586364061
transform 1 0 12604 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_137
timestamp 1586364061
transform 1 0 13708 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_64_149
timestamp 1586364061
transform 1 0 14812 0 -1 37536
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_556
timestamp 1586364061
transform 1 0 15364 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_156
timestamp 1586364061
transform 1 0 15456 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_168
timestamp 1586364061
transform 1 0 16560 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_557
timestamp 1586364061
transform 1 0 18216 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_180
timestamp 1586364061
transform 1 0 17664 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_187
timestamp 1586364061
transform 1 0 18308 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_558
timestamp 1586364061
transform 1 0 21068 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_199
timestamp 1586364061
transform 1 0 19412 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_64_211
timestamp 1586364061
transform 1 0 20516 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_218
timestamp 1586364061
transform 1 0 21160 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_559
timestamp 1586364061
transform 1 0 23920 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_230
timestamp 1586364061
transform 1 0 22264 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_64_242
timestamp 1586364061
transform 1 0 23368 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_249
timestamp 1586364061
transform 1 0 24012 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_261
timestamp 1586364061
transform 1 0 25116 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_64_273
timestamp 1586364061
transform 1 0 26220 0 -1 37536
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_560
timestamp 1586364061
transform 1 0 26772 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_280
timestamp 1586364061
transform 1 0 26864 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_292
timestamp 1586364061
transform 1 0 27968 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_561
timestamp 1586364061
transform 1 0 29624 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_304
timestamp 1586364061
transform 1 0 29072 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_311
timestamp 1586364061
transform 1 0 29716 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_562
timestamp 1586364061
transform 1 0 32476 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_323
timestamp 1586364061
transform 1 0 30820 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_64_335
timestamp 1586364061
transform 1 0 31924 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_342
timestamp 1586364061
transform 1 0 32568 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_563
timestamp 1586364061
transform 1 0 35328 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_354
timestamp 1586364061
transform 1 0 33672 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_64_366
timestamp 1586364061
transform 1 0 34776 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_373
timestamp 1586364061
transform 1 0 35420 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_385
timestamp 1586364061
transform 1 0 36524 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_64_397
timestamp 1586364061
transform 1 0 37628 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_3  PHY_129
timestamp 1586364061
transform -1 0 38824 0 -1 37536
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_564
timestamp 1586364061
transform 1 0 38180 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_3  FILLER_64_404
timestamp 1586364061
transform 1 0 38272 0 -1 37536
box -38 -48 314 592
<< labels >>
rlabel metal2 s 38290 0 38346 480 6 Test_en
port 0 nsew default input
rlabel metal2 s 9402 0 9458 480 6 bottom_width_0_height_0__pin_16_
port 1 nsew default input
rlabel metal2 s 10506 0 10562 480 6 bottom_width_0_height_0__pin_17_
port 2 nsew default input
rlabel metal2 s 11610 0 11666 480 6 bottom_width_0_height_0__pin_18_
port 3 nsew default input
rlabel metal2 s 12714 0 12770 480 6 bottom_width_0_height_0__pin_19_
port 4 nsew default input
rlabel metal2 s 13910 0 13966 480 6 bottom_width_0_height_0__pin_20_
port 5 nsew default input
rlabel metal2 s 15014 0 15070 480 6 bottom_width_0_height_0__pin_21_
port 6 nsew default input
rlabel metal2 s 16118 0 16174 480 6 bottom_width_0_height_0__pin_22_
port 7 nsew default input
rlabel metal2 s 17222 0 17278 480 6 bottom_width_0_height_0__pin_23_
port 8 nsew default input
rlabel metal2 s 18326 0 18382 480 6 bottom_width_0_height_0__pin_24_
port 9 nsew default input
rlabel metal2 s 19430 0 19486 480 6 bottom_width_0_height_0__pin_25_
port 10 nsew default input
rlabel metal2 s 20534 0 20590 480 6 bottom_width_0_height_0__pin_26_
port 11 nsew default input
rlabel metal2 s 21638 0 21694 480 6 bottom_width_0_height_0__pin_27_
port 12 nsew default input
rlabel metal2 s 22742 0 22798 480 6 bottom_width_0_height_0__pin_28_
port 13 nsew default input
rlabel metal2 s 23846 0 23902 480 6 bottom_width_0_height_0__pin_29_
port 14 nsew default input
rlabel metal2 s 24950 0 25006 480 6 bottom_width_0_height_0__pin_30_
port 15 nsew default input
rlabel metal2 s 26054 0 26110 480 6 bottom_width_0_height_0__pin_31_
port 16 nsew default input
rlabel metal2 s 29458 0 29514 480 6 bottom_width_0_height_0__pin_42_lower
port 17 nsew default tristate
rlabel metal2 s 570 0 626 480 6 bottom_width_0_height_0__pin_42_upper
port 18 nsew default tristate
rlabel metal2 s 30562 0 30618 480 6 bottom_width_0_height_0__pin_43_lower
port 19 nsew default tristate
rlabel metal2 s 1674 0 1730 480 6 bottom_width_0_height_0__pin_43_upper
port 20 nsew default tristate
rlabel metal2 s 31666 0 31722 480 6 bottom_width_0_height_0__pin_44_lower
port 21 nsew default tristate
rlabel metal2 s 2778 0 2834 480 6 bottom_width_0_height_0__pin_44_upper
port 22 nsew default tristate
rlabel metal2 s 32770 0 32826 480 6 bottom_width_0_height_0__pin_45_lower
port 23 nsew default tristate
rlabel metal2 s 3882 0 3938 480 6 bottom_width_0_height_0__pin_45_upper
port 24 nsew default tristate
rlabel metal2 s 33874 0 33930 480 6 bottom_width_0_height_0__pin_46_lower
port 25 nsew default tristate
rlabel metal2 s 4986 0 5042 480 6 bottom_width_0_height_0__pin_46_upper
port 26 nsew default tristate
rlabel metal2 s 34978 0 35034 480 6 bottom_width_0_height_0__pin_47_lower
port 27 nsew default tristate
rlabel metal2 s 6090 0 6146 480 6 bottom_width_0_height_0__pin_47_upper
port 28 nsew default tristate
rlabel metal2 s 36082 0 36138 480 6 bottom_width_0_height_0__pin_48_lower
port 29 nsew default tristate
rlabel metal2 s 7194 0 7250 480 6 bottom_width_0_height_0__pin_48_upper
port 30 nsew default tristate
rlabel metal2 s 37186 0 37242 480 6 bottom_width_0_height_0__pin_49_lower
port 31 nsew default tristate
rlabel metal2 s 8298 0 8354 480 6 bottom_width_0_height_0__pin_49_upper
port 32 nsew default tristate
rlabel metal2 s 27250 0 27306 480 6 bottom_width_0_height_0__pin_50_
port 33 nsew default tristate
rlabel metal2 s 28354 0 28410 480 6 bottom_width_0_height_0__pin_51_
port 34 nsew default tristate
rlabel metal3 s 0 20000 480 20120 6 ccff_head
port 35 nsew default input
rlabel metal3 s 39520 11976 40000 12096 6 ccff_tail
port 36 nsew default tristate
rlabel metal2 s 39394 0 39450 480 6 clk
port 37 nsew default input
rlabel metal3 s 0 33328 480 33448 6 left_width_0_height_0__pin_52_
port 38 nsew default input
rlabel metal3 s 0 6672 480 6792 6 prog_clk
port 39 nsew default input
rlabel metal3 s 39520 13064 40000 13184 6 right_width_0_height_0__pin_0_
port 40 nsew default input
rlabel metal3 s 39520 24488 40000 24608 6 right_width_0_height_0__pin_10_
port 41 nsew default input
rlabel metal3 s 39520 25576 40000 25696 6 right_width_0_height_0__pin_11_
port 42 nsew default input
rlabel metal3 s 39520 26800 40000 26920 6 right_width_0_height_0__pin_12_
port 43 nsew default input
rlabel metal3 s 39520 27888 40000 28008 6 right_width_0_height_0__pin_13_
port 44 nsew default input
rlabel metal3 s 39520 29112 40000 29232 6 right_width_0_height_0__pin_14_
port 45 nsew default input
rlabel metal3 s 39520 30200 40000 30320 6 right_width_0_height_0__pin_15_
port 46 nsew default input
rlabel metal3 s 39520 14152 40000 14272 6 right_width_0_height_0__pin_1_
port 47 nsew default input
rlabel metal3 s 39520 15376 40000 15496 6 right_width_0_height_0__pin_2_
port 48 nsew default input
rlabel metal3 s 39520 5040 40000 5160 6 right_width_0_height_0__pin_34_lower
port 49 nsew default tristate
rlabel metal3 s 39520 31288 40000 31408 6 right_width_0_height_0__pin_34_upper
port 50 nsew default tristate
rlabel metal3 s 39520 6264 40000 6384 6 right_width_0_height_0__pin_35_lower
port 51 nsew default tristate
rlabel metal3 s 39520 32512 40000 32632 6 right_width_0_height_0__pin_35_upper
port 52 nsew default tristate
rlabel metal3 s 39520 7352 40000 7472 6 right_width_0_height_0__pin_36_lower
port 53 nsew default tristate
rlabel metal3 s 39520 33600 40000 33720 6 right_width_0_height_0__pin_36_upper
port 54 nsew default tristate
rlabel metal3 s 39520 8440 40000 8560 6 right_width_0_height_0__pin_37_lower
port 55 nsew default tristate
rlabel metal3 s 39520 34824 40000 34944 6 right_width_0_height_0__pin_37_upper
port 56 nsew default tristate
rlabel metal3 s 39520 9664 40000 9784 6 right_width_0_height_0__pin_38_lower
port 57 nsew default tristate
rlabel metal3 s 39520 35912 40000 36032 6 right_width_0_height_0__pin_38_upper
port 58 nsew default tristate
rlabel metal3 s 39520 10752 40000 10872 6 right_width_0_height_0__pin_39_lower
port 59 nsew default tristate
rlabel metal3 s 39520 37000 40000 37120 6 right_width_0_height_0__pin_39_upper
port 60 nsew default tristate
rlabel metal3 s 39520 16464 40000 16584 6 right_width_0_height_0__pin_3_
port 61 nsew default input
rlabel metal3 s 39520 2728 40000 2848 6 right_width_0_height_0__pin_40_lower
port 62 nsew default tristate
rlabel metal3 s 39520 38224 40000 38344 6 right_width_0_height_0__pin_40_upper
port 63 nsew default tristate
rlabel metal3 s 39520 3952 40000 4072 6 right_width_0_height_0__pin_41_lower
port 64 nsew default tristate
rlabel metal3 s 39520 39312 40000 39432 6 right_width_0_height_0__pin_41_upper
port 65 nsew default tristate
rlabel metal3 s 39520 17688 40000 17808 6 right_width_0_height_0__pin_4_
port 66 nsew default input
rlabel metal3 s 39520 18776 40000 18896 6 right_width_0_height_0__pin_5_
port 67 nsew default input
rlabel metal3 s 39520 19864 40000 19984 6 right_width_0_height_0__pin_6_
port 68 nsew default input
rlabel metal3 s 39520 21088 40000 21208 6 right_width_0_height_0__pin_7_
port 69 nsew default input
rlabel metal3 s 39520 22176 40000 22296 6 right_width_0_height_0__pin_8_
port 70 nsew default input
rlabel metal3 s 39520 23400 40000 23520 6 right_width_0_height_0__pin_9_
port 71 nsew default input
rlabel metal3 s 39520 552 40000 672 6 top_width_0_height_0__pin_32_
port 72 nsew default input
rlabel metal3 s 39520 1640 40000 1760 6 top_width_0_height_0__pin_33_
port 73 nsew default input
rlabel metal4 s 4208 2128 4528 37584 6 vpwr
port 74 nsew default input
rlabel metal4 s 19568 2128 19888 37584 6 vgnd
port 75 nsew default input
<< properties >>
string FIXED_BBOX 0 0 40000 39432
<< end >>
