magic
tech sky130A
magscale 1 2
timestamp 1609018222
<< locali >>
rect 22017 16779 22051 17561
rect 19901 15963 19935 16065
rect 9689 12087 9723 12257
rect 22017 11339 22051 11985
rect 17785 11067 17819 11237
rect 17325 9979 17359 10149
rect 7849 8891 7883 9129
rect 10793 8347 10827 8449
rect 13277 8279 13311 8585
rect 6653 7259 6687 7429
rect 11713 7259 11747 7497
rect 22017 5559 22051 6613
rect 16221 2295 16255 2465
rect 6193 1819 6227 2057
<< viali >>
rect 4813 20553 4847 20587
rect 18981 20553 19015 20587
rect 19165 20553 19199 20587
rect 21373 20553 21407 20587
rect 6929 20485 6963 20519
rect 21189 20485 21223 20519
rect 7481 20417 7515 20451
rect 20821 20417 20855 20451
rect 4629 20349 4663 20383
rect 19993 20349 20027 20383
rect 20545 20349 20579 20383
rect 7389 20281 7423 20315
rect 20269 20281 20303 20315
rect 7297 20213 7331 20247
rect 19717 20213 19751 20247
rect 19901 20213 19935 20247
rect 7297 20009 7331 20043
rect 9965 20009 9999 20043
rect 11069 20009 11103 20043
rect 11989 20009 12023 20043
rect 13277 20009 13311 20043
rect 14749 20009 14783 20043
rect 15485 20009 15519 20043
rect 17325 20009 17359 20043
rect 18705 19941 18739 19975
rect 19349 19941 19383 19975
rect 19993 19941 20027 19975
rect 20545 19941 20579 19975
rect 21189 19941 21223 19975
rect 4344 19873 4378 19907
rect 6092 19873 6126 19907
rect 8033 19873 8067 19907
rect 9781 19873 9815 19907
rect 10333 19873 10367 19907
rect 10885 19873 10919 19907
rect 11437 19873 11471 19907
rect 11805 19873 11839 19907
rect 12173 19873 12207 19907
rect 13093 19873 13127 19907
rect 14565 19873 14599 19907
rect 15301 19873 15335 19907
rect 15669 19873 15703 19907
rect 17049 19873 17083 19907
rect 17141 19873 17175 19907
rect 18429 19873 18463 19907
rect 19073 19873 19107 19907
rect 19717 19873 19751 19907
rect 20269 19873 20303 19907
rect 20913 19873 20947 19907
rect 4077 19805 4111 19839
rect 5825 19805 5859 19839
rect 8125 19805 8159 19839
rect 8309 19805 8343 19839
rect 10609 19805 10643 19839
rect 21465 19805 21499 19839
rect 7573 19737 7607 19771
rect 8585 19737 8619 19771
rect 11621 19737 11655 19771
rect 5457 19669 5491 19703
rect 7205 19669 7239 19703
rect 7665 19669 7699 19703
rect 8769 19669 8803 19703
rect 1961 19465 1995 19499
rect 6653 19465 6687 19499
rect 15117 19465 15151 19499
rect 12081 19397 12115 19431
rect 3801 19329 3835 19363
rect 8953 19329 8987 19363
rect 10057 19329 10091 19363
rect 10977 19329 11011 19363
rect 11897 19329 11931 19363
rect 12725 19329 12759 19363
rect 21281 19329 21315 19363
rect 1777 19261 1811 19295
rect 3249 19261 3283 19295
rect 5273 19261 5307 19295
rect 6929 19261 6963 19295
rect 7196 19261 7230 19295
rect 8769 19261 8803 19295
rect 9229 19261 9263 19295
rect 9505 19261 9539 19295
rect 9781 19261 9815 19295
rect 10793 19261 10827 19295
rect 11621 19261 11655 19295
rect 12449 19261 12483 19295
rect 13001 19261 13035 19295
rect 13369 19261 13403 19295
rect 13737 19261 13771 19295
rect 14197 19261 14231 19295
rect 14565 19261 14599 19295
rect 14933 19261 14967 19295
rect 15577 19261 15611 19295
rect 16129 19261 16163 19295
rect 16497 19261 16531 19295
rect 17141 19261 17175 19295
rect 17601 19261 17635 19295
rect 18061 19261 18095 19295
rect 18245 19261 18279 19295
rect 18521 19261 18555 19295
rect 18889 19261 18923 19295
rect 19993 19261 20027 19295
rect 20177 19261 20211 19295
rect 20453 19261 20487 19295
rect 20729 19261 20763 19295
rect 21005 19261 21039 19295
rect 3525 19193 3559 19227
rect 4068 19193 4102 19227
rect 5540 19193 5574 19227
rect 15853 19193 15887 19227
rect 19717 19193 19751 19227
rect 21465 19193 21499 19227
rect 2237 19125 2271 19159
rect 5181 19125 5215 19159
rect 8309 19125 8343 19159
rect 8401 19125 8435 19159
rect 8861 19125 8895 19159
rect 10425 19125 10459 19159
rect 10885 19125 10919 19159
rect 11253 19125 11287 19159
rect 11713 19125 11747 19159
rect 13185 19125 13219 19159
rect 13553 19125 13587 19159
rect 13921 19125 13955 19159
rect 14381 19125 14415 19159
rect 14749 19125 14783 19159
rect 15301 19125 15335 19159
rect 16313 19125 16347 19159
rect 16681 19125 16715 19159
rect 16957 19125 16991 19159
rect 17325 19125 17359 19159
rect 17785 19125 17819 19159
rect 1961 18921 1995 18955
rect 3801 18921 3835 18955
rect 4721 18921 4755 18955
rect 5457 18921 5491 18955
rect 5917 18921 5951 18955
rect 6285 18921 6319 18955
rect 7205 18921 7239 18955
rect 7573 18921 7607 18955
rect 10149 18921 10183 18955
rect 16221 18921 16255 18955
rect 19809 18921 19843 18955
rect 19993 18921 20027 18955
rect 21465 18921 21499 18955
rect 5365 18853 5399 18887
rect 8033 18853 8067 18887
rect 8677 18853 8711 18887
rect 17049 18853 17083 18887
rect 17969 18853 18003 18887
rect 20545 18853 20579 18887
rect 21189 18853 21223 18887
rect 1777 18785 1811 18819
rect 2145 18785 2179 18819
rect 3065 18785 3099 18819
rect 5825 18785 5859 18819
rect 6653 18785 6687 18819
rect 7665 18785 7699 18819
rect 8585 18785 8619 18819
rect 10876 18785 10910 18819
rect 18061 18785 18095 18819
rect 18613 18785 18647 18819
rect 19165 18785 19199 18819
rect 20269 18785 20303 18819
rect 20913 18785 20947 18819
rect 2973 18717 3007 18751
rect 4169 18717 4203 18751
rect 4813 18717 4847 18751
rect 4997 18717 5031 18751
rect 6101 18717 6135 18751
rect 6745 18717 6779 18751
rect 6929 18717 6963 18751
rect 7757 18717 7791 18751
rect 8861 18717 8895 18751
rect 10241 18717 10275 18751
rect 10425 18717 10459 18751
rect 10609 18717 10643 18751
rect 12817 18717 12851 18751
rect 18245 18717 18279 18751
rect 18797 18717 18831 18751
rect 19349 18717 19383 18751
rect 9781 18649 9815 18683
rect 13185 18649 13219 18683
rect 2697 18581 2731 18615
rect 4353 18581 4387 18615
rect 8217 18581 8251 18615
rect 11989 18581 12023 18615
rect 13645 18581 13679 18615
rect 14105 18581 14139 18615
rect 14473 18581 14507 18615
rect 15945 18581 15979 18615
rect 2329 18377 2363 18411
rect 4905 18377 4939 18411
rect 7389 18377 7423 18411
rect 8217 18377 8251 18411
rect 16681 18377 16715 18411
rect 18705 18377 18739 18411
rect 19717 18377 19751 18411
rect 19993 18377 20027 18411
rect 20269 18377 20303 18411
rect 21465 18377 21499 18411
rect 10057 18309 10091 18343
rect 20361 18309 20395 18343
rect 3709 18241 3743 18275
rect 4537 18241 4571 18275
rect 6377 18241 6411 18275
rect 6561 18241 6595 18275
rect 6837 18241 6871 18275
rect 7941 18241 7975 18275
rect 12449 18241 12483 18275
rect 14197 18241 14231 18275
rect 1777 18173 1811 18207
rect 2145 18173 2179 18207
rect 2513 18173 2547 18207
rect 3433 18173 3467 18207
rect 4353 18173 4387 18207
rect 6285 18173 6319 18207
rect 8677 18173 8711 18207
rect 10149 18173 10183 18207
rect 10416 18173 10450 18207
rect 11621 18173 11655 18207
rect 13921 18173 13955 18207
rect 16497 18173 16531 18207
rect 18429 18173 18463 18207
rect 18521 18173 18555 18207
rect 19533 18173 19567 18207
rect 20729 18173 20763 18207
rect 21281 18173 21315 18207
rect 3525 18105 3559 18139
rect 4261 18105 4295 18139
rect 5089 18105 5123 18139
rect 7849 18105 7883 18139
rect 8922 18105 8956 18139
rect 12694 18105 12728 18139
rect 21005 18105 21039 18139
rect 1961 18037 1995 18071
rect 2697 18037 2731 18071
rect 2881 18037 2915 18071
rect 3065 18037 3099 18071
rect 3893 18037 3927 18071
rect 4721 18037 4755 18071
rect 5917 18037 5951 18071
rect 7757 18037 7791 18071
rect 11529 18037 11563 18071
rect 13829 18037 13863 18071
rect 19349 18037 19383 18071
rect 20545 18037 20579 18071
rect 1593 17833 1627 17867
rect 2789 17833 2823 17867
rect 3617 17833 3651 17867
rect 4077 17833 4111 17867
rect 4445 17833 4479 17867
rect 4905 17833 4939 17867
rect 6469 17833 6503 17867
rect 6929 17833 6963 17867
rect 9965 17833 9999 17867
rect 10425 17833 10459 17867
rect 10793 17833 10827 17867
rect 11621 17833 11655 17867
rect 11989 17833 12023 17867
rect 13553 17833 13587 17867
rect 14197 17833 14231 17867
rect 20085 17833 20119 17867
rect 21465 17833 21499 17867
rect 2053 17765 2087 17799
rect 3525 17765 3559 17799
rect 5273 17765 5307 17799
rect 8217 17765 8251 17799
rect 10333 17765 10367 17799
rect 11161 17765 11195 17799
rect 15117 17765 15151 17799
rect 16405 17765 16439 17799
rect 1409 17697 1443 17731
rect 1777 17697 1811 17731
rect 2697 17697 2731 17731
rect 4537 17697 4571 17731
rect 6377 17697 6411 17731
rect 6837 17697 6871 17731
rect 8309 17697 8343 17731
rect 9873 17697 9907 17731
rect 11253 17697 11287 17731
rect 12449 17697 12483 17731
rect 13461 17697 13495 17731
rect 14105 17697 14139 17731
rect 15669 17697 15703 17731
rect 16129 17697 16163 17731
rect 19901 17697 19935 17731
rect 20269 17697 20303 17731
rect 20913 17697 20947 17731
rect 2973 17629 3007 17663
rect 3709 17629 3743 17663
rect 4629 17629 4663 17663
rect 5365 17629 5399 17663
rect 5457 17629 5491 17663
rect 7113 17629 7147 17663
rect 8493 17629 8527 17663
rect 10609 17629 10643 17663
rect 11345 17629 11379 17663
rect 12081 17629 12115 17663
rect 12173 17629 12207 17663
rect 14381 17629 14415 17663
rect 15761 17629 15795 17663
rect 15945 17629 15979 17663
rect 20545 17629 20579 17663
rect 21189 17629 21223 17663
rect 8677 17561 8711 17595
rect 13737 17561 13771 17595
rect 19717 17561 19751 17595
rect 22017 17561 22051 17595
rect 2329 17493 2363 17527
rect 3157 17493 3191 17527
rect 7389 17493 7423 17527
rect 7665 17493 7699 17527
rect 7849 17493 7883 17527
rect 15301 17493 15335 17527
rect 1869 17289 1903 17323
rect 6009 17289 6043 17323
rect 6929 17289 6963 17323
rect 9873 17289 9907 17323
rect 10701 17289 10735 17323
rect 15393 17289 15427 17323
rect 16221 17289 16255 17323
rect 20637 17289 20671 17323
rect 21465 17289 21499 17323
rect 4077 17221 4111 17255
rect 4169 17221 4203 17255
rect 5181 17221 5215 17255
rect 6193 17221 6227 17255
rect 7757 17221 7791 17255
rect 15301 17221 15335 17255
rect 2329 17153 2363 17187
rect 2513 17153 2547 17187
rect 4629 17153 4663 17187
rect 4813 17153 4847 17187
rect 5641 17153 5675 17187
rect 5825 17153 5859 17187
rect 6469 17153 6503 17187
rect 7389 17153 7423 17187
rect 7573 17153 7607 17187
rect 8309 17153 8343 17187
rect 8677 17153 8711 17187
rect 10517 17153 10551 17187
rect 11253 17153 11287 17187
rect 11621 17153 11655 17187
rect 15945 17153 15979 17187
rect 16773 17153 16807 17187
rect 20177 17153 20211 17187
rect 2237 17085 2271 17119
rect 2697 17085 2731 17119
rect 5549 17085 5583 17119
rect 9689 17085 9723 17119
rect 10333 17085 10367 17119
rect 11069 17085 11103 17119
rect 11161 17085 11195 17119
rect 12449 17085 12483 17119
rect 13921 17085 13955 17119
rect 15853 17085 15887 17119
rect 16589 17085 16623 17119
rect 19901 17085 19935 17119
rect 20729 17085 20763 17119
rect 21281 17085 21315 17119
rect 2964 17017 2998 17051
rect 6653 17017 6687 17051
rect 7297 17017 7331 17051
rect 12716 17017 12750 17051
rect 14166 17017 14200 17051
rect 21005 17017 21039 17051
rect 1777 16949 1811 16983
rect 4537 16949 4571 16983
rect 4997 16949 5031 16983
rect 8125 16949 8159 16983
rect 8217 16949 8251 16983
rect 8769 16949 8803 16983
rect 9505 16949 9539 16983
rect 10241 16949 10275 16983
rect 13829 16949 13863 16983
rect 15761 16949 15795 16983
rect 16681 16949 16715 16983
rect 3525 16745 3559 16779
rect 5549 16745 5583 16779
rect 6469 16745 6503 16779
rect 8769 16745 8803 16779
rect 9689 16745 9723 16779
rect 11069 16745 11103 16779
rect 11253 16745 11287 16779
rect 12541 16745 12575 16779
rect 12909 16745 12943 16779
rect 14197 16745 14231 16779
rect 16773 16745 16807 16779
rect 17233 16745 17267 16779
rect 21097 16745 21131 16779
rect 22017 16745 22051 16779
rect 4414 16677 4448 16711
rect 6101 16677 6135 16711
rect 6929 16677 6963 16711
rect 9229 16677 9263 16711
rect 10701 16677 10735 16711
rect 11621 16677 11655 16711
rect 13369 16677 13403 16711
rect 14105 16677 14139 16711
rect 21465 16677 21499 16711
rect 1501 16609 1535 16643
rect 2136 16609 2170 16643
rect 6009 16609 6043 16643
rect 6837 16609 6871 16643
rect 7564 16609 7598 16643
rect 9137 16609 9171 16643
rect 10057 16609 10091 16643
rect 10149 16609 10183 16643
rect 11713 16609 11747 16643
rect 12449 16609 12483 16643
rect 13277 16609 13311 16643
rect 15025 16609 15059 16643
rect 15568 16609 15602 16643
rect 17141 16609 17175 16643
rect 20913 16609 20947 16643
rect 21281 16609 21315 16643
rect 1869 16541 1903 16575
rect 4169 16541 4203 16575
rect 6285 16541 6319 16575
rect 7113 16541 7147 16575
rect 7297 16541 7331 16575
rect 9321 16541 9355 16575
rect 10241 16541 10275 16575
rect 11897 16541 11931 16575
rect 12725 16541 12759 16575
rect 13461 16541 13495 16575
rect 14289 16541 14323 16575
rect 15301 16541 15335 16575
rect 17325 16541 17359 16575
rect 1685 16473 1719 16507
rect 3801 16473 3835 16507
rect 8677 16473 8711 16507
rect 10609 16473 10643 16507
rect 12081 16473 12115 16507
rect 13737 16473 13771 16507
rect 16681 16473 16715 16507
rect 3249 16405 3283 16439
rect 3433 16405 3467 16439
rect 5641 16405 5675 16439
rect 10885 16405 10919 16439
rect 1593 16201 1627 16235
rect 2329 16201 2363 16235
rect 2697 16201 2731 16235
rect 2881 16201 2915 16235
rect 4813 16201 4847 16235
rect 4997 16201 5031 16235
rect 8217 16201 8251 16235
rect 11069 16201 11103 16235
rect 15669 16201 15703 16235
rect 20637 16201 20671 16235
rect 21005 16201 21039 16235
rect 21373 16201 21407 16235
rect 8309 16133 8343 16167
rect 17325 16133 17359 16167
rect 3433 16065 3467 16099
rect 4261 16065 4295 16099
rect 5273 16065 5307 16099
rect 6837 16065 6871 16099
rect 8861 16065 8895 16099
rect 9597 16065 9631 16099
rect 11621 16065 11655 16099
rect 12449 16065 12483 16099
rect 19901 16065 19935 16099
rect 1409 15997 1443 16031
rect 1777 15997 1811 16031
rect 2145 15997 2179 16031
rect 2513 15997 2547 16031
rect 7104 15997 7138 16031
rect 12716 15997 12750 16031
rect 14289 15997 14323 16031
rect 14556 15997 14590 16031
rect 15945 15997 15979 16031
rect 16212 15997 16246 16031
rect 20269 15997 20303 16031
rect 20453 15997 20487 16031
rect 20821 15997 20855 16031
rect 21189 15997 21223 16031
rect 4169 15929 4203 15963
rect 4629 15929 4663 15963
rect 5540 15929 5574 15963
rect 9864 15929 9898 15963
rect 11437 15929 11471 15963
rect 11989 15929 12023 15963
rect 14105 15929 14139 15963
rect 19901 15929 19935 15963
rect 20177 15929 20211 15963
rect 1961 15861 1995 15895
rect 3249 15861 3283 15895
rect 3341 15861 3375 15895
rect 3709 15861 3743 15895
rect 4077 15861 4111 15895
rect 5181 15861 5215 15895
rect 6653 15861 6687 15895
rect 8677 15861 8711 15895
rect 8769 15861 8803 15895
rect 10977 15861 11011 15895
rect 11529 15861 11563 15895
rect 12081 15861 12115 15895
rect 13829 15861 13863 15895
rect 14013 15861 14047 15895
rect 17417 15861 17451 15895
rect 1777 15657 1811 15691
rect 3801 15657 3835 15691
rect 4445 15657 4479 15691
rect 5273 15657 5307 15691
rect 5733 15657 5767 15691
rect 6101 15657 6135 15691
rect 6469 15657 6503 15691
rect 6929 15657 6963 15691
rect 9229 15657 9263 15691
rect 11069 15657 11103 15691
rect 11437 15657 11471 15691
rect 12265 15657 12299 15691
rect 13093 15657 13127 15691
rect 13553 15657 13587 15691
rect 13921 15657 13955 15691
rect 14381 15657 14415 15691
rect 15301 15657 15335 15691
rect 16129 15657 16163 15691
rect 16497 15657 16531 15691
rect 20545 15657 20579 15691
rect 21097 15657 21131 15691
rect 21465 15657 21499 15691
rect 2145 15589 2179 15623
rect 9137 15589 9171 15623
rect 11805 15589 11839 15623
rect 13461 15589 13495 15623
rect 17233 15589 17267 15623
rect 1869 15521 1903 15555
rect 2421 15521 2455 15555
rect 2688 15521 2722 15555
rect 4813 15521 4847 15555
rect 5641 15521 5675 15555
rect 6561 15521 6595 15555
rect 7297 15521 7331 15555
rect 7757 15521 7791 15555
rect 8125 15521 8159 15555
rect 9956 15521 9990 15555
rect 12633 15521 12667 15555
rect 14289 15521 14323 15555
rect 15669 15521 15703 15555
rect 15761 15521 15795 15555
rect 18153 15521 18187 15555
rect 20913 15521 20947 15555
rect 21281 15521 21315 15555
rect 4905 15453 4939 15487
rect 4997 15453 5031 15487
rect 5917 15453 5951 15487
rect 6745 15453 6779 15487
rect 7389 15453 7423 15487
rect 7481 15453 7515 15487
rect 9321 15453 9355 15487
rect 9689 15453 9723 15487
rect 11897 15453 11931 15487
rect 12081 15453 12115 15487
rect 12725 15453 12759 15487
rect 12909 15453 12943 15487
rect 13737 15453 13771 15487
rect 14473 15453 14507 15487
rect 15945 15453 15979 15487
rect 16589 15453 16623 15487
rect 16681 15453 16715 15487
rect 18245 15453 18279 15487
rect 18337 15453 18371 15487
rect 14749 15385 14783 15419
rect 16957 15385 16991 15419
rect 20729 15385 20763 15419
rect 1593 15317 1627 15351
rect 8769 15317 8803 15351
rect 11253 15317 11287 15351
rect 17785 15317 17819 15351
rect 1961 15113 1995 15147
rect 3985 15113 4019 15147
rect 6377 15113 6411 15147
rect 9873 15113 9907 15147
rect 11529 15113 11563 15147
rect 15669 15113 15703 15147
rect 19441 15113 19475 15147
rect 21005 15113 21039 15147
rect 1777 15045 1811 15079
rect 2789 15045 2823 15079
rect 6193 15045 6227 15079
rect 8125 15045 8159 15079
rect 13829 15045 13863 15079
rect 16037 15045 16071 15079
rect 2421 14977 2455 15011
rect 2605 14977 2639 15011
rect 3433 14977 3467 15011
rect 4629 14977 4663 15011
rect 4813 14977 4847 15011
rect 7757 14977 7791 15011
rect 7941 14977 7975 15011
rect 10609 14977 10643 15011
rect 12173 14977 12207 15011
rect 13921 14977 13955 15011
rect 15393 14977 15427 15011
rect 18061 14977 18095 15011
rect 20177 14977 20211 15011
rect 1593 14909 1627 14943
rect 4353 14909 4387 14943
rect 5080 14909 5114 14943
rect 8309 14909 8343 14943
rect 8493 14909 8527 14943
rect 10425 14909 10459 14943
rect 11253 14909 11287 14943
rect 11897 14909 11931 14943
rect 12449 14909 12483 14943
rect 15853 14909 15887 14943
rect 16313 14909 16347 14943
rect 16580 14909 16614 14943
rect 19901 14909 19935 14943
rect 20821 14909 20855 14943
rect 1501 14841 1535 14875
rect 7205 14841 7239 14875
rect 7665 14841 7699 14875
rect 8760 14841 8794 14875
rect 11437 14841 11471 14875
rect 12716 14841 12750 14875
rect 15209 14841 15243 14875
rect 18328 14841 18362 14875
rect 2329 14773 2363 14807
rect 3157 14773 3191 14807
rect 3249 14773 3283 14807
rect 3617 14773 3651 14807
rect 4445 14773 4479 14807
rect 6837 14773 6871 14807
rect 7297 14773 7331 14807
rect 10057 14773 10091 14807
rect 10517 14773 10551 14807
rect 10885 14773 10919 14807
rect 11989 14773 12023 14807
rect 14841 14773 14875 14807
rect 15301 14773 15335 14807
rect 17693 14773 17727 14807
rect 19533 14773 19567 14807
rect 21189 14773 21223 14807
rect 1869 14569 1903 14603
rect 2697 14569 2731 14603
rect 3157 14569 3191 14603
rect 3801 14569 3835 14603
rect 4077 14569 4111 14603
rect 4905 14569 4939 14603
rect 6561 14569 6595 14603
rect 6745 14569 6779 14603
rect 7113 14569 7147 14603
rect 9873 14569 9907 14603
rect 10241 14569 10275 14603
rect 10701 14569 10735 14603
rect 11069 14569 11103 14603
rect 11529 14569 11563 14603
rect 12265 14569 12299 14603
rect 12541 14569 12575 14603
rect 19349 14569 19383 14603
rect 20453 14569 20487 14603
rect 21097 14569 21131 14603
rect 21465 14569 21499 14603
rect 5917 14501 5951 14535
rect 6469 14501 6503 14535
rect 10609 14501 10643 14535
rect 13912 14501 13946 14535
rect 15568 14501 15602 14535
rect 19441 14501 19475 14535
rect 20177 14501 20211 14535
rect 1685 14433 1719 14467
rect 2053 14433 2087 14467
rect 3617 14433 3651 14467
rect 4445 14433 4479 14467
rect 4537 14433 4571 14467
rect 7573 14433 7607 14467
rect 7840 14433 7874 14467
rect 9229 14433 9263 14467
rect 11437 14433 11471 14467
rect 12449 14433 12483 14467
rect 12909 14433 12943 14467
rect 13645 14433 13679 14467
rect 15301 14433 15335 14467
rect 17776 14433 17810 14467
rect 19901 14433 19935 14467
rect 20913 14433 20947 14467
rect 21281 14433 21315 14467
rect 2329 14365 2363 14399
rect 3249 14365 3283 14399
rect 3433 14365 3467 14399
rect 4721 14365 4755 14399
rect 6009 14365 6043 14399
rect 6193 14365 6227 14399
rect 7205 14365 7239 14399
rect 7389 14365 7423 14399
rect 9965 14365 9999 14399
rect 10885 14365 10919 14399
rect 11621 14365 11655 14399
rect 13001 14365 13035 14399
rect 13093 14365 13127 14399
rect 17509 14365 17543 14399
rect 19533 14365 19567 14399
rect 2789 14297 2823 14331
rect 8953 14297 8987 14331
rect 11989 14297 12023 14331
rect 13369 14297 13403 14331
rect 18889 14297 18923 14331
rect 1501 14229 1535 14263
rect 5181 14229 5215 14263
rect 5549 14229 5583 14263
rect 9137 14229 9171 14263
rect 12081 14229 12115 14263
rect 15025 14229 15059 14263
rect 16681 14229 16715 14263
rect 18981 14229 19015 14263
rect 20729 14229 20763 14263
rect 1777 14025 1811 14059
rect 5825 14025 5859 14059
rect 7665 14025 7699 14059
rect 9689 14025 9723 14059
rect 12725 14025 12759 14059
rect 15853 14025 15887 14059
rect 17141 14025 17175 14059
rect 17601 14025 17635 14059
rect 18061 14025 18095 14059
rect 18889 14025 18923 14059
rect 21005 14025 21039 14059
rect 3985 13957 4019 13991
rect 8861 13957 8895 13991
rect 10517 13957 10551 13991
rect 11437 13957 11471 13991
rect 14933 13957 14967 13991
rect 21373 13957 21407 13991
rect 2237 13889 2271 13923
rect 6469 13889 6503 13923
rect 7389 13889 7423 13923
rect 8217 13889 8251 13923
rect 9505 13889 9539 13923
rect 10149 13889 10183 13923
rect 10333 13889 10367 13923
rect 11069 13889 11103 13923
rect 13369 13889 13403 13923
rect 15577 13889 15611 13923
rect 16405 13889 16439 13923
rect 18613 13889 18647 13923
rect 19441 13889 19475 13923
rect 1501 13821 1535 13855
rect 1593 13821 1627 13855
rect 1961 13821 1995 13855
rect 2605 13821 2639 13855
rect 4445 13821 4479 13855
rect 7297 13821 7331 13855
rect 8125 13821 8159 13855
rect 8769 13821 8803 13855
rect 9321 13821 9355 13855
rect 10885 13821 10919 13855
rect 10977 13821 11011 13855
rect 13553 13821 13587 13855
rect 16221 13821 16255 13855
rect 16957 13821 16991 13855
rect 18429 13821 18463 13855
rect 19257 13821 19291 13855
rect 20269 13821 20303 13855
rect 20545 13821 20579 13855
rect 20821 13821 20855 13855
rect 21281 13821 21315 13855
rect 2872 13753 2906 13787
rect 4690 13753 4724 13787
rect 7205 13753 7239 13787
rect 11621 13753 11655 13787
rect 13093 13753 13127 13787
rect 13820 13753 13854 13787
rect 17785 13753 17819 13787
rect 19349 13753 19383 13787
rect 5917 13685 5951 13719
rect 6285 13685 6319 13719
rect 6377 13685 6411 13719
rect 6837 13685 6871 13719
rect 8033 13685 8067 13719
rect 8585 13685 8619 13719
rect 9229 13685 9263 13719
rect 10057 13685 10091 13719
rect 12449 13685 12483 13719
rect 13185 13685 13219 13719
rect 15025 13685 15059 13719
rect 15393 13685 15427 13719
rect 15485 13685 15519 13719
rect 16313 13685 16347 13719
rect 16681 13685 16715 13719
rect 18521 13685 18555 13719
rect 2421 13481 2455 13515
rect 2789 13481 2823 13515
rect 3157 13481 3191 13515
rect 5457 13481 5491 13515
rect 6101 13481 6135 13515
rect 6469 13481 6503 13515
rect 8401 13481 8435 13515
rect 9505 13481 9539 13515
rect 9689 13481 9723 13515
rect 10057 13481 10091 13515
rect 13553 13481 13587 13515
rect 13921 13481 13955 13515
rect 14381 13481 14415 13515
rect 14749 13481 14783 13515
rect 15301 13481 15335 13515
rect 16129 13481 16163 13515
rect 16497 13481 16531 13515
rect 17049 13481 17083 13515
rect 17509 13481 17543 13515
rect 17877 13481 17911 13515
rect 21097 13481 21131 13515
rect 7174 13413 7208 13447
rect 10149 13413 10183 13447
rect 10609 13413 10643 13447
rect 11069 13413 11103 13447
rect 14013 13413 14047 13447
rect 15669 13413 15703 13447
rect 16589 13413 16623 13447
rect 1685 13345 1719 13379
rect 2237 13345 2271 13379
rect 2605 13345 2639 13379
rect 3525 13345 3559 13379
rect 4344 13345 4378 13379
rect 5733 13345 5767 13379
rect 6009 13345 6043 13379
rect 6929 13345 6963 13379
rect 8769 13345 8803 13379
rect 11161 13345 11195 13379
rect 11529 13345 11563 13379
rect 11796 13345 11830 13379
rect 17417 13345 17451 13379
rect 18245 13345 18279 13379
rect 20913 13345 20947 13379
rect 21281 13345 21315 13379
rect 1869 13277 1903 13311
rect 3617 13277 3651 13311
rect 3709 13277 3743 13311
rect 4077 13277 4111 13311
rect 6561 13277 6595 13311
rect 6745 13277 6779 13311
rect 8861 13277 8895 13311
rect 8953 13277 8987 13311
rect 10333 13277 10367 13311
rect 11253 13277 11287 13311
rect 14197 13277 14231 13311
rect 14841 13277 14875 13311
rect 14933 13277 14967 13311
rect 15761 13277 15795 13311
rect 15945 13277 15979 13311
rect 16681 13277 16715 13311
rect 17601 13277 17635 13311
rect 18337 13277 18371 13311
rect 18521 13277 18555 13311
rect 3065 13209 3099 13243
rect 5549 13141 5583 13175
rect 8309 13141 8343 13175
rect 9321 13141 9355 13175
rect 10701 13141 10735 13175
rect 12909 13141 12943 13175
rect 19441 13141 19475 13175
rect 3249 12937 3283 12971
rect 3801 12937 3835 12971
rect 4813 12937 4847 12971
rect 5917 12937 5951 12971
rect 6837 12937 6871 12971
rect 11805 12937 11839 12971
rect 14381 12937 14415 12971
rect 14657 12937 14691 12971
rect 14933 12937 14967 12971
rect 16037 12937 16071 12971
rect 17141 12937 17175 12971
rect 19533 12937 19567 12971
rect 21005 12937 21039 12971
rect 13277 12869 13311 12903
rect 14105 12869 14139 12903
rect 19441 12869 19475 12903
rect 4353 12801 4387 12835
rect 5365 12801 5399 12835
rect 6561 12801 6595 12835
rect 7389 12801 7423 12835
rect 8401 12801 8435 12835
rect 9045 12801 9079 12835
rect 9137 12801 9171 12835
rect 10241 12801 10275 12835
rect 13001 12801 13035 12835
rect 13829 12801 13863 12835
rect 15577 12801 15611 12835
rect 16589 12801 16623 12835
rect 17785 12801 17819 12835
rect 20085 12801 20119 12835
rect 1869 12733 1903 12767
rect 7205 12733 7239 12767
rect 8953 12733 8987 12767
rect 9965 12733 9999 12767
rect 10425 12733 10459 12767
rect 13737 12733 13771 12767
rect 14289 12733 14323 12767
rect 16497 12733 16531 12767
rect 16865 12733 16899 12767
rect 18061 12733 18095 12767
rect 19901 12733 19935 12767
rect 20821 12733 20855 12767
rect 2136 12665 2170 12699
rect 3709 12665 3743 12699
rect 4261 12665 4295 12699
rect 5273 12665 5307 12699
rect 6377 12665 6411 12699
rect 8125 12665 8159 12699
rect 10692 12665 10726 12699
rect 12173 12665 12207 12699
rect 13645 12665 13679 12699
rect 14749 12665 14783 12699
rect 15301 12665 15335 12699
rect 15393 12665 15427 12699
rect 16405 12665 16439 12699
rect 17601 12665 17635 12699
rect 18328 12665 18362 12699
rect 19993 12665 20027 12699
rect 4169 12597 4203 12631
rect 5181 12597 5215 12631
rect 5733 12597 5767 12631
rect 6285 12597 6319 12631
rect 7297 12597 7331 12631
rect 7757 12597 7791 12631
rect 8217 12597 8251 12631
rect 8585 12597 8619 12631
rect 9413 12597 9447 12631
rect 9597 12597 9631 12631
rect 10057 12597 10091 12631
rect 11897 12597 11931 12631
rect 12449 12597 12483 12631
rect 12817 12597 12851 12631
rect 12909 12597 12943 12631
rect 15853 12597 15887 12631
rect 17509 12597 17543 12631
rect 1685 12393 1719 12427
rect 1869 12393 1903 12427
rect 2329 12393 2363 12427
rect 2789 12393 2823 12427
rect 4077 12393 4111 12427
rect 4537 12393 4571 12427
rect 4997 12393 5031 12427
rect 5457 12393 5491 12427
rect 7297 12393 7331 12427
rect 9413 12393 9447 12427
rect 10149 12393 10183 12427
rect 11437 12393 11471 12427
rect 11805 12393 11839 12427
rect 12173 12393 12207 12427
rect 16773 12393 16807 12427
rect 16957 12393 16991 12427
rect 17233 12393 17267 12427
rect 18797 12393 18831 12427
rect 19257 12393 19291 12427
rect 8300 12325 8334 12359
rect 9873 12325 9907 12359
rect 12970 12325 13004 12359
rect 15546 12325 15580 12359
rect 20269 12325 20303 12359
rect 1501 12257 1535 12291
rect 2237 12257 2271 12291
rect 3157 12257 3191 12291
rect 4905 12257 4939 12291
rect 6092 12257 6126 12291
rect 7481 12257 7515 12291
rect 7941 12257 7975 12291
rect 9689 12257 9723 12291
rect 10517 12257 10551 12291
rect 11345 12257 11379 12291
rect 12725 12257 12759 12291
rect 17325 12257 17359 12291
rect 17592 12257 17626 12291
rect 19165 12257 19199 12291
rect 19993 12257 20027 12291
rect 2513 12189 2547 12223
rect 3249 12189 3283 12223
rect 3341 12189 3375 12223
rect 5089 12189 5123 12223
rect 5825 12189 5859 12223
rect 8033 12189 8067 12223
rect 10609 12189 10643 12223
rect 10793 12189 10827 12223
rect 11529 12189 11563 12223
rect 12265 12189 12299 12223
rect 12449 12189 12483 12223
rect 14197 12189 14231 12223
rect 15301 12189 15335 12223
rect 19349 12189 19383 12223
rect 18705 12121 18739 12155
rect 4353 12053 4387 12087
rect 5641 12053 5675 12087
rect 7205 12053 7239 12087
rect 7757 12053 7791 12087
rect 9689 12053 9723 12087
rect 9965 12053 9999 12087
rect 10977 12053 11011 12087
rect 14105 12053 14139 12087
rect 14841 12053 14875 12087
rect 15025 12053 15059 12087
rect 16681 12053 16715 12087
rect 19717 12053 19751 12087
rect 22017 11985 22051 12019
rect 2881 11849 2915 11883
rect 3157 11849 3191 11883
rect 3433 11849 3467 11883
rect 4261 11849 4295 11883
rect 6929 11849 6963 11883
rect 7113 11849 7147 11883
rect 8769 11849 8803 11883
rect 10149 11849 10183 11883
rect 12449 11849 12483 11883
rect 15393 11849 15427 11883
rect 17601 11849 17635 11883
rect 18153 11849 18187 11883
rect 21005 11849 21039 11883
rect 21373 11849 21407 11883
rect 11713 11781 11747 11815
rect 18981 11781 19015 11815
rect 1501 11713 1535 11747
rect 4077 11713 4111 11747
rect 4813 11713 4847 11747
rect 7573 11713 7607 11747
rect 7665 11713 7699 11747
rect 8493 11713 8527 11747
rect 9413 11713 9447 11747
rect 9965 11713 9999 11747
rect 10333 11713 10367 11747
rect 12909 11713 12943 11747
rect 13001 11713 13035 11747
rect 16037 11713 16071 11747
rect 18705 11713 18739 11747
rect 2973 11645 3007 11679
rect 5273 11645 5307 11679
rect 5540 11645 5574 11679
rect 8401 11645 8435 11679
rect 9137 11645 9171 11679
rect 9229 11645 9263 11679
rect 13277 11645 13311 11679
rect 13461 11645 13495 11679
rect 16221 11645 16255 11679
rect 20821 11645 20855 11679
rect 21189 11645 21223 11679
rect 1768 11577 1802 11611
rect 10600 11577 10634 11611
rect 11805 11577 11839 11611
rect 12173 11577 12207 11611
rect 13728 11577 13762 11611
rect 16488 11577 16522 11611
rect 18613 11577 18647 11611
rect 19165 11577 19199 11611
rect 3801 11509 3835 11543
rect 3893 11509 3927 11543
rect 4629 11509 4663 11543
rect 4721 11509 4755 11543
rect 5089 11509 5123 11543
rect 6653 11509 6687 11543
rect 7481 11509 7515 11543
rect 7941 11509 7975 11543
rect 8309 11509 8343 11543
rect 9689 11509 9723 11543
rect 9781 11509 9815 11543
rect 12817 11509 12851 11543
rect 14841 11509 14875 11543
rect 15025 11509 15059 11543
rect 15761 11509 15795 11543
rect 15853 11509 15887 11543
rect 17785 11509 17819 11543
rect 18521 11509 18555 11543
rect 1593 11305 1627 11339
rect 3157 11305 3191 11339
rect 4169 11305 4203 11339
rect 4997 11305 5031 11339
rect 6561 11305 6595 11339
rect 7389 11305 7423 11339
rect 7941 11305 7975 11339
rect 8401 11305 8435 11339
rect 12265 11305 12299 11339
rect 13093 11305 13127 11339
rect 14381 11305 14415 11339
rect 15669 11305 15703 11339
rect 16129 11305 16163 11339
rect 17417 11305 17451 11339
rect 17877 11305 17911 11339
rect 19073 11305 19107 11339
rect 21097 11305 21131 11339
rect 22017 11305 22051 11339
rect 5641 11237 5675 11271
rect 6929 11237 6963 11271
rect 10425 11237 10459 11271
rect 12725 11237 12759 11271
rect 13461 11237 13495 11271
rect 13921 11237 13955 11271
rect 14841 11237 14875 11271
rect 17785 11237 17819 11271
rect 18337 11237 18371 11271
rect 1409 11169 1443 11203
rect 1777 11169 1811 11203
rect 2044 11169 2078 11203
rect 4537 11169 4571 11203
rect 4629 11169 4663 11203
rect 6469 11169 6503 11203
rect 7297 11169 7331 11203
rect 8309 11169 8343 11203
rect 8953 11169 8987 11203
rect 9781 11169 9815 11203
rect 12633 11169 12667 11203
rect 13277 11169 13311 11203
rect 14749 11169 14783 11203
rect 16497 11169 16531 11203
rect 17325 11169 17359 11203
rect 3801 11101 3835 11135
rect 4813 11101 4847 11135
rect 5733 11101 5767 11135
rect 5917 11101 5951 11135
rect 6653 11101 6687 11135
rect 7573 11101 7607 11135
rect 8585 11101 8619 11135
rect 9505 11101 9539 11135
rect 12817 11101 12851 11135
rect 14013 11101 14047 11135
rect 14197 11101 14231 11135
rect 14933 11101 14967 11135
rect 15761 11101 15795 11135
rect 15945 11101 15979 11135
rect 16589 11101 16623 11135
rect 16773 11101 16807 11135
rect 17601 11101 17635 11135
rect 18245 11169 18279 11203
rect 20913 11169 20947 11203
rect 18521 11101 18555 11135
rect 19165 11101 19199 11135
rect 19257 11101 19291 11135
rect 3709 11033 3743 11067
rect 5273 11033 5307 11067
rect 8769 11033 8803 11067
rect 11713 11033 11747 11067
rect 13553 11033 13587 11067
rect 15301 11033 15335 11067
rect 16957 11033 16991 11067
rect 17785 11033 17819 11067
rect 18705 11033 18739 11067
rect 6101 10965 6135 10999
rect 7849 10965 7883 10999
rect 9045 10965 9079 10999
rect 9229 10965 9263 10999
rect 1501 10761 1535 10795
rect 3709 10761 3743 10795
rect 3893 10761 3927 10795
rect 4721 10761 4755 10795
rect 5733 10761 5767 10795
rect 8309 10761 8343 10795
rect 11345 10761 11379 10795
rect 11437 10761 11471 10795
rect 13921 10761 13955 10795
rect 15117 10761 15151 10795
rect 17785 10761 17819 10795
rect 8217 10693 8251 10727
rect 14841 10693 14875 10727
rect 18061 10693 18095 10727
rect 19349 10693 19383 10727
rect 2145 10625 2179 10659
rect 4353 10625 4387 10659
rect 4537 10625 4571 10659
rect 5365 10625 5399 10659
rect 5641 10625 5675 10659
rect 6193 10625 6227 10659
rect 6377 10625 6411 10659
rect 8861 10625 8895 10659
rect 9689 10625 9723 10659
rect 9965 10625 9999 10659
rect 11989 10625 12023 10659
rect 14565 10625 14599 10659
rect 15761 10625 15795 10659
rect 18521 10625 18555 10659
rect 18705 10625 18739 10659
rect 18889 10625 18923 10659
rect 19901 10625 19935 10659
rect 20453 10625 20487 10659
rect 21005 10625 21039 10659
rect 2329 10557 2363 10591
rect 4261 10557 4295 10591
rect 6837 10557 6871 10591
rect 8769 10557 8803 10591
rect 10221 10557 10255 10591
rect 11897 10557 11931 10591
rect 12541 10557 12575 10591
rect 15485 10557 15519 10591
rect 15945 10557 15979 10591
rect 16212 10557 16246 10591
rect 17509 10557 17543 10591
rect 18429 10557 18463 10591
rect 19165 10557 19199 10591
rect 20177 10557 20211 10591
rect 20729 10557 20763 10591
rect 2596 10489 2630 10523
rect 5181 10489 5215 10523
rect 6101 10489 6135 10523
rect 7082 10489 7116 10523
rect 8677 10489 8711 10523
rect 9505 10489 9539 10523
rect 11805 10489 11839 10523
rect 12808 10489 12842 10523
rect 14381 10489 14415 10523
rect 1869 10421 1903 10455
rect 1961 10421 1995 10455
rect 5089 10421 5123 10455
rect 6561 10421 6595 10455
rect 9137 10421 9171 10455
rect 9597 10421 9631 10455
rect 14013 10421 14047 10455
rect 14473 10421 14507 10455
rect 15577 10421 15611 10455
rect 17325 10421 17359 10455
rect 19717 10421 19751 10455
rect 19809 10421 19843 10455
rect 2053 10217 2087 10251
rect 3157 10217 3191 10251
rect 4353 10217 4387 10251
rect 5273 10217 5307 10251
rect 6101 10217 6135 10251
rect 6745 10217 6779 10251
rect 7113 10217 7147 10251
rect 11345 10217 11379 10251
rect 11805 10217 11839 10251
rect 11897 10217 11931 10251
rect 13645 10217 13679 10251
rect 13921 10217 13955 10251
rect 14289 10217 14323 10251
rect 14657 10217 14691 10251
rect 15301 10217 15335 10251
rect 16129 10217 16163 10251
rect 16497 10217 16531 10251
rect 18797 10217 18831 10251
rect 20637 10217 20671 10251
rect 4261 10149 4295 10183
rect 4721 10149 4755 10183
rect 6653 10149 6687 10183
rect 9137 10149 9171 10183
rect 9934 10149 9968 10183
rect 14749 10149 14783 10183
rect 15761 10149 15795 10183
rect 17141 10149 17175 10183
rect 17325 10149 17359 10183
rect 17662 10149 17696 10183
rect 2421 10081 2455 10115
rect 5641 10081 5675 10115
rect 5733 10081 5767 10115
rect 7481 10081 7515 10115
rect 7573 10081 7607 10115
rect 8309 10081 8343 10115
rect 12265 10081 12299 10115
rect 12532 10081 12566 10115
rect 15669 10081 15703 10115
rect 16589 10081 16623 10115
rect 2513 10013 2547 10047
rect 2697 10013 2731 10047
rect 4813 10013 4847 10047
rect 4997 10013 5031 10047
rect 5917 10013 5951 10047
rect 6837 10013 6871 10047
rect 7757 10013 7791 10047
rect 8401 10013 8435 10047
rect 8585 10013 8619 10047
rect 9229 10013 9263 10047
rect 9413 10013 9447 10047
rect 9689 10013 9723 10047
rect 12081 10013 12115 10047
rect 13737 10013 13771 10047
rect 14933 10013 14967 10047
rect 15853 10013 15887 10047
rect 16773 10013 16807 10047
rect 19524 10081 19558 10115
rect 17417 10013 17451 10047
rect 18889 10013 18923 10047
rect 19257 10013 19291 10047
rect 2973 9945 3007 9979
rect 8769 9945 8803 9979
rect 14197 9945 14231 9979
rect 17325 9945 17359 9979
rect 3249 9877 3283 9911
rect 6285 9877 6319 9911
rect 7941 9877 7975 9911
rect 11069 9877 11103 9911
rect 11437 9877 11471 9911
rect 16957 9877 16991 9911
rect 19165 9877 19199 9911
rect 1593 9673 1627 9707
rect 2421 9673 2455 9707
rect 4261 9673 4295 9707
rect 10149 9673 10183 9707
rect 12265 9673 12299 9707
rect 12541 9673 12575 9707
rect 14657 9673 14691 9707
rect 17509 9673 17543 9707
rect 20453 9673 20487 9707
rect 3249 9605 3283 9639
rect 4169 9605 4203 9639
rect 5089 9605 5123 9639
rect 14197 9605 14231 9639
rect 14841 9605 14875 9639
rect 15669 9605 15703 9639
rect 20361 9605 20395 9639
rect 2053 9537 2087 9571
rect 2237 9537 2271 9571
rect 3065 9537 3099 9571
rect 3893 9537 3927 9571
rect 4813 9537 4847 9571
rect 5641 9537 5675 9571
rect 6561 9537 6595 9571
rect 8769 9537 8803 9571
rect 10241 9537 10275 9571
rect 13185 9537 13219 9571
rect 14013 9537 14047 9571
rect 15301 9537 15335 9571
rect 15485 9537 15519 9571
rect 16313 9537 16347 9571
rect 17049 9537 17083 9571
rect 18797 9537 18831 9571
rect 21005 9537 21039 9571
rect 3709 9469 3743 9503
rect 7021 9469 7055 9503
rect 7277 9469 7311 9503
rect 9036 9469 9070 9503
rect 10885 9469 10919 9503
rect 11152 9469 11186 9503
rect 13001 9469 13035 9503
rect 13737 9469 13771 9503
rect 14381 9469 14415 9503
rect 18981 9469 19015 9503
rect 19248 9469 19282 9503
rect 2881 9401 2915 9435
rect 13829 9401 13863 9435
rect 14473 9401 14507 9435
rect 15209 9401 15243 9435
rect 17693 9401 17727 9435
rect 1409 9333 1443 9367
rect 1961 9333 1995 9367
rect 2789 9333 2823 9367
rect 3617 9333 3651 9367
rect 4629 9333 4663 9367
rect 4721 9333 4755 9367
rect 5457 9333 5491 9367
rect 5549 9333 5583 9367
rect 5917 9333 5951 9367
rect 6285 9333 6319 9367
rect 6377 9333 6411 9367
rect 6929 9333 6963 9367
rect 8401 9333 8435 9367
rect 8585 9333 8619 9367
rect 12909 9333 12943 9367
rect 13369 9333 13403 9367
rect 16037 9333 16071 9367
rect 16129 9333 16163 9367
rect 16497 9333 16531 9367
rect 16865 9333 16899 9367
rect 16957 9333 16991 9367
rect 17417 9333 17451 9367
rect 18153 9333 18187 9367
rect 18521 9333 18555 9367
rect 18613 9333 18647 9367
rect 20821 9333 20855 9367
rect 20913 9333 20947 9367
rect 1593 9129 1627 9163
rect 2421 9129 2455 9163
rect 2881 9129 2915 9163
rect 5457 9129 5491 9163
rect 7849 9129 7883 9163
rect 8309 9129 8343 9163
rect 8401 9129 8435 9163
rect 8769 9129 8803 9163
rect 9137 9129 9171 9163
rect 9689 9129 9723 9163
rect 13185 9129 13219 9163
rect 13553 9129 13587 9163
rect 15301 9129 15335 9163
rect 17141 9129 17175 9163
rect 17601 9129 17635 9163
rect 17969 9129 18003 9163
rect 20177 9129 20211 9163
rect 1961 9061 1995 9095
rect 3249 9061 3283 9095
rect 4333 9061 4367 9095
rect 1409 8993 1443 9027
rect 2789 8993 2823 9027
rect 4077 8993 4111 9027
rect 5733 8993 5767 9027
rect 6000 8993 6034 9027
rect 7389 8993 7423 9027
rect 7757 8993 7791 9027
rect 2053 8925 2087 8959
rect 2237 8925 2271 8959
rect 3065 8925 3099 8959
rect 10701 9061 10735 9095
rect 11253 9061 11287 9095
rect 13093 9061 13127 9095
rect 14289 9061 14323 9095
rect 14657 9061 14691 9095
rect 17509 9061 17543 9095
rect 18337 9061 18371 9095
rect 9229 8993 9263 9027
rect 10057 8993 10091 9027
rect 13645 8993 13679 9027
rect 15485 8993 15519 9027
rect 15669 8993 15703 9027
rect 15936 8993 15970 9027
rect 19064 8993 19098 9027
rect 8585 8925 8619 8959
rect 9413 8925 9447 8959
rect 10149 8925 10183 8959
rect 10241 8925 10275 8959
rect 11345 8925 11379 8959
rect 11529 8925 11563 8959
rect 13737 8925 13771 8959
rect 14933 8925 14967 8959
rect 17693 8925 17727 8959
rect 18429 8925 18463 8959
rect 18613 8925 18647 8959
rect 18797 8925 18831 8959
rect 7205 8857 7239 8891
rect 7573 8857 7607 8891
rect 7849 8857 7883 8891
rect 10517 8857 10551 8891
rect 14841 8857 14875 8891
rect 3617 8789 3651 8823
rect 5641 8789 5675 8823
rect 7113 8789 7147 8823
rect 7941 8789 7975 8823
rect 10885 8789 10919 8823
rect 14197 8789 14231 8823
rect 17049 8789 17083 8823
rect 20361 8789 20395 8823
rect 4261 8585 4295 8619
rect 6193 8585 6227 8619
rect 7205 8585 7239 8619
rect 9965 8585 9999 8619
rect 12449 8585 12483 8619
rect 13277 8585 13311 8619
rect 16589 8585 16623 8619
rect 18889 8585 18923 8619
rect 19717 8585 19751 8619
rect 1961 8517 1995 8551
rect 9873 8517 9907 8551
rect 1685 8449 1719 8483
rect 2605 8449 2639 8483
rect 7849 8449 7883 8483
rect 8033 8449 8067 8483
rect 8493 8449 8527 8483
rect 10517 8449 10551 8483
rect 10793 8449 10827 8483
rect 10885 8449 10919 8483
rect 13093 8449 13127 8483
rect 1409 8381 1443 8415
rect 2421 8381 2455 8415
rect 2881 8381 2915 8415
rect 4813 8381 4847 8415
rect 7021 8381 7055 8415
rect 10425 8381 10459 8415
rect 11141 8381 11175 8415
rect 12817 8381 12851 8415
rect 2329 8313 2363 8347
rect 3126 8313 3160 8347
rect 5080 8313 5114 8347
rect 8760 8313 8794 8347
rect 10333 8313 10367 8347
rect 10793 8313 10827 8347
rect 20545 8517 20579 8551
rect 13553 8449 13587 8483
rect 15209 8449 15243 8483
rect 17233 8449 17267 8483
rect 18613 8449 18647 8483
rect 19441 8449 19475 8483
rect 20269 8449 20303 8483
rect 21097 8449 21131 8483
rect 13737 8381 13771 8415
rect 14004 8381 14038 8415
rect 17141 8381 17175 8415
rect 17785 8381 17819 8415
rect 18521 8381 18555 8415
rect 20177 8381 20211 8415
rect 15476 8313 15510 8347
rect 17049 8313 17083 8347
rect 17509 8313 17543 8347
rect 18429 8313 18463 8347
rect 19257 8313 19291 8347
rect 6285 8245 6319 8279
rect 6837 8245 6871 8279
rect 7389 8245 7423 8279
rect 7757 8245 7791 8279
rect 8309 8245 8343 8279
rect 12265 8245 12299 8279
rect 12909 8245 12943 8279
rect 13277 8245 13311 8279
rect 13461 8245 13495 8279
rect 15117 8245 15151 8279
rect 16681 8245 16715 8279
rect 18061 8245 18095 8279
rect 19349 8245 19383 8279
rect 20085 8245 20119 8279
rect 20913 8245 20947 8279
rect 21005 8245 21039 8279
rect 21465 8245 21499 8279
rect 1501 8041 1535 8075
rect 3525 8041 3559 8075
rect 5089 8041 5123 8075
rect 5457 8041 5491 8075
rect 6745 8041 6779 8075
rect 7113 8041 7147 8075
rect 7941 8041 7975 8075
rect 8401 8041 8435 8075
rect 8769 8041 8803 8075
rect 9229 8041 9263 8075
rect 10149 8041 10183 8075
rect 12449 8041 12483 8075
rect 12725 8041 12759 8075
rect 13185 8041 13219 8075
rect 13553 8041 13587 8075
rect 14381 8041 14415 8075
rect 14749 8041 14783 8075
rect 16589 8041 16623 8075
rect 17141 8041 17175 8075
rect 19441 8041 19475 8075
rect 19993 8041 20027 8075
rect 20361 8041 20395 8075
rect 21097 8041 21131 8075
rect 7205 7973 7239 8007
rect 9137 7973 9171 8007
rect 10609 7973 10643 8007
rect 13093 7973 13127 8007
rect 14841 7973 14875 8007
rect 16681 7973 16715 8007
rect 17509 7973 17543 8007
rect 1952 7905 1986 7939
rect 6285 7905 6319 7939
rect 6377 7905 6411 7939
rect 7849 7905 7883 7939
rect 8309 7905 8343 7939
rect 10517 7905 10551 7939
rect 11244 7905 11278 7939
rect 12633 7905 12667 7939
rect 13921 7905 13955 7939
rect 15669 7905 15703 7939
rect 17969 7905 18003 7939
rect 18236 7905 18270 7939
rect 21005 7905 21039 7939
rect 1685 7837 1719 7871
rect 3617 7837 3651 7871
rect 3709 7837 3743 7871
rect 5549 7837 5583 7871
rect 5733 7837 5767 7871
rect 6561 7837 6595 7871
rect 7297 7837 7331 7871
rect 8585 7837 8619 7871
rect 9413 7837 9447 7871
rect 10793 7837 10827 7871
rect 10977 7837 11011 7871
rect 13369 7837 13403 7871
rect 14013 7837 14047 7871
rect 14105 7837 14139 7871
rect 14933 7837 14967 7871
rect 15761 7837 15795 7871
rect 15945 7837 15979 7871
rect 16773 7837 16807 7871
rect 17601 7837 17635 7871
rect 17693 7837 17727 7871
rect 20453 7837 20487 7871
rect 20637 7837 20671 7871
rect 3065 7769 3099 7803
rect 5917 7769 5951 7803
rect 7665 7769 7699 7803
rect 9965 7769 9999 7803
rect 16221 7769 16255 7803
rect 19625 7769 19659 7803
rect 21465 7769 21499 7803
rect 3157 7701 3191 7735
rect 4721 7701 4755 7735
rect 4997 7701 5031 7735
rect 9781 7701 9815 7735
rect 12357 7701 12391 7735
rect 15301 7701 15335 7735
rect 19349 7701 19383 7735
rect 3709 7497 3743 7531
rect 5825 7497 5859 7531
rect 9137 7497 9171 7531
rect 10701 7497 10735 7531
rect 10885 7497 10919 7531
rect 11713 7497 11747 7531
rect 15025 7497 15059 7531
rect 17141 7497 17175 7531
rect 17693 7497 17727 7531
rect 18061 7497 18095 7531
rect 20361 7497 20395 7531
rect 6653 7429 6687 7463
rect 6837 7429 6871 7463
rect 9045 7429 9079 7463
rect 4169 7361 4203 7395
rect 4261 7361 4295 7395
rect 5549 7361 5583 7395
rect 6377 7361 6411 7395
rect 1869 7293 1903 7327
rect 4721 7293 4755 7327
rect 5365 7293 5399 7327
rect 6285 7293 6319 7327
rect 7389 7361 7423 7395
rect 9689 7361 9723 7395
rect 10241 7361 10275 7395
rect 11529 7361 11563 7395
rect 7205 7293 7239 7327
rect 7665 7293 7699 7327
rect 9597 7293 9631 7327
rect 10609 7293 10643 7327
rect 12173 7429 12207 7463
rect 12449 7429 12483 7463
rect 15209 7429 15243 7463
rect 16037 7429 16071 7463
rect 13093 7361 13127 7395
rect 13737 7361 13771 7395
rect 13921 7361 13955 7395
rect 14657 7361 14691 7395
rect 15669 7361 15703 7395
rect 15853 7361 15887 7395
rect 16589 7361 16623 7395
rect 16865 7361 16899 7395
rect 18613 7361 18647 7395
rect 20177 7361 20211 7395
rect 20913 7361 20947 7395
rect 18521 7293 18555 7327
rect 18981 7293 19015 7327
rect 19901 7293 19935 7327
rect 2136 7225 2170 7259
rect 4077 7225 4111 7259
rect 4905 7225 4939 7259
rect 6193 7225 6227 7259
rect 6653 7225 6687 7259
rect 7910 7225 7944 7259
rect 9505 7225 9539 7259
rect 10425 7225 10459 7259
rect 11345 7225 11379 7259
rect 11713 7225 11747 7259
rect 14565 7225 14599 7259
rect 15577 7225 15611 7259
rect 17877 7225 17911 7259
rect 18429 7225 18463 7259
rect 19257 7225 19291 7259
rect 21373 7225 21407 7259
rect 3249 7157 3283 7191
rect 4997 7157 5031 7191
rect 5457 7157 5491 7191
rect 7297 7157 7331 7191
rect 9965 7157 9999 7191
rect 11253 7157 11287 7191
rect 11805 7157 11839 7191
rect 12081 7157 12115 7191
rect 12817 7157 12851 7191
rect 12909 7157 12943 7191
rect 13277 7157 13311 7191
rect 13645 7157 13679 7191
rect 14105 7157 14139 7191
rect 14473 7157 14507 7191
rect 16405 7157 16439 7191
rect 16497 7157 16531 7191
rect 19533 7157 19567 7191
rect 19993 7157 20027 7191
rect 20729 7157 20763 7191
rect 20821 7157 20855 7191
rect 21189 7157 21223 7191
rect 7021 6953 7055 6987
rect 10333 6953 10367 6987
rect 11529 6953 11563 6987
rect 14565 6953 14599 6987
rect 15025 6953 15059 6987
rect 15393 6953 15427 6987
rect 16589 6953 16623 6987
rect 19257 6953 19291 6987
rect 19349 6953 19383 6987
rect 20085 6953 20119 6987
rect 9781 6885 9815 6919
rect 13461 6885 13495 6919
rect 18429 6885 18463 6919
rect 2329 6817 2363 6851
rect 3157 6817 3191 6851
rect 4333 6817 4367 6851
rect 5816 6817 5850 6851
rect 7389 6817 7423 6851
rect 8309 6817 8343 6851
rect 8953 6817 8987 6851
rect 10241 6817 10275 6851
rect 10701 6817 10735 6851
rect 11888 6817 11922 6851
rect 13921 6817 13955 6851
rect 14657 6817 14691 6851
rect 17417 6817 17451 6851
rect 20545 6817 20579 6851
rect 1685 6749 1719 6783
rect 2421 6749 2455 6783
rect 2605 6749 2639 6783
rect 3249 6749 3283 6783
rect 3433 6749 3467 6783
rect 4077 6749 4111 6783
rect 5549 6749 5583 6783
rect 7481 6749 7515 6783
rect 7573 6749 7607 6783
rect 7849 6749 7883 6783
rect 8033 6749 8067 6783
rect 8401 6749 8435 6783
rect 10517 6749 10551 6783
rect 11621 6749 11655 6783
rect 13553 6749 13587 6783
rect 13645 6749 13679 6783
rect 14841 6749 14875 6783
rect 16681 6749 16715 6783
rect 16865 6749 16899 6783
rect 17509 6749 17543 6783
rect 17601 6749 17635 6783
rect 18521 6749 18555 6783
rect 18705 6749 18739 6783
rect 19441 6749 19475 6783
rect 20177 6749 20211 6783
rect 20361 6749 20395 6783
rect 1961 6681 1995 6715
rect 2789 6681 2823 6715
rect 8677 6681 8711 6715
rect 13093 6681 13127 6715
rect 16037 6681 16071 6715
rect 18061 6681 18095 6715
rect 18889 6681 18923 6715
rect 19717 6681 19751 6715
rect 21097 6681 21131 6715
rect 1501 6613 1535 6647
rect 5457 6613 5491 6647
rect 6929 6613 6963 6647
rect 8769 6613 8803 6647
rect 9413 6613 9447 6647
rect 9873 6613 9907 6647
rect 13001 6613 13035 6647
rect 14197 6613 14231 6647
rect 15577 6613 15611 6647
rect 16221 6613 16255 6647
rect 17049 6613 17083 6647
rect 17969 6613 18003 6647
rect 21005 6613 21039 6647
rect 22017 6613 22051 6647
rect 2053 6409 2087 6443
rect 4721 6409 4755 6443
rect 10701 6409 10735 6443
rect 11989 6409 12023 6443
rect 13369 6409 13403 6443
rect 15577 6409 15611 6443
rect 18153 6409 18187 6443
rect 20637 6409 20671 6443
rect 5825 6341 5859 6375
rect 12449 6341 12483 6375
rect 15761 6341 15795 6375
rect 2697 6273 2731 6307
rect 3801 6273 3835 6307
rect 5181 6273 5215 6307
rect 5273 6273 5307 6307
rect 6561 6273 6595 6307
rect 7389 6273 7423 6307
rect 8309 6273 8343 6307
rect 9137 6273 9171 6307
rect 10241 6273 10275 6307
rect 11529 6273 11563 6307
rect 11713 6273 11747 6307
rect 12909 6273 12943 6307
rect 13001 6273 13035 6307
rect 16221 6273 16255 6307
rect 16405 6273 16439 6307
rect 17233 6273 17267 6307
rect 17417 6273 17451 6307
rect 18797 6273 18831 6307
rect 19257 6273 19291 6307
rect 2421 6205 2455 6239
rect 5549 6205 5583 6239
rect 6377 6205 6411 6239
rect 7297 6205 7331 6239
rect 9045 6205 9079 6239
rect 10977 6205 11011 6239
rect 11437 6205 11471 6239
rect 14197 6205 14231 6239
rect 14464 6205 14498 6239
rect 16129 6205 16163 6239
rect 1593 6137 1627 6171
rect 2973 6137 3007 6171
rect 5089 6137 5123 6171
rect 7205 6137 7239 6171
rect 8125 6137 8159 6171
rect 9965 6137 9999 6171
rect 10517 6137 10551 6171
rect 12817 6137 12851 6171
rect 13829 6137 13863 6171
rect 16957 6137 16991 6171
rect 17785 6137 17819 6171
rect 18613 6137 18647 6171
rect 19524 6137 19558 6171
rect 1777 6069 1811 6103
rect 2513 6069 2547 6103
rect 3157 6069 3191 6103
rect 3525 6069 3559 6103
rect 3617 6069 3651 6103
rect 5917 6069 5951 6103
rect 6285 6069 6319 6103
rect 6837 6069 6871 6103
rect 7665 6069 7699 6103
rect 8033 6069 8067 6103
rect 8585 6069 8619 6103
rect 8953 6069 8987 6103
rect 9413 6069 9447 6103
rect 9597 6069 9631 6103
rect 10057 6069 10091 6103
rect 11069 6069 11103 6103
rect 13645 6069 13679 6103
rect 14105 6069 14139 6103
rect 16589 6069 16623 6103
rect 17049 6069 17083 6103
rect 18521 6069 18555 6103
rect 2329 5865 2363 5899
rect 2697 5865 2731 5899
rect 6193 5865 6227 5899
rect 6745 5865 6779 5899
rect 7481 5865 7515 5899
rect 8585 5865 8619 5899
rect 11621 5865 11655 5899
rect 12081 5865 12115 5899
rect 12357 5865 12391 5899
rect 15761 5865 15795 5899
rect 16221 5865 16255 5899
rect 16589 5865 16623 5899
rect 16773 5865 16807 5899
rect 17233 5865 17267 5899
rect 17601 5865 17635 5899
rect 17969 5865 18003 5899
rect 18429 5865 18463 5899
rect 20085 5865 20119 5899
rect 1961 5797 1995 5831
rect 2789 5797 2823 5831
rect 7113 5797 7147 5831
rect 8125 5797 8159 5831
rect 11529 5797 11563 5831
rect 12808 5797 12842 5831
rect 20453 5797 20487 5831
rect 1685 5729 1719 5763
rect 3525 5729 3559 5763
rect 4436 5729 4470 5763
rect 6653 5729 6687 5763
rect 8953 5729 8987 5763
rect 9956 5729 9990 5763
rect 12541 5729 12575 5763
rect 14013 5729 14047 5763
rect 14749 5729 14783 5763
rect 16129 5729 16163 5763
rect 17141 5729 17175 5763
rect 18705 5729 18739 5763
rect 18972 5729 19006 5763
rect 20177 5729 20211 5763
rect 2881 5661 2915 5695
rect 3617 5661 3651 5695
rect 3801 5661 3835 5695
rect 4169 5661 4203 5695
rect 6837 5661 6871 5695
rect 7297 5661 7331 5695
rect 8217 5661 8251 5695
rect 8401 5661 8435 5695
rect 9045 5661 9079 5695
rect 9137 5661 9171 5695
rect 9689 5661 9723 5695
rect 11713 5661 11747 5695
rect 14841 5661 14875 5695
rect 15025 5661 15059 5695
rect 16405 5661 16439 5695
rect 17325 5661 17359 5695
rect 18061 5661 18095 5695
rect 18153 5661 18187 5695
rect 3157 5593 3191 5627
rect 5549 5593 5583 5627
rect 11161 5593 11195 5627
rect 14197 5593 14231 5627
rect 5733 5525 5767 5559
rect 6285 5525 6319 5559
rect 7757 5525 7791 5559
rect 9505 5525 9539 5559
rect 11069 5525 11103 5559
rect 13921 5525 13955 5559
rect 14381 5525 14415 5559
rect 15301 5525 15335 5559
rect 15577 5525 15611 5559
rect 22017 5525 22051 5559
rect 4721 5321 4755 5355
rect 5549 5321 5583 5355
rect 7021 5321 7055 5355
rect 7205 5321 7239 5355
rect 8309 5321 8343 5355
rect 14197 5321 14231 5355
rect 16589 5321 16623 5355
rect 17877 5321 17911 5355
rect 19533 5321 19567 5355
rect 19625 5321 19659 5355
rect 4629 5253 4663 5287
rect 16497 5253 16531 5287
rect 5365 5185 5399 5219
rect 6009 5185 6043 5219
rect 6193 5185 6227 5219
rect 6469 5185 6503 5219
rect 7849 5185 7883 5219
rect 7941 5185 7975 5219
rect 8861 5185 8895 5219
rect 9137 5185 9171 5219
rect 11069 5185 11103 5219
rect 11161 5185 11195 5219
rect 11989 5185 12023 5219
rect 13093 5185 13127 5219
rect 14013 5185 14047 5219
rect 14841 5185 14875 5219
rect 17049 5185 17083 5219
rect 17233 5185 17267 5219
rect 20177 5185 20211 5219
rect 1777 5117 1811 5151
rect 3249 5117 3283 5151
rect 3516 5117 3550 5151
rect 9404 5117 9438 5151
rect 11805 5117 11839 5151
rect 11897 5117 11931 5151
rect 13829 5117 13863 5151
rect 14657 5117 14691 5151
rect 15117 5117 15151 5151
rect 16957 5117 16991 5151
rect 17693 5117 17727 5151
rect 18153 5117 18187 5151
rect 2044 5049 2078 5083
rect 5089 5049 5123 5083
rect 5917 5049 5951 5083
rect 6653 5049 6687 5083
rect 7757 5049 7791 5083
rect 8677 5049 8711 5083
rect 8769 5049 8803 5083
rect 10977 5049 11011 5083
rect 12817 5049 12851 5083
rect 15362 5049 15396 5083
rect 18398 5049 18432 5083
rect 20085 5049 20119 5083
rect 3157 4981 3191 5015
rect 5181 4981 5215 5015
rect 7389 4981 7423 5015
rect 10517 4981 10551 5015
rect 10609 4981 10643 5015
rect 11437 4981 11471 5015
rect 12449 4981 12483 5015
rect 12909 4981 12943 5015
rect 13369 4981 13403 5015
rect 13737 4981 13771 5015
rect 14565 4981 14599 5015
rect 19993 4981 20027 5015
rect 2789 4777 2823 4811
rect 4077 4777 4111 4811
rect 5273 4777 5307 4811
rect 7573 4777 7607 4811
rect 7941 4777 7975 4811
rect 8401 4777 8435 4811
rect 8769 4777 8803 4811
rect 9137 4777 9171 4811
rect 9689 4777 9723 4811
rect 10609 4777 10643 4811
rect 11989 4777 12023 4811
rect 12265 4777 12299 4811
rect 12449 4777 12483 4811
rect 15301 4777 15335 4811
rect 16865 4777 16899 4811
rect 17693 4777 17727 4811
rect 18521 4777 18555 4811
rect 19809 4777 19843 4811
rect 1676 4709 1710 4743
rect 5908 4709 5942 4743
rect 12992 4709 13026 4743
rect 14657 4709 14691 4743
rect 15025 4709 15059 4743
rect 15752 4709 15786 4743
rect 18981 4709 19015 4743
rect 1409 4641 1443 4675
rect 3525 4641 3559 4675
rect 5181 4641 5215 4675
rect 7481 4641 7515 4675
rect 8309 4641 8343 4675
rect 10057 4641 10091 4675
rect 10149 4641 10183 4675
rect 10885 4641 10919 4675
rect 11529 4641 11563 4675
rect 14565 4641 14599 4675
rect 18061 4641 18095 4675
rect 18889 4641 18923 4675
rect 19717 4641 19751 4675
rect 3617 4573 3651 4607
rect 3709 4573 3743 4607
rect 5365 4573 5399 4607
rect 5641 4573 5675 4607
rect 7665 4573 7699 4607
rect 8493 4573 8527 4607
rect 9229 4573 9263 4607
rect 9321 4573 9355 4607
rect 10333 4573 10367 4607
rect 11621 4573 11655 4607
rect 11805 4573 11839 4607
rect 12725 4573 12759 4607
rect 14749 4573 14783 4607
rect 15485 4573 15519 4607
rect 18153 4573 18187 4607
rect 18337 4573 18371 4607
rect 19165 4573 19199 4607
rect 19901 4573 19935 4607
rect 3157 4505 3191 4539
rect 17601 4505 17635 4539
rect 19349 4505 19383 4539
rect 2973 4437 3007 4471
rect 4537 4437 4571 4471
rect 4813 4437 4847 4471
rect 7021 4437 7055 4471
rect 7113 4437 7147 4471
rect 10977 4437 11011 4471
rect 11161 4437 11195 4471
rect 14105 4437 14139 4471
rect 14197 4437 14231 4471
rect 16957 4437 16991 4471
rect 4169 4233 4203 4267
rect 4813 4233 4847 4267
rect 15117 4233 15151 4267
rect 17509 4233 17543 4267
rect 19441 4233 19475 4267
rect 19533 4233 19567 4267
rect 9689 4165 9723 4199
rect 12909 4165 12943 4199
rect 14933 4165 14967 4199
rect 2421 4097 2455 4131
rect 2605 4097 2639 4131
rect 4629 4097 4663 4131
rect 5549 4097 5583 4131
rect 6285 4097 6319 4131
rect 6377 4097 6411 4131
rect 8493 4097 8527 4131
rect 9137 4097 9171 4131
rect 9229 4097 9263 4131
rect 10425 4097 10459 4131
rect 11805 4097 11839 4131
rect 11897 4097 11931 4131
rect 12173 4097 12207 4131
rect 13645 4097 13679 4131
rect 14473 4097 14507 4131
rect 15577 4097 15611 4131
rect 15761 4097 15795 4131
rect 16129 4097 16163 4131
rect 20085 4097 20119 4131
rect 2789 4029 2823 4063
rect 6929 4029 6963 4063
rect 9597 4029 9631 4063
rect 10241 4029 10275 4063
rect 10333 4029 10367 4063
rect 11713 4029 11747 4063
rect 13369 4029 13403 4063
rect 13461 4029 13495 4063
rect 14749 4029 14783 4063
rect 16396 4029 16430 4063
rect 18068 4029 18102 4063
rect 3056 3961 3090 3995
rect 5457 3961 5491 3995
rect 7196 3961 7230 3995
rect 9045 3961 9079 3995
rect 12633 3961 12667 3995
rect 14289 3961 14323 3995
rect 15945 3961 15979 3995
rect 17877 3961 17911 3995
rect 18306 3961 18340 3995
rect 1961 3893 1995 3927
rect 2329 3893 2363 3927
rect 4997 3893 5031 3927
rect 5365 3893 5399 3927
rect 5825 3893 5859 3927
rect 6193 3893 6227 3927
rect 8309 3893 8343 3927
rect 8677 3893 8711 3927
rect 9873 3893 9907 3927
rect 11345 3893 11379 3927
rect 12541 3893 12575 3927
rect 13001 3893 13035 3927
rect 13829 3893 13863 3927
rect 14197 3893 14231 3927
rect 15485 3893 15519 3927
rect 17601 3893 17635 3927
rect 19901 3893 19935 3927
rect 19993 3893 20027 3927
rect 20361 3893 20395 3927
rect 2329 3689 2363 3723
rect 3157 3689 3191 3723
rect 3617 3689 3651 3723
rect 5457 3689 5491 3723
rect 5917 3689 5951 3723
rect 6285 3689 6319 3723
rect 8125 3689 8159 3723
rect 8769 3689 8803 3723
rect 12909 3689 12943 3723
rect 13461 3689 13495 3723
rect 14289 3689 14323 3723
rect 15025 3689 15059 3723
rect 16313 3689 16347 3723
rect 18981 3689 19015 3723
rect 19809 3689 19843 3723
rect 20177 3689 20211 3723
rect 2789 3621 2823 3655
rect 4322 3621 4356 3655
rect 6990 3621 7024 3655
rect 8585 3621 8619 3655
rect 9229 3621 9263 3655
rect 19441 3621 19475 3655
rect 2697 3553 2731 3587
rect 3525 3553 3559 3587
rect 4077 3553 4111 3587
rect 8493 3553 8527 3587
rect 9137 3553 9171 3587
rect 9956 3553 9990 3587
rect 11529 3553 11563 3587
rect 11796 3553 11830 3587
rect 13369 3553 13403 3587
rect 14197 3553 14231 3587
rect 14657 3553 14691 3587
rect 15669 3553 15703 3587
rect 16129 3553 16163 3587
rect 16948 3553 16982 3587
rect 18521 3553 18555 3587
rect 19349 3553 19383 3587
rect 2973 3485 3007 3519
rect 3801 3485 3835 3519
rect 6377 3485 6411 3519
rect 6561 3485 6595 3519
rect 6745 3485 6779 3519
rect 9413 3485 9447 3519
rect 9689 3485 9723 3519
rect 11161 3485 11195 3519
rect 13645 3485 13679 3519
rect 14381 3485 14415 3519
rect 15761 3485 15795 3519
rect 15853 3485 15887 3519
rect 16681 3485 16715 3519
rect 18613 3485 18647 3519
rect 18797 3485 18831 3519
rect 19533 3485 19567 3519
rect 5825 3349 5859 3383
rect 8309 3349 8343 3383
rect 11069 3349 11103 3383
rect 13001 3349 13035 3383
rect 13829 3349 13863 3383
rect 14841 3349 14875 3383
rect 15301 3349 15335 3383
rect 16497 3349 16531 3383
rect 18061 3349 18095 3383
rect 18153 3349 18187 3383
rect 20361 3349 20395 3383
rect 2513 3145 2547 3179
rect 3341 3145 3375 3179
rect 5917 3145 5951 3179
rect 8401 3145 8435 3179
rect 9045 3145 9079 3179
rect 13829 3145 13863 3179
rect 16865 3145 16899 3179
rect 17141 3145 17175 3179
rect 18153 3145 18187 3179
rect 11253 3077 11287 3111
rect 3157 3009 3191 3043
rect 3893 3009 3927 3043
rect 4353 3009 4387 3043
rect 6561 3009 6595 3043
rect 9597 3009 9631 3043
rect 12081 3009 12115 3043
rect 15117 3009 15151 3043
rect 15669 3009 15703 3043
rect 17785 3009 17819 3043
rect 18797 3009 18831 3043
rect 19533 3009 19567 3043
rect 2421 2941 2455 2975
rect 2973 2941 3007 2975
rect 3709 2941 3743 2975
rect 3801 2941 3835 2975
rect 6377 2941 6411 2975
rect 7021 2941 7055 2975
rect 8493 2941 8527 2975
rect 8769 2941 8803 2975
rect 9505 2941 9539 2975
rect 9873 2941 9907 2975
rect 10140 2941 10174 2975
rect 12449 2941 12483 2975
rect 13921 2941 13955 2975
rect 14565 2941 14599 2975
rect 15393 2941 15427 2975
rect 15945 2941 15979 2975
rect 16497 2941 16531 2975
rect 17509 2941 17543 2975
rect 18521 2941 18555 2975
rect 19349 2941 19383 2975
rect 19809 2941 19843 2975
rect 20177 2941 20211 2975
rect 20545 2941 20579 2975
rect 20913 2941 20947 2975
rect 4261 2873 4295 2907
rect 4620 2873 4654 2907
rect 6285 2873 6319 2907
rect 6929 2873 6963 2907
rect 7288 2873 7322 2907
rect 11897 2873 11931 2907
rect 12716 2873 12750 2907
rect 14197 2873 14231 2907
rect 14841 2873 14875 2907
rect 16221 2873 16255 2907
rect 17601 2873 17635 2907
rect 19441 2873 19475 2907
rect 2881 2805 2915 2839
rect 5733 2805 5767 2839
rect 9413 2805 9447 2839
rect 11529 2805 11563 2839
rect 11989 2805 12023 2839
rect 16681 2805 16715 2839
rect 18613 2805 18647 2839
rect 18981 2805 19015 2839
rect 19993 2805 20027 2839
rect 20361 2805 20395 2839
rect 20729 2805 20763 2839
rect 3341 2601 3375 2635
rect 4169 2601 4203 2635
rect 4997 2601 5031 2635
rect 5365 2601 5399 2635
rect 6009 2601 6043 2635
rect 7389 2601 7423 2635
rect 9321 2601 9355 2635
rect 9781 2601 9815 2635
rect 11437 2601 11471 2635
rect 12633 2601 12667 2635
rect 13093 2601 13127 2635
rect 16313 2601 16347 2635
rect 17049 2601 17083 2635
rect 19625 2601 19659 2635
rect 20085 2601 20119 2635
rect 6469 2533 6503 2567
rect 8585 2533 8619 2567
rect 10241 2533 10275 2567
rect 12265 2533 12299 2567
rect 19257 2533 19291 2567
rect 4537 2465 4571 2499
rect 5457 2465 5491 2499
rect 5917 2465 5951 2499
rect 6377 2465 6411 2499
rect 7021 2465 7055 2499
rect 7757 2465 7791 2499
rect 10149 2465 10183 2499
rect 10609 2465 10643 2499
rect 11621 2465 11655 2499
rect 11989 2465 12023 2499
rect 13001 2465 13035 2499
rect 13461 2465 13495 2499
rect 13829 2465 13863 2499
rect 14197 2465 14231 2499
rect 14565 2465 14599 2499
rect 15025 2465 15059 2499
rect 15485 2465 15519 2499
rect 15853 2465 15887 2499
rect 16221 2465 16255 2499
rect 16497 2465 16531 2499
rect 16865 2465 16899 2499
rect 17233 2465 17267 2499
rect 18337 2465 18371 2499
rect 18705 2465 18739 2499
rect 19073 2465 19107 2499
rect 4629 2397 4663 2431
rect 4813 2397 4847 2431
rect 5549 2397 5583 2431
rect 6561 2397 6595 2431
rect 7849 2397 7883 2431
rect 8033 2397 8067 2431
rect 8677 2397 8711 2431
rect 8861 2397 8895 2431
rect 10425 2397 10459 2431
rect 10885 2397 10919 2431
rect 13185 2397 13219 2431
rect 8217 2329 8251 2363
rect 14013 2329 14047 2363
rect 17785 2397 17819 2431
rect 17969 2397 18003 2431
rect 16681 2329 16715 2363
rect 17417 2329 17451 2363
rect 3157 2261 3191 2295
rect 3617 2261 3651 2295
rect 3801 2261 3835 2295
rect 7205 2261 7239 2295
rect 9045 2261 9079 2295
rect 9597 2261 9631 2295
rect 11161 2261 11195 2295
rect 11805 2261 11839 2295
rect 13645 2261 13679 2295
rect 14381 2261 14415 2295
rect 14749 2261 14783 2295
rect 15209 2261 15243 2295
rect 15669 2261 15703 2295
rect 16037 2261 16071 2295
rect 16221 2261 16255 2295
rect 17601 2261 17635 2295
rect 18521 2261 18555 2295
rect 18889 2261 18923 2295
rect 19533 2261 19567 2295
rect 19901 2261 19935 2295
rect 6193 2057 6227 2091
rect 6193 1785 6227 1819
<< metal1 >>
rect 1104 20698 21896 20720
rect 1104 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 4575 20698
rect 4627 20646 4639 20698
rect 4691 20646 11378 20698
rect 11430 20646 11442 20698
rect 11494 20646 11506 20698
rect 11558 20646 11570 20698
rect 11622 20646 18308 20698
rect 18360 20646 18372 20698
rect 18424 20646 18436 20698
rect 18488 20646 18500 20698
rect 18552 20646 21896 20698
rect 1104 20624 21896 20646
rect 4801 20587 4859 20593
rect 4801 20553 4813 20587
rect 4847 20584 4859 20587
rect 11698 20584 11704 20596
rect 4847 20556 11704 20584
rect 4847 20553 4859 20556
rect 4801 20547 4859 20553
rect 11698 20544 11704 20556
rect 11756 20544 11762 20596
rect 18966 20584 18972 20596
rect 18927 20556 18972 20584
rect 18966 20544 18972 20556
rect 19024 20544 19030 20596
rect 19153 20587 19211 20593
rect 19153 20553 19165 20587
rect 19199 20584 19211 20587
rect 19334 20584 19340 20596
rect 19199 20556 19340 20584
rect 19199 20553 19211 20556
rect 19153 20547 19211 20553
rect 19334 20544 19340 20556
rect 19392 20544 19398 20596
rect 20898 20544 20904 20596
rect 20956 20584 20962 20596
rect 21361 20587 21419 20593
rect 21361 20584 21373 20587
rect 20956 20556 21373 20584
rect 20956 20544 20962 20556
rect 21361 20553 21373 20556
rect 21407 20553 21419 20587
rect 21361 20547 21419 20553
rect 4338 20476 4344 20528
rect 4396 20516 4402 20528
rect 5350 20516 5356 20528
rect 4396 20488 5356 20516
rect 4396 20476 4402 20488
rect 5350 20476 5356 20488
rect 5408 20476 5414 20528
rect 6917 20519 6975 20525
rect 6917 20485 6929 20519
rect 6963 20516 6975 20519
rect 9858 20516 9864 20528
rect 6963 20488 9864 20516
rect 6963 20485 6975 20488
rect 6917 20479 6975 20485
rect 9858 20476 9864 20488
rect 9916 20476 9922 20528
rect 20622 20476 20628 20528
rect 20680 20516 20686 20528
rect 21177 20519 21235 20525
rect 21177 20516 21189 20519
rect 20680 20488 21189 20516
rect 20680 20476 20686 20488
rect 21177 20485 21189 20488
rect 21223 20485 21235 20519
rect 21177 20479 21235 20485
rect 6638 20408 6644 20460
rect 6696 20448 6702 20460
rect 7469 20451 7527 20457
rect 7469 20448 7481 20451
rect 6696 20420 7481 20448
rect 6696 20408 6702 20420
rect 7469 20417 7481 20420
rect 7515 20417 7527 20451
rect 7469 20411 7527 20417
rect 20809 20451 20867 20457
rect 20809 20417 20821 20451
rect 20855 20448 20867 20451
rect 22370 20448 22376 20460
rect 20855 20420 22376 20448
rect 20855 20417 20867 20420
rect 20809 20411 20867 20417
rect 22370 20408 22376 20420
rect 22428 20408 22434 20460
rect 4338 20340 4344 20392
rect 4396 20380 4402 20392
rect 4617 20383 4675 20389
rect 4617 20380 4629 20383
rect 4396 20352 4629 20380
rect 4396 20340 4402 20352
rect 4617 20349 4629 20352
rect 4663 20349 4675 20383
rect 4617 20343 4675 20349
rect 19981 20383 20039 20389
rect 19981 20349 19993 20383
rect 20027 20349 20039 20383
rect 19981 20343 20039 20349
rect 20533 20383 20591 20389
rect 20533 20349 20545 20383
rect 20579 20380 20591 20383
rect 20714 20380 20720 20392
rect 20579 20352 20720 20380
rect 20579 20349 20591 20352
rect 20533 20343 20591 20349
rect 5442 20272 5448 20324
rect 5500 20312 5506 20324
rect 7377 20315 7435 20321
rect 7377 20312 7389 20315
rect 5500 20284 7389 20312
rect 5500 20272 5506 20284
rect 7377 20281 7389 20284
rect 7423 20281 7435 20315
rect 7377 20275 7435 20281
rect 7834 20272 7840 20324
rect 7892 20312 7898 20324
rect 13446 20312 13452 20324
rect 7892 20284 13452 20312
rect 7892 20272 7898 20284
rect 13446 20272 13452 20284
rect 13504 20272 13510 20324
rect 7282 20244 7288 20256
rect 7243 20216 7288 20244
rect 7282 20204 7288 20216
rect 7340 20204 7346 20256
rect 19610 20204 19616 20256
rect 19668 20244 19674 20256
rect 19705 20247 19763 20253
rect 19705 20244 19717 20247
rect 19668 20216 19717 20244
rect 19668 20204 19674 20216
rect 19705 20213 19717 20216
rect 19751 20244 19763 20247
rect 19889 20247 19947 20253
rect 19889 20244 19901 20247
rect 19751 20216 19901 20244
rect 19751 20213 19763 20216
rect 19705 20207 19763 20213
rect 19889 20213 19901 20216
rect 19935 20244 19947 20247
rect 19996 20244 20024 20343
rect 20714 20340 20720 20352
rect 20772 20380 20778 20392
rect 20898 20380 20904 20392
rect 20772 20352 20904 20380
rect 20772 20340 20778 20352
rect 20898 20340 20904 20352
rect 20956 20340 20962 20392
rect 20257 20315 20315 20321
rect 20257 20281 20269 20315
rect 20303 20312 20315 20315
rect 22738 20312 22744 20324
rect 20303 20284 22744 20312
rect 20303 20281 20315 20284
rect 20257 20275 20315 20281
rect 22738 20272 22744 20284
rect 22796 20272 22802 20324
rect 21266 20244 21272 20256
rect 19935 20216 21272 20244
rect 19935 20213 19947 20216
rect 19889 20207 19947 20213
rect 21266 20204 21272 20216
rect 21324 20204 21330 20256
rect 1104 20154 21896 20176
rect 1104 20102 7912 20154
rect 7964 20102 7976 20154
rect 8028 20102 8040 20154
rect 8092 20102 8104 20154
rect 8156 20102 14843 20154
rect 14895 20102 14907 20154
rect 14959 20102 14971 20154
rect 15023 20102 15035 20154
rect 15087 20102 21896 20154
rect 1104 20080 21896 20102
rect 2866 20000 2872 20052
rect 2924 20040 2930 20052
rect 3326 20040 3332 20052
rect 2924 20012 3332 20040
rect 2924 20000 2930 20012
rect 3326 20000 3332 20012
rect 3384 20040 3390 20052
rect 7285 20043 7343 20049
rect 7285 20040 7297 20043
rect 3384 20012 7297 20040
rect 3384 20000 3390 20012
rect 7285 20009 7297 20012
rect 7331 20040 7343 20043
rect 7374 20040 7380 20052
rect 7331 20012 7380 20040
rect 7331 20009 7343 20012
rect 7285 20003 7343 20009
rect 7374 20000 7380 20012
rect 7432 20000 7438 20052
rect 7558 20000 7564 20052
rect 7616 20040 7622 20052
rect 9030 20040 9036 20052
rect 7616 20012 9036 20040
rect 7616 20000 7622 20012
rect 9030 20000 9036 20012
rect 9088 20000 9094 20052
rect 9953 20043 10011 20049
rect 9953 20009 9965 20043
rect 9999 20040 10011 20043
rect 10870 20040 10876 20052
rect 9999 20012 10876 20040
rect 9999 20009 10011 20012
rect 9953 20003 10011 20009
rect 10870 20000 10876 20012
rect 10928 20000 10934 20052
rect 11057 20043 11115 20049
rect 11057 20009 11069 20043
rect 11103 20040 11115 20043
rect 11238 20040 11244 20052
rect 11103 20012 11244 20040
rect 11103 20009 11115 20012
rect 11057 20003 11115 20009
rect 11238 20000 11244 20012
rect 11296 20000 11302 20052
rect 11977 20043 12035 20049
rect 11977 20009 11989 20043
rect 12023 20040 12035 20043
rect 12066 20040 12072 20052
rect 12023 20012 12072 20040
rect 12023 20009 12035 20012
rect 11977 20003 12035 20009
rect 12066 20000 12072 20012
rect 12124 20000 12130 20052
rect 13265 20043 13323 20049
rect 13265 20009 13277 20043
rect 13311 20040 13323 20043
rect 13998 20040 14004 20052
rect 13311 20012 14004 20040
rect 13311 20009 13323 20012
rect 13265 20003 13323 20009
rect 13998 20000 14004 20012
rect 14056 20000 14062 20052
rect 14737 20043 14795 20049
rect 14737 20009 14749 20043
rect 14783 20040 14795 20043
rect 15378 20040 15384 20052
rect 14783 20012 15384 20040
rect 14783 20009 14795 20012
rect 14737 20003 14795 20009
rect 15378 20000 15384 20012
rect 15436 20000 15442 20052
rect 15473 20043 15531 20049
rect 15473 20009 15485 20043
rect 15519 20040 15531 20043
rect 15838 20040 15844 20052
rect 15519 20012 15844 20040
rect 15519 20009 15531 20012
rect 15473 20003 15531 20009
rect 15838 20000 15844 20012
rect 15896 20000 15902 20052
rect 17313 20043 17371 20049
rect 17313 20009 17325 20043
rect 17359 20040 17371 20043
rect 18138 20040 18144 20052
rect 17359 20012 18144 20040
rect 17359 20009 17371 20012
rect 17313 20003 17371 20009
rect 18138 20000 18144 20012
rect 18196 20000 18202 20052
rect 4062 19932 4068 19984
rect 4120 19972 4126 19984
rect 18693 19975 18751 19981
rect 18693 19972 18705 19975
rect 4120 19944 18705 19972
rect 4120 19932 4126 19944
rect 18693 19941 18705 19944
rect 18739 19941 18751 19975
rect 18693 19935 18751 19941
rect 19242 19932 19248 19984
rect 19300 19972 19306 19984
rect 19337 19975 19395 19981
rect 19337 19972 19349 19975
rect 19300 19944 19349 19972
rect 19300 19932 19306 19944
rect 19337 19941 19349 19944
rect 19383 19941 19395 19975
rect 19337 19935 19395 19941
rect 19426 19932 19432 19984
rect 19484 19972 19490 19984
rect 19978 19972 19984 19984
rect 19484 19944 19840 19972
rect 19939 19944 19984 19972
rect 19484 19932 19490 19944
rect 4332 19907 4390 19913
rect 4332 19873 4344 19907
rect 4378 19904 4390 19907
rect 5534 19904 5540 19916
rect 4378 19876 5540 19904
rect 4378 19873 4390 19876
rect 4332 19867 4390 19873
rect 5534 19864 5540 19876
rect 5592 19864 5598 19916
rect 6080 19907 6138 19913
rect 6080 19873 6092 19907
rect 6126 19904 6138 19907
rect 6822 19904 6828 19916
rect 6126 19876 6828 19904
rect 6126 19873 6138 19876
rect 6080 19867 6138 19873
rect 6822 19864 6828 19876
rect 6880 19864 6886 19916
rect 7374 19864 7380 19916
rect 7432 19904 7438 19916
rect 8021 19907 8079 19913
rect 8021 19904 8033 19907
rect 7432 19876 8033 19904
rect 7432 19864 7438 19876
rect 8021 19873 8033 19876
rect 8067 19904 8079 19907
rect 8067 19876 9628 19904
rect 8067 19873 8079 19876
rect 8021 19867 8079 19873
rect 4062 19836 4068 19848
rect 4023 19808 4068 19836
rect 4062 19796 4068 19808
rect 4120 19796 4126 19848
rect 5258 19796 5264 19848
rect 5316 19836 5322 19848
rect 5813 19839 5871 19845
rect 5813 19836 5825 19839
rect 5316 19808 5825 19836
rect 5316 19796 5322 19808
rect 5813 19805 5825 19808
rect 5859 19805 5871 19839
rect 5813 19799 5871 19805
rect 8113 19839 8171 19845
rect 8113 19805 8125 19839
rect 8159 19805 8171 19839
rect 8294 19836 8300 19848
rect 8255 19808 8300 19836
rect 8113 19799 8171 19805
rect 7558 19768 7564 19780
rect 7519 19740 7564 19768
rect 7558 19728 7564 19740
rect 7616 19768 7622 19780
rect 8128 19768 8156 19799
rect 8294 19796 8300 19808
rect 8352 19796 8358 19848
rect 7616 19740 8156 19768
rect 8573 19771 8631 19777
rect 7616 19728 7622 19740
rect 8573 19737 8585 19771
rect 8619 19768 8631 19771
rect 8846 19768 8852 19780
rect 8619 19740 8852 19768
rect 8619 19737 8631 19740
rect 8573 19731 8631 19737
rect 8846 19728 8852 19740
rect 8904 19728 8910 19780
rect 4982 19660 4988 19712
rect 5040 19700 5046 19712
rect 5445 19703 5503 19709
rect 5445 19700 5457 19703
rect 5040 19672 5457 19700
rect 5040 19660 5046 19672
rect 5445 19669 5457 19672
rect 5491 19669 5503 19703
rect 7190 19700 7196 19712
rect 7151 19672 7196 19700
rect 5445 19663 5503 19669
rect 7190 19660 7196 19672
rect 7248 19660 7254 19712
rect 7650 19700 7656 19712
rect 7611 19672 7656 19700
rect 7650 19660 7656 19672
rect 7708 19660 7714 19712
rect 8754 19700 8760 19712
rect 8715 19672 8760 19700
rect 8754 19660 8760 19672
rect 8812 19660 8818 19712
rect 9600 19700 9628 19876
rect 9674 19864 9680 19916
rect 9732 19904 9738 19916
rect 9769 19907 9827 19913
rect 9769 19904 9781 19907
rect 9732 19876 9781 19904
rect 9732 19864 9738 19876
rect 9769 19873 9781 19876
rect 9815 19873 9827 19907
rect 9769 19867 9827 19873
rect 9950 19864 9956 19916
rect 10008 19904 10014 19916
rect 10321 19907 10379 19913
rect 10321 19904 10333 19907
rect 10008 19876 10333 19904
rect 10008 19864 10014 19876
rect 10321 19873 10333 19876
rect 10367 19873 10379 19907
rect 10870 19904 10876 19916
rect 10831 19876 10876 19904
rect 10321 19867 10379 19873
rect 10870 19864 10876 19876
rect 10928 19864 10934 19916
rect 11425 19907 11483 19913
rect 11425 19873 11437 19907
rect 11471 19873 11483 19907
rect 11425 19867 11483 19873
rect 11793 19907 11851 19913
rect 11793 19873 11805 19907
rect 11839 19904 11851 19907
rect 12158 19904 12164 19916
rect 11839 19876 12164 19904
rect 11839 19873 11851 19876
rect 11793 19867 11851 19873
rect 10597 19839 10655 19845
rect 10597 19805 10609 19839
rect 10643 19836 10655 19839
rect 11440 19836 11468 19867
rect 12158 19864 12164 19876
rect 12216 19864 12222 19916
rect 13078 19904 13084 19916
rect 13039 19876 13084 19904
rect 13078 19864 13084 19876
rect 13136 19864 13142 19916
rect 14550 19904 14556 19916
rect 14511 19876 14556 19904
rect 14550 19864 14556 19876
rect 14608 19864 14614 19916
rect 15194 19864 15200 19916
rect 15252 19904 15258 19916
rect 15289 19907 15347 19913
rect 15289 19904 15301 19907
rect 15252 19876 15301 19904
rect 15252 19864 15258 19876
rect 15289 19873 15301 19876
rect 15335 19904 15347 19907
rect 15657 19907 15715 19913
rect 15657 19904 15669 19907
rect 15335 19876 15669 19904
rect 15335 19873 15347 19876
rect 15289 19867 15347 19873
rect 15657 19873 15669 19876
rect 15703 19873 15715 19907
rect 15657 19867 15715 19873
rect 16114 19864 16120 19916
rect 16172 19904 16178 19916
rect 17037 19907 17095 19913
rect 17037 19904 17049 19907
rect 16172 19876 17049 19904
rect 16172 19864 16178 19876
rect 17037 19873 17049 19876
rect 17083 19904 17095 19907
rect 17129 19907 17187 19913
rect 17129 19904 17141 19907
rect 17083 19876 17141 19904
rect 17083 19873 17095 19876
rect 17037 19867 17095 19873
rect 17129 19873 17141 19876
rect 17175 19873 17187 19907
rect 17129 19867 17187 19873
rect 18417 19907 18475 19913
rect 18417 19873 18429 19907
rect 18463 19873 18475 19907
rect 18417 19867 18475 19873
rect 10643 19808 11468 19836
rect 18432 19836 18460 19867
rect 18966 19864 18972 19916
rect 19024 19904 19030 19916
rect 19061 19907 19119 19913
rect 19061 19904 19073 19907
rect 19024 19876 19073 19904
rect 19024 19864 19030 19876
rect 19061 19873 19073 19876
rect 19107 19873 19119 19907
rect 19061 19867 19119 19873
rect 19610 19864 19616 19916
rect 19668 19904 19674 19916
rect 19705 19907 19763 19913
rect 19705 19904 19717 19907
rect 19668 19876 19717 19904
rect 19668 19864 19674 19876
rect 19705 19873 19717 19876
rect 19751 19873 19763 19907
rect 19812 19904 19840 19944
rect 19978 19932 19984 19944
rect 20036 19932 20042 19984
rect 20530 19972 20536 19984
rect 20491 19944 20536 19972
rect 20530 19932 20536 19944
rect 20588 19932 20594 19984
rect 20622 19932 20628 19984
rect 20680 19932 20686 19984
rect 21177 19975 21235 19981
rect 21177 19941 21189 19975
rect 21223 19972 21235 19975
rect 21634 19972 21640 19984
rect 21223 19944 21640 19972
rect 21223 19941 21235 19944
rect 21177 19935 21235 19941
rect 21634 19932 21640 19944
rect 21692 19932 21698 19984
rect 20257 19907 20315 19913
rect 20257 19904 20269 19907
rect 19812 19876 20269 19904
rect 19705 19867 19763 19873
rect 20257 19873 20269 19876
rect 20303 19904 20315 19907
rect 20640 19904 20668 19932
rect 20303 19876 20668 19904
rect 20901 19907 20959 19913
rect 20303 19873 20315 19876
rect 20257 19867 20315 19873
rect 20901 19873 20913 19907
rect 20947 19873 20959 19907
rect 20901 19867 20959 19873
rect 19334 19836 19340 19848
rect 18432 19808 19340 19836
rect 10643 19805 10655 19808
rect 10597 19799 10655 19805
rect 19334 19796 19340 19808
rect 19392 19836 19398 19848
rect 20622 19836 20628 19848
rect 19392 19808 20628 19836
rect 19392 19796 19398 19808
rect 20622 19796 20628 19808
rect 20680 19836 20686 19848
rect 20916 19836 20944 19867
rect 21453 19839 21511 19845
rect 21453 19836 21465 19839
rect 20680 19808 21465 19836
rect 20680 19796 20686 19808
rect 21453 19805 21465 19808
rect 21499 19805 21511 19839
rect 21453 19799 21511 19805
rect 11609 19771 11667 19777
rect 11609 19737 11621 19771
rect 11655 19768 11667 19771
rect 12434 19768 12440 19780
rect 11655 19740 12440 19768
rect 11655 19737 11667 19740
rect 11609 19731 11667 19737
rect 12434 19728 12440 19740
rect 12492 19728 12498 19780
rect 12250 19700 12256 19712
rect 9600 19672 12256 19700
rect 12250 19660 12256 19672
rect 12308 19660 12314 19712
rect 1104 19610 21896 19632
rect 1104 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 4575 19610
rect 4627 19558 4639 19610
rect 4691 19558 11378 19610
rect 11430 19558 11442 19610
rect 11494 19558 11506 19610
rect 11558 19558 11570 19610
rect 11622 19558 18308 19610
rect 18360 19558 18372 19610
rect 18424 19558 18436 19610
rect 18488 19558 18500 19610
rect 18552 19558 21896 19610
rect 1104 19536 21896 19558
rect 1946 19496 1952 19508
rect 1907 19468 1952 19496
rect 1946 19456 1952 19468
rect 2004 19456 2010 19508
rect 4154 19496 4160 19508
rect 3804 19468 4160 19496
rect 3804 19369 3832 19468
rect 4154 19456 4160 19468
rect 4212 19496 4218 19508
rect 5258 19496 5264 19508
rect 4212 19468 5264 19496
rect 4212 19456 4218 19468
rect 5258 19456 5264 19468
rect 5316 19456 5322 19508
rect 5534 19456 5540 19508
rect 5592 19496 5598 19508
rect 6638 19496 6644 19508
rect 5592 19468 6644 19496
rect 5592 19456 5598 19468
rect 6638 19456 6644 19468
rect 6696 19456 6702 19508
rect 9122 19496 9128 19508
rect 6840 19468 9128 19496
rect 3789 19363 3847 19369
rect 3789 19329 3801 19363
rect 3835 19329 3847 19363
rect 3789 19323 3847 19329
rect 1765 19295 1823 19301
rect 1765 19261 1777 19295
rect 1811 19292 1823 19295
rect 3237 19295 3295 19301
rect 1811 19264 2268 19292
rect 1811 19261 1823 19264
rect 1765 19255 1823 19261
rect 198 19184 204 19236
rect 256 19224 262 19236
rect 2130 19224 2136 19236
rect 256 19196 2136 19224
rect 256 19184 262 19196
rect 2130 19184 2136 19196
rect 2188 19184 2194 19236
rect 2240 19165 2268 19264
rect 3237 19261 3249 19295
rect 3283 19261 3295 19295
rect 4338 19292 4344 19304
rect 3237 19255 3295 19261
rect 3988 19264 4344 19292
rect 2225 19159 2283 19165
rect 2225 19125 2237 19159
rect 2271 19156 2283 19159
rect 3050 19156 3056 19168
rect 2271 19128 3056 19156
rect 2271 19125 2283 19128
rect 2225 19119 2283 19125
rect 3050 19116 3056 19128
rect 3108 19116 3114 19168
rect 3252 19156 3280 19255
rect 3513 19227 3571 19233
rect 3513 19193 3525 19227
rect 3559 19224 3571 19227
rect 3988 19224 4016 19264
rect 4338 19252 4344 19264
rect 4396 19252 4402 19304
rect 5276 19301 5304 19456
rect 5261 19295 5319 19301
rect 5261 19261 5273 19295
rect 5307 19261 5319 19295
rect 5261 19255 5319 19261
rect 5902 19252 5908 19304
rect 5960 19292 5966 19304
rect 6840 19292 6868 19468
rect 9122 19456 9128 19468
rect 9180 19456 9186 19508
rect 15102 19496 15108 19508
rect 15063 19468 15108 19496
rect 15102 19456 15108 19468
rect 15160 19456 15166 19508
rect 10134 19388 10140 19440
rect 10192 19428 10198 19440
rect 10594 19428 10600 19440
rect 10192 19400 10600 19428
rect 10192 19388 10198 19400
rect 10594 19388 10600 19400
rect 10652 19388 10658 19440
rect 12069 19431 12127 19437
rect 12069 19428 12081 19431
rect 11532 19400 12081 19428
rect 8941 19363 8999 19369
rect 8941 19360 8953 19363
rect 8312 19332 8953 19360
rect 8312 19304 8340 19332
rect 8941 19329 8953 19332
rect 8987 19329 8999 19363
rect 10045 19363 10103 19369
rect 8941 19323 8999 19329
rect 9048 19332 9352 19360
rect 5960 19264 6868 19292
rect 5960 19252 5966 19264
rect 6914 19252 6920 19304
rect 6972 19292 6978 19304
rect 7184 19295 7242 19301
rect 6972 19264 7017 19292
rect 6972 19252 6978 19264
rect 7184 19261 7196 19295
rect 7230 19292 7242 19295
rect 8294 19292 8300 19304
rect 7230 19264 8300 19292
rect 7230 19261 7242 19264
rect 7184 19255 7242 19261
rect 8294 19252 8300 19264
rect 8352 19252 8358 19304
rect 8754 19292 8760 19304
rect 8715 19264 8760 19292
rect 8754 19252 8760 19264
rect 8812 19292 8818 19304
rect 9048 19292 9076 19332
rect 8812 19264 9076 19292
rect 9217 19295 9275 19301
rect 8812 19252 8818 19264
rect 9217 19261 9229 19295
rect 9263 19261 9275 19295
rect 9217 19255 9275 19261
rect 3559 19196 4016 19224
rect 4056 19227 4114 19233
rect 3559 19193 3571 19196
rect 3513 19187 3571 19193
rect 4056 19193 4068 19227
rect 4102 19224 4114 19227
rect 4982 19224 4988 19236
rect 4102 19196 4988 19224
rect 4102 19193 4114 19196
rect 4056 19187 4114 19193
rect 4982 19184 4988 19196
rect 5040 19184 5046 19236
rect 5528 19227 5586 19233
rect 5528 19193 5540 19227
rect 5574 19224 5586 19227
rect 7006 19224 7012 19236
rect 5574 19196 7012 19224
rect 5574 19193 5586 19196
rect 5528 19187 5586 19193
rect 7006 19184 7012 19196
rect 7064 19184 7070 19236
rect 7374 19184 7380 19236
rect 7432 19224 7438 19236
rect 9232 19224 9260 19255
rect 7432 19196 9260 19224
rect 9324 19224 9352 19332
rect 10045 19329 10057 19363
rect 10091 19360 10103 19363
rect 10870 19360 10876 19372
rect 10091 19332 10876 19360
rect 10091 19329 10103 19332
rect 10045 19323 10103 19329
rect 10870 19320 10876 19332
rect 10928 19320 10934 19372
rect 10962 19320 10968 19372
rect 11020 19360 11026 19372
rect 11020 19332 11065 19360
rect 11020 19320 11026 19332
rect 9493 19295 9551 19301
rect 9493 19261 9505 19295
rect 9539 19292 9551 19295
rect 9674 19292 9680 19304
rect 9539 19264 9680 19292
rect 9539 19261 9551 19264
rect 9493 19255 9551 19261
rect 9674 19252 9680 19264
rect 9732 19252 9738 19304
rect 9769 19295 9827 19301
rect 9769 19261 9781 19295
rect 9815 19292 9827 19295
rect 9858 19292 9864 19304
rect 9815 19264 9864 19292
rect 9815 19261 9827 19264
rect 9769 19255 9827 19261
rect 9858 19252 9864 19264
rect 9916 19252 9922 19304
rect 10781 19295 10839 19301
rect 10781 19261 10793 19295
rect 10827 19292 10839 19295
rect 11532 19292 11560 19400
rect 12069 19397 12081 19400
rect 12115 19397 12127 19431
rect 12069 19391 12127 19397
rect 11885 19363 11943 19369
rect 11885 19329 11897 19363
rect 11931 19360 11943 19363
rect 11974 19360 11980 19372
rect 11931 19332 11980 19360
rect 11931 19329 11943 19332
rect 11885 19323 11943 19329
rect 11974 19320 11980 19332
rect 12032 19320 12038 19372
rect 12084 19304 12112 19391
rect 12713 19363 12771 19369
rect 12713 19329 12725 19363
rect 12759 19360 12771 19363
rect 13078 19360 13084 19372
rect 12759 19332 13084 19360
rect 12759 19329 12771 19332
rect 12713 19323 12771 19329
rect 13078 19320 13084 19332
rect 13136 19320 13142 19372
rect 18966 19360 18972 19372
rect 18248 19332 18972 19360
rect 10827 19264 11560 19292
rect 11609 19295 11667 19301
rect 10827 19261 10839 19264
rect 10781 19255 10839 19261
rect 11609 19261 11621 19295
rect 11655 19292 11667 19295
rect 11698 19292 11704 19304
rect 11655 19264 11704 19292
rect 11655 19261 11667 19264
rect 11609 19255 11667 19261
rect 11698 19252 11704 19264
rect 11756 19252 11762 19304
rect 12066 19252 12072 19304
rect 12124 19252 12130 19304
rect 12437 19295 12495 19301
rect 12437 19261 12449 19295
rect 12483 19261 12495 19295
rect 12986 19292 12992 19304
rect 12947 19264 12992 19292
rect 12437 19255 12495 19261
rect 11146 19224 11152 19236
rect 9324 19196 11152 19224
rect 7432 19184 7438 19196
rect 11146 19184 11152 19196
rect 11204 19184 11210 19236
rect 12452 19224 12480 19255
rect 12986 19252 12992 19264
rect 13044 19252 13050 19304
rect 13354 19292 13360 19304
rect 13315 19264 13360 19292
rect 13354 19252 13360 19264
rect 13412 19252 13418 19304
rect 13722 19292 13728 19304
rect 13683 19264 13728 19292
rect 13722 19252 13728 19264
rect 13780 19252 13786 19304
rect 14182 19292 14188 19304
rect 14143 19264 14188 19292
rect 14182 19252 14188 19264
rect 14240 19252 14246 19304
rect 14458 19252 14464 19304
rect 14516 19292 14522 19304
rect 14553 19295 14611 19301
rect 14553 19292 14565 19295
rect 14516 19264 14565 19292
rect 14516 19252 14522 19264
rect 14553 19261 14565 19264
rect 14599 19261 14611 19295
rect 14553 19255 14611 19261
rect 14921 19295 14979 19301
rect 14921 19261 14933 19295
rect 14967 19292 14979 19295
rect 15562 19292 15568 19304
rect 14967 19264 15332 19292
rect 15523 19264 15568 19292
rect 14967 19261 14979 19264
rect 14921 19255 14979 19261
rect 11256 19196 12480 19224
rect 4890 19156 4896 19168
rect 3252 19128 4896 19156
rect 4890 19116 4896 19128
rect 4948 19116 4954 19168
rect 5074 19116 5080 19168
rect 5132 19156 5138 19168
rect 5169 19159 5227 19165
rect 5169 19156 5181 19159
rect 5132 19128 5181 19156
rect 5132 19116 5138 19128
rect 5169 19125 5181 19128
rect 5215 19125 5227 19159
rect 5169 19119 5227 19125
rect 5258 19116 5264 19168
rect 5316 19156 5322 19168
rect 6730 19156 6736 19168
rect 5316 19128 6736 19156
rect 5316 19116 5322 19128
rect 6730 19116 6736 19128
rect 6788 19116 6794 19168
rect 6822 19116 6828 19168
rect 6880 19156 6886 19168
rect 8297 19159 8355 19165
rect 8297 19156 8309 19159
rect 6880 19128 8309 19156
rect 6880 19116 6886 19128
rect 8297 19125 8309 19128
rect 8343 19125 8355 19159
rect 8297 19119 8355 19125
rect 8386 19116 8392 19168
rect 8444 19156 8450 19168
rect 8846 19156 8852 19168
rect 8444 19128 8489 19156
rect 8807 19128 8852 19156
rect 8444 19116 8450 19128
rect 8846 19116 8852 19128
rect 8904 19116 8910 19168
rect 10134 19116 10140 19168
rect 10192 19156 10198 19168
rect 10413 19159 10471 19165
rect 10413 19156 10425 19159
rect 10192 19128 10425 19156
rect 10192 19116 10198 19128
rect 10413 19125 10425 19128
rect 10459 19125 10471 19159
rect 10413 19119 10471 19125
rect 10870 19116 10876 19168
rect 10928 19156 10934 19168
rect 11256 19165 11284 19196
rect 15304 19168 15332 19264
rect 15562 19252 15568 19264
rect 15620 19252 15626 19304
rect 16022 19252 16028 19304
rect 16080 19292 16086 19304
rect 16117 19295 16175 19301
rect 16117 19292 16129 19295
rect 16080 19264 16129 19292
rect 16080 19252 16086 19264
rect 16117 19261 16129 19264
rect 16163 19261 16175 19295
rect 16117 19255 16175 19261
rect 16485 19295 16543 19301
rect 16485 19261 16497 19295
rect 16531 19292 16543 19295
rect 17126 19292 17132 19304
rect 16531 19264 16988 19292
rect 17087 19264 17132 19292
rect 16531 19261 16543 19264
rect 16485 19255 16543 19261
rect 15838 19224 15844 19236
rect 15799 19196 15844 19224
rect 15838 19184 15844 19196
rect 15896 19184 15902 19236
rect 16960 19168 16988 19264
rect 17126 19252 17132 19264
rect 17184 19252 17190 19304
rect 17586 19292 17592 19304
rect 17547 19264 17592 19292
rect 17586 19252 17592 19264
rect 17644 19292 17650 19304
rect 18248 19301 18276 19332
rect 18966 19320 18972 19332
rect 19024 19320 19030 19372
rect 21266 19360 21272 19372
rect 20732 19332 21272 19360
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 17644 19264 18061 19292
rect 17644 19252 17650 19264
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18049 19255 18107 19261
rect 18233 19295 18291 19301
rect 18233 19261 18245 19295
rect 18279 19261 18291 19295
rect 18506 19292 18512 19304
rect 18467 19264 18512 19292
rect 18233 19255 18291 19261
rect 18506 19252 18512 19264
rect 18564 19252 18570 19304
rect 18877 19295 18935 19301
rect 18877 19261 18889 19295
rect 18923 19261 18935 19295
rect 18984 19292 19012 19320
rect 19981 19295 20039 19301
rect 19981 19292 19993 19295
rect 18984 19264 19993 19292
rect 18877 19255 18935 19261
rect 19981 19261 19993 19264
rect 20027 19261 20039 19295
rect 20162 19292 20168 19304
rect 20123 19264 20168 19292
rect 19981 19255 20039 19261
rect 11241 19159 11299 19165
rect 10928 19128 10973 19156
rect 10928 19116 10934 19128
rect 11241 19125 11253 19159
rect 11287 19125 11299 19159
rect 11241 19119 11299 19125
rect 11330 19116 11336 19168
rect 11388 19156 11394 19168
rect 11701 19159 11759 19165
rect 11701 19156 11713 19159
rect 11388 19128 11713 19156
rect 11388 19116 11394 19128
rect 11701 19125 11713 19128
rect 11747 19125 11759 19159
rect 11701 19119 11759 19125
rect 12802 19116 12808 19168
rect 12860 19156 12866 19168
rect 13173 19159 13231 19165
rect 13173 19156 13185 19159
rect 12860 19128 13185 19156
rect 12860 19116 12866 19128
rect 13173 19125 13185 19128
rect 13219 19125 13231 19159
rect 13173 19119 13231 19125
rect 13262 19116 13268 19168
rect 13320 19156 13326 19168
rect 13541 19159 13599 19165
rect 13541 19156 13553 19159
rect 13320 19128 13553 19156
rect 13320 19116 13326 19128
rect 13541 19125 13553 19128
rect 13587 19125 13599 19159
rect 13541 19119 13599 19125
rect 13630 19116 13636 19168
rect 13688 19156 13694 19168
rect 13909 19159 13967 19165
rect 13909 19156 13921 19159
rect 13688 19128 13921 19156
rect 13688 19116 13694 19128
rect 13909 19125 13921 19128
rect 13955 19125 13967 19159
rect 14366 19156 14372 19168
rect 14327 19128 14372 19156
rect 13909 19119 13967 19125
rect 14366 19116 14372 19128
rect 14424 19116 14430 19168
rect 14734 19156 14740 19168
rect 14695 19128 14740 19156
rect 14734 19116 14740 19128
rect 14792 19116 14798 19168
rect 15286 19156 15292 19168
rect 15247 19128 15292 19156
rect 15286 19116 15292 19128
rect 15344 19116 15350 19168
rect 16298 19156 16304 19168
rect 16259 19128 16304 19156
rect 16298 19116 16304 19128
rect 16356 19116 16362 19168
rect 16666 19156 16672 19168
rect 16627 19128 16672 19156
rect 16666 19116 16672 19128
rect 16724 19116 16730 19168
rect 16942 19156 16948 19168
rect 16903 19128 16948 19156
rect 16942 19116 16948 19128
rect 17000 19116 17006 19168
rect 17313 19159 17371 19165
rect 17313 19125 17325 19159
rect 17359 19156 17371 19159
rect 17402 19156 17408 19168
rect 17359 19128 17408 19156
rect 17359 19125 17371 19128
rect 17313 19119 17371 19125
rect 17402 19116 17408 19128
rect 17460 19116 17466 19168
rect 17770 19156 17776 19168
rect 17731 19128 17776 19156
rect 17770 19116 17776 19128
rect 17828 19116 17834 19168
rect 18892 19156 18920 19255
rect 20162 19252 20168 19264
rect 20220 19252 20226 19304
rect 20438 19292 20444 19304
rect 20399 19264 20444 19292
rect 20438 19252 20444 19264
rect 20496 19252 20502 19304
rect 20622 19252 20628 19304
rect 20680 19292 20686 19304
rect 20732 19301 20760 19332
rect 21266 19320 21272 19332
rect 21324 19320 21330 19372
rect 20717 19295 20775 19301
rect 20717 19292 20729 19295
rect 20680 19264 20729 19292
rect 20680 19252 20686 19264
rect 20717 19261 20729 19264
rect 20763 19261 20775 19295
rect 20990 19292 20996 19304
rect 20951 19264 20996 19292
rect 20717 19255 20775 19261
rect 20990 19252 20996 19264
rect 21048 19252 21054 19304
rect 18966 19184 18972 19236
rect 19024 19224 19030 19236
rect 19518 19224 19524 19236
rect 19024 19196 19524 19224
rect 19024 19184 19030 19196
rect 19518 19184 19524 19196
rect 19576 19184 19582 19236
rect 19610 19184 19616 19236
rect 19668 19224 19674 19236
rect 19705 19227 19763 19233
rect 19705 19224 19717 19227
rect 19668 19196 19717 19224
rect 19668 19184 19674 19196
rect 19705 19193 19717 19196
rect 19751 19193 19763 19227
rect 21453 19227 21511 19233
rect 21453 19224 21465 19227
rect 19705 19187 19763 19193
rect 20088 19196 21465 19224
rect 20088 19168 20116 19196
rect 21453 19193 21465 19196
rect 21499 19193 21511 19227
rect 21453 19187 21511 19193
rect 20070 19156 20076 19168
rect 18892 19128 20076 19156
rect 20070 19116 20076 19128
rect 20128 19116 20134 19168
rect 1104 19066 21896 19088
rect 1104 19014 7912 19066
rect 7964 19014 7976 19066
rect 8028 19014 8040 19066
rect 8092 19014 8104 19066
rect 8156 19014 14843 19066
rect 14895 19014 14907 19066
rect 14959 19014 14971 19066
rect 15023 19014 15035 19066
rect 15087 19014 21896 19066
rect 1104 18992 21896 19014
rect 1854 18912 1860 18964
rect 1912 18952 1918 18964
rect 1949 18955 2007 18961
rect 1949 18952 1961 18955
rect 1912 18924 1961 18952
rect 1912 18912 1918 18924
rect 1949 18921 1961 18924
rect 1995 18921 2007 18955
rect 3789 18955 3847 18961
rect 3789 18952 3801 18955
rect 1949 18915 2007 18921
rect 3068 18924 3801 18952
rect 566 18844 572 18896
rect 624 18884 630 18896
rect 3068 18884 3096 18924
rect 3789 18921 3801 18924
rect 3835 18952 3847 18955
rect 4709 18955 4767 18961
rect 4709 18952 4721 18955
rect 3835 18924 4721 18952
rect 3835 18921 3847 18924
rect 3789 18915 3847 18921
rect 4709 18921 4721 18924
rect 4755 18952 4767 18955
rect 5258 18952 5264 18964
rect 4755 18924 5264 18952
rect 4755 18921 4767 18924
rect 4709 18915 4767 18921
rect 5258 18912 5264 18924
rect 5316 18912 5322 18964
rect 5442 18952 5448 18964
rect 5403 18924 5448 18952
rect 5442 18912 5448 18924
rect 5500 18912 5506 18964
rect 5902 18952 5908 18964
rect 5863 18924 5908 18952
rect 5902 18912 5908 18924
rect 5960 18912 5966 18964
rect 6273 18955 6331 18961
rect 6273 18921 6285 18955
rect 6319 18952 6331 18955
rect 6362 18952 6368 18964
rect 6319 18924 6368 18952
rect 6319 18921 6331 18924
rect 6273 18915 6331 18921
rect 6362 18912 6368 18924
rect 6420 18912 6426 18964
rect 7098 18912 7104 18964
rect 7156 18952 7162 18964
rect 7193 18955 7251 18961
rect 7193 18952 7205 18955
rect 7156 18924 7205 18952
rect 7156 18912 7162 18924
rect 7193 18921 7205 18924
rect 7239 18921 7251 18955
rect 7193 18915 7251 18921
rect 7561 18955 7619 18961
rect 7561 18921 7573 18955
rect 7607 18952 7619 18955
rect 7650 18952 7656 18964
rect 7607 18924 7656 18952
rect 7607 18921 7619 18924
rect 7561 18915 7619 18921
rect 7650 18912 7656 18924
rect 7708 18912 7714 18964
rect 10134 18952 10140 18964
rect 10095 18924 10140 18952
rect 10134 18912 10140 18924
rect 10192 18912 10198 18964
rect 11606 18912 11612 18964
rect 11664 18952 11670 18964
rect 13538 18952 13544 18964
rect 11664 18924 13544 18952
rect 11664 18912 11670 18924
rect 13538 18912 13544 18924
rect 13596 18912 13602 18964
rect 15562 18912 15568 18964
rect 15620 18952 15626 18964
rect 16209 18955 16267 18961
rect 16209 18952 16221 18955
rect 15620 18924 16221 18952
rect 15620 18912 15626 18924
rect 16209 18921 16221 18924
rect 16255 18952 16267 18955
rect 19426 18952 19432 18964
rect 16255 18924 19432 18952
rect 16255 18921 16267 18924
rect 16209 18915 16267 18921
rect 19426 18912 19432 18924
rect 19484 18912 19490 18964
rect 19794 18952 19800 18964
rect 19755 18924 19800 18952
rect 19794 18912 19800 18924
rect 19852 18952 19858 18964
rect 19981 18955 20039 18961
rect 19981 18952 19993 18955
rect 19852 18924 19993 18952
rect 19852 18912 19858 18924
rect 19981 18921 19993 18924
rect 20027 18952 20039 18955
rect 20162 18952 20168 18964
rect 20027 18924 20168 18952
rect 20027 18921 20039 18924
rect 19981 18915 20039 18921
rect 20162 18912 20168 18924
rect 20220 18952 20226 18964
rect 21453 18955 21511 18961
rect 21453 18952 21465 18955
rect 20220 18924 21465 18952
rect 20220 18912 20226 18924
rect 624 18856 3096 18884
rect 5353 18887 5411 18893
rect 624 18844 630 18856
rect 5353 18853 5365 18887
rect 5399 18884 5411 18887
rect 5399 18856 6224 18884
rect 5399 18853 5411 18856
rect 5353 18847 5411 18853
rect 1765 18819 1823 18825
rect 1765 18785 1777 18819
rect 1811 18816 1823 18819
rect 2133 18819 2191 18825
rect 2133 18816 2145 18819
rect 1811 18788 2145 18816
rect 1811 18785 1823 18788
rect 1765 18779 1823 18785
rect 2133 18785 2145 18788
rect 2179 18785 2191 18819
rect 2133 18779 2191 18785
rect 2148 18748 2176 18779
rect 2222 18776 2228 18828
rect 2280 18816 2286 18828
rect 2866 18816 2872 18828
rect 2280 18788 2872 18816
rect 2280 18776 2286 18788
rect 2866 18776 2872 18788
rect 2924 18816 2930 18828
rect 3053 18819 3111 18825
rect 3053 18816 3065 18819
rect 2924 18788 3065 18816
rect 2924 18776 2930 18788
rect 3053 18785 3065 18788
rect 3099 18785 3111 18819
rect 5810 18816 5816 18828
rect 5771 18788 5816 18816
rect 3053 18779 3111 18785
rect 5810 18776 5816 18788
rect 5868 18776 5874 18828
rect 6196 18760 6224 18856
rect 6730 18844 6736 18896
rect 6788 18884 6794 18896
rect 8021 18887 8079 18893
rect 8021 18884 8033 18887
rect 6788 18856 8033 18884
rect 6788 18844 6794 18856
rect 8021 18853 8033 18856
rect 8067 18884 8079 18887
rect 8665 18887 8723 18893
rect 8665 18884 8677 18887
rect 8067 18856 8677 18884
rect 8067 18853 8079 18856
rect 8021 18847 8079 18853
rect 8665 18853 8677 18856
rect 8711 18884 8723 18887
rect 8846 18884 8852 18896
rect 8711 18856 8852 18884
rect 8711 18853 8723 18856
rect 8665 18847 8723 18853
rect 8846 18844 8852 18856
rect 8904 18844 8910 18896
rect 17037 18887 17095 18893
rect 17037 18853 17049 18887
rect 17083 18884 17095 18887
rect 17126 18884 17132 18896
rect 17083 18856 17132 18884
rect 17083 18853 17095 18856
rect 17037 18847 17095 18853
rect 17126 18844 17132 18856
rect 17184 18884 17190 18896
rect 17862 18884 17868 18896
rect 17184 18856 17868 18884
rect 17184 18844 17190 18856
rect 17862 18844 17868 18856
rect 17920 18844 17926 18896
rect 17957 18887 18015 18893
rect 17957 18853 17969 18887
rect 18003 18884 18015 18887
rect 18966 18884 18972 18896
rect 18003 18856 18972 18884
rect 18003 18853 18015 18856
rect 17957 18847 18015 18853
rect 6638 18816 6644 18828
rect 6599 18788 6644 18816
rect 6638 18776 6644 18788
rect 6696 18776 6702 18828
rect 7653 18819 7711 18825
rect 7653 18785 7665 18819
rect 7699 18816 7711 18819
rect 8386 18816 8392 18828
rect 7699 18788 8392 18816
rect 7699 18785 7711 18788
rect 7653 18779 7711 18785
rect 8386 18776 8392 18788
rect 8444 18776 8450 18828
rect 8573 18819 8631 18825
rect 8573 18785 8585 18819
rect 8619 18785 8631 18819
rect 10864 18819 10922 18825
rect 10864 18816 10876 18819
rect 8573 18779 8631 18785
rect 10428 18788 10876 18816
rect 2406 18748 2412 18760
rect 2148 18720 2412 18748
rect 2406 18708 2412 18720
rect 2464 18708 2470 18760
rect 2682 18708 2688 18760
rect 2740 18748 2746 18760
rect 2961 18751 3019 18757
rect 2961 18748 2973 18751
rect 2740 18720 2973 18748
rect 2740 18708 2746 18720
rect 2961 18717 2973 18720
rect 3007 18717 3019 18751
rect 4154 18748 4160 18760
rect 4115 18720 4160 18748
rect 2961 18711 3019 18717
rect 4154 18708 4160 18720
rect 4212 18748 4218 18760
rect 4801 18751 4859 18757
rect 4801 18748 4813 18751
rect 4212 18720 4813 18748
rect 4212 18708 4218 18720
rect 4801 18717 4813 18720
rect 4847 18717 4859 18751
rect 4982 18748 4988 18760
rect 4943 18720 4988 18748
rect 4801 18711 4859 18717
rect 1670 18640 1676 18692
rect 1728 18680 1734 18692
rect 4062 18680 4068 18692
rect 1728 18652 4068 18680
rect 1728 18640 1734 18652
rect 4062 18640 4068 18652
rect 4120 18640 4126 18692
rect 4816 18680 4844 18711
rect 4982 18708 4988 18720
rect 5040 18708 5046 18760
rect 6089 18751 6147 18757
rect 6089 18717 6101 18751
rect 6135 18717 6147 18751
rect 6089 18711 6147 18717
rect 5902 18680 5908 18692
rect 4816 18652 5908 18680
rect 5902 18640 5908 18652
rect 5960 18640 5966 18692
rect 6104 18680 6132 18711
rect 6178 18708 6184 18760
rect 6236 18748 6242 18760
rect 6733 18751 6791 18757
rect 6733 18748 6745 18751
rect 6236 18720 6745 18748
rect 6236 18708 6242 18720
rect 6733 18717 6745 18720
rect 6779 18717 6791 18751
rect 6733 18711 6791 18717
rect 6914 18708 6920 18760
rect 6972 18748 6978 18760
rect 7745 18751 7803 18757
rect 7745 18748 7757 18751
rect 6972 18720 7757 18748
rect 6972 18708 6978 18720
rect 7745 18717 7757 18720
rect 7791 18717 7803 18751
rect 7745 18711 7803 18717
rect 8110 18708 8116 18760
rect 8168 18748 8174 18760
rect 8588 18748 8616 18779
rect 8846 18748 8852 18760
rect 8168 18720 8616 18748
rect 8807 18720 8852 18748
rect 8168 18708 8174 18720
rect 8846 18708 8852 18720
rect 8904 18708 8910 18760
rect 10226 18748 10232 18760
rect 10187 18720 10232 18748
rect 10226 18708 10232 18720
rect 10284 18708 10290 18760
rect 10428 18757 10456 18788
rect 10864 18785 10876 18788
rect 10910 18816 10922 18819
rect 11146 18816 11152 18828
rect 10910 18788 11152 18816
rect 10910 18785 10922 18788
rect 10864 18779 10922 18785
rect 11146 18776 11152 18788
rect 11204 18776 11210 18828
rect 11238 18776 11244 18828
rect 11296 18816 11302 18828
rect 11296 18788 11652 18816
rect 11296 18776 11302 18788
rect 10413 18751 10471 18757
rect 10413 18717 10425 18751
rect 10459 18717 10471 18751
rect 10413 18711 10471 18717
rect 10597 18751 10655 18757
rect 10597 18717 10609 18751
rect 10643 18717 10655 18751
rect 11624 18748 11652 18788
rect 12066 18776 12072 18828
rect 12124 18816 12130 18828
rect 17586 18816 17592 18828
rect 12124 18788 17592 18816
rect 12124 18776 12130 18788
rect 17586 18776 17592 18788
rect 17644 18776 17650 18828
rect 18064 18825 18092 18856
rect 18966 18844 18972 18856
rect 19024 18844 19030 18896
rect 19242 18844 19248 18896
rect 19300 18884 19306 18896
rect 20533 18887 20591 18893
rect 20533 18884 20545 18887
rect 19300 18856 20545 18884
rect 19300 18844 19306 18856
rect 20533 18853 20545 18856
rect 20579 18853 20591 18887
rect 20533 18847 20591 18853
rect 18049 18819 18107 18825
rect 18049 18785 18061 18819
rect 18095 18816 18107 18819
rect 18601 18819 18659 18825
rect 18095 18788 18129 18816
rect 18095 18785 18107 18788
rect 18049 18779 18107 18785
rect 18601 18785 18613 18819
rect 18647 18785 18659 18819
rect 18601 18779 18659 18785
rect 19153 18819 19211 18825
rect 19153 18785 19165 18819
rect 19199 18816 19211 18819
rect 20257 18819 20315 18825
rect 20257 18816 20269 18819
rect 19199 18788 20269 18816
rect 19199 18785 19211 18788
rect 19153 18779 19211 18785
rect 20257 18785 20269 18788
rect 20303 18816 20315 18819
rect 20714 18816 20720 18828
rect 20303 18788 20720 18816
rect 20303 18785 20315 18788
rect 20257 18779 20315 18785
rect 12805 18751 12863 18757
rect 12805 18748 12817 18751
rect 11624 18720 12817 18748
rect 10597 18711 10655 18717
rect 12805 18717 12817 18720
rect 12851 18748 12863 18751
rect 12986 18748 12992 18760
rect 12851 18720 12992 18748
rect 12851 18717 12863 18720
rect 12805 18711 12863 18717
rect 7190 18680 7196 18692
rect 6104 18652 7196 18680
rect 7190 18640 7196 18652
rect 7248 18640 7254 18692
rect 8754 18680 8760 18692
rect 8128 18652 8760 18680
rect 2498 18572 2504 18624
rect 2556 18612 2562 18624
rect 2685 18615 2743 18621
rect 2685 18612 2697 18615
rect 2556 18584 2697 18612
rect 2556 18572 2562 18584
rect 2685 18581 2697 18584
rect 2731 18581 2743 18615
rect 2685 18575 2743 18581
rect 3326 18572 3332 18624
rect 3384 18612 3390 18624
rect 3786 18612 3792 18624
rect 3384 18584 3792 18612
rect 3384 18572 3390 18584
rect 3786 18572 3792 18584
rect 3844 18572 3850 18624
rect 4338 18612 4344 18624
rect 4299 18584 4344 18612
rect 4338 18572 4344 18584
rect 4396 18572 4402 18624
rect 4982 18572 4988 18624
rect 5040 18612 5046 18624
rect 8128 18612 8156 18652
rect 8754 18640 8760 18652
rect 8812 18640 8818 18692
rect 9769 18683 9827 18689
rect 9769 18649 9781 18683
rect 9815 18680 9827 18683
rect 9858 18680 9864 18692
rect 9815 18652 9864 18680
rect 9815 18649 9827 18652
rect 9769 18643 9827 18649
rect 9858 18640 9864 18652
rect 9916 18640 9922 18692
rect 5040 18584 8156 18612
rect 8205 18615 8263 18621
rect 5040 18572 5046 18584
rect 8205 18581 8217 18615
rect 8251 18612 8263 18615
rect 10410 18612 10416 18624
rect 8251 18584 10416 18612
rect 8251 18581 8263 18584
rect 8205 18575 8263 18581
rect 10410 18572 10416 18584
rect 10468 18572 10474 18624
rect 10612 18612 10640 18711
rect 12986 18708 12992 18720
rect 13044 18708 13050 18760
rect 18230 18748 18236 18760
rect 18191 18720 18236 18748
rect 18230 18708 18236 18720
rect 18288 18708 18294 18760
rect 12066 18640 12072 18692
rect 12124 18680 12130 18692
rect 13173 18683 13231 18689
rect 13173 18680 13185 18683
rect 12124 18652 13185 18680
rect 12124 18640 12130 18652
rect 13173 18649 13185 18652
rect 13219 18680 13231 18683
rect 13354 18680 13360 18692
rect 13219 18652 13360 18680
rect 13219 18649 13231 18652
rect 13173 18643 13231 18649
rect 13354 18640 13360 18652
rect 13412 18640 13418 18692
rect 18616 18680 18644 18779
rect 20714 18776 20720 18788
rect 20772 18776 20778 18828
rect 20916 18825 20944 18924
rect 21453 18921 21465 18924
rect 21499 18921 21511 18955
rect 21453 18915 21511 18921
rect 21177 18887 21235 18893
rect 21177 18853 21189 18887
rect 21223 18884 21235 18887
rect 22002 18884 22008 18896
rect 21223 18856 22008 18884
rect 21223 18853 21235 18856
rect 21177 18847 21235 18853
rect 22002 18844 22008 18856
rect 22060 18844 22066 18896
rect 20901 18819 20959 18825
rect 20901 18785 20913 18819
rect 20947 18785 20959 18819
rect 20901 18779 20959 18785
rect 18782 18748 18788 18760
rect 18743 18720 18788 18748
rect 18782 18708 18788 18720
rect 18840 18708 18846 18760
rect 19334 18748 19340 18760
rect 19295 18720 19340 18748
rect 19334 18708 19340 18720
rect 19392 18708 19398 18760
rect 19794 18680 19800 18692
rect 18616 18652 19800 18680
rect 19794 18640 19800 18652
rect 19852 18640 19858 18692
rect 11790 18612 11796 18624
rect 10612 18584 11796 18612
rect 11790 18572 11796 18584
rect 11848 18572 11854 18624
rect 11974 18612 11980 18624
rect 11935 18584 11980 18612
rect 11974 18572 11980 18584
rect 12032 18572 12038 18624
rect 13630 18612 13636 18624
rect 13591 18584 13636 18612
rect 13630 18572 13636 18584
rect 13688 18572 13694 18624
rect 14093 18615 14151 18621
rect 14093 18581 14105 18615
rect 14139 18612 14151 18615
rect 14182 18612 14188 18624
rect 14139 18584 14188 18612
rect 14139 18581 14151 18584
rect 14093 18575 14151 18581
rect 14182 18572 14188 18584
rect 14240 18572 14246 18624
rect 14458 18612 14464 18624
rect 14419 18584 14464 18612
rect 14458 18572 14464 18584
rect 14516 18572 14522 18624
rect 15562 18572 15568 18624
rect 15620 18612 15626 18624
rect 15933 18615 15991 18621
rect 15933 18612 15945 18615
rect 15620 18584 15945 18612
rect 15620 18572 15626 18584
rect 15933 18581 15945 18584
rect 15979 18612 15991 18615
rect 16022 18612 16028 18624
rect 15979 18584 16028 18612
rect 15979 18581 15991 18584
rect 15933 18575 15991 18581
rect 16022 18572 16028 18584
rect 16080 18572 16086 18624
rect 18598 18572 18604 18624
rect 18656 18612 18662 18624
rect 20530 18612 20536 18624
rect 18656 18584 20536 18612
rect 18656 18572 18662 18584
rect 20530 18572 20536 18584
rect 20588 18572 20594 18624
rect 1104 18522 21896 18544
rect 1104 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 4575 18522
rect 4627 18470 4639 18522
rect 4691 18470 11378 18522
rect 11430 18470 11442 18522
rect 11494 18470 11506 18522
rect 11558 18470 11570 18522
rect 11622 18470 18308 18522
rect 18360 18470 18372 18522
rect 18424 18470 18436 18522
rect 18488 18470 18500 18522
rect 18552 18470 21896 18522
rect 1104 18448 21896 18470
rect 2317 18411 2375 18417
rect 2317 18377 2329 18411
rect 2363 18408 2375 18411
rect 2774 18408 2780 18420
rect 2363 18380 2780 18408
rect 2363 18377 2375 18380
rect 2317 18371 2375 18377
rect 2774 18368 2780 18380
rect 2832 18368 2838 18420
rect 4154 18368 4160 18420
rect 4212 18408 4218 18420
rect 4893 18411 4951 18417
rect 4893 18408 4905 18411
rect 4212 18380 4905 18408
rect 4212 18368 4218 18380
rect 4893 18377 4905 18380
rect 4939 18408 4951 18411
rect 4982 18408 4988 18420
rect 4939 18380 4988 18408
rect 4939 18377 4951 18380
rect 4893 18371 4951 18377
rect 4982 18368 4988 18380
rect 5040 18368 5046 18420
rect 5810 18368 5816 18420
rect 5868 18408 5874 18420
rect 7377 18411 7435 18417
rect 7377 18408 7389 18411
rect 5868 18380 7389 18408
rect 5868 18368 5874 18380
rect 7377 18377 7389 18380
rect 7423 18377 7435 18411
rect 7377 18371 7435 18377
rect 7558 18368 7564 18420
rect 7616 18408 7622 18420
rect 8110 18408 8116 18420
rect 7616 18380 8116 18408
rect 7616 18368 7622 18380
rect 8110 18368 8116 18380
rect 8168 18408 8174 18420
rect 8205 18411 8263 18417
rect 8205 18408 8217 18411
rect 8168 18380 8217 18408
rect 8168 18368 8174 18380
rect 8205 18377 8217 18380
rect 8251 18377 8263 18411
rect 8205 18371 8263 18377
rect 8846 18368 8852 18420
rect 8904 18408 8910 18420
rect 16669 18411 16727 18417
rect 8904 18380 11284 18408
rect 8904 18368 8910 18380
rect 3050 18300 3056 18352
rect 3108 18340 3114 18352
rect 7190 18340 7196 18352
rect 3108 18312 6500 18340
rect 3108 18300 3114 18312
rect 934 18232 940 18284
rect 992 18272 998 18284
rect 3697 18275 3755 18281
rect 992 18244 3648 18272
rect 992 18232 998 18244
rect 1765 18207 1823 18213
rect 1765 18173 1777 18207
rect 1811 18173 1823 18207
rect 2130 18204 2136 18216
rect 2091 18176 2136 18204
rect 1765 18167 1823 18173
rect 1780 18136 1808 18167
rect 2130 18164 2136 18176
rect 2188 18164 2194 18216
rect 2501 18207 2559 18213
rect 2501 18173 2513 18207
rect 2547 18204 2559 18207
rect 2682 18204 2688 18216
rect 2547 18176 2688 18204
rect 2547 18173 2559 18176
rect 2501 18167 2559 18173
rect 2682 18164 2688 18176
rect 2740 18164 2746 18216
rect 3142 18164 3148 18216
rect 3200 18204 3206 18216
rect 3421 18207 3479 18213
rect 3421 18204 3433 18207
rect 3200 18176 3433 18204
rect 3200 18164 3206 18176
rect 3421 18173 3433 18176
rect 3467 18173 3479 18207
rect 3421 18167 3479 18173
rect 1780 18108 2912 18136
rect 2884 18080 2912 18108
rect 2958 18096 2964 18148
rect 3016 18136 3022 18148
rect 3513 18139 3571 18145
rect 3513 18136 3525 18139
rect 3016 18108 3525 18136
rect 3016 18096 3022 18108
rect 3513 18105 3525 18108
rect 3559 18105 3571 18139
rect 3620 18136 3648 18244
rect 3697 18241 3709 18275
rect 3743 18272 3755 18275
rect 4525 18275 4583 18281
rect 4525 18272 4537 18275
rect 3743 18244 4537 18272
rect 3743 18241 3755 18244
rect 3697 18235 3755 18241
rect 4525 18241 4537 18244
rect 4571 18272 4583 18275
rect 4614 18272 4620 18284
rect 4571 18244 4620 18272
rect 4571 18241 4583 18244
rect 4525 18235 4583 18241
rect 4614 18232 4620 18244
rect 4672 18272 4678 18284
rect 5074 18272 5080 18284
rect 4672 18244 5080 18272
rect 4672 18232 4678 18244
rect 5074 18232 5080 18244
rect 5132 18232 5138 18284
rect 6086 18232 6092 18284
rect 6144 18272 6150 18284
rect 6365 18275 6423 18281
rect 6365 18272 6377 18275
rect 6144 18244 6377 18272
rect 6144 18232 6150 18244
rect 6365 18241 6377 18244
rect 6411 18241 6423 18275
rect 6365 18235 6423 18241
rect 4338 18204 4344 18216
rect 4299 18176 4344 18204
rect 4338 18164 4344 18176
rect 4396 18164 4402 18216
rect 6270 18204 6276 18216
rect 6231 18176 6276 18204
rect 6270 18164 6276 18176
rect 6328 18164 6334 18216
rect 6472 18204 6500 18312
rect 6564 18312 7196 18340
rect 6564 18281 6592 18312
rect 7190 18300 7196 18312
rect 7248 18300 7254 18352
rect 10045 18343 10103 18349
rect 10045 18309 10057 18343
rect 10091 18309 10103 18343
rect 11256 18340 11284 18380
rect 16669 18377 16681 18411
rect 16715 18408 16727 18411
rect 17034 18408 17040 18420
rect 16715 18380 17040 18408
rect 16715 18377 16727 18380
rect 16669 18371 16727 18377
rect 17034 18368 17040 18380
rect 17092 18368 17098 18420
rect 18690 18408 18696 18420
rect 18651 18380 18696 18408
rect 18690 18368 18696 18380
rect 18748 18368 18754 18420
rect 19702 18408 19708 18420
rect 19663 18380 19708 18408
rect 19702 18368 19708 18380
rect 19760 18368 19766 18420
rect 19981 18411 20039 18417
rect 19981 18377 19993 18411
rect 20027 18408 20039 18411
rect 20257 18411 20315 18417
rect 20257 18408 20269 18411
rect 20027 18380 20269 18408
rect 20027 18377 20039 18380
rect 19981 18371 20039 18377
rect 20257 18377 20269 18380
rect 20303 18408 20315 18411
rect 20714 18408 20720 18420
rect 20303 18380 20720 18408
rect 20303 18377 20315 18380
rect 20257 18371 20315 18377
rect 20714 18368 20720 18380
rect 20772 18368 20778 18420
rect 21450 18408 21456 18420
rect 21411 18380 21456 18408
rect 21450 18368 21456 18380
rect 21508 18368 21514 18420
rect 11330 18340 11336 18352
rect 11256 18312 11336 18340
rect 10045 18303 10103 18309
rect 6549 18275 6607 18281
rect 6549 18241 6561 18275
rect 6595 18241 6607 18275
rect 6549 18235 6607 18241
rect 6638 18232 6644 18284
rect 6696 18272 6702 18284
rect 6825 18275 6883 18281
rect 6825 18272 6837 18275
rect 6696 18244 6837 18272
rect 6696 18232 6702 18244
rect 6825 18241 6837 18244
rect 6871 18241 6883 18275
rect 6825 18235 6883 18241
rect 6914 18232 6920 18284
rect 6972 18272 6978 18284
rect 7929 18275 7987 18281
rect 7929 18272 7941 18275
rect 6972 18244 7941 18272
rect 6972 18232 6978 18244
rect 7929 18241 7941 18244
rect 7975 18241 7987 18275
rect 10060 18272 10088 18303
rect 11330 18300 11336 18312
rect 11388 18300 11394 18352
rect 20162 18300 20168 18352
rect 20220 18340 20226 18352
rect 20349 18343 20407 18349
rect 20349 18340 20361 18343
rect 20220 18312 20361 18340
rect 20220 18300 20226 18312
rect 20349 18309 20361 18312
rect 20395 18309 20407 18343
rect 20349 18303 20407 18309
rect 7929 18235 7987 18241
rect 8036 18244 8791 18272
rect 10060 18244 10272 18272
rect 8036 18204 8064 18244
rect 8662 18204 8668 18216
rect 6472 18176 8064 18204
rect 8623 18176 8668 18204
rect 8662 18164 8668 18176
rect 8720 18164 8726 18216
rect 8763 18204 8791 18244
rect 9858 18204 9864 18216
rect 8763 18176 9864 18204
rect 9858 18164 9864 18176
rect 9916 18164 9922 18216
rect 10134 18204 10140 18216
rect 10095 18176 10140 18204
rect 10134 18164 10140 18176
rect 10192 18164 10198 18216
rect 10244 18204 10272 18244
rect 11790 18232 11796 18284
rect 11848 18272 11854 18284
rect 12434 18272 12440 18284
rect 11848 18244 12440 18272
rect 11848 18232 11854 18244
rect 12434 18232 12440 18244
rect 12492 18232 12498 18284
rect 14185 18275 14243 18281
rect 14185 18241 14197 18275
rect 14231 18272 14243 18275
rect 14550 18272 14556 18284
rect 14231 18244 14556 18272
rect 14231 18241 14243 18244
rect 14185 18235 14243 18241
rect 14550 18232 14556 18244
rect 14608 18232 14614 18284
rect 10404 18207 10462 18213
rect 10404 18204 10416 18207
rect 10244 18176 10416 18204
rect 10404 18173 10416 18176
rect 10450 18204 10462 18207
rect 10778 18204 10784 18216
rect 10450 18176 10784 18204
rect 10450 18173 10462 18176
rect 10404 18167 10462 18173
rect 10778 18164 10784 18176
rect 10836 18204 10842 18216
rect 10962 18204 10968 18216
rect 10836 18176 10968 18204
rect 10836 18164 10842 18176
rect 10962 18164 10968 18176
rect 11020 18164 11026 18216
rect 11514 18164 11520 18216
rect 11572 18204 11578 18216
rect 11609 18207 11667 18213
rect 11609 18204 11621 18207
rect 11572 18176 11621 18204
rect 11572 18164 11578 18176
rect 11609 18173 11621 18176
rect 11655 18173 11667 18207
rect 12158 18204 12164 18216
rect 11609 18167 11667 18173
rect 11716 18176 12164 18204
rect 4249 18139 4307 18145
rect 4249 18136 4261 18139
rect 3620 18108 4261 18136
rect 3513 18099 3571 18105
rect 4249 18105 4261 18108
rect 4295 18105 4307 18139
rect 4249 18099 4307 18105
rect 1946 18068 1952 18080
rect 1907 18040 1952 18068
rect 1946 18028 1952 18040
rect 2004 18028 2010 18080
rect 2590 18028 2596 18080
rect 2648 18068 2654 18080
rect 2685 18071 2743 18077
rect 2685 18068 2697 18071
rect 2648 18040 2697 18068
rect 2648 18028 2654 18040
rect 2685 18037 2697 18040
rect 2731 18037 2743 18071
rect 2866 18068 2872 18080
rect 2827 18040 2872 18068
rect 2685 18031 2743 18037
rect 2866 18028 2872 18040
rect 2924 18028 2930 18080
rect 3050 18068 3056 18080
rect 3011 18040 3056 18068
rect 3050 18028 3056 18040
rect 3108 18028 3114 18080
rect 3878 18068 3884 18080
rect 3839 18040 3884 18068
rect 3878 18028 3884 18040
rect 3936 18028 3942 18080
rect 4264 18068 4292 18099
rect 4430 18096 4436 18148
rect 4488 18136 4494 18148
rect 5077 18139 5135 18145
rect 5077 18136 5089 18139
rect 4488 18108 5089 18136
rect 4488 18096 4494 18108
rect 5077 18105 5089 18108
rect 5123 18136 5135 18139
rect 5626 18136 5632 18148
rect 5123 18108 5632 18136
rect 5123 18105 5135 18108
rect 5077 18099 5135 18105
rect 5626 18096 5632 18108
rect 5684 18096 5690 18148
rect 7837 18139 7895 18145
rect 7837 18105 7849 18139
rect 7883 18136 7895 18139
rect 8754 18136 8760 18148
rect 7883 18108 8760 18136
rect 7883 18105 7895 18108
rect 7837 18099 7895 18105
rect 8754 18096 8760 18108
rect 8812 18096 8818 18148
rect 8846 18096 8852 18148
rect 8904 18145 8910 18148
rect 8904 18139 8968 18145
rect 8904 18105 8922 18139
rect 8956 18105 8968 18139
rect 8904 18099 8968 18105
rect 8904 18096 8910 18099
rect 10318 18096 10324 18148
rect 10376 18136 10382 18148
rect 11716 18136 11744 18176
rect 12158 18164 12164 18176
rect 12216 18164 12222 18216
rect 13906 18204 13912 18216
rect 13867 18176 13912 18204
rect 13906 18164 13912 18176
rect 13964 18164 13970 18216
rect 16482 18204 16488 18216
rect 16443 18176 16488 18204
rect 16482 18164 16488 18176
rect 16540 18164 16546 18216
rect 18046 18164 18052 18216
rect 18104 18204 18110 18216
rect 18417 18207 18475 18213
rect 18417 18204 18429 18207
rect 18104 18176 18429 18204
rect 18104 18164 18110 18176
rect 18417 18173 18429 18176
rect 18463 18204 18475 18207
rect 18509 18207 18567 18213
rect 18509 18204 18521 18207
rect 18463 18176 18521 18204
rect 18463 18173 18475 18176
rect 18417 18167 18475 18173
rect 18509 18173 18521 18176
rect 18555 18173 18567 18207
rect 19521 18207 19579 18213
rect 19521 18204 19533 18207
rect 18509 18167 18567 18173
rect 19352 18176 19533 18204
rect 10376 18108 11744 18136
rect 10376 18096 10382 18108
rect 11974 18096 11980 18148
rect 12032 18136 12038 18148
rect 12682 18139 12740 18145
rect 12682 18136 12694 18139
rect 12032 18108 12694 18136
rect 12032 18096 12038 18108
rect 12682 18105 12694 18108
rect 12728 18105 12740 18139
rect 12682 18099 12740 18105
rect 19352 18080 19380 18176
rect 19521 18173 19533 18176
rect 19567 18173 19579 18207
rect 20364 18204 20392 18303
rect 20717 18207 20775 18213
rect 20717 18204 20729 18207
rect 20364 18176 20729 18204
rect 19521 18167 19579 18173
rect 20717 18173 20729 18176
rect 20763 18173 20775 18207
rect 20717 18167 20775 18173
rect 21269 18207 21327 18213
rect 21269 18173 21281 18207
rect 21315 18173 21327 18207
rect 21269 18167 21327 18173
rect 20898 18096 20904 18148
rect 20956 18136 20962 18148
rect 20993 18139 21051 18145
rect 20993 18136 21005 18139
rect 20956 18108 21005 18136
rect 20956 18096 20962 18108
rect 20993 18105 21005 18108
rect 21039 18105 21051 18139
rect 20993 18099 21051 18105
rect 4709 18071 4767 18077
rect 4709 18068 4721 18071
rect 4264 18040 4721 18068
rect 4709 18037 4721 18040
rect 4755 18068 4767 18071
rect 5258 18068 5264 18080
rect 4755 18040 5264 18068
rect 4755 18037 4767 18040
rect 4709 18031 4767 18037
rect 5258 18028 5264 18040
rect 5316 18028 5322 18080
rect 5905 18071 5963 18077
rect 5905 18037 5917 18071
rect 5951 18068 5963 18071
rect 7282 18068 7288 18080
rect 5951 18040 7288 18068
rect 5951 18037 5963 18040
rect 5905 18031 5963 18037
rect 7282 18028 7288 18040
rect 7340 18028 7346 18080
rect 7742 18068 7748 18080
rect 7703 18040 7748 18068
rect 7742 18028 7748 18040
rect 7800 18028 7806 18080
rect 8662 18028 8668 18080
rect 8720 18068 8726 18080
rect 9306 18068 9312 18080
rect 8720 18040 9312 18068
rect 8720 18028 8726 18040
rect 9306 18028 9312 18040
rect 9364 18068 9370 18080
rect 10134 18068 10140 18080
rect 9364 18040 10140 18068
rect 9364 18028 9370 18040
rect 10134 18028 10140 18040
rect 10192 18028 10198 18080
rect 11146 18028 11152 18080
rect 11204 18068 11210 18080
rect 11517 18071 11575 18077
rect 11517 18068 11529 18071
rect 11204 18040 11529 18068
rect 11204 18028 11210 18040
rect 11517 18037 11529 18040
rect 11563 18068 11575 18071
rect 12158 18068 12164 18080
rect 11563 18040 12164 18068
rect 11563 18037 11575 18040
rect 11517 18031 11575 18037
rect 12158 18028 12164 18040
rect 12216 18028 12222 18080
rect 12802 18028 12808 18080
rect 12860 18068 12866 18080
rect 13817 18071 13875 18077
rect 13817 18068 13829 18071
rect 12860 18040 13829 18068
rect 12860 18028 12866 18040
rect 13817 18037 13829 18040
rect 13863 18037 13875 18071
rect 19334 18068 19340 18080
rect 19295 18040 19340 18068
rect 13817 18031 13875 18037
rect 19334 18028 19340 18040
rect 19392 18028 19398 18080
rect 19978 18028 19984 18080
rect 20036 18068 20042 18080
rect 20533 18071 20591 18077
rect 20533 18068 20545 18071
rect 20036 18040 20545 18068
rect 20036 18028 20042 18040
rect 20533 18037 20545 18040
rect 20579 18068 20591 18071
rect 21284 18068 21312 18167
rect 20579 18040 21312 18068
rect 20579 18037 20591 18040
rect 20533 18031 20591 18037
rect 1104 17978 21896 18000
rect 1104 17926 7912 17978
rect 7964 17926 7976 17978
rect 8028 17926 8040 17978
rect 8092 17926 8104 17978
rect 8156 17926 14843 17978
rect 14895 17926 14907 17978
rect 14959 17926 14971 17978
rect 15023 17926 15035 17978
rect 15087 17926 21896 17978
rect 1104 17904 21896 17926
rect 1578 17864 1584 17876
rect 1539 17836 1584 17864
rect 1578 17824 1584 17836
rect 1636 17824 1642 17876
rect 2777 17867 2835 17873
rect 2777 17833 2789 17867
rect 2823 17864 2835 17867
rect 3050 17864 3056 17876
rect 2823 17836 3056 17864
rect 2823 17833 2835 17836
rect 2777 17827 2835 17833
rect 3050 17824 3056 17836
rect 3108 17824 3114 17876
rect 3605 17867 3663 17873
rect 3605 17833 3617 17867
rect 3651 17864 3663 17867
rect 3878 17864 3884 17876
rect 3651 17836 3884 17864
rect 3651 17833 3663 17836
rect 3605 17827 3663 17833
rect 3878 17824 3884 17836
rect 3936 17824 3942 17876
rect 4065 17867 4123 17873
rect 4065 17833 4077 17867
rect 4111 17833 4123 17867
rect 4065 17827 4123 17833
rect 2041 17799 2099 17805
rect 2041 17765 2053 17799
rect 2087 17796 2099 17799
rect 2130 17796 2136 17808
rect 2087 17768 2136 17796
rect 2087 17765 2099 17768
rect 2041 17759 2099 17765
rect 2130 17756 2136 17768
rect 2188 17756 2194 17808
rect 3513 17799 3571 17805
rect 3513 17765 3525 17799
rect 3559 17796 3571 17799
rect 4080 17796 4108 17827
rect 4154 17824 4160 17876
rect 4212 17864 4218 17876
rect 4430 17864 4436 17876
rect 4212 17836 4436 17864
rect 4212 17824 4218 17836
rect 4430 17824 4436 17836
rect 4488 17824 4494 17876
rect 4890 17864 4896 17876
rect 4851 17836 4896 17864
rect 4890 17824 4896 17836
rect 4948 17824 4954 17876
rect 6086 17824 6092 17876
rect 6144 17864 6150 17876
rect 6457 17867 6515 17873
rect 6457 17864 6469 17867
rect 6144 17836 6469 17864
rect 6144 17824 6150 17836
rect 6457 17833 6469 17836
rect 6503 17833 6515 17867
rect 6457 17827 6515 17833
rect 6822 17824 6828 17876
rect 6880 17824 6886 17876
rect 6914 17824 6920 17876
rect 6972 17864 6978 17876
rect 6972 17836 7017 17864
rect 6972 17824 6978 17836
rect 8386 17824 8392 17876
rect 8444 17824 8450 17876
rect 8846 17824 8852 17876
rect 8904 17864 8910 17876
rect 9122 17864 9128 17876
rect 8904 17836 9128 17864
rect 8904 17824 8910 17836
rect 9122 17824 9128 17836
rect 9180 17824 9186 17876
rect 9953 17867 10011 17873
rect 9953 17833 9965 17867
rect 9999 17864 10011 17867
rect 10226 17864 10232 17876
rect 9999 17836 10232 17864
rect 9999 17833 10011 17836
rect 9953 17827 10011 17833
rect 10226 17824 10232 17836
rect 10284 17824 10290 17876
rect 10410 17864 10416 17876
rect 10371 17836 10416 17864
rect 10410 17824 10416 17836
rect 10468 17824 10474 17876
rect 10781 17867 10839 17873
rect 10781 17833 10793 17867
rect 10827 17864 10839 17867
rect 10870 17864 10876 17876
rect 10827 17836 10876 17864
rect 10827 17833 10839 17836
rect 10781 17827 10839 17833
rect 10870 17824 10876 17836
rect 10928 17824 10934 17876
rect 11054 17824 11060 17876
rect 11112 17864 11118 17876
rect 11514 17864 11520 17876
rect 11112 17836 11520 17864
rect 11112 17824 11118 17836
rect 11514 17824 11520 17836
rect 11572 17824 11578 17876
rect 11609 17867 11667 17873
rect 11609 17833 11621 17867
rect 11655 17864 11667 17867
rect 11698 17864 11704 17876
rect 11655 17836 11704 17864
rect 11655 17833 11667 17836
rect 11609 17827 11667 17833
rect 11698 17824 11704 17836
rect 11756 17824 11762 17876
rect 11974 17864 11980 17876
rect 11935 17836 11980 17864
rect 11974 17824 11980 17836
rect 12032 17824 12038 17876
rect 13538 17864 13544 17876
rect 13499 17836 13544 17864
rect 13538 17824 13544 17836
rect 13596 17864 13602 17876
rect 14185 17867 14243 17873
rect 14185 17864 14197 17867
rect 13596 17836 14197 17864
rect 13596 17824 13602 17836
rect 14185 17833 14197 17836
rect 14231 17833 14243 17867
rect 20070 17864 20076 17876
rect 20031 17836 20076 17864
rect 14185 17827 14243 17833
rect 20070 17824 20076 17836
rect 20128 17824 20134 17876
rect 21266 17824 21272 17876
rect 21324 17864 21330 17876
rect 21453 17867 21511 17873
rect 21453 17864 21465 17867
rect 21324 17836 21465 17864
rect 21324 17824 21330 17836
rect 21453 17833 21465 17836
rect 21499 17833 21511 17867
rect 21453 17827 21511 17833
rect 5261 17799 5319 17805
rect 5261 17796 5273 17799
rect 3559 17768 4108 17796
rect 4264 17768 5273 17796
rect 3559 17765 3571 17768
rect 3513 17759 3571 17765
rect 1394 17728 1400 17740
rect 1355 17700 1400 17728
rect 1394 17688 1400 17700
rect 1452 17688 1458 17740
rect 1765 17731 1823 17737
rect 1765 17697 1777 17731
rect 1811 17697 1823 17731
rect 1765 17691 1823 17697
rect 2685 17731 2743 17737
rect 2685 17697 2697 17731
rect 2731 17728 2743 17731
rect 4154 17728 4160 17740
rect 2731 17700 4160 17728
rect 2731 17697 2743 17700
rect 2685 17691 2743 17697
rect 1780 17660 1808 17691
rect 4154 17688 4160 17700
rect 4212 17688 4218 17740
rect 2130 17660 2136 17672
rect 1780 17632 2136 17660
rect 2130 17620 2136 17632
rect 2188 17620 2194 17672
rect 2590 17620 2596 17672
rect 2648 17660 2654 17672
rect 2961 17663 3019 17669
rect 2961 17660 2973 17663
rect 2648 17632 2973 17660
rect 2648 17620 2654 17632
rect 2961 17629 2973 17632
rect 3007 17660 3019 17663
rect 3697 17663 3755 17669
rect 3697 17660 3709 17663
rect 3007 17632 3709 17660
rect 3007 17629 3019 17632
rect 2961 17623 3019 17629
rect 3697 17629 3709 17632
rect 3743 17629 3755 17663
rect 4264 17660 4292 17768
rect 5261 17765 5273 17768
rect 5307 17765 5319 17799
rect 6840 17796 6868 17824
rect 6840 17768 7144 17796
rect 5261 17759 5319 17765
rect 4525 17731 4583 17737
rect 4525 17697 4537 17731
rect 4571 17728 4583 17731
rect 4890 17728 4896 17740
rect 4571 17700 4896 17728
rect 4571 17697 4583 17700
rect 4525 17691 4583 17697
rect 4890 17688 4896 17700
rect 4948 17688 4954 17740
rect 6365 17731 6423 17737
rect 6365 17697 6377 17731
rect 6411 17728 6423 17731
rect 6546 17728 6552 17740
rect 6411 17700 6552 17728
rect 6411 17697 6423 17700
rect 6365 17691 6423 17697
rect 6546 17688 6552 17700
rect 6604 17728 6610 17740
rect 6825 17731 6883 17737
rect 6825 17728 6837 17731
rect 6604 17700 6837 17728
rect 6604 17688 6610 17700
rect 6825 17697 6837 17700
rect 6871 17697 6883 17731
rect 6825 17691 6883 17697
rect 4614 17660 4620 17672
rect 3697 17623 3755 17629
rect 3804 17632 4292 17660
rect 4575 17632 4620 17660
rect 2866 17552 2872 17604
rect 2924 17592 2930 17604
rect 3804 17592 3832 17632
rect 4614 17620 4620 17632
rect 4672 17660 4678 17672
rect 4982 17660 4988 17672
rect 4672 17632 4988 17660
rect 4672 17620 4678 17632
rect 4982 17620 4988 17632
rect 5040 17620 5046 17672
rect 5350 17660 5356 17672
rect 5311 17632 5356 17660
rect 5350 17620 5356 17632
rect 5408 17620 5414 17672
rect 7116 17669 7144 17768
rect 7650 17756 7656 17808
rect 7708 17796 7714 17808
rect 8205 17799 8263 17805
rect 8205 17796 8217 17799
rect 7708 17768 8217 17796
rect 7708 17756 7714 17768
rect 8205 17765 8217 17768
rect 8251 17765 8263 17799
rect 8404 17796 8432 17824
rect 10321 17799 10379 17805
rect 8404 17768 8524 17796
rect 8205 17759 8263 17765
rect 7558 17688 7564 17740
rect 7616 17728 7622 17740
rect 8297 17731 8355 17737
rect 8297 17728 8309 17731
rect 7616 17700 8309 17728
rect 7616 17688 7622 17700
rect 8297 17697 8309 17700
rect 8343 17728 8355 17731
rect 8343 17700 8432 17728
rect 8343 17697 8355 17700
rect 8297 17691 8355 17697
rect 5445 17663 5503 17669
rect 5445 17629 5457 17663
rect 5491 17629 5503 17663
rect 5445 17623 5503 17629
rect 7101 17663 7159 17669
rect 7101 17629 7113 17663
rect 7147 17629 7159 17663
rect 7101 17623 7159 17629
rect 2924 17564 3832 17592
rect 2924 17552 2930 17564
rect 4062 17552 4068 17604
rect 4120 17592 4126 17604
rect 5460 17592 5488 17623
rect 8404 17604 8432 17700
rect 8496 17672 8524 17768
rect 10321 17765 10333 17799
rect 10367 17796 10379 17799
rect 10686 17796 10692 17808
rect 10367 17768 10692 17796
rect 10367 17765 10379 17768
rect 10321 17759 10379 17765
rect 10686 17756 10692 17768
rect 10744 17756 10750 17808
rect 11149 17799 11207 17805
rect 11149 17796 11161 17799
rect 11072 17768 11161 17796
rect 9861 17731 9919 17737
rect 9861 17697 9873 17731
rect 9907 17728 9919 17731
rect 11072 17728 11100 17768
rect 11149 17765 11161 17768
rect 11195 17796 11207 17799
rect 15105 17799 15163 17805
rect 11195 17768 14228 17796
rect 11195 17765 11207 17768
rect 11149 17759 11207 17765
rect 14200 17740 14228 17768
rect 15105 17765 15117 17799
rect 15151 17796 15163 17799
rect 15286 17796 15292 17808
rect 15151 17768 15292 17796
rect 15151 17765 15163 17768
rect 15105 17759 15163 17765
rect 15286 17756 15292 17768
rect 15344 17796 15350 17808
rect 15746 17796 15752 17808
rect 15344 17768 15752 17796
rect 15344 17756 15350 17768
rect 15746 17756 15752 17768
rect 15804 17756 15810 17808
rect 16393 17799 16451 17805
rect 16393 17765 16405 17799
rect 16439 17796 16451 17799
rect 16482 17796 16488 17808
rect 16439 17768 16488 17796
rect 16439 17765 16451 17768
rect 16393 17759 16451 17765
rect 16482 17756 16488 17768
rect 16540 17756 16546 17808
rect 11238 17728 11244 17740
rect 9907 17700 11100 17728
rect 11151 17700 11244 17728
rect 9907 17697 9919 17700
rect 9861 17691 9919 17697
rect 11238 17688 11244 17700
rect 11296 17728 11302 17740
rect 11790 17728 11796 17740
rect 11296 17700 11796 17728
rect 11296 17688 11302 17700
rect 11790 17688 11796 17700
rect 11848 17728 11854 17740
rect 12437 17731 12495 17737
rect 12437 17728 12449 17731
rect 11848 17700 12449 17728
rect 11848 17688 11854 17700
rect 12437 17697 12449 17700
rect 12483 17697 12495 17731
rect 12437 17691 12495 17697
rect 13262 17688 13268 17740
rect 13320 17728 13326 17740
rect 13449 17731 13507 17737
rect 13449 17728 13461 17731
rect 13320 17700 13461 17728
rect 13320 17688 13326 17700
rect 13449 17697 13461 17700
rect 13495 17728 13507 17731
rect 14093 17731 14151 17737
rect 14093 17728 14105 17731
rect 13495 17700 14105 17728
rect 13495 17697 13507 17700
rect 13449 17691 13507 17697
rect 14093 17697 14105 17700
rect 14139 17697 14151 17731
rect 14093 17691 14151 17697
rect 14182 17688 14188 17740
rect 14240 17688 14246 17740
rect 15654 17728 15660 17740
rect 15615 17700 15660 17728
rect 15654 17688 15660 17700
rect 15712 17688 15718 17740
rect 16117 17731 16175 17737
rect 16117 17697 16129 17731
rect 16163 17728 16175 17731
rect 16206 17728 16212 17740
rect 16163 17700 16212 17728
rect 16163 17697 16175 17700
rect 16117 17691 16175 17697
rect 16206 17688 16212 17700
rect 16264 17688 16270 17740
rect 19889 17731 19947 17737
rect 19889 17728 19901 17731
rect 19720 17700 19901 17728
rect 8478 17620 8484 17672
rect 8536 17660 8542 17672
rect 10597 17663 10655 17669
rect 8536 17632 8581 17660
rect 8536 17620 8542 17632
rect 10597 17629 10609 17663
rect 10643 17660 10655 17663
rect 10778 17660 10784 17672
rect 10643 17632 10784 17660
rect 10643 17629 10655 17632
rect 10597 17623 10655 17629
rect 10778 17620 10784 17632
rect 10836 17620 10842 17672
rect 11330 17620 11336 17672
rect 11388 17660 11394 17672
rect 12069 17663 12127 17669
rect 11388 17632 11433 17660
rect 11388 17620 11394 17632
rect 12069 17629 12081 17663
rect 12115 17629 12127 17663
rect 12069 17623 12127 17629
rect 4120 17564 5488 17592
rect 4120 17552 4126 17564
rect 6822 17552 6828 17604
rect 6880 17592 6886 17604
rect 8202 17592 8208 17604
rect 6880 17564 8208 17592
rect 6880 17552 6886 17564
rect 8202 17552 8208 17564
rect 8260 17552 8266 17604
rect 8386 17592 8392 17604
rect 8299 17564 8392 17592
rect 8386 17552 8392 17564
rect 8444 17592 8450 17604
rect 8665 17595 8723 17601
rect 8665 17592 8677 17595
rect 8444 17564 8677 17592
rect 8444 17552 8450 17564
rect 8665 17561 8677 17564
rect 8711 17561 8723 17595
rect 8665 17555 8723 17561
rect 9858 17552 9864 17604
rect 9916 17592 9922 17604
rect 12084 17592 12112 17623
rect 12158 17620 12164 17672
rect 12216 17660 12222 17672
rect 14369 17663 14427 17669
rect 12216 17632 12261 17660
rect 12216 17620 12222 17632
rect 14369 17629 14381 17663
rect 14415 17660 14427 17663
rect 15286 17660 15292 17672
rect 14415 17632 15292 17660
rect 14415 17629 14427 17632
rect 14369 17623 14427 17629
rect 15286 17620 15292 17632
rect 15344 17620 15350 17672
rect 15378 17620 15384 17672
rect 15436 17660 15442 17672
rect 15749 17663 15807 17669
rect 15749 17660 15761 17663
rect 15436 17632 15761 17660
rect 15436 17620 15442 17632
rect 15749 17629 15761 17632
rect 15795 17629 15807 17663
rect 15930 17660 15936 17672
rect 15891 17632 15936 17660
rect 15749 17623 15807 17629
rect 15930 17620 15936 17632
rect 15988 17620 15994 17672
rect 19720 17604 19748 17700
rect 19889 17697 19901 17700
rect 19935 17697 19947 17731
rect 19889 17691 19947 17697
rect 20257 17731 20315 17737
rect 20257 17697 20269 17731
rect 20303 17728 20315 17731
rect 20714 17728 20720 17740
rect 20303 17700 20720 17728
rect 20303 17697 20315 17700
rect 20257 17691 20315 17697
rect 20714 17688 20720 17700
rect 20772 17688 20778 17740
rect 20901 17731 20959 17737
rect 20901 17697 20913 17731
rect 20947 17728 20959 17731
rect 21284 17728 21312 17824
rect 20947 17700 21312 17728
rect 20947 17697 20959 17700
rect 20901 17691 20959 17697
rect 20533 17663 20591 17669
rect 20533 17629 20545 17663
rect 20579 17660 20591 17663
rect 20622 17660 20628 17672
rect 20579 17632 20628 17660
rect 20579 17629 20591 17632
rect 20533 17623 20591 17629
rect 20622 17620 20628 17632
rect 20680 17620 20686 17672
rect 21177 17663 21235 17669
rect 21177 17629 21189 17663
rect 21223 17660 21235 17663
rect 21542 17660 21548 17672
rect 21223 17632 21548 17660
rect 21223 17629 21235 17632
rect 21177 17623 21235 17629
rect 21542 17620 21548 17632
rect 21600 17620 21606 17672
rect 9916 17564 12112 17592
rect 13725 17595 13783 17601
rect 9916 17552 9922 17564
rect 13725 17561 13737 17595
rect 13771 17592 13783 17595
rect 17218 17592 17224 17604
rect 13771 17564 17224 17592
rect 13771 17561 13783 17564
rect 13725 17555 13783 17561
rect 17218 17552 17224 17564
rect 17276 17552 17282 17604
rect 19702 17592 19708 17604
rect 19663 17564 19708 17592
rect 19702 17552 19708 17564
rect 19760 17552 19766 17604
rect 22002 17592 22008 17604
rect 21963 17564 22008 17592
rect 22002 17552 22008 17564
rect 22060 17552 22066 17604
rect 2222 17484 2228 17536
rect 2280 17524 2286 17536
rect 2317 17527 2375 17533
rect 2317 17524 2329 17527
rect 2280 17496 2329 17524
rect 2280 17484 2286 17496
rect 2317 17493 2329 17496
rect 2363 17493 2375 17527
rect 2317 17487 2375 17493
rect 2406 17484 2412 17536
rect 2464 17524 2470 17536
rect 3145 17527 3203 17533
rect 3145 17524 3157 17527
rect 2464 17496 3157 17524
rect 2464 17484 2470 17496
rect 3145 17493 3157 17496
rect 3191 17493 3203 17527
rect 3145 17487 3203 17493
rect 3234 17484 3240 17536
rect 3292 17524 3298 17536
rect 3878 17524 3884 17536
rect 3292 17496 3884 17524
rect 3292 17484 3298 17496
rect 3878 17484 3884 17496
rect 3936 17484 3942 17536
rect 6730 17484 6736 17536
rect 6788 17524 6794 17536
rect 7098 17524 7104 17536
rect 6788 17496 7104 17524
rect 6788 17484 6794 17496
rect 7098 17484 7104 17496
rect 7156 17524 7162 17536
rect 7377 17527 7435 17533
rect 7377 17524 7389 17527
rect 7156 17496 7389 17524
rect 7156 17484 7162 17496
rect 7377 17493 7389 17496
rect 7423 17493 7435 17527
rect 7650 17524 7656 17536
rect 7611 17496 7656 17524
rect 7377 17487 7435 17493
rect 7650 17484 7656 17496
rect 7708 17484 7714 17536
rect 7742 17484 7748 17536
rect 7800 17524 7806 17536
rect 7837 17527 7895 17533
rect 7837 17524 7849 17527
rect 7800 17496 7849 17524
rect 7800 17484 7806 17496
rect 7837 17493 7849 17496
rect 7883 17493 7895 17527
rect 7837 17487 7895 17493
rect 10134 17484 10140 17536
rect 10192 17524 10198 17536
rect 10594 17524 10600 17536
rect 10192 17496 10600 17524
rect 10192 17484 10198 17496
rect 10594 17484 10600 17496
rect 10652 17484 10658 17536
rect 12250 17484 12256 17536
rect 12308 17524 12314 17536
rect 13262 17524 13268 17536
rect 12308 17496 13268 17524
rect 12308 17484 12314 17496
rect 13262 17484 13268 17496
rect 13320 17484 13326 17536
rect 15289 17527 15347 17533
rect 15289 17493 15301 17527
rect 15335 17524 15347 17527
rect 16574 17524 16580 17536
rect 15335 17496 16580 17524
rect 15335 17493 15347 17496
rect 15289 17487 15347 17493
rect 16574 17484 16580 17496
rect 16632 17484 16638 17536
rect 1104 17434 21896 17456
rect 1104 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 4575 17434
rect 4627 17382 4639 17434
rect 4691 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 18308 17434
rect 18360 17382 18372 17434
rect 18424 17382 18436 17434
rect 18488 17382 18500 17434
rect 18552 17382 21896 17434
rect 1104 17360 21896 17382
rect 1857 17323 1915 17329
rect 1857 17289 1869 17323
rect 1903 17320 1915 17323
rect 5350 17320 5356 17332
rect 1903 17292 5356 17320
rect 1903 17289 1915 17292
rect 1857 17283 1915 17289
rect 5350 17280 5356 17292
rect 5408 17280 5414 17332
rect 5902 17280 5908 17332
rect 5960 17320 5966 17332
rect 5997 17323 6055 17329
rect 5997 17320 6009 17323
rect 5960 17292 6009 17320
rect 5960 17280 5966 17292
rect 5997 17289 6009 17292
rect 6043 17320 6055 17323
rect 6086 17320 6092 17332
rect 6043 17292 6092 17320
rect 6043 17289 6055 17292
rect 5997 17283 6055 17289
rect 6086 17280 6092 17292
rect 6144 17280 6150 17332
rect 6730 17320 6736 17332
rect 6196 17292 6736 17320
rect 4062 17252 4068 17264
rect 4023 17224 4068 17252
rect 4062 17212 4068 17224
rect 4120 17212 4126 17264
rect 4154 17212 4160 17264
rect 4212 17252 4218 17264
rect 5169 17255 5227 17261
rect 4212 17224 4257 17252
rect 4212 17212 4218 17224
rect 5169 17221 5181 17255
rect 5215 17252 5227 17255
rect 5534 17252 5540 17264
rect 5215 17224 5540 17252
rect 5215 17221 5227 17224
rect 5169 17215 5227 17221
rect 5534 17212 5540 17224
rect 5592 17212 5598 17264
rect 6196 17261 6224 17292
rect 6730 17280 6736 17292
rect 6788 17280 6794 17332
rect 6914 17280 6920 17332
rect 6972 17320 6978 17332
rect 6972 17292 7017 17320
rect 6972 17280 6978 17292
rect 7282 17280 7288 17332
rect 7340 17320 7346 17332
rect 8662 17320 8668 17332
rect 7340 17292 8668 17320
rect 7340 17280 7346 17292
rect 8662 17280 8668 17292
rect 8720 17280 8726 17332
rect 9858 17320 9864 17332
rect 9819 17292 9864 17320
rect 9858 17280 9864 17292
rect 9916 17280 9922 17332
rect 10689 17323 10747 17329
rect 9968 17292 10180 17320
rect 6181 17255 6239 17261
rect 6181 17252 6193 17255
rect 5644 17224 6193 17252
rect 5644 17196 5672 17224
rect 6181 17221 6193 17224
rect 6227 17221 6239 17255
rect 6181 17215 6239 17221
rect 6362 17212 6368 17264
rect 6420 17252 6426 17264
rect 7745 17255 7803 17261
rect 6420 17224 7696 17252
rect 6420 17212 6426 17224
rect 2317 17187 2375 17193
rect 2317 17153 2329 17187
rect 2363 17184 2375 17187
rect 2406 17184 2412 17196
rect 2363 17156 2412 17184
rect 2363 17153 2375 17156
rect 2317 17147 2375 17153
rect 2406 17144 2412 17156
rect 2464 17144 2470 17196
rect 2501 17187 2559 17193
rect 2501 17153 2513 17187
rect 2547 17153 2559 17187
rect 2501 17147 2559 17153
rect 2222 17116 2228 17128
rect 2183 17088 2228 17116
rect 2222 17076 2228 17088
rect 2280 17076 2286 17128
rect 2516 17048 2544 17147
rect 3786 17144 3792 17196
rect 3844 17184 3850 17196
rect 4617 17187 4675 17193
rect 4617 17184 4629 17187
rect 3844 17156 4629 17184
rect 3844 17144 3850 17156
rect 4617 17153 4629 17156
rect 4663 17184 4675 17187
rect 4706 17184 4712 17196
rect 4663 17156 4712 17184
rect 4663 17153 4675 17156
rect 4617 17147 4675 17153
rect 4706 17144 4712 17156
rect 4764 17144 4770 17196
rect 4801 17187 4859 17193
rect 4801 17153 4813 17187
rect 4847 17184 4859 17187
rect 4982 17184 4988 17196
rect 4847 17156 4988 17184
rect 4847 17153 4859 17156
rect 4801 17147 4859 17153
rect 4982 17144 4988 17156
rect 5040 17144 5046 17196
rect 5626 17184 5632 17196
rect 5587 17156 5632 17184
rect 5626 17144 5632 17156
rect 5684 17144 5690 17196
rect 5813 17187 5871 17193
rect 5813 17153 5825 17187
rect 5859 17184 5871 17187
rect 6270 17184 6276 17196
rect 5859 17156 6276 17184
rect 5859 17153 5871 17156
rect 5813 17147 5871 17153
rect 6270 17144 6276 17156
rect 6328 17144 6334 17196
rect 6457 17187 6515 17193
rect 6457 17153 6469 17187
rect 6503 17184 6515 17187
rect 6546 17184 6552 17196
rect 6503 17156 6552 17184
rect 6503 17153 6515 17156
rect 6457 17147 6515 17153
rect 6546 17144 6552 17156
rect 6604 17144 6610 17196
rect 7282 17144 7288 17196
rect 7340 17184 7346 17196
rect 7377 17187 7435 17193
rect 7377 17184 7389 17187
rect 7340 17156 7389 17184
rect 7340 17144 7346 17156
rect 7377 17153 7389 17156
rect 7423 17153 7435 17187
rect 7377 17147 7435 17153
rect 7561 17187 7619 17193
rect 7561 17153 7573 17187
rect 7607 17153 7619 17187
rect 7668 17184 7696 17224
rect 7745 17221 7757 17255
rect 7791 17252 7803 17255
rect 9214 17252 9220 17264
rect 7791 17224 9220 17252
rect 7791 17221 7803 17224
rect 7745 17215 7803 17221
rect 9214 17212 9220 17224
rect 9272 17212 9278 17264
rect 9490 17212 9496 17264
rect 9548 17252 9554 17264
rect 9968 17252 9996 17292
rect 9548 17224 9996 17252
rect 10152 17252 10180 17292
rect 10689 17289 10701 17323
rect 10735 17320 10747 17323
rect 11974 17320 11980 17332
rect 10735 17292 11980 17320
rect 10735 17289 10747 17292
rect 10689 17283 10747 17289
rect 11974 17280 11980 17292
rect 12032 17280 12038 17332
rect 15378 17320 15384 17332
rect 12452 17292 14964 17320
rect 15339 17292 15384 17320
rect 10152 17224 11652 17252
rect 9548 17212 9554 17224
rect 11624 17196 11652 17224
rect 7834 17184 7840 17196
rect 7668 17156 7840 17184
rect 7561 17147 7619 17153
rect 2682 17116 2688 17128
rect 2643 17088 2688 17116
rect 2682 17076 2688 17088
rect 2740 17076 2746 17128
rect 3418 17076 3424 17128
rect 3476 17116 3482 17128
rect 3970 17116 3976 17128
rect 3476 17088 3976 17116
rect 3476 17076 3482 17088
rect 3970 17076 3976 17088
rect 4028 17076 4034 17128
rect 5537 17119 5595 17125
rect 5537 17085 5549 17119
rect 5583 17116 5595 17119
rect 5902 17116 5908 17128
rect 5583 17088 5908 17116
rect 5583 17085 5595 17088
rect 5537 17079 5595 17085
rect 5902 17076 5908 17088
rect 5960 17076 5966 17128
rect 6178 17076 6184 17128
rect 6236 17116 6242 17128
rect 6730 17116 6736 17128
rect 6236 17088 6736 17116
rect 6236 17076 6242 17088
rect 6730 17076 6736 17088
rect 6788 17076 6794 17128
rect 7576 17116 7604 17147
rect 7834 17144 7840 17156
rect 7892 17184 7898 17196
rect 8297 17187 8355 17193
rect 8297 17184 8309 17187
rect 7892 17156 8309 17184
rect 7892 17144 7898 17156
rect 8297 17153 8309 17156
rect 8343 17153 8355 17187
rect 8662 17184 8668 17196
rect 8575 17156 8668 17184
rect 8297 17147 8355 17153
rect 8662 17144 8668 17156
rect 8720 17184 8726 17196
rect 9582 17184 9588 17196
rect 8720 17156 9588 17184
rect 8720 17144 8726 17156
rect 9582 17144 9588 17156
rect 9640 17184 9646 17196
rect 9858 17184 9864 17196
rect 9640 17156 9864 17184
rect 9640 17144 9646 17156
rect 9858 17144 9864 17156
rect 9916 17144 9922 17196
rect 10505 17187 10563 17193
rect 10505 17153 10517 17187
rect 10551 17184 10563 17187
rect 10778 17184 10784 17196
rect 10551 17156 10784 17184
rect 10551 17153 10563 17156
rect 10505 17147 10563 17153
rect 10778 17144 10784 17156
rect 10836 17184 10842 17196
rect 11241 17187 11299 17193
rect 11241 17184 11253 17187
rect 10836 17156 11253 17184
rect 10836 17144 10842 17156
rect 11241 17153 11253 17156
rect 11287 17153 11299 17187
rect 11606 17184 11612 17196
rect 11567 17156 11612 17184
rect 11241 17147 11299 17153
rect 11606 17144 11612 17156
rect 11664 17144 11670 17196
rect 12452 17184 12480 17292
rect 12360 17156 12480 17184
rect 14936 17184 14964 17292
rect 15378 17280 15384 17292
rect 15436 17280 15442 17332
rect 16206 17320 16212 17332
rect 16167 17292 16212 17320
rect 16206 17280 16212 17292
rect 16264 17280 16270 17332
rect 20625 17323 20683 17329
rect 20625 17289 20637 17323
rect 20671 17320 20683 17323
rect 20714 17320 20720 17332
rect 20671 17292 20720 17320
rect 20671 17289 20683 17292
rect 20625 17283 20683 17289
rect 20714 17280 20720 17292
rect 20772 17280 20778 17332
rect 21453 17323 21511 17329
rect 21453 17289 21465 17323
rect 21499 17320 21511 17323
rect 21634 17320 21640 17332
rect 21499 17292 21640 17320
rect 21499 17289 21511 17292
rect 21453 17283 21511 17289
rect 21634 17280 21640 17292
rect 21692 17280 21698 17332
rect 15286 17252 15292 17264
rect 15247 17224 15292 17252
rect 15286 17212 15292 17224
rect 15344 17252 15350 17264
rect 15344 17224 15976 17252
rect 15344 17212 15350 17224
rect 15948 17193 15976 17224
rect 15933 17187 15991 17193
rect 14936 17156 15700 17184
rect 8478 17116 8484 17128
rect 7576 17088 8484 17116
rect 8478 17076 8484 17088
rect 8536 17076 8542 17128
rect 9674 17076 9680 17128
rect 9732 17116 9738 17128
rect 10321 17119 10379 17125
rect 10321 17116 10333 17119
rect 9732 17088 10333 17116
rect 9732 17076 9738 17088
rect 10321 17085 10333 17088
rect 10367 17085 10379 17119
rect 11054 17116 11060 17128
rect 11015 17088 11060 17116
rect 10321 17079 10379 17085
rect 11054 17076 11060 17088
rect 11112 17076 11118 17128
rect 11149 17119 11207 17125
rect 11149 17085 11161 17119
rect 11195 17116 11207 17119
rect 11330 17116 11336 17128
rect 11195 17088 11336 17116
rect 11195 17085 11207 17088
rect 11149 17079 11207 17085
rect 11330 17076 11336 17088
rect 11388 17116 11394 17128
rect 12360 17116 12388 17156
rect 11388 17088 12388 17116
rect 11388 17076 11394 17088
rect 12434 17076 12440 17128
rect 12492 17116 12498 17128
rect 12492 17088 12537 17116
rect 12492 17076 12498 17088
rect 13814 17076 13820 17128
rect 13872 17116 13878 17128
rect 13909 17119 13967 17125
rect 13909 17116 13921 17119
rect 13872 17088 13921 17116
rect 13872 17076 13878 17088
rect 13909 17085 13921 17088
rect 13955 17085 13967 17119
rect 13909 17079 13967 17085
rect 2952 17051 3010 17057
rect 2952 17048 2964 17051
rect 2516 17020 2964 17048
rect 2952 17017 2964 17020
rect 2998 17048 3010 17051
rect 3234 17048 3240 17060
rect 2998 17020 3240 17048
rect 2998 17017 3010 17020
rect 2952 17011 3010 17017
rect 3234 17008 3240 17020
rect 3292 17008 3298 17060
rect 3510 17008 3516 17060
rect 3568 17048 3574 17060
rect 6641 17051 6699 17057
rect 3568 17020 4568 17048
rect 3568 17008 3574 17020
rect 1394 16940 1400 16992
rect 1452 16980 1458 16992
rect 1765 16983 1823 16989
rect 1765 16980 1777 16983
rect 1452 16952 1777 16980
rect 1452 16940 1458 16952
rect 1765 16949 1777 16952
rect 1811 16980 1823 16983
rect 4338 16980 4344 16992
rect 1811 16952 4344 16980
rect 1811 16949 1823 16952
rect 1765 16943 1823 16949
rect 4338 16940 4344 16952
rect 4396 16940 4402 16992
rect 4540 16989 4568 17020
rect 6641 17017 6653 17051
rect 6687 17048 6699 17051
rect 7285 17051 7343 17057
rect 7285 17048 7297 17051
rect 6687 17020 7297 17048
rect 6687 17017 6699 17020
rect 6641 17011 6699 17017
rect 7285 17017 7297 17020
rect 7331 17048 7343 17051
rect 11698 17048 11704 17060
rect 7331 17020 11704 17048
rect 7331 17017 7343 17020
rect 7285 17011 7343 17017
rect 11698 17008 11704 17020
rect 11756 17008 11762 17060
rect 12704 17051 12762 17057
rect 12704 17017 12716 17051
rect 12750 17048 12762 17051
rect 13354 17048 13360 17060
rect 12750 17020 13360 17048
rect 12750 17017 12762 17020
rect 12704 17011 12762 17017
rect 13354 17008 13360 17020
rect 13412 17008 13418 17060
rect 14154 17051 14212 17057
rect 14154 17048 14166 17051
rect 13832 17020 14166 17048
rect 4525 16983 4583 16989
rect 4525 16949 4537 16983
rect 4571 16980 4583 16983
rect 4985 16983 5043 16989
rect 4985 16980 4997 16983
rect 4571 16952 4997 16980
rect 4571 16949 4583 16952
rect 4525 16943 4583 16949
rect 4985 16949 4997 16952
rect 5031 16949 5043 16983
rect 4985 16943 5043 16949
rect 7098 16940 7104 16992
rect 7156 16980 7162 16992
rect 8113 16983 8171 16989
rect 8113 16980 8125 16983
rect 7156 16952 8125 16980
rect 7156 16940 7162 16952
rect 8113 16949 8125 16952
rect 8159 16949 8171 16983
rect 8113 16943 8171 16949
rect 8202 16940 8208 16992
rect 8260 16980 8266 16992
rect 8757 16983 8815 16989
rect 8757 16980 8769 16983
rect 8260 16952 8769 16980
rect 8260 16940 8266 16952
rect 8757 16949 8769 16952
rect 8803 16949 8815 16983
rect 9490 16980 9496 16992
rect 9451 16952 9496 16980
rect 8757 16943 8815 16949
rect 9490 16940 9496 16952
rect 9548 16980 9554 16992
rect 13832 16989 13860 17020
rect 14154 17017 14166 17020
rect 14200 17048 14212 17051
rect 14274 17048 14280 17060
rect 14200 17020 14280 17048
rect 14200 17017 14212 17020
rect 14154 17011 14212 17017
rect 14274 17008 14280 17020
rect 14332 17008 14338 17060
rect 15672 17048 15700 17156
rect 15933 17153 15945 17187
rect 15979 17153 15991 17187
rect 15933 17147 15991 17153
rect 16666 17144 16672 17196
rect 16724 17184 16730 17196
rect 16761 17187 16819 17193
rect 16761 17184 16773 17187
rect 16724 17156 16773 17184
rect 16724 17144 16730 17156
rect 16761 17153 16773 17156
rect 16807 17153 16819 17187
rect 16761 17147 16819 17153
rect 19518 17144 19524 17196
rect 19576 17184 19582 17196
rect 20165 17187 20223 17193
rect 19576 17156 20024 17184
rect 19576 17144 19582 17156
rect 15746 17076 15752 17128
rect 15804 17116 15810 17128
rect 15841 17119 15899 17125
rect 15841 17116 15853 17119
rect 15804 17088 15853 17116
rect 15804 17076 15810 17088
rect 15841 17085 15853 17088
rect 15887 17085 15899 17119
rect 16574 17116 16580 17128
rect 16535 17088 16580 17116
rect 15841 17079 15899 17085
rect 16574 17076 16580 17088
rect 16632 17076 16638 17128
rect 19702 17076 19708 17128
rect 19760 17116 19766 17128
rect 19889 17119 19947 17125
rect 19889 17116 19901 17119
rect 19760 17088 19901 17116
rect 19760 17076 19766 17088
rect 19889 17085 19901 17088
rect 19935 17085 19947 17119
rect 19996 17116 20024 17156
rect 20165 17153 20177 17187
rect 20211 17184 20223 17187
rect 20211 17156 21312 17184
rect 20211 17153 20223 17156
rect 20165 17147 20223 17153
rect 20438 17116 20444 17128
rect 19996 17088 20444 17116
rect 19889 17079 19947 17085
rect 20438 17076 20444 17088
rect 20496 17116 20502 17128
rect 21284 17125 21312 17156
rect 20717 17119 20775 17125
rect 20717 17116 20729 17119
rect 20496 17088 20729 17116
rect 20496 17076 20502 17088
rect 20717 17085 20729 17088
rect 20763 17085 20775 17119
rect 20717 17079 20775 17085
rect 21269 17119 21327 17125
rect 21269 17085 21281 17119
rect 21315 17085 21327 17119
rect 21269 17079 21327 17085
rect 19334 17048 19340 17060
rect 15672 17020 19340 17048
rect 19334 17008 19340 17020
rect 19392 17008 19398 17060
rect 20993 17051 21051 17057
rect 20993 17017 21005 17051
rect 21039 17017 21051 17051
rect 20993 17011 21051 17017
rect 10229 16983 10287 16989
rect 10229 16980 10241 16983
rect 9548 16952 10241 16980
rect 9548 16940 9554 16952
rect 10229 16949 10241 16952
rect 10275 16949 10287 16983
rect 10229 16943 10287 16949
rect 13817 16983 13875 16989
rect 13817 16949 13829 16983
rect 13863 16949 13875 16983
rect 13817 16943 13875 16949
rect 14458 16940 14464 16992
rect 14516 16980 14522 16992
rect 15749 16983 15807 16989
rect 15749 16980 15761 16983
rect 14516 16952 15761 16980
rect 14516 16940 14522 16952
rect 15749 16949 15761 16952
rect 15795 16949 15807 16983
rect 15749 16943 15807 16949
rect 16669 16983 16727 16989
rect 16669 16949 16681 16983
rect 16715 16980 16727 16983
rect 16758 16980 16764 16992
rect 16715 16952 16764 16980
rect 16715 16949 16727 16952
rect 16669 16943 16727 16949
rect 16758 16940 16764 16952
rect 16816 16940 16822 16992
rect 21008 16980 21036 17011
rect 21266 16980 21272 16992
rect 21008 16952 21272 16980
rect 21266 16940 21272 16952
rect 21324 16940 21330 16992
rect 1104 16890 21896 16912
rect 1104 16838 7912 16890
rect 7964 16838 7976 16890
rect 8028 16838 8040 16890
rect 8092 16838 8104 16890
rect 8156 16838 14843 16890
rect 14895 16838 14907 16890
rect 14959 16838 14971 16890
rect 15023 16838 15035 16890
rect 15087 16838 21896 16890
rect 1104 16816 21896 16838
rect 3513 16779 3571 16785
rect 3513 16776 3525 16779
rect 1504 16748 3525 16776
rect 1504 16649 1532 16748
rect 3513 16745 3525 16748
rect 3559 16776 3571 16779
rect 3694 16776 3700 16788
rect 3559 16748 3700 16776
rect 3559 16745 3571 16748
rect 3513 16739 3571 16745
rect 3694 16736 3700 16748
rect 3752 16736 3758 16788
rect 5537 16779 5595 16785
rect 5537 16745 5549 16779
rect 5583 16776 5595 16779
rect 6362 16776 6368 16788
rect 5583 16748 6368 16776
rect 5583 16745 5595 16748
rect 5537 16739 5595 16745
rect 6362 16736 6368 16748
rect 6420 16736 6426 16788
rect 6457 16779 6515 16785
rect 6457 16745 6469 16779
rect 6503 16776 6515 16779
rect 7374 16776 7380 16788
rect 6503 16748 7380 16776
rect 6503 16745 6515 16748
rect 6457 16739 6515 16745
rect 7374 16736 7380 16748
rect 7432 16736 7438 16788
rect 8754 16776 8760 16788
rect 8715 16748 8760 16776
rect 8754 16736 8760 16748
rect 8812 16736 8818 16788
rect 9677 16779 9735 16785
rect 9677 16745 9689 16779
rect 9723 16776 9735 16779
rect 9950 16776 9956 16788
rect 9723 16748 9956 16776
rect 9723 16745 9735 16748
rect 9677 16739 9735 16745
rect 9950 16736 9956 16748
rect 10008 16736 10014 16788
rect 10962 16736 10968 16788
rect 11020 16776 11026 16788
rect 11057 16779 11115 16785
rect 11057 16776 11069 16779
rect 11020 16748 11069 16776
rect 11020 16736 11026 16748
rect 11057 16745 11069 16748
rect 11103 16745 11115 16779
rect 11057 16739 11115 16745
rect 11241 16779 11299 16785
rect 11241 16745 11253 16779
rect 11287 16776 11299 16779
rect 12529 16779 12587 16785
rect 12529 16776 12541 16779
rect 11287 16748 12541 16776
rect 11287 16745 11299 16748
rect 11241 16739 11299 16745
rect 12529 16745 12541 16748
rect 12575 16745 12587 16779
rect 12529 16739 12587 16745
rect 12897 16779 12955 16785
rect 12897 16745 12909 16779
rect 12943 16776 12955 16779
rect 14185 16779 14243 16785
rect 14185 16776 14197 16779
rect 12943 16748 14197 16776
rect 12943 16745 12955 16748
rect 12897 16739 12955 16745
rect 14185 16745 14197 16748
rect 14231 16745 14243 16779
rect 16758 16776 16764 16788
rect 16719 16748 16764 16776
rect 14185 16739 14243 16745
rect 2498 16668 2504 16720
rect 2556 16708 2562 16720
rect 2682 16708 2688 16720
rect 2556 16680 2688 16708
rect 2556 16668 2562 16680
rect 2682 16668 2688 16680
rect 2740 16668 2746 16720
rect 4062 16668 4068 16720
rect 4120 16708 4126 16720
rect 4402 16711 4460 16717
rect 4402 16708 4414 16711
rect 4120 16680 4414 16708
rect 4120 16668 4126 16680
rect 4402 16677 4414 16680
rect 4448 16677 4460 16711
rect 6086 16708 6092 16720
rect 6047 16680 6092 16708
rect 4402 16671 4460 16677
rect 6086 16668 6092 16680
rect 6144 16668 6150 16720
rect 6638 16708 6644 16720
rect 6288 16680 6644 16708
rect 1489 16643 1547 16649
rect 1489 16609 1501 16643
rect 1535 16609 1547 16643
rect 1489 16603 1547 16609
rect 1670 16600 1676 16652
rect 1728 16600 1734 16652
rect 2124 16643 2182 16649
rect 2124 16609 2136 16643
rect 2170 16640 2182 16643
rect 2590 16640 2596 16652
rect 2170 16612 2596 16640
rect 2170 16609 2182 16612
rect 2124 16603 2182 16609
rect 2590 16600 2596 16612
rect 2648 16600 2654 16652
rect 5258 16600 5264 16652
rect 5316 16640 5322 16652
rect 5997 16643 6055 16649
rect 5997 16640 6009 16643
rect 5316 16612 6009 16640
rect 5316 16600 5322 16612
rect 5997 16609 6009 16612
rect 6043 16640 6055 16643
rect 6288 16640 6316 16680
rect 6638 16668 6644 16680
rect 6696 16668 6702 16720
rect 6917 16711 6975 16717
rect 6917 16677 6929 16711
rect 6963 16708 6975 16711
rect 8110 16708 8116 16720
rect 6963 16680 8116 16708
rect 6963 16677 6975 16680
rect 6917 16671 6975 16677
rect 8110 16668 8116 16680
rect 8168 16668 8174 16720
rect 9217 16711 9275 16717
rect 9217 16677 9229 16711
rect 9263 16708 9275 16711
rect 10502 16708 10508 16720
rect 9263 16680 10508 16708
rect 9263 16677 9275 16680
rect 9217 16671 9275 16677
rect 10502 16668 10508 16680
rect 10560 16708 10566 16720
rect 10689 16711 10747 16717
rect 10689 16708 10701 16711
rect 10560 16680 10701 16708
rect 10560 16668 10566 16680
rect 10689 16677 10701 16680
rect 10735 16677 10747 16711
rect 11072 16708 11100 16739
rect 16758 16736 16764 16748
rect 16816 16736 16822 16788
rect 17218 16776 17224 16788
rect 17179 16748 17224 16776
rect 17218 16736 17224 16748
rect 17276 16736 17282 16788
rect 21085 16779 21143 16785
rect 21085 16745 21097 16779
rect 21131 16776 21143 16779
rect 22005 16779 22063 16785
rect 22005 16776 22017 16779
rect 21131 16748 22017 16776
rect 21131 16745 21143 16748
rect 21085 16739 21143 16745
rect 22005 16745 22017 16748
rect 22051 16745 22063 16779
rect 22005 16739 22063 16745
rect 11606 16708 11612 16720
rect 11072 16680 11192 16708
rect 11567 16680 11612 16708
rect 10689 16671 10747 16677
rect 6043 16612 6316 16640
rect 6043 16609 6055 16612
rect 5997 16603 6055 16609
rect 6362 16600 6368 16652
rect 6420 16640 6426 16652
rect 7558 16649 7564 16652
rect 6825 16643 6883 16649
rect 6825 16640 6837 16643
rect 6420 16612 6837 16640
rect 6420 16600 6426 16612
rect 6825 16609 6837 16612
rect 6871 16609 6883 16643
rect 7552 16640 7564 16649
rect 6825 16603 6883 16609
rect 7116 16612 7564 16640
rect 1688 16513 1716 16600
rect 1857 16575 1915 16581
rect 1857 16541 1869 16575
rect 1903 16541 1915 16575
rect 1857 16535 1915 16541
rect 1673 16507 1731 16513
rect 1673 16473 1685 16507
rect 1719 16473 1731 16507
rect 1673 16467 1731 16473
rect 1872 16436 1900 16535
rect 4062 16532 4068 16584
rect 4120 16572 4126 16584
rect 4157 16575 4215 16581
rect 4157 16572 4169 16575
rect 4120 16544 4169 16572
rect 4120 16532 4126 16544
rect 4157 16541 4169 16544
rect 4203 16541 4215 16575
rect 6270 16572 6276 16584
rect 6231 16544 6276 16572
rect 4157 16535 4215 16541
rect 6270 16532 6276 16544
rect 6328 16532 6334 16584
rect 7116 16581 7144 16612
rect 7552 16603 7564 16612
rect 7558 16600 7564 16603
rect 7616 16600 7622 16652
rect 9122 16640 9128 16652
rect 9035 16612 9128 16640
rect 9122 16600 9128 16612
rect 9180 16640 9186 16652
rect 9180 16612 9444 16640
rect 9180 16600 9186 16612
rect 7101 16575 7159 16581
rect 7101 16541 7113 16575
rect 7147 16541 7159 16575
rect 7101 16535 7159 16541
rect 7190 16532 7196 16584
rect 7248 16572 7254 16584
rect 7285 16575 7343 16581
rect 7285 16572 7297 16575
rect 7248 16544 7297 16572
rect 7248 16532 7254 16544
rect 7285 16541 7297 16544
rect 7331 16541 7343 16575
rect 7285 16535 7343 16541
rect 8478 16532 8484 16584
rect 8536 16572 8542 16584
rect 9309 16575 9367 16581
rect 9309 16572 9321 16575
rect 8536 16544 9321 16572
rect 8536 16532 8542 16544
rect 3786 16504 3792 16516
rect 3747 16476 3792 16504
rect 3786 16464 3792 16476
rect 3844 16464 3850 16516
rect 8680 16513 8708 16544
rect 9309 16541 9321 16544
rect 9355 16541 9367 16575
rect 9416 16572 9444 16612
rect 9674 16600 9680 16652
rect 9732 16640 9738 16652
rect 10045 16643 10103 16649
rect 10045 16640 10057 16643
rect 9732 16612 10057 16640
rect 9732 16600 9738 16612
rect 10045 16609 10057 16612
rect 10091 16609 10103 16643
rect 10045 16603 10103 16609
rect 10137 16643 10195 16649
rect 10137 16609 10149 16643
rect 10183 16640 10195 16643
rect 11054 16640 11060 16652
rect 10183 16612 11060 16640
rect 10183 16609 10195 16612
rect 10137 16603 10195 16609
rect 11054 16600 11060 16612
rect 11112 16600 11118 16652
rect 11164 16640 11192 16680
rect 11606 16668 11612 16680
rect 11664 16668 11670 16720
rect 13357 16711 13415 16717
rect 13357 16708 13369 16711
rect 12084 16680 13369 16708
rect 11701 16643 11759 16649
rect 11701 16640 11713 16643
rect 11164 16612 11713 16640
rect 11701 16609 11713 16612
rect 11747 16609 11759 16643
rect 11701 16603 11759 16609
rect 10229 16575 10287 16581
rect 9416 16544 9812 16572
rect 9309 16535 9367 16541
rect 8665 16507 8723 16513
rect 5552 16476 6224 16504
rect 2498 16436 2504 16448
rect 1872 16408 2504 16436
rect 2498 16396 2504 16408
rect 2556 16396 2562 16448
rect 3234 16436 3240 16448
rect 3195 16408 3240 16436
rect 3234 16396 3240 16408
rect 3292 16396 3298 16448
rect 3326 16396 3332 16448
rect 3384 16436 3390 16448
rect 3421 16439 3479 16445
rect 3421 16436 3433 16439
rect 3384 16408 3433 16436
rect 3384 16396 3390 16408
rect 3421 16405 3433 16408
rect 3467 16436 3479 16439
rect 5552 16436 5580 16476
rect 3467 16408 5580 16436
rect 3467 16405 3479 16408
rect 3421 16399 3479 16405
rect 5626 16396 5632 16448
rect 5684 16436 5690 16448
rect 6196 16436 6224 16476
rect 8665 16473 8677 16507
rect 8711 16473 8723 16507
rect 8665 16467 8723 16473
rect 8754 16436 8760 16448
rect 5684 16408 5729 16436
rect 6196 16408 8760 16436
rect 5684 16396 5690 16408
rect 8754 16396 8760 16408
rect 8812 16396 8818 16448
rect 9784 16436 9812 16544
rect 10229 16541 10241 16575
rect 10275 16541 10287 16575
rect 10229 16535 10287 16541
rect 11885 16575 11943 16581
rect 11885 16541 11897 16575
rect 11931 16572 11943 16575
rect 11931 16544 12020 16572
rect 11931 16541 11943 16544
rect 11885 16535 11943 16541
rect 9858 16464 9864 16516
rect 9916 16504 9922 16516
rect 10244 16504 10272 16535
rect 9916 16476 10272 16504
rect 10597 16507 10655 16513
rect 9916 16464 9922 16476
rect 10597 16473 10609 16507
rect 10643 16504 10655 16507
rect 11330 16504 11336 16516
rect 10643 16476 11336 16504
rect 10643 16473 10655 16476
rect 10597 16467 10655 16473
rect 11330 16464 11336 16476
rect 11388 16464 11394 16516
rect 10873 16439 10931 16445
rect 10873 16436 10885 16439
rect 9784 16408 10885 16436
rect 10873 16405 10885 16408
rect 10919 16405 10931 16439
rect 11992 16436 12020 16544
rect 12084 16513 12112 16680
rect 13357 16677 13369 16680
rect 13403 16677 13415 16711
rect 14093 16711 14151 16717
rect 14093 16708 14105 16711
rect 13357 16671 13415 16677
rect 13556 16680 14105 16708
rect 12434 16600 12440 16652
rect 12492 16640 12498 16652
rect 13262 16640 13268 16652
rect 12492 16612 12537 16640
rect 13223 16612 13268 16640
rect 12492 16600 12498 16612
rect 13262 16600 13268 16612
rect 13320 16600 13326 16652
rect 12710 16572 12716 16584
rect 12671 16544 12716 16572
rect 12710 16532 12716 16544
rect 12768 16532 12774 16584
rect 13354 16532 13360 16584
rect 13412 16572 13418 16584
rect 13449 16575 13507 16581
rect 13449 16572 13461 16575
rect 13412 16544 13461 16572
rect 13412 16532 13418 16544
rect 13449 16541 13461 16544
rect 13495 16541 13507 16575
rect 13449 16535 13507 16541
rect 12069 16507 12127 16513
rect 12069 16473 12081 16507
rect 12115 16473 12127 16507
rect 12069 16467 12127 16473
rect 12250 16464 12256 16516
rect 12308 16504 12314 16516
rect 13556 16504 13584 16680
rect 14093 16677 14105 16680
rect 14139 16677 14151 16711
rect 14093 16671 14151 16677
rect 20438 16668 20444 16720
rect 20496 16708 20502 16720
rect 21453 16711 21511 16717
rect 21453 16708 21465 16711
rect 20496 16680 21465 16708
rect 20496 16668 20502 16680
rect 21453 16677 21465 16680
rect 21499 16677 21511 16711
rect 21453 16671 21511 16677
rect 13906 16640 13912 16652
rect 13740 16612 13912 16640
rect 13740 16513 13768 16612
rect 13906 16600 13912 16612
rect 13964 16600 13970 16652
rect 14458 16600 14464 16652
rect 14516 16640 14522 16652
rect 15562 16649 15568 16652
rect 15013 16643 15071 16649
rect 15013 16640 15025 16643
rect 14516 16612 15025 16640
rect 14516 16600 14522 16612
rect 15013 16609 15025 16612
rect 15059 16609 15071 16643
rect 15556 16640 15568 16649
rect 15475 16612 15568 16640
rect 15013 16603 15071 16609
rect 15556 16603 15568 16612
rect 15620 16640 15626 16652
rect 15930 16640 15936 16652
rect 15620 16612 15936 16640
rect 15562 16600 15568 16603
rect 15620 16600 15626 16612
rect 15930 16600 15936 16612
rect 15988 16640 15994 16652
rect 17126 16640 17132 16652
rect 15988 16612 16344 16640
rect 17087 16612 17132 16640
rect 15988 16600 15994 16612
rect 14274 16572 14280 16584
rect 14235 16544 14280 16572
rect 14274 16532 14280 16544
rect 14332 16532 14338 16584
rect 15289 16575 15347 16581
rect 15289 16541 15301 16575
rect 15335 16541 15347 16575
rect 16316 16572 16344 16612
rect 17126 16600 17132 16612
rect 17184 16600 17190 16652
rect 20806 16600 20812 16652
rect 20864 16640 20870 16652
rect 20901 16643 20959 16649
rect 20901 16640 20913 16643
rect 20864 16612 20913 16640
rect 20864 16600 20870 16612
rect 20901 16609 20913 16612
rect 20947 16640 20959 16643
rect 21269 16643 21327 16649
rect 21269 16640 21281 16643
rect 20947 16612 21281 16640
rect 20947 16609 20959 16612
rect 20901 16603 20959 16609
rect 21269 16609 21281 16612
rect 21315 16609 21327 16643
rect 21269 16603 21327 16609
rect 17313 16575 17371 16581
rect 16316 16544 16804 16572
rect 15289 16535 15347 16541
rect 12308 16476 13584 16504
rect 13725 16507 13783 16513
rect 12308 16464 12314 16476
rect 13725 16473 13737 16507
rect 13771 16473 13783 16507
rect 13725 16467 13783 16473
rect 12802 16436 12808 16448
rect 11992 16408 12808 16436
rect 10873 16399 10931 16405
rect 12802 16396 12808 16408
rect 12860 16396 12866 16448
rect 15304 16436 15332 16535
rect 16666 16504 16672 16516
rect 16627 16476 16672 16504
rect 16666 16464 16672 16476
rect 16724 16464 16730 16516
rect 16776 16504 16804 16544
rect 17313 16541 17325 16575
rect 17359 16541 17371 16575
rect 17313 16535 17371 16541
rect 17328 16504 17356 16535
rect 16776 16476 17356 16504
rect 15930 16436 15936 16448
rect 15304 16408 15936 16436
rect 15930 16396 15936 16408
rect 15988 16396 15994 16448
rect 1104 16346 21896 16368
rect 1104 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 4575 16346
rect 4627 16294 4639 16346
rect 4691 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 18308 16346
rect 18360 16294 18372 16346
rect 18424 16294 18436 16346
rect 18488 16294 18500 16346
rect 18552 16294 21896 16346
rect 1104 16272 21896 16294
rect 1578 16232 1584 16244
rect 1539 16204 1584 16232
rect 1578 16192 1584 16204
rect 1636 16192 1642 16244
rect 2314 16232 2320 16244
rect 2275 16204 2320 16232
rect 2314 16192 2320 16204
rect 2372 16192 2378 16244
rect 2685 16235 2743 16241
rect 2685 16201 2697 16235
rect 2731 16232 2743 16235
rect 2774 16232 2780 16244
rect 2731 16204 2780 16232
rect 2731 16201 2743 16204
rect 2685 16195 2743 16201
rect 2774 16192 2780 16204
rect 2832 16192 2838 16244
rect 2866 16192 2872 16244
rect 2924 16232 2930 16244
rect 2924 16204 2969 16232
rect 2924 16192 2930 16204
rect 3050 16192 3056 16244
rect 3108 16232 3114 16244
rect 4246 16232 4252 16244
rect 3108 16204 4252 16232
rect 3108 16192 3114 16204
rect 4246 16192 4252 16204
rect 4304 16192 4310 16244
rect 4798 16232 4804 16244
rect 4759 16204 4804 16232
rect 4798 16192 4804 16204
rect 4856 16192 4862 16244
rect 4985 16235 5043 16241
rect 4985 16201 4997 16235
rect 5031 16232 5043 16235
rect 5258 16232 5264 16244
rect 5031 16204 5264 16232
rect 5031 16201 5043 16204
rect 4985 16195 5043 16201
rect 5258 16192 5264 16204
rect 5316 16192 5322 16244
rect 7190 16232 7196 16244
rect 6840 16204 7196 16232
rect 2590 16124 2596 16176
rect 2648 16164 2654 16176
rect 2648 16136 3556 16164
rect 2648 16124 2654 16136
rect 3234 16056 3240 16108
rect 3292 16096 3298 16108
rect 3421 16099 3479 16105
rect 3421 16096 3433 16099
rect 3292 16068 3433 16096
rect 3292 16056 3298 16068
rect 3421 16065 3433 16068
rect 3467 16065 3479 16099
rect 3528 16096 3556 16136
rect 4062 16124 4068 16176
rect 4120 16164 4126 16176
rect 4120 16136 5304 16164
rect 4120 16124 4126 16136
rect 5276 16105 5304 16136
rect 6840 16105 6868 16204
rect 7190 16192 7196 16204
rect 7248 16192 7254 16244
rect 7558 16192 7564 16244
rect 7616 16232 7622 16244
rect 8205 16235 8263 16241
rect 8205 16232 8217 16235
rect 7616 16204 8217 16232
rect 7616 16192 7622 16204
rect 8205 16201 8217 16204
rect 8251 16201 8263 16235
rect 8205 16195 8263 16201
rect 8754 16192 8760 16244
rect 8812 16232 8818 16244
rect 8812 16204 10640 16232
rect 8812 16192 8818 16204
rect 8110 16124 8116 16176
rect 8168 16164 8174 16176
rect 8297 16167 8355 16173
rect 8297 16164 8309 16167
rect 8168 16136 8309 16164
rect 8168 16124 8174 16136
rect 8297 16133 8309 16136
rect 8343 16133 8355 16167
rect 10612 16164 10640 16204
rect 10686 16192 10692 16244
rect 10744 16232 10750 16244
rect 11057 16235 11115 16241
rect 11057 16232 11069 16235
rect 10744 16204 11069 16232
rect 10744 16192 10750 16204
rect 11057 16201 11069 16204
rect 11103 16201 11115 16235
rect 15470 16232 15476 16244
rect 11057 16195 11115 16201
rect 12452 16204 15476 16232
rect 12452 16164 12480 16204
rect 15470 16192 15476 16204
rect 15528 16192 15534 16244
rect 15562 16192 15568 16244
rect 15620 16232 15626 16244
rect 15657 16235 15715 16241
rect 15657 16232 15669 16235
rect 15620 16204 15669 16232
rect 15620 16192 15626 16204
rect 15657 16201 15669 16204
rect 15703 16201 15715 16235
rect 15657 16195 15715 16201
rect 19058 16192 19064 16244
rect 19116 16232 19122 16244
rect 20625 16235 20683 16241
rect 20625 16232 20637 16235
rect 19116 16204 20637 16232
rect 19116 16192 19122 16204
rect 20625 16201 20637 16204
rect 20671 16201 20683 16235
rect 20990 16232 20996 16244
rect 20951 16204 20996 16232
rect 20625 16195 20683 16201
rect 20990 16192 20996 16204
rect 21048 16192 21054 16244
rect 21358 16232 21364 16244
rect 21319 16204 21364 16232
rect 21358 16192 21364 16204
rect 21416 16192 21422 16244
rect 10612 16136 12480 16164
rect 17313 16167 17371 16173
rect 8297 16127 8355 16133
rect 17313 16133 17325 16167
rect 17359 16164 17371 16167
rect 17494 16164 17500 16176
rect 17359 16136 17500 16164
rect 17359 16133 17371 16136
rect 17313 16127 17371 16133
rect 17494 16124 17500 16136
rect 17552 16124 17558 16176
rect 20162 16124 20168 16176
rect 20220 16164 20226 16176
rect 20220 16136 21220 16164
rect 20220 16124 20226 16136
rect 4249 16099 4307 16105
rect 4249 16096 4261 16099
rect 3528 16068 4261 16096
rect 3421 16059 3479 16065
rect 4249 16065 4261 16068
rect 4295 16065 4307 16099
rect 4249 16059 4307 16065
rect 5261 16099 5319 16105
rect 5261 16065 5273 16099
rect 5307 16065 5319 16099
rect 5261 16059 5319 16065
rect 6825 16099 6883 16105
rect 6825 16065 6837 16099
rect 6871 16065 6883 16099
rect 6825 16059 6883 16065
rect 8849 16099 8907 16105
rect 8849 16065 8861 16099
rect 8895 16065 8907 16099
rect 8849 16059 8907 16065
rect 1394 16028 1400 16040
rect 1355 16000 1400 16028
rect 1394 15988 1400 16000
rect 1452 15988 1458 16040
rect 1762 16028 1768 16040
rect 1723 16000 1768 16028
rect 1762 15988 1768 16000
rect 1820 15988 1826 16040
rect 2133 16031 2191 16037
rect 2133 15997 2145 16031
rect 2179 15997 2191 16031
rect 2133 15991 2191 15997
rect 2501 16031 2559 16037
rect 2501 15997 2513 16031
rect 2547 16028 2559 16031
rect 3326 16028 3332 16040
rect 2547 16000 3332 16028
rect 2547 15997 2559 16000
rect 2501 15991 2559 15997
rect 2148 15960 2176 15991
rect 3326 15988 3332 16000
rect 3384 15988 3390 16040
rect 4798 15988 4804 16040
rect 4856 16028 4862 16040
rect 6840 16028 6868 16059
rect 4856 16000 6868 16028
rect 7092 16031 7150 16037
rect 4856 15988 4862 16000
rect 7092 15997 7104 16031
rect 7138 16028 7150 16031
rect 8864 16028 8892 16059
rect 9122 16056 9128 16108
rect 9180 16096 9186 16108
rect 9306 16096 9312 16108
rect 9180 16068 9312 16096
rect 9180 16056 9186 16068
rect 9306 16056 9312 16068
rect 9364 16096 9370 16108
rect 9585 16099 9643 16105
rect 9585 16096 9597 16099
rect 9364 16068 9597 16096
rect 9364 16056 9370 16068
rect 9585 16065 9597 16068
rect 9631 16065 9643 16099
rect 9585 16059 9643 16065
rect 11146 16056 11152 16108
rect 11204 16096 11210 16108
rect 11609 16099 11667 16105
rect 11609 16096 11621 16099
rect 11204 16068 11621 16096
rect 11204 16056 11210 16068
rect 11609 16065 11621 16068
rect 11655 16065 11667 16099
rect 11609 16059 11667 16065
rect 12342 16056 12348 16108
rect 12400 16096 12406 16108
rect 12437 16099 12495 16105
rect 12437 16096 12449 16099
rect 12400 16068 12449 16096
rect 12400 16056 12406 16068
rect 12437 16065 12449 16068
rect 12483 16065 12495 16099
rect 12437 16059 12495 16065
rect 12066 16028 12072 16040
rect 7138 16000 8892 16028
rect 9692 16000 12072 16028
rect 7138 15997 7150 16000
rect 7092 15991 7150 15997
rect 3050 15960 3056 15972
rect 2148 15932 3056 15960
rect 3050 15920 3056 15932
rect 3108 15920 3114 15972
rect 3970 15920 3976 15972
rect 4028 15960 4034 15972
rect 4157 15963 4215 15969
rect 4157 15960 4169 15963
rect 4028 15932 4169 15960
rect 4028 15920 4034 15932
rect 4157 15929 4169 15932
rect 4203 15929 4215 15963
rect 4157 15923 4215 15929
rect 4246 15920 4252 15972
rect 4304 15960 4310 15972
rect 4617 15963 4675 15969
rect 4617 15960 4629 15963
rect 4304 15932 4629 15960
rect 4304 15920 4310 15932
rect 4617 15929 4629 15932
rect 4663 15960 4675 15963
rect 5350 15960 5356 15972
rect 4663 15932 5356 15960
rect 4663 15929 4675 15932
rect 4617 15923 4675 15929
rect 5350 15920 5356 15932
rect 5408 15920 5414 15972
rect 5528 15963 5586 15969
rect 5528 15929 5540 15963
rect 5574 15960 5586 15963
rect 5902 15960 5908 15972
rect 5574 15932 5908 15960
rect 5574 15929 5586 15932
rect 5528 15923 5586 15929
rect 5902 15920 5908 15932
rect 5960 15920 5966 15972
rect 6730 15960 6736 15972
rect 6643 15932 6736 15960
rect 1946 15892 1952 15904
rect 1907 15864 1952 15892
rect 1946 15852 1952 15864
rect 2004 15852 2010 15904
rect 3234 15892 3240 15904
rect 3195 15864 3240 15892
rect 3234 15852 3240 15864
rect 3292 15852 3298 15904
rect 3329 15895 3387 15901
rect 3329 15861 3341 15895
rect 3375 15892 3387 15895
rect 3697 15895 3755 15901
rect 3697 15892 3709 15895
rect 3375 15864 3709 15892
rect 3375 15861 3387 15864
rect 3329 15855 3387 15861
rect 3697 15861 3709 15864
rect 3743 15861 3755 15895
rect 3697 15855 3755 15861
rect 4065 15895 4123 15901
rect 4065 15861 4077 15895
rect 4111 15892 4123 15895
rect 4430 15892 4436 15904
rect 4111 15864 4436 15892
rect 4111 15861 4123 15864
rect 4065 15855 4123 15861
rect 4430 15852 4436 15864
rect 4488 15852 4494 15904
rect 5169 15895 5227 15901
rect 5169 15861 5181 15895
rect 5215 15892 5227 15895
rect 5258 15892 5264 15904
rect 5215 15864 5264 15892
rect 5215 15861 5227 15864
rect 5169 15855 5227 15861
rect 5258 15852 5264 15864
rect 5316 15852 5322 15904
rect 6656 15901 6684 15932
rect 6730 15920 6736 15932
rect 6788 15960 6794 15972
rect 7107 15960 7135 15991
rect 6788 15932 7135 15960
rect 6788 15920 6794 15932
rect 8202 15920 8208 15972
rect 8260 15960 8266 15972
rect 9692 15960 9720 16000
rect 12066 15988 12072 16000
rect 12124 15988 12130 16040
rect 12452 16028 12480 16059
rect 17034 16056 17040 16108
rect 17092 16096 17098 16108
rect 19889 16099 19947 16105
rect 19889 16096 19901 16099
rect 17092 16068 19901 16096
rect 17092 16056 17098 16068
rect 19889 16065 19901 16068
rect 19935 16065 19947 16099
rect 19889 16059 19947 16065
rect 20272 16068 20852 16096
rect 12526 16028 12532 16040
rect 12452 16000 12532 16028
rect 12526 15988 12532 16000
rect 12584 15988 12590 16040
rect 12710 16037 12716 16040
rect 12704 16028 12716 16037
rect 12671 16000 12716 16028
rect 12704 15991 12716 16000
rect 12710 15988 12716 15991
rect 12768 15988 12774 16040
rect 13906 15988 13912 16040
rect 13964 16028 13970 16040
rect 14277 16031 14335 16037
rect 14277 16028 14289 16031
rect 13964 16000 14289 16028
rect 13964 15988 13970 16000
rect 14277 15997 14289 16000
rect 14323 15997 14335 16031
rect 14277 15991 14335 15997
rect 14544 16031 14602 16037
rect 14544 15997 14556 16031
rect 14590 16028 14602 16031
rect 15286 16028 15292 16040
rect 14590 16000 15292 16028
rect 14590 15997 14602 16000
rect 14544 15991 14602 15997
rect 9858 15969 9864 15972
rect 9852 15960 9864 15969
rect 8260 15932 9720 15960
rect 9819 15932 9864 15960
rect 8260 15920 8266 15932
rect 9852 15923 9864 15932
rect 9858 15920 9864 15923
rect 9916 15920 9922 15972
rect 11425 15963 11483 15969
rect 10060 15932 11376 15960
rect 10060 15904 10088 15932
rect 6641 15895 6699 15901
rect 6641 15861 6653 15895
rect 6687 15861 6699 15895
rect 6641 15855 6699 15861
rect 7098 15852 7104 15904
rect 7156 15892 7162 15904
rect 8665 15895 8723 15901
rect 8665 15892 8677 15895
rect 7156 15864 8677 15892
rect 7156 15852 7162 15864
rect 8665 15861 8677 15864
rect 8711 15861 8723 15895
rect 8665 15855 8723 15861
rect 8754 15852 8760 15904
rect 8812 15892 8818 15904
rect 8812 15864 8857 15892
rect 8812 15852 8818 15864
rect 8938 15852 8944 15904
rect 8996 15892 9002 15904
rect 10042 15892 10048 15904
rect 8996 15864 10048 15892
rect 8996 15852 9002 15864
rect 10042 15852 10048 15864
rect 10100 15852 10106 15904
rect 10965 15895 11023 15901
rect 10965 15861 10977 15895
rect 11011 15892 11023 15895
rect 11146 15892 11152 15904
rect 11011 15864 11152 15892
rect 11011 15861 11023 15864
rect 10965 15855 11023 15861
rect 11146 15852 11152 15864
rect 11204 15852 11210 15904
rect 11348 15892 11376 15932
rect 11425 15929 11437 15963
rect 11471 15960 11483 15963
rect 11977 15963 12035 15969
rect 11977 15960 11989 15963
rect 11471 15932 11989 15960
rect 11471 15929 11483 15932
rect 11425 15923 11483 15929
rect 11977 15929 11989 15932
rect 12023 15960 12035 15963
rect 12342 15960 12348 15972
rect 12023 15932 12348 15960
rect 12023 15929 12035 15932
rect 11977 15923 12035 15929
rect 12342 15920 12348 15932
rect 12400 15920 12406 15972
rect 12802 15920 12808 15972
rect 12860 15960 12866 15972
rect 14093 15963 14151 15969
rect 14093 15960 14105 15963
rect 12860 15932 14105 15960
rect 12860 15920 12866 15932
rect 14093 15929 14105 15932
rect 14139 15929 14151 15963
rect 14292 15960 14320 15991
rect 15286 15988 15292 16000
rect 15344 15988 15350 16040
rect 15930 16028 15936 16040
rect 15891 16000 15936 16028
rect 15930 15988 15936 16000
rect 15988 15988 15994 16040
rect 16200 16031 16258 16037
rect 16200 15997 16212 16031
rect 16246 16028 16258 16031
rect 16666 16028 16672 16040
rect 16246 16000 16672 16028
rect 16246 15997 16258 16000
rect 16200 15991 16258 15997
rect 16666 15988 16672 16000
rect 16724 15988 16730 16040
rect 20272 16037 20300 16068
rect 20824 16037 20852 16068
rect 21192 16037 21220 16136
rect 20257 16031 20315 16037
rect 20257 16028 20269 16031
rect 19260 16000 20269 16028
rect 15948 15960 15976 15988
rect 14292 15932 15976 15960
rect 14093 15923 14151 15929
rect 16298 15920 16304 15972
rect 16356 15960 16362 15972
rect 19260 15960 19288 16000
rect 20257 15997 20269 16000
rect 20303 15997 20315 16031
rect 20257 15991 20315 15997
rect 20441 16031 20499 16037
rect 20441 15997 20453 16031
rect 20487 15997 20499 16031
rect 20441 15991 20499 15997
rect 20809 16031 20867 16037
rect 20809 15997 20821 16031
rect 20855 15997 20867 16031
rect 20809 15991 20867 15997
rect 21177 16031 21235 16037
rect 21177 15997 21189 16031
rect 21223 15997 21235 16031
rect 21177 15991 21235 15997
rect 16356 15932 19288 15960
rect 19889 15963 19947 15969
rect 16356 15920 16362 15932
rect 19889 15929 19901 15963
rect 19935 15960 19947 15963
rect 20165 15963 20223 15969
rect 20165 15960 20177 15963
rect 19935 15932 20177 15960
rect 19935 15929 19947 15932
rect 19889 15923 19947 15929
rect 20165 15929 20177 15932
rect 20211 15960 20223 15963
rect 20456 15960 20484 15991
rect 20211 15932 20484 15960
rect 20211 15929 20223 15932
rect 20165 15923 20223 15929
rect 11517 15895 11575 15901
rect 11517 15892 11529 15895
rect 11348 15864 11529 15892
rect 11517 15861 11529 15864
rect 11563 15892 11575 15895
rect 12069 15895 12127 15901
rect 12069 15892 12081 15895
rect 11563 15864 12081 15892
rect 11563 15861 11575 15864
rect 11517 15855 11575 15861
rect 12069 15861 12081 15864
rect 12115 15861 12127 15895
rect 12069 15855 12127 15861
rect 13354 15852 13360 15904
rect 13412 15892 13418 15904
rect 13814 15892 13820 15904
rect 13412 15864 13820 15892
rect 13412 15852 13418 15864
rect 13814 15852 13820 15864
rect 13872 15852 13878 15904
rect 13998 15892 14004 15904
rect 13959 15864 14004 15892
rect 13998 15852 14004 15864
rect 14056 15892 14062 15904
rect 17034 15892 17040 15904
rect 14056 15864 17040 15892
rect 14056 15852 14062 15864
rect 17034 15852 17040 15864
rect 17092 15852 17098 15904
rect 17402 15852 17408 15904
rect 17460 15892 17466 15904
rect 17460 15864 17505 15892
rect 17460 15852 17466 15864
rect 1104 15802 21896 15824
rect 1104 15750 7912 15802
rect 7964 15750 7976 15802
rect 8028 15750 8040 15802
rect 8092 15750 8104 15802
rect 8156 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 15035 15802
rect 15087 15750 21896 15802
rect 1104 15728 21896 15750
rect 1670 15648 1676 15700
rect 1728 15688 1734 15700
rect 1765 15691 1823 15697
rect 1765 15688 1777 15691
rect 1728 15660 1777 15688
rect 1728 15648 1734 15660
rect 1765 15657 1777 15660
rect 1811 15688 1823 15691
rect 1811 15660 2544 15688
rect 1811 15657 1823 15660
rect 1765 15651 1823 15657
rect 1394 15580 1400 15632
rect 1452 15620 1458 15632
rect 2133 15623 2191 15629
rect 2133 15620 2145 15623
rect 1452 15592 2145 15620
rect 1452 15580 1458 15592
rect 2133 15589 2145 15592
rect 2179 15589 2191 15623
rect 2516 15620 2544 15660
rect 2590 15648 2596 15700
rect 2648 15688 2654 15700
rect 3789 15691 3847 15697
rect 3789 15688 3801 15691
rect 2648 15660 3801 15688
rect 2648 15648 2654 15660
rect 3789 15657 3801 15660
rect 3835 15657 3847 15691
rect 4430 15688 4436 15700
rect 4391 15660 4436 15688
rect 3789 15651 3847 15657
rect 4430 15648 4436 15660
rect 4488 15648 4494 15700
rect 5261 15691 5319 15697
rect 5261 15657 5273 15691
rect 5307 15657 5319 15691
rect 5261 15651 5319 15657
rect 3510 15620 3516 15632
rect 2516 15592 3516 15620
rect 2133 15583 2191 15589
rect 3510 15580 3516 15592
rect 3568 15580 3574 15632
rect 5276 15620 5304 15651
rect 5626 15648 5632 15700
rect 5684 15688 5690 15700
rect 5721 15691 5779 15697
rect 5721 15688 5733 15691
rect 5684 15660 5733 15688
rect 5684 15648 5690 15660
rect 5721 15657 5733 15660
rect 5767 15657 5779 15691
rect 5721 15651 5779 15657
rect 6089 15691 6147 15697
rect 6089 15657 6101 15691
rect 6135 15688 6147 15691
rect 6362 15688 6368 15700
rect 6135 15660 6368 15688
rect 6135 15657 6147 15660
rect 6089 15651 6147 15657
rect 6362 15648 6368 15660
rect 6420 15648 6426 15700
rect 6457 15691 6515 15697
rect 6457 15657 6469 15691
rect 6503 15688 6515 15691
rect 6917 15691 6975 15697
rect 6917 15688 6929 15691
rect 6503 15660 6929 15688
rect 6503 15657 6515 15660
rect 6457 15651 6515 15657
rect 6917 15657 6929 15660
rect 6963 15657 6975 15691
rect 6917 15651 6975 15657
rect 7374 15648 7380 15700
rect 7432 15688 7438 15700
rect 9214 15688 9220 15700
rect 7432 15660 9076 15688
rect 9175 15660 9220 15688
rect 7432 15648 7438 15660
rect 8754 15620 8760 15632
rect 5276 15592 8760 15620
rect 8754 15580 8760 15592
rect 8812 15580 8818 15632
rect 1857 15555 1915 15561
rect 1857 15521 1869 15555
rect 1903 15521 1915 15555
rect 1857 15515 1915 15521
rect 2409 15555 2467 15561
rect 2409 15521 2421 15555
rect 2455 15552 2467 15555
rect 2498 15552 2504 15564
rect 2455 15524 2504 15552
rect 2455 15521 2467 15524
rect 2409 15515 2467 15521
rect 1578 15348 1584 15360
rect 1539 15320 1584 15348
rect 1578 15308 1584 15320
rect 1636 15308 1642 15360
rect 1872 15348 1900 15515
rect 2498 15512 2504 15524
rect 2556 15512 2562 15564
rect 2676 15555 2734 15561
rect 2676 15521 2688 15555
rect 2722 15552 2734 15555
rect 4154 15552 4160 15564
rect 2722 15524 4160 15552
rect 2722 15521 2734 15524
rect 2676 15515 2734 15521
rect 4154 15512 4160 15524
rect 4212 15512 4218 15564
rect 4801 15555 4859 15561
rect 4801 15521 4813 15555
rect 4847 15552 4859 15555
rect 5258 15552 5264 15564
rect 4847 15524 5264 15552
rect 4847 15521 4859 15524
rect 4801 15515 4859 15521
rect 5258 15512 5264 15524
rect 5316 15512 5322 15564
rect 5534 15512 5540 15564
rect 5592 15552 5598 15564
rect 5629 15555 5687 15561
rect 5629 15552 5641 15555
rect 5592 15524 5641 15552
rect 5592 15512 5598 15524
rect 5629 15521 5641 15524
rect 5675 15521 5687 15555
rect 5629 15515 5687 15521
rect 6549 15555 6607 15561
rect 6549 15521 6561 15555
rect 6595 15552 6607 15555
rect 7098 15552 7104 15564
rect 6595 15524 7104 15552
rect 6595 15521 6607 15524
rect 6549 15515 6607 15521
rect 7098 15512 7104 15524
rect 7156 15512 7162 15564
rect 7285 15555 7343 15561
rect 7285 15521 7297 15555
rect 7331 15552 7343 15555
rect 7745 15555 7803 15561
rect 7745 15552 7757 15555
rect 7331 15524 7757 15552
rect 7331 15521 7343 15524
rect 7285 15515 7343 15521
rect 7745 15521 7757 15524
rect 7791 15521 7803 15555
rect 8110 15552 8116 15564
rect 8071 15524 8116 15552
rect 7745 15515 7803 15521
rect 8110 15512 8116 15524
rect 8168 15512 8174 15564
rect 9048 15552 9076 15660
rect 9214 15648 9220 15660
rect 9272 15648 9278 15700
rect 9858 15648 9864 15700
rect 9916 15688 9922 15700
rect 11057 15691 11115 15697
rect 11057 15688 11069 15691
rect 9916 15660 11069 15688
rect 9916 15648 9922 15660
rect 11057 15657 11069 15660
rect 11103 15657 11115 15691
rect 11057 15651 11115 15657
rect 11425 15691 11483 15697
rect 11425 15657 11437 15691
rect 11471 15688 11483 15691
rect 12158 15688 12164 15700
rect 11471 15660 12164 15688
rect 11471 15657 11483 15660
rect 11425 15651 11483 15657
rect 12158 15648 12164 15660
rect 12216 15648 12222 15700
rect 12253 15691 12311 15697
rect 12253 15657 12265 15691
rect 12299 15688 12311 15691
rect 12434 15688 12440 15700
rect 12299 15660 12440 15688
rect 12299 15657 12311 15660
rect 12253 15651 12311 15657
rect 12434 15648 12440 15660
rect 12492 15648 12498 15700
rect 13081 15691 13139 15697
rect 13081 15657 13093 15691
rect 13127 15688 13139 15691
rect 13262 15688 13268 15700
rect 13127 15660 13268 15688
rect 13127 15657 13139 15660
rect 13081 15651 13139 15657
rect 13262 15648 13268 15660
rect 13320 15648 13326 15700
rect 13538 15688 13544 15700
rect 13499 15660 13544 15688
rect 13538 15648 13544 15660
rect 13596 15648 13602 15700
rect 13722 15648 13728 15700
rect 13780 15688 13786 15700
rect 13909 15691 13967 15697
rect 13909 15688 13921 15691
rect 13780 15660 13921 15688
rect 13780 15648 13786 15660
rect 13909 15657 13921 15660
rect 13955 15657 13967 15691
rect 13909 15651 13967 15657
rect 14090 15648 14096 15700
rect 14148 15688 14154 15700
rect 14369 15691 14427 15697
rect 14369 15688 14381 15691
rect 14148 15660 14381 15688
rect 14148 15648 14154 15660
rect 14369 15657 14381 15660
rect 14415 15657 14427 15691
rect 14369 15651 14427 15657
rect 15289 15691 15347 15697
rect 15289 15657 15301 15691
rect 15335 15657 15347 15691
rect 15289 15651 15347 15657
rect 9125 15623 9183 15629
rect 9125 15589 9137 15623
rect 9171 15620 9183 15623
rect 9306 15620 9312 15632
rect 9171 15592 9312 15620
rect 9171 15589 9183 15592
rect 9125 15583 9183 15589
rect 9306 15580 9312 15592
rect 9364 15580 9370 15632
rect 11793 15623 11851 15629
rect 9876 15592 10171 15620
rect 9876 15552 9904 15592
rect 9950 15561 9956 15564
rect 9048 15524 9904 15552
rect 9944 15515 9956 15561
rect 10008 15552 10014 15564
rect 10143 15552 10171 15592
rect 11793 15589 11805 15623
rect 11839 15620 11851 15623
rect 11974 15620 11980 15632
rect 11839 15592 11980 15620
rect 11839 15589 11851 15592
rect 11793 15583 11851 15589
rect 11974 15580 11980 15592
rect 12032 15580 12038 15632
rect 12066 15580 12072 15632
rect 12124 15620 12130 15632
rect 13449 15623 13507 15629
rect 13449 15620 13461 15623
rect 12124 15592 13461 15620
rect 12124 15580 12130 15592
rect 13449 15589 13461 15592
rect 13495 15620 13507 15623
rect 15304 15620 15332 15651
rect 15654 15648 15660 15700
rect 15712 15688 15718 15700
rect 16117 15691 16175 15697
rect 16117 15688 16129 15691
rect 15712 15660 16129 15688
rect 15712 15648 15718 15660
rect 16117 15657 16129 15660
rect 16163 15657 16175 15691
rect 16117 15651 16175 15657
rect 16485 15691 16543 15697
rect 16485 15657 16497 15691
rect 16531 15688 16543 15691
rect 17402 15688 17408 15700
rect 16531 15660 17408 15688
rect 16531 15657 16543 15660
rect 16485 15651 16543 15657
rect 17402 15648 17408 15660
rect 17460 15648 17466 15700
rect 19334 15648 19340 15700
rect 19392 15688 19398 15700
rect 20533 15691 20591 15697
rect 20533 15688 20545 15691
rect 19392 15660 20545 15688
rect 19392 15648 19398 15660
rect 20533 15657 20545 15660
rect 20579 15688 20591 15691
rect 21082 15688 21088 15700
rect 20579 15660 20944 15688
rect 21043 15660 21088 15688
rect 20579 15657 20591 15660
rect 20533 15651 20591 15657
rect 17126 15620 17132 15632
rect 13495 15592 14964 15620
rect 15304 15592 17132 15620
rect 13495 15589 13507 15592
rect 13449 15583 13507 15589
rect 12618 15552 12624 15564
rect 10008 15524 10044 15552
rect 10143 15524 11652 15552
rect 12579 15524 12624 15552
rect 9950 15512 9956 15515
rect 10008 15512 10014 15524
rect 4893 15487 4951 15493
rect 4893 15453 4905 15487
rect 4939 15453 4951 15487
rect 4893 15447 4951 15453
rect 4908 15416 4936 15447
rect 4982 15444 4988 15496
rect 5040 15484 5046 15496
rect 5902 15484 5908 15496
rect 5040 15456 5085 15484
rect 5863 15456 5908 15484
rect 5040 15444 5046 15456
rect 5902 15444 5908 15456
rect 5960 15444 5966 15496
rect 6730 15484 6736 15496
rect 6691 15456 6736 15484
rect 6730 15444 6736 15456
rect 6788 15444 6794 15496
rect 6822 15444 6828 15496
rect 6880 15484 6886 15496
rect 7374 15484 7380 15496
rect 6880 15456 7380 15484
rect 6880 15444 6886 15456
rect 7374 15444 7380 15456
rect 7432 15444 7438 15496
rect 7466 15444 7472 15496
rect 7524 15484 7530 15496
rect 7524 15456 7569 15484
rect 7524 15444 7530 15456
rect 8754 15444 8760 15496
rect 8812 15444 8818 15496
rect 8938 15444 8944 15496
rect 8996 15484 9002 15496
rect 9309 15487 9367 15493
rect 9309 15484 9321 15487
rect 8996 15456 9321 15484
rect 8996 15444 9002 15456
rect 9309 15453 9321 15456
rect 9355 15453 9367 15487
rect 9309 15447 9367 15453
rect 9677 15487 9735 15493
rect 9677 15453 9689 15487
rect 9723 15453 9735 15487
rect 9677 15447 9735 15453
rect 6362 15416 6368 15428
rect 4908 15388 6368 15416
rect 6362 15376 6368 15388
rect 6420 15376 6426 15428
rect 8772 15416 8800 15444
rect 6656 15388 8800 15416
rect 4982 15348 4988 15360
rect 1872 15320 4988 15348
rect 4982 15308 4988 15320
rect 5040 15308 5046 15360
rect 5350 15308 5356 15360
rect 5408 15348 5414 15360
rect 6656 15348 6684 15388
rect 9122 15376 9128 15428
rect 9180 15416 9186 15428
rect 9692 15416 9720 15447
rect 11146 15416 11152 15428
rect 9180 15388 9720 15416
rect 11072 15388 11152 15416
rect 9180 15376 9186 15388
rect 5408 15320 6684 15348
rect 5408 15308 5414 15320
rect 6730 15308 6736 15360
rect 6788 15348 6794 15360
rect 8202 15348 8208 15360
rect 6788 15320 8208 15348
rect 6788 15308 6794 15320
rect 8202 15308 8208 15320
rect 8260 15308 8266 15360
rect 8757 15351 8815 15357
rect 8757 15317 8769 15351
rect 8803 15348 8815 15351
rect 11072 15348 11100 15388
rect 11146 15376 11152 15388
rect 11204 15376 11210 15428
rect 11238 15348 11244 15360
rect 8803 15320 11100 15348
rect 11199 15320 11244 15348
rect 8803 15317 8815 15320
rect 8757 15311 8815 15317
rect 11238 15308 11244 15320
rect 11296 15308 11302 15360
rect 11624 15348 11652 15524
rect 12618 15512 12624 15524
rect 12676 15552 12682 15564
rect 13998 15552 14004 15564
rect 12676 15524 14004 15552
rect 12676 15512 12682 15524
rect 13998 15512 14004 15524
rect 14056 15512 14062 15564
rect 14274 15552 14280 15564
rect 14235 15524 14280 15552
rect 14274 15512 14280 15524
rect 14332 15512 14338 15564
rect 11882 15484 11888 15496
rect 11843 15456 11888 15484
rect 11882 15444 11888 15456
rect 11940 15444 11946 15496
rect 12069 15487 12127 15493
rect 12069 15453 12081 15487
rect 12115 15453 12127 15487
rect 12710 15484 12716 15496
rect 12671 15456 12716 15484
rect 12069 15447 12127 15453
rect 12084 15416 12112 15447
rect 12710 15444 12716 15456
rect 12768 15444 12774 15496
rect 12894 15444 12900 15496
rect 12952 15484 12958 15496
rect 13722 15484 13728 15496
rect 12952 15456 12997 15484
rect 13683 15456 13728 15484
rect 12952 15444 12958 15456
rect 13722 15444 13728 15456
rect 13780 15484 13786 15496
rect 14461 15487 14519 15493
rect 14461 15484 14473 15487
rect 13780 15456 14473 15484
rect 13780 15444 13786 15456
rect 14461 15453 14473 15456
rect 14507 15453 14519 15487
rect 14936 15484 14964 15592
rect 17126 15580 17132 15592
rect 17184 15580 17190 15632
rect 17218 15580 17224 15632
rect 17276 15620 17282 15632
rect 20806 15620 20812 15632
rect 17276 15592 17321 15620
rect 17420 15592 20812 15620
rect 17276 15580 17282 15592
rect 15470 15512 15476 15564
rect 15528 15552 15534 15564
rect 15657 15555 15715 15561
rect 15657 15552 15669 15555
rect 15528 15524 15669 15552
rect 15528 15512 15534 15524
rect 15657 15521 15669 15524
rect 15703 15521 15715 15555
rect 15657 15515 15715 15521
rect 15749 15555 15807 15561
rect 15749 15521 15761 15555
rect 15795 15552 15807 15555
rect 16850 15552 16856 15564
rect 15795 15524 16856 15552
rect 15795 15521 15807 15524
rect 15749 15515 15807 15521
rect 16850 15512 16856 15524
rect 16908 15512 16914 15564
rect 17420 15552 17448 15592
rect 20806 15580 20812 15592
rect 20864 15580 20870 15632
rect 20916 15620 20944 15660
rect 21082 15648 21088 15660
rect 21140 15648 21146 15700
rect 21450 15688 21456 15700
rect 21411 15660 21456 15688
rect 21450 15648 21456 15660
rect 21508 15648 21514 15700
rect 20916 15592 21312 15620
rect 18138 15552 18144 15564
rect 16960 15524 17448 15552
rect 18099 15524 18144 15552
rect 15838 15484 15844 15496
rect 14936 15456 15844 15484
rect 14461 15447 14519 15453
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 15933 15487 15991 15493
rect 15933 15453 15945 15487
rect 15979 15453 15991 15487
rect 15933 15447 15991 15453
rect 13814 15416 13820 15428
rect 12084 15388 13820 15416
rect 13814 15376 13820 15388
rect 13872 15376 13878 15428
rect 13998 15376 14004 15428
rect 14056 15416 14062 15428
rect 14737 15419 14795 15425
rect 14737 15416 14749 15419
rect 14056 15388 14749 15416
rect 14056 15376 14062 15388
rect 14737 15385 14749 15388
rect 14783 15385 14795 15419
rect 14737 15379 14795 15385
rect 15286 15376 15292 15428
rect 15344 15416 15350 15428
rect 15948 15416 15976 15447
rect 16298 15444 16304 15496
rect 16356 15484 16362 15496
rect 16577 15487 16635 15493
rect 16577 15484 16589 15487
rect 16356 15456 16589 15484
rect 16356 15444 16362 15456
rect 16577 15453 16589 15456
rect 16623 15453 16635 15487
rect 16577 15447 16635 15453
rect 16669 15487 16727 15493
rect 16669 15453 16681 15487
rect 16715 15453 16727 15487
rect 16960 15484 16988 15524
rect 18138 15512 18144 15524
rect 18196 15512 18202 15564
rect 21284 15561 21312 15592
rect 20901 15555 20959 15561
rect 20901 15552 20913 15555
rect 20732 15524 20913 15552
rect 16669 15447 16727 15453
rect 16776 15456 16988 15484
rect 16684 15416 16712 15447
rect 15344 15388 16712 15416
rect 15344 15376 15350 15388
rect 16776 15348 16804 15456
rect 17034 15444 17040 15496
rect 17092 15484 17098 15496
rect 18233 15487 18291 15493
rect 18233 15484 18245 15487
rect 17092 15456 18245 15484
rect 17092 15444 17098 15456
rect 18233 15453 18245 15456
rect 18279 15453 18291 15487
rect 18233 15447 18291 15453
rect 18325 15487 18383 15493
rect 18325 15453 18337 15487
rect 18371 15453 18383 15487
rect 18325 15447 18383 15453
rect 16850 15376 16856 15428
rect 16908 15416 16914 15428
rect 16945 15419 17003 15425
rect 16945 15416 16957 15419
rect 16908 15388 16957 15416
rect 16908 15376 16914 15388
rect 16945 15385 16957 15388
rect 16991 15385 17003 15419
rect 16945 15379 17003 15385
rect 17954 15376 17960 15428
rect 18012 15416 18018 15428
rect 18340 15416 18368 15447
rect 18012 15388 18368 15416
rect 18012 15376 18018 15388
rect 18690 15376 18696 15428
rect 18748 15416 18754 15428
rect 20732 15425 20760 15524
rect 20901 15521 20913 15524
rect 20947 15521 20959 15555
rect 20901 15515 20959 15521
rect 21269 15555 21327 15561
rect 21269 15521 21281 15555
rect 21315 15521 21327 15555
rect 21269 15515 21327 15521
rect 20717 15419 20775 15425
rect 20717 15416 20729 15419
rect 18748 15388 20729 15416
rect 18748 15376 18754 15388
rect 20717 15385 20729 15388
rect 20763 15385 20775 15419
rect 20717 15379 20775 15385
rect 11624 15320 16804 15348
rect 17773 15351 17831 15357
rect 17773 15317 17785 15351
rect 17819 15348 17831 15351
rect 19150 15348 19156 15360
rect 17819 15320 19156 15348
rect 17819 15317 17831 15320
rect 17773 15311 17831 15317
rect 19150 15308 19156 15320
rect 19208 15308 19214 15360
rect 1104 15258 21896 15280
rect 1104 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 4575 15258
rect 4627 15206 4639 15258
rect 4691 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 18308 15258
rect 18360 15206 18372 15258
rect 18424 15206 18436 15258
rect 18488 15206 18500 15258
rect 18552 15206 21896 15258
rect 1104 15184 21896 15206
rect 1949 15147 2007 15153
rect 1949 15113 1961 15147
rect 1995 15144 2007 15147
rect 3234 15144 3240 15156
rect 1995 15116 3240 15144
rect 1995 15113 2007 15116
rect 1949 15107 2007 15113
rect 3234 15104 3240 15116
rect 3292 15104 3298 15156
rect 3970 15144 3976 15156
rect 3931 15116 3976 15144
rect 3970 15104 3976 15116
rect 4028 15104 4034 15156
rect 5074 15144 5080 15156
rect 4632 15116 5080 15144
rect 1762 15076 1768 15088
rect 1723 15048 1768 15076
rect 1762 15036 1768 15048
rect 1820 15036 1826 15088
rect 2777 15079 2835 15085
rect 2777 15076 2789 15079
rect 2424 15048 2789 15076
rect 2424 15017 2452 15048
rect 2777 15045 2789 15048
rect 2823 15045 2835 15079
rect 2777 15039 2835 15045
rect 2409 15011 2467 15017
rect 2409 14977 2421 15011
rect 2455 14977 2467 15011
rect 2590 15008 2596 15020
rect 2551 14980 2596 15008
rect 2409 14971 2467 14977
rect 2590 14968 2596 14980
rect 2648 14968 2654 15020
rect 3421 15011 3479 15017
rect 3421 14977 3433 15011
rect 3467 15008 3479 15011
rect 4154 15008 4160 15020
rect 3467 14980 4160 15008
rect 3467 14977 3479 14980
rect 3421 14971 3479 14977
rect 4154 14968 4160 14980
rect 4212 15008 4218 15020
rect 4632 15017 4660 15116
rect 5074 15104 5080 15116
rect 5132 15104 5138 15156
rect 6362 15144 6368 15156
rect 6275 15116 6368 15144
rect 6362 15104 6368 15116
rect 6420 15144 6426 15156
rect 6730 15144 6736 15156
rect 6420 15116 6736 15144
rect 6420 15104 6426 15116
rect 6730 15104 6736 15116
rect 6788 15104 6794 15156
rect 7742 15104 7748 15156
rect 7800 15144 7806 15156
rect 9861 15147 9919 15153
rect 7800 15116 9812 15144
rect 7800 15104 7806 15116
rect 5902 15036 5908 15088
rect 5960 15076 5966 15088
rect 6181 15079 6239 15085
rect 6181 15076 6193 15079
rect 5960 15048 6193 15076
rect 5960 15036 5966 15048
rect 6181 15045 6193 15048
rect 6227 15076 6239 15079
rect 7466 15076 7472 15088
rect 6227 15048 7472 15076
rect 6227 15045 6239 15048
rect 6181 15039 6239 15045
rect 7466 15036 7472 15048
rect 7524 15036 7530 15088
rect 8018 15076 8024 15088
rect 7760 15048 8024 15076
rect 4617 15011 4675 15017
rect 4617 15008 4629 15011
rect 4212 14980 4629 15008
rect 4212 14968 4218 14980
rect 4617 14977 4629 14980
rect 4663 14977 4675 15011
rect 4798 15008 4804 15020
rect 4759 14980 4804 15008
rect 4617 14971 4675 14977
rect 4798 14968 4804 14980
rect 4856 14968 4862 15020
rect 7760 15017 7788 15048
rect 8018 15036 8024 15048
rect 8076 15036 8082 15088
rect 8113 15079 8171 15085
rect 8113 15045 8125 15079
rect 8159 15076 8171 15079
rect 8202 15076 8208 15088
rect 8159 15048 8208 15076
rect 8159 15045 8171 15048
rect 8113 15039 8171 15045
rect 8202 15036 8208 15048
rect 8260 15076 8266 15088
rect 8260 15048 8524 15076
rect 8260 15036 8266 15048
rect 7745 15011 7803 15017
rect 7745 14977 7757 15011
rect 7791 14977 7803 15011
rect 7926 15008 7932 15020
rect 7839 14980 7932 15008
rect 7745 14971 7803 14977
rect 7926 14968 7932 14980
rect 7984 15008 7990 15020
rect 8386 15008 8392 15020
rect 7984 14980 8392 15008
rect 7984 14968 7990 14980
rect 8386 14968 8392 14980
rect 8444 14968 8450 15020
rect 1578 14940 1584 14952
rect 1491 14912 1584 14940
rect 1578 14900 1584 14912
rect 1636 14940 1642 14952
rect 4338 14940 4344 14952
rect 1636 14912 3924 14940
rect 4299 14912 4344 14940
rect 1636 14900 1642 14912
rect 1489 14875 1547 14881
rect 1489 14841 1501 14875
rect 1535 14872 1547 14875
rect 3896 14872 3924 14912
rect 4338 14900 4344 14912
rect 4396 14900 4402 14952
rect 5068 14943 5126 14949
rect 5068 14909 5080 14943
rect 5114 14940 5126 14943
rect 5350 14940 5356 14952
rect 5114 14912 5356 14940
rect 5114 14909 5126 14912
rect 5068 14903 5126 14909
rect 5350 14900 5356 14912
rect 5408 14900 5414 14952
rect 7558 14900 7564 14952
rect 7616 14940 7622 14952
rect 8496 14949 8524 15048
rect 9784 15008 9812 15116
rect 9861 15113 9873 15147
rect 9907 15144 9919 15147
rect 9950 15144 9956 15156
rect 9907 15116 9956 15144
rect 9907 15113 9919 15116
rect 9861 15107 9919 15113
rect 9950 15104 9956 15116
rect 10008 15144 10014 15156
rect 10594 15144 10600 15156
rect 10008 15116 10600 15144
rect 10008 15104 10014 15116
rect 10594 15104 10600 15116
rect 10652 15104 10658 15156
rect 11517 15147 11575 15153
rect 11517 15113 11529 15147
rect 11563 15144 11575 15147
rect 11882 15144 11888 15156
rect 11563 15116 11888 15144
rect 11563 15113 11575 15116
rect 11517 15107 11575 15113
rect 11882 15104 11888 15116
rect 11940 15104 11946 15156
rect 15657 15147 15715 15153
rect 15657 15113 15669 15147
rect 15703 15144 15715 15147
rect 15930 15144 15936 15156
rect 15703 15116 15936 15144
rect 15703 15113 15715 15116
rect 15657 15107 15715 15113
rect 15930 15104 15936 15116
rect 15988 15144 15994 15156
rect 16574 15144 16580 15156
rect 15988 15116 16580 15144
rect 15988 15104 15994 15116
rect 16574 15104 16580 15116
rect 16632 15104 16638 15156
rect 17954 15104 17960 15156
rect 18012 15144 18018 15156
rect 19429 15147 19487 15153
rect 19429 15144 19441 15147
rect 18012 15116 19441 15144
rect 18012 15104 18018 15116
rect 19429 15113 19441 15116
rect 19475 15113 19487 15147
rect 20990 15144 20996 15156
rect 20951 15116 20996 15144
rect 19429 15107 19487 15113
rect 20990 15104 20996 15116
rect 21048 15104 21054 15156
rect 11238 15036 11244 15088
rect 11296 15076 11302 15088
rect 12066 15076 12072 15088
rect 11296 15048 12072 15076
rect 11296 15036 11302 15048
rect 12066 15036 12072 15048
rect 12124 15036 12130 15088
rect 13722 15036 13728 15088
rect 13780 15076 13786 15088
rect 13817 15079 13875 15085
rect 13817 15076 13829 15079
rect 13780 15048 13829 15076
rect 13780 15036 13786 15048
rect 13817 15045 13829 15048
rect 13863 15045 13875 15079
rect 13817 15039 13875 15045
rect 16025 15079 16083 15085
rect 16025 15045 16037 15079
rect 16071 15076 16083 15079
rect 16298 15076 16304 15088
rect 16071 15048 16304 15076
rect 16071 15045 16083 15048
rect 16025 15039 16083 15045
rect 16298 15036 16304 15048
rect 16356 15036 16362 15088
rect 10597 15011 10655 15017
rect 10597 15008 10609 15011
rect 9784 14980 10609 15008
rect 10597 14977 10609 14980
rect 10643 15008 10655 15011
rect 10870 15008 10876 15020
rect 10643 14980 10876 15008
rect 10643 14977 10655 14980
rect 10597 14971 10655 14977
rect 10870 14968 10876 14980
rect 10928 14968 10934 15020
rect 12158 15008 12164 15020
rect 12119 14980 12164 15008
rect 12158 14968 12164 14980
rect 12216 14968 12222 15020
rect 13909 15011 13967 15017
rect 13909 14977 13921 15011
rect 13955 15008 13967 15011
rect 14274 15008 14280 15020
rect 13955 14980 14280 15008
rect 13955 14977 13967 14980
rect 13909 14971 13967 14977
rect 14274 14968 14280 14980
rect 14332 14968 14338 15020
rect 15378 15008 15384 15020
rect 15339 14980 15384 15008
rect 15378 14968 15384 14980
rect 15436 14968 15442 15020
rect 15488 14980 16252 15008
rect 8297 14943 8355 14949
rect 8297 14940 8309 14943
rect 7616 14912 8309 14940
rect 7616 14900 7622 14912
rect 8297 14909 8309 14912
rect 8343 14909 8355 14943
rect 8297 14903 8355 14909
rect 8481 14943 8539 14949
rect 8481 14909 8493 14943
rect 8527 14940 8539 14943
rect 9122 14940 9128 14952
rect 8527 14912 9128 14940
rect 8527 14909 8539 14912
rect 8481 14903 8539 14909
rect 9122 14900 9128 14912
rect 9180 14900 9186 14952
rect 9858 14900 9864 14952
rect 9916 14940 9922 14952
rect 10413 14943 10471 14949
rect 10413 14940 10425 14943
rect 9916 14912 10425 14940
rect 9916 14900 9922 14912
rect 10413 14909 10425 14912
rect 10459 14940 10471 14943
rect 11241 14943 11299 14949
rect 10459 14912 11100 14940
rect 10459 14909 10471 14912
rect 10413 14903 10471 14909
rect 6086 14872 6092 14884
rect 1535 14844 3280 14872
rect 3896 14844 6092 14872
rect 1535 14841 1547 14844
rect 1489 14835 1547 14841
rect 2317 14807 2375 14813
rect 2317 14773 2329 14807
rect 2363 14804 2375 14807
rect 2590 14804 2596 14816
rect 2363 14776 2596 14804
rect 2363 14773 2375 14776
rect 2317 14767 2375 14773
rect 2590 14764 2596 14776
rect 2648 14764 2654 14816
rect 3050 14764 3056 14816
rect 3108 14804 3114 14816
rect 3252 14813 3280 14844
rect 6086 14832 6092 14844
rect 6144 14832 6150 14884
rect 7193 14875 7251 14881
rect 7193 14841 7205 14875
rect 7239 14872 7251 14875
rect 7653 14875 7711 14881
rect 7653 14872 7665 14875
rect 7239 14844 7665 14872
rect 7239 14841 7251 14844
rect 7193 14835 7251 14841
rect 7653 14841 7665 14844
rect 7699 14872 7711 14875
rect 8748 14875 8806 14881
rect 7699 14844 8708 14872
rect 7699 14841 7711 14844
rect 7653 14835 7711 14841
rect 8680 14816 8708 14844
rect 8748 14841 8760 14875
rect 8794 14872 8806 14875
rect 8938 14872 8944 14884
rect 8794 14844 8944 14872
rect 8794 14841 8806 14844
rect 8748 14835 8806 14841
rect 8938 14832 8944 14844
rect 8996 14832 9002 14884
rect 11072 14872 11100 14912
rect 11241 14909 11253 14943
rect 11287 14940 11299 14943
rect 11885 14943 11943 14949
rect 11885 14940 11897 14943
rect 11287 14912 11897 14940
rect 11287 14909 11299 14912
rect 11241 14903 11299 14909
rect 11885 14909 11897 14912
rect 11931 14940 11943 14943
rect 12066 14940 12072 14952
rect 11931 14912 12072 14940
rect 11931 14909 11943 14912
rect 11885 14903 11943 14909
rect 12066 14900 12072 14912
rect 12124 14900 12130 14952
rect 12437 14943 12495 14949
rect 12437 14909 12449 14943
rect 12483 14940 12495 14943
rect 12526 14940 12532 14952
rect 12483 14912 12532 14940
rect 12483 14909 12495 14912
rect 12437 14903 12495 14909
rect 12526 14900 12532 14912
rect 12584 14900 12590 14952
rect 13170 14900 13176 14952
rect 13228 14940 13234 14952
rect 15488 14940 15516 14980
rect 15838 14940 15844 14952
rect 13228 14912 15516 14940
rect 15799 14912 15844 14940
rect 13228 14900 13234 14912
rect 15838 14900 15844 14912
rect 15896 14900 15902 14952
rect 11330 14872 11336 14884
rect 11072 14844 11336 14872
rect 11330 14832 11336 14844
rect 11388 14832 11394 14884
rect 11425 14875 11483 14881
rect 11425 14841 11437 14875
rect 11471 14872 11483 14875
rect 12704 14875 12762 14881
rect 11471 14844 12020 14872
rect 11471 14841 11483 14844
rect 11425 14835 11483 14841
rect 11992 14816 12020 14844
rect 12704 14841 12716 14875
rect 12750 14872 12762 14875
rect 12802 14872 12808 14884
rect 12750 14844 12808 14872
rect 12750 14841 12762 14844
rect 12704 14835 12762 14841
rect 12802 14832 12808 14844
rect 12860 14832 12866 14884
rect 15197 14875 15255 14881
rect 15197 14841 15209 14875
rect 15243 14872 15255 14875
rect 16114 14872 16120 14884
rect 15243 14844 16120 14872
rect 15243 14841 15255 14844
rect 15197 14835 15255 14841
rect 16114 14832 16120 14844
rect 16172 14832 16178 14884
rect 16224 14872 16252 14980
rect 17310 14968 17316 15020
rect 17368 15008 17374 15020
rect 18049 15011 18107 15017
rect 18049 15008 18061 15011
rect 17368 14980 18061 15008
rect 17368 14968 17374 14980
rect 18049 14977 18061 14980
rect 18095 14977 18107 15011
rect 20162 15008 20168 15020
rect 20123 14980 20168 15008
rect 18049 14971 18107 14977
rect 20162 14968 20168 14980
rect 20220 14968 20226 15020
rect 16301 14943 16359 14949
rect 16301 14909 16313 14943
rect 16347 14940 16359 14943
rect 16390 14940 16396 14952
rect 16347 14912 16396 14940
rect 16347 14909 16359 14912
rect 16301 14903 16359 14909
rect 16390 14900 16396 14912
rect 16448 14900 16454 14952
rect 16568 14943 16626 14949
rect 16568 14909 16580 14943
rect 16614 14940 16626 14943
rect 17954 14940 17960 14952
rect 16614 14912 17960 14940
rect 16614 14909 16626 14912
rect 16568 14903 16626 14909
rect 17954 14900 17960 14912
rect 18012 14900 18018 14952
rect 19889 14943 19947 14949
rect 19889 14940 19901 14943
rect 18156 14912 19901 14940
rect 18156 14872 18184 14912
rect 19889 14909 19901 14912
rect 19935 14909 19947 14943
rect 20806 14940 20812 14952
rect 20767 14912 20812 14940
rect 19889 14903 19947 14909
rect 20806 14900 20812 14912
rect 20864 14900 20870 14952
rect 16224 14844 18184 14872
rect 18316 14875 18374 14881
rect 18316 14841 18328 14875
rect 18362 14872 18374 14875
rect 18874 14872 18880 14884
rect 18362 14844 18880 14872
rect 18362 14841 18374 14844
rect 18316 14835 18374 14841
rect 18874 14832 18880 14844
rect 18932 14832 18938 14884
rect 3145 14807 3203 14813
rect 3145 14804 3157 14807
rect 3108 14776 3157 14804
rect 3108 14764 3114 14776
rect 3145 14773 3157 14776
rect 3191 14773 3203 14807
rect 3145 14767 3203 14773
rect 3237 14807 3295 14813
rect 3237 14773 3249 14807
rect 3283 14804 3295 14807
rect 3418 14804 3424 14816
rect 3283 14776 3424 14804
rect 3283 14773 3295 14776
rect 3237 14767 3295 14773
rect 3418 14764 3424 14776
rect 3476 14764 3482 14816
rect 3602 14804 3608 14816
rect 3563 14776 3608 14804
rect 3602 14764 3608 14776
rect 3660 14764 3666 14816
rect 4433 14807 4491 14813
rect 4433 14773 4445 14807
rect 4479 14804 4491 14807
rect 5166 14804 5172 14816
rect 4479 14776 5172 14804
rect 4479 14773 4491 14776
rect 4433 14767 4491 14773
rect 5166 14764 5172 14776
rect 5224 14764 5230 14816
rect 6730 14764 6736 14816
rect 6788 14804 6794 14816
rect 6825 14807 6883 14813
rect 6825 14804 6837 14807
rect 6788 14776 6837 14804
rect 6788 14764 6794 14776
rect 6825 14773 6837 14776
rect 6871 14773 6883 14807
rect 7282 14804 7288 14816
rect 7243 14776 7288 14804
rect 6825 14767 6883 14773
rect 7282 14764 7288 14776
rect 7340 14764 7346 14816
rect 8662 14764 8668 14816
rect 8720 14764 8726 14816
rect 10045 14807 10103 14813
rect 10045 14773 10057 14807
rect 10091 14804 10103 14807
rect 10134 14804 10140 14816
rect 10091 14776 10140 14804
rect 10091 14773 10103 14776
rect 10045 14767 10103 14773
rect 10134 14764 10140 14776
rect 10192 14764 10198 14816
rect 10410 14764 10416 14816
rect 10468 14804 10474 14816
rect 10505 14807 10563 14813
rect 10505 14804 10517 14807
rect 10468 14776 10517 14804
rect 10468 14764 10474 14776
rect 10505 14773 10517 14776
rect 10551 14804 10563 14807
rect 10873 14807 10931 14813
rect 10873 14804 10885 14807
rect 10551 14776 10885 14804
rect 10551 14773 10563 14776
rect 10505 14767 10563 14773
rect 10873 14773 10885 14776
rect 10919 14773 10931 14807
rect 11974 14804 11980 14816
rect 11935 14776 11980 14804
rect 10873 14767 10931 14773
rect 11974 14764 11980 14776
rect 12032 14764 12038 14816
rect 14090 14764 14096 14816
rect 14148 14804 14154 14816
rect 14829 14807 14887 14813
rect 14829 14804 14841 14807
rect 14148 14776 14841 14804
rect 14148 14764 14154 14776
rect 14829 14773 14841 14776
rect 14875 14773 14887 14807
rect 15286 14804 15292 14816
rect 15247 14776 15292 14804
rect 14829 14767 14887 14773
rect 15286 14764 15292 14776
rect 15344 14764 15350 14816
rect 16022 14764 16028 14816
rect 16080 14804 16086 14816
rect 17681 14807 17739 14813
rect 17681 14804 17693 14807
rect 16080 14776 17693 14804
rect 16080 14764 16086 14776
rect 17681 14773 17693 14776
rect 17727 14773 17739 14807
rect 17681 14767 17739 14773
rect 19518 14764 19524 14816
rect 19576 14804 19582 14816
rect 21174 14804 21180 14816
rect 19576 14776 19621 14804
rect 21135 14776 21180 14804
rect 19576 14764 19582 14776
rect 21174 14764 21180 14776
rect 21232 14764 21238 14816
rect 1104 14714 21896 14736
rect 1104 14662 7912 14714
rect 7964 14662 7976 14714
rect 8028 14662 8040 14714
rect 8092 14662 8104 14714
rect 8156 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 15035 14714
rect 15087 14662 21896 14714
rect 1104 14640 21896 14662
rect 1854 14600 1860 14612
rect 1815 14572 1860 14600
rect 1854 14560 1860 14572
rect 1912 14560 1918 14612
rect 2685 14603 2743 14609
rect 2685 14569 2697 14603
rect 2731 14600 2743 14603
rect 3050 14600 3056 14612
rect 2731 14572 3056 14600
rect 2731 14569 2743 14572
rect 2685 14563 2743 14569
rect 3050 14560 3056 14572
rect 3108 14560 3114 14612
rect 3145 14603 3203 14609
rect 3145 14569 3157 14603
rect 3191 14600 3203 14603
rect 3602 14600 3608 14612
rect 3191 14572 3608 14600
rect 3191 14569 3203 14572
rect 3145 14563 3203 14569
rect 3602 14560 3608 14572
rect 3660 14560 3666 14612
rect 3786 14600 3792 14612
rect 3747 14572 3792 14600
rect 3786 14560 3792 14572
rect 3844 14560 3850 14612
rect 3970 14560 3976 14612
rect 4028 14600 4034 14612
rect 4065 14603 4123 14609
rect 4065 14600 4077 14603
rect 4028 14572 4077 14600
rect 4028 14560 4034 14572
rect 4065 14569 4077 14572
rect 4111 14569 4123 14603
rect 4065 14563 4123 14569
rect 4338 14560 4344 14612
rect 4396 14600 4402 14612
rect 4893 14603 4951 14609
rect 4893 14600 4905 14603
rect 4396 14572 4905 14600
rect 4396 14560 4402 14572
rect 4893 14569 4905 14572
rect 4939 14600 4951 14603
rect 5718 14600 5724 14612
rect 4939 14572 5724 14600
rect 4939 14569 4951 14572
rect 4893 14563 4951 14569
rect 5718 14560 5724 14572
rect 5776 14560 5782 14612
rect 5810 14560 5816 14612
rect 5868 14600 5874 14612
rect 6546 14600 6552 14612
rect 5868 14572 6552 14600
rect 5868 14560 5874 14572
rect 6546 14560 6552 14572
rect 6604 14560 6610 14612
rect 6733 14603 6791 14609
rect 6733 14569 6745 14603
rect 6779 14600 6791 14603
rect 7006 14600 7012 14612
rect 6779 14572 7012 14600
rect 6779 14569 6791 14572
rect 6733 14563 6791 14569
rect 7006 14560 7012 14572
rect 7064 14560 7070 14612
rect 7101 14603 7159 14609
rect 7101 14569 7113 14603
rect 7147 14600 7159 14603
rect 7282 14600 7288 14612
rect 7147 14572 7288 14600
rect 7147 14569 7159 14572
rect 7101 14563 7159 14569
rect 7282 14560 7288 14572
rect 7340 14560 7346 14612
rect 9858 14600 9864 14612
rect 7576 14572 9864 14600
rect 5905 14535 5963 14541
rect 3068 14504 3648 14532
rect 1670 14464 1676 14476
rect 1631 14436 1676 14464
rect 1670 14424 1676 14436
rect 1728 14424 1734 14476
rect 2038 14464 2044 14476
rect 1999 14436 2044 14464
rect 2038 14424 2044 14436
rect 2096 14424 2102 14476
rect 2682 14424 2688 14476
rect 2740 14464 2746 14476
rect 3068 14464 3096 14504
rect 3620 14473 3648 14504
rect 5905 14501 5917 14535
rect 5951 14532 5963 14535
rect 6457 14535 6515 14541
rect 6457 14532 6469 14535
rect 5951 14504 6469 14532
rect 5951 14501 5963 14504
rect 5905 14495 5963 14501
rect 6457 14501 6469 14504
rect 6503 14532 6515 14535
rect 6822 14532 6828 14544
rect 6503 14504 6828 14532
rect 6503 14501 6515 14504
rect 6457 14495 6515 14501
rect 6822 14492 6828 14504
rect 6880 14532 6886 14544
rect 7576 14532 7604 14572
rect 9858 14560 9864 14572
rect 9916 14560 9922 14612
rect 10226 14600 10232 14612
rect 10187 14572 10232 14600
rect 10226 14560 10232 14572
rect 10284 14560 10290 14612
rect 10689 14603 10747 14609
rect 10689 14600 10701 14603
rect 10520 14572 10701 14600
rect 8202 14532 8208 14544
rect 6880 14504 7604 14532
rect 7760 14504 8208 14532
rect 6880 14492 6886 14504
rect 2740 14436 3096 14464
rect 3605 14467 3663 14473
rect 2740 14424 2746 14436
rect 3605 14433 3617 14467
rect 3651 14433 3663 14467
rect 3605 14427 3663 14433
rect 3786 14424 3792 14476
rect 3844 14464 3850 14476
rect 4433 14467 4491 14473
rect 4433 14464 4445 14467
rect 3844 14436 4445 14464
rect 3844 14424 3850 14436
rect 4433 14433 4445 14436
rect 4479 14433 4491 14467
rect 4433 14427 4491 14433
rect 4525 14467 4583 14473
rect 4525 14433 4537 14467
rect 4571 14464 4583 14467
rect 4798 14464 4804 14476
rect 4571 14436 4804 14464
rect 4571 14433 4583 14436
rect 4525 14427 4583 14433
rect 4798 14424 4804 14436
rect 4856 14424 4862 14476
rect 7561 14467 7619 14473
rect 7561 14433 7573 14467
rect 7607 14464 7619 14467
rect 7760 14464 7788 14504
rect 8202 14492 8208 14504
rect 8260 14492 8266 14544
rect 10520 14532 10548 14572
rect 10689 14569 10701 14572
rect 10735 14600 10747 14603
rect 10778 14600 10784 14612
rect 10735 14572 10784 14600
rect 10735 14569 10747 14572
rect 10689 14563 10747 14569
rect 10778 14560 10784 14572
rect 10836 14560 10842 14612
rect 11054 14600 11060 14612
rect 11015 14572 11060 14600
rect 11054 14560 11060 14572
rect 11112 14560 11118 14612
rect 11146 14560 11152 14612
rect 11204 14600 11210 14612
rect 11517 14603 11575 14609
rect 11517 14600 11529 14603
rect 11204 14572 11529 14600
rect 11204 14560 11210 14572
rect 11517 14569 11529 14572
rect 11563 14569 11575 14603
rect 11517 14563 11575 14569
rect 11790 14560 11796 14612
rect 11848 14600 11854 14612
rect 12253 14603 12311 14609
rect 12253 14600 12265 14603
rect 11848 14572 12265 14600
rect 11848 14560 11854 14572
rect 12253 14569 12265 14572
rect 12299 14600 12311 14603
rect 12434 14600 12440 14612
rect 12299 14572 12440 14600
rect 12299 14569 12311 14572
rect 12253 14563 12311 14569
rect 12434 14560 12440 14572
rect 12492 14560 12498 14612
rect 12529 14603 12587 14609
rect 12529 14569 12541 14603
rect 12575 14600 12587 14603
rect 13538 14600 13544 14612
rect 12575 14572 13544 14600
rect 12575 14569 12587 14572
rect 12529 14563 12587 14569
rect 13538 14560 13544 14572
rect 13596 14560 13602 14612
rect 14274 14600 14280 14612
rect 13648 14572 14280 14600
rect 8588 14504 10548 14532
rect 10597 14535 10655 14541
rect 7834 14473 7840 14476
rect 7607 14436 7788 14464
rect 7607 14433 7619 14436
rect 7561 14427 7619 14433
rect 7828 14427 7840 14473
rect 7892 14464 7898 14476
rect 7892 14436 7928 14464
rect 7834 14424 7840 14427
rect 7892 14424 7898 14436
rect 8110 14424 8116 14476
rect 8168 14464 8174 14476
rect 8588 14464 8616 14504
rect 10597 14501 10609 14535
rect 10643 14532 10655 14535
rect 13648 14532 13676 14572
rect 14274 14560 14280 14572
rect 14332 14600 14338 14612
rect 15838 14600 15844 14612
rect 14332 14572 15844 14600
rect 14332 14560 14338 14572
rect 15838 14560 15844 14572
rect 15896 14560 15902 14612
rect 19337 14603 19395 14609
rect 19337 14569 19349 14603
rect 19383 14600 19395 14603
rect 19518 14600 19524 14612
rect 19383 14572 19524 14600
rect 19383 14569 19395 14572
rect 19337 14563 19395 14569
rect 19518 14560 19524 14572
rect 19576 14560 19582 14612
rect 20441 14603 20499 14609
rect 20441 14600 20453 14603
rect 19628 14572 20453 14600
rect 10643 14504 12020 14532
rect 10643 14501 10655 14504
rect 10597 14495 10655 14501
rect 8168 14436 8616 14464
rect 8168 14424 8174 14436
rect 9030 14424 9036 14476
rect 9088 14464 9094 14476
rect 9217 14467 9275 14473
rect 9217 14464 9229 14467
rect 9088 14436 9229 14464
rect 9088 14424 9094 14436
rect 9217 14433 9229 14436
rect 9263 14433 9275 14467
rect 11425 14467 11483 14473
rect 11425 14464 11437 14467
rect 9217 14427 9275 14433
rect 10980 14436 11437 14464
rect 10980 14408 11008 14436
rect 11425 14433 11437 14436
rect 11471 14433 11483 14467
rect 11425 14427 11483 14433
rect 2314 14396 2320 14408
rect 2275 14368 2320 14396
rect 2314 14356 2320 14368
rect 2372 14356 2378 14408
rect 3237 14399 3295 14405
rect 3237 14396 3249 14399
rect 2976 14368 3249 14396
rect 2590 14288 2596 14340
rect 2648 14328 2654 14340
rect 2777 14331 2835 14337
rect 2777 14328 2789 14331
rect 2648 14300 2789 14328
rect 2648 14288 2654 14300
rect 2777 14297 2789 14300
rect 2823 14297 2835 14331
rect 2777 14291 2835 14297
rect 1394 14220 1400 14272
rect 1452 14260 1458 14272
rect 1489 14263 1547 14269
rect 1489 14260 1501 14263
rect 1452 14232 1501 14260
rect 1452 14220 1458 14232
rect 1489 14229 1501 14232
rect 1535 14260 1547 14263
rect 2976 14260 3004 14368
rect 3237 14365 3249 14368
rect 3283 14365 3295 14399
rect 3237 14359 3295 14365
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14396 3479 14399
rect 4154 14396 4160 14408
rect 3467 14368 4160 14396
rect 3467 14365 3479 14368
rect 3421 14359 3479 14365
rect 3252 14328 3280 14359
rect 4154 14356 4160 14368
rect 4212 14356 4218 14408
rect 4709 14399 4767 14405
rect 4709 14365 4721 14399
rect 4755 14396 4767 14399
rect 5810 14396 5816 14408
rect 4755 14368 5816 14396
rect 4755 14365 4767 14368
rect 4709 14359 4767 14365
rect 5810 14356 5816 14368
rect 5868 14356 5874 14408
rect 5994 14396 6000 14408
rect 5955 14368 6000 14396
rect 5994 14356 6000 14368
rect 6052 14356 6058 14408
rect 6178 14396 6184 14408
rect 6139 14368 6184 14396
rect 6178 14356 6184 14368
rect 6236 14356 6242 14408
rect 7190 14396 7196 14408
rect 7151 14368 7196 14396
rect 7190 14356 7196 14368
rect 7248 14356 7254 14408
rect 7377 14399 7435 14405
rect 7377 14365 7389 14399
rect 7423 14396 7435 14399
rect 7466 14396 7472 14408
rect 7423 14368 7472 14396
rect 7423 14365 7435 14368
rect 7377 14359 7435 14365
rect 7466 14356 7472 14368
rect 7524 14356 7530 14408
rect 9950 14396 9956 14408
rect 9911 14368 9956 14396
rect 9950 14356 9956 14368
rect 10008 14356 10014 14408
rect 10870 14396 10876 14408
rect 10831 14368 10876 14396
rect 10870 14356 10876 14368
rect 10928 14356 10934 14408
rect 10962 14356 10968 14408
rect 11020 14356 11026 14408
rect 11609 14399 11667 14405
rect 11609 14365 11621 14399
rect 11655 14365 11667 14399
rect 11609 14359 11667 14365
rect 5902 14328 5908 14340
rect 3252 14300 5908 14328
rect 5902 14288 5908 14300
rect 5960 14288 5966 14340
rect 8938 14328 8944 14340
rect 8851 14300 8944 14328
rect 8938 14288 8944 14300
rect 8996 14328 9002 14340
rect 9398 14328 9404 14340
rect 8996 14300 9404 14328
rect 8996 14288 9002 14300
rect 9398 14288 9404 14300
rect 9456 14288 9462 14340
rect 10594 14288 10600 14340
rect 10652 14328 10658 14340
rect 11624 14328 11652 14359
rect 11992 14337 12020 14504
rect 12452 14504 13676 14532
rect 13900 14535 13958 14541
rect 12452 14473 12480 14504
rect 13900 14501 13912 14535
rect 13946 14532 13958 14535
rect 15378 14532 15384 14544
rect 13946 14504 15384 14532
rect 13946 14501 13958 14504
rect 13900 14495 13958 14501
rect 15378 14492 15384 14504
rect 15436 14492 15442 14544
rect 15556 14535 15614 14541
rect 15556 14501 15568 14535
rect 15602 14532 15614 14535
rect 16022 14532 16028 14544
rect 15602 14504 16028 14532
rect 15602 14501 15614 14504
rect 15556 14495 15614 14501
rect 16022 14492 16028 14504
rect 16080 14492 16086 14544
rect 19426 14532 19432 14544
rect 19387 14504 19432 14532
rect 19426 14492 19432 14504
rect 19484 14532 19490 14544
rect 19628 14532 19656 14572
rect 20441 14569 20453 14572
rect 20487 14569 20499 14603
rect 21082 14600 21088 14612
rect 21043 14572 21088 14600
rect 20441 14563 20499 14569
rect 21082 14560 21088 14572
rect 21140 14560 21146 14612
rect 21450 14600 21456 14612
rect 21411 14572 21456 14600
rect 21450 14560 21456 14572
rect 21508 14560 21514 14612
rect 19484 14504 19656 14532
rect 20165 14535 20223 14541
rect 19484 14492 19490 14504
rect 20165 14501 20177 14535
rect 20211 14532 20223 14535
rect 20806 14532 20812 14544
rect 20211 14504 20812 14532
rect 20211 14501 20223 14504
rect 20165 14495 20223 14501
rect 20806 14492 20812 14504
rect 20864 14492 20870 14544
rect 21174 14492 21180 14544
rect 21232 14532 21238 14544
rect 21232 14504 21312 14532
rect 21232 14492 21238 14504
rect 12437 14467 12495 14473
rect 12437 14433 12449 14467
rect 12483 14433 12495 14467
rect 12437 14427 12495 14433
rect 12526 14424 12532 14476
rect 12584 14464 12590 14476
rect 12897 14467 12955 14473
rect 12897 14464 12909 14467
rect 12584 14436 12909 14464
rect 12584 14424 12590 14436
rect 12897 14433 12909 14436
rect 12943 14433 12955 14467
rect 12897 14427 12955 14433
rect 13633 14467 13691 14473
rect 13633 14433 13645 14467
rect 13679 14464 13691 14467
rect 13722 14464 13728 14476
rect 13679 14436 13728 14464
rect 13679 14433 13691 14436
rect 13633 14427 13691 14433
rect 13722 14424 13728 14436
rect 13780 14424 13786 14476
rect 15289 14467 15347 14473
rect 15289 14433 15301 14467
rect 15335 14464 15347 14467
rect 15335 14436 16620 14464
rect 15335 14433 15347 14436
rect 15289 14427 15347 14433
rect 16592 14408 16620 14436
rect 16666 14424 16672 14476
rect 16724 14464 16730 14476
rect 17586 14464 17592 14476
rect 16724 14436 17592 14464
rect 16724 14424 16730 14436
rect 17586 14424 17592 14436
rect 17644 14424 17650 14476
rect 17764 14467 17822 14473
rect 17764 14433 17776 14467
rect 17810 14464 17822 14467
rect 18598 14464 18604 14476
rect 17810 14436 18604 14464
rect 17810 14433 17822 14436
rect 17764 14427 17822 14433
rect 18598 14424 18604 14436
rect 18656 14424 18662 14476
rect 19150 14424 19156 14476
rect 19208 14464 19214 14476
rect 19889 14467 19947 14473
rect 19889 14464 19901 14467
rect 19208 14436 19901 14464
rect 19208 14424 19214 14436
rect 19889 14433 19901 14436
rect 19935 14433 19947 14467
rect 19889 14427 19947 14433
rect 20901 14467 20959 14473
rect 20901 14433 20913 14467
rect 20947 14464 20959 14467
rect 21082 14464 21088 14476
rect 20947 14436 21088 14464
rect 20947 14433 20959 14436
rect 20901 14427 20959 14433
rect 21082 14424 21088 14436
rect 21140 14424 21146 14476
rect 21284 14473 21312 14504
rect 21269 14467 21327 14473
rect 21269 14433 21281 14467
rect 21315 14433 21327 14467
rect 21269 14427 21327 14433
rect 12986 14396 12992 14408
rect 12947 14368 12992 14396
rect 12986 14356 12992 14368
rect 13044 14356 13050 14408
rect 13078 14356 13084 14408
rect 13136 14396 13142 14408
rect 13136 14368 13181 14396
rect 13136 14356 13142 14368
rect 16574 14356 16580 14408
rect 16632 14396 16638 14408
rect 17310 14396 17316 14408
rect 16632 14368 17316 14396
rect 16632 14356 16638 14368
rect 17310 14356 17316 14368
rect 17368 14396 17374 14408
rect 17497 14399 17555 14405
rect 17497 14396 17509 14399
rect 17368 14368 17509 14396
rect 17368 14356 17374 14368
rect 17497 14365 17509 14368
rect 17543 14365 17555 14399
rect 18616 14396 18644 14424
rect 19521 14399 19579 14405
rect 18616 14368 19380 14396
rect 17497 14359 17555 14365
rect 10652 14300 11652 14328
rect 11977 14331 12035 14337
rect 10652 14288 10658 14300
rect 11977 14297 11989 14331
rect 12023 14328 12035 14331
rect 12618 14328 12624 14340
rect 12023 14300 12624 14328
rect 12023 14297 12035 14300
rect 11977 14291 12035 14297
rect 12618 14288 12624 14300
rect 12676 14288 12682 14340
rect 13004 14328 13032 14356
rect 13357 14331 13415 14337
rect 13357 14328 13369 14331
rect 13004 14300 13369 14328
rect 13357 14297 13369 14300
rect 13403 14297 13415 14331
rect 18874 14328 18880 14340
rect 18835 14300 18880 14328
rect 13357 14291 13415 14297
rect 18874 14288 18880 14300
rect 18932 14288 18938 14340
rect 19352 14328 19380 14368
rect 19521 14365 19533 14399
rect 19567 14365 19579 14399
rect 19521 14359 19579 14365
rect 19536 14328 19564 14359
rect 20346 14356 20352 14408
rect 20404 14396 20410 14408
rect 21284 14396 21312 14427
rect 20404 14368 21312 14396
rect 20404 14356 20410 14368
rect 19352 14300 19564 14328
rect 1535 14232 3004 14260
rect 1535 14229 1547 14232
rect 1489 14223 1547 14229
rect 3050 14220 3056 14272
rect 3108 14260 3114 14272
rect 3602 14260 3608 14272
rect 3108 14232 3608 14260
rect 3108 14220 3114 14232
rect 3602 14220 3608 14232
rect 3660 14220 3666 14272
rect 5166 14260 5172 14272
rect 5127 14232 5172 14260
rect 5166 14220 5172 14232
rect 5224 14220 5230 14272
rect 5534 14260 5540 14272
rect 5495 14232 5540 14260
rect 5534 14220 5540 14232
rect 5592 14220 5598 14272
rect 9125 14263 9183 14269
rect 9125 14229 9137 14263
rect 9171 14260 9183 14263
rect 9214 14260 9220 14272
rect 9171 14232 9220 14260
rect 9171 14229 9183 14232
rect 9125 14223 9183 14229
rect 9214 14220 9220 14232
rect 9272 14220 9278 14272
rect 10778 14220 10784 14272
rect 10836 14260 10842 14272
rect 12069 14263 12127 14269
rect 12069 14260 12081 14263
rect 10836 14232 12081 14260
rect 10836 14220 10842 14232
rect 12069 14229 12081 14232
rect 12115 14229 12127 14263
rect 12069 14223 12127 14229
rect 13814 14220 13820 14272
rect 13872 14260 13878 14272
rect 14366 14260 14372 14272
rect 13872 14232 14372 14260
rect 13872 14220 13878 14232
rect 14366 14220 14372 14232
rect 14424 14260 14430 14272
rect 15013 14263 15071 14269
rect 15013 14260 15025 14263
rect 14424 14232 15025 14260
rect 14424 14220 14430 14232
rect 15013 14229 15025 14232
rect 15059 14229 15071 14263
rect 15013 14223 15071 14229
rect 16390 14220 16396 14272
rect 16448 14260 16454 14272
rect 16669 14263 16727 14269
rect 16669 14260 16681 14263
rect 16448 14232 16681 14260
rect 16448 14220 16454 14232
rect 16669 14229 16681 14232
rect 16715 14229 16727 14263
rect 16669 14223 16727 14229
rect 16942 14220 16948 14272
rect 17000 14260 17006 14272
rect 17770 14260 17776 14272
rect 17000 14232 17776 14260
rect 17000 14220 17006 14232
rect 17770 14220 17776 14232
rect 17828 14220 17834 14272
rect 18966 14260 18972 14272
rect 18927 14232 18972 14260
rect 18966 14220 18972 14232
rect 19024 14220 19030 14272
rect 20717 14263 20775 14269
rect 20717 14229 20729 14263
rect 20763 14260 20775 14263
rect 21082 14260 21088 14272
rect 20763 14232 21088 14260
rect 20763 14229 20775 14232
rect 20717 14223 20775 14229
rect 21082 14220 21088 14232
rect 21140 14260 21146 14272
rect 21450 14260 21456 14272
rect 21140 14232 21456 14260
rect 21140 14220 21146 14232
rect 21450 14220 21456 14232
rect 21508 14220 21514 14272
rect 1104 14170 21896 14192
rect 1104 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 4575 14170
rect 4627 14118 4639 14170
rect 4691 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 18308 14170
rect 18360 14118 18372 14170
rect 18424 14118 18436 14170
rect 18488 14118 18500 14170
rect 18552 14118 21896 14170
rect 1104 14096 21896 14118
rect 1762 14056 1768 14068
rect 1723 14028 1768 14056
rect 1762 14016 1768 14028
rect 1820 14016 1826 14068
rect 5626 14056 5632 14068
rect 1964 14028 5632 14056
rect 1489 13855 1547 13861
rect 1489 13821 1501 13855
rect 1535 13852 1547 13855
rect 1578 13852 1584 13864
rect 1535 13824 1584 13852
rect 1535 13821 1547 13824
rect 1489 13815 1547 13821
rect 1578 13812 1584 13824
rect 1636 13812 1642 13864
rect 1964 13861 1992 14028
rect 5626 14016 5632 14028
rect 5684 14016 5690 14068
rect 5810 14056 5816 14068
rect 5771 14028 5816 14056
rect 5810 14016 5816 14028
rect 5868 14056 5874 14068
rect 7006 14056 7012 14068
rect 5868 14028 7012 14056
rect 5868 14016 5874 14028
rect 7006 14016 7012 14028
rect 7064 14016 7070 14068
rect 7098 14016 7104 14068
rect 7156 14056 7162 14068
rect 7653 14059 7711 14065
rect 7653 14056 7665 14059
rect 7156 14028 7665 14056
rect 7156 14016 7162 14028
rect 7653 14025 7665 14028
rect 7699 14025 7711 14059
rect 8938 14056 8944 14068
rect 7653 14019 7711 14025
rect 8772 14028 8944 14056
rect 2590 13988 2596 14000
rect 2240 13960 2596 13988
rect 2240 13929 2268 13960
rect 2590 13948 2596 13960
rect 2648 13948 2654 14000
rect 3973 13991 4031 13997
rect 3973 13957 3985 13991
rect 4019 13957 4031 13991
rect 3973 13951 4031 13957
rect 2225 13923 2283 13929
rect 2225 13889 2237 13923
rect 2271 13889 2283 13923
rect 3988 13920 4016 13951
rect 5902 13948 5908 14000
rect 5960 13988 5966 14000
rect 8772 13988 8800 14028
rect 8938 14016 8944 14028
rect 8996 14016 9002 14068
rect 9677 14059 9735 14065
rect 9677 14025 9689 14059
rect 9723 14056 9735 14059
rect 10962 14056 10968 14068
rect 9723 14028 10968 14056
rect 9723 14025 9735 14028
rect 9677 14019 9735 14025
rect 10962 14016 10968 14028
rect 11020 14016 11026 14068
rect 12713 14059 12771 14065
rect 12713 14025 12725 14059
rect 12759 14056 12771 14059
rect 13170 14056 13176 14068
rect 12759 14028 13176 14056
rect 12759 14025 12771 14028
rect 12713 14019 12771 14025
rect 13170 14016 13176 14028
rect 13228 14016 13234 14068
rect 13814 14056 13820 14068
rect 13372 14028 13820 14056
rect 5960 13960 8800 13988
rect 8849 13991 8907 13997
rect 5960 13948 5966 13960
rect 8849 13957 8861 13991
rect 8895 13988 8907 13991
rect 10502 13988 10508 14000
rect 8895 13960 9904 13988
rect 8895 13957 8907 13960
rect 8849 13951 8907 13957
rect 9876 13932 9904 13960
rect 9968 13960 10364 13988
rect 10463 13960 10508 13988
rect 3988 13892 4568 13920
rect 2225 13883 2283 13889
rect 4540 13864 4568 13892
rect 6178 13880 6184 13932
rect 6236 13920 6242 13932
rect 6457 13923 6515 13929
rect 6457 13920 6469 13923
rect 6236 13892 6469 13920
rect 6236 13880 6242 13892
rect 6457 13889 6469 13892
rect 6503 13889 6515 13923
rect 7374 13920 7380 13932
rect 7335 13892 7380 13920
rect 6457 13883 6515 13889
rect 7374 13880 7380 13892
rect 7432 13880 7438 13932
rect 7466 13880 7472 13932
rect 7524 13920 7530 13932
rect 8205 13923 8263 13929
rect 8205 13920 8217 13923
rect 7524 13892 8217 13920
rect 7524 13880 7530 13892
rect 8205 13889 8217 13892
rect 8251 13889 8263 13923
rect 9030 13920 9036 13932
rect 8205 13883 8263 13889
rect 8680 13892 9036 13920
rect 1949 13855 2007 13861
rect 1949 13821 1961 13855
rect 1995 13821 2007 13855
rect 2590 13852 2596 13864
rect 2503 13824 2596 13852
rect 1949 13815 2007 13821
rect 2590 13812 2596 13824
rect 2648 13852 2654 13864
rect 3970 13852 3976 13864
rect 2648 13824 3976 13852
rect 2648 13812 2654 13824
rect 3970 13812 3976 13824
rect 4028 13852 4034 13864
rect 4433 13855 4491 13861
rect 4433 13852 4445 13855
rect 4028 13824 4445 13852
rect 4028 13812 4034 13824
rect 4433 13821 4445 13824
rect 4479 13821 4491 13855
rect 4433 13815 4491 13821
rect 4522 13812 4528 13864
rect 4580 13852 4586 13864
rect 6196 13852 6224 13880
rect 4580 13824 6224 13852
rect 4580 13812 4586 13824
rect 6546 13812 6552 13864
rect 6604 13852 6610 13864
rect 7098 13852 7104 13864
rect 6604 13824 7104 13852
rect 6604 13812 6610 13824
rect 7098 13812 7104 13824
rect 7156 13852 7162 13864
rect 7285 13855 7343 13861
rect 7285 13852 7297 13855
rect 7156 13824 7297 13852
rect 7156 13812 7162 13824
rect 7285 13821 7297 13824
rect 7331 13821 7343 13855
rect 8110 13852 8116 13864
rect 8071 13824 8116 13852
rect 7285 13815 7343 13821
rect 8110 13812 8116 13824
rect 8168 13812 8174 13864
rect 2860 13787 2918 13793
rect 2860 13753 2872 13787
rect 2906 13784 2918 13787
rect 3234 13784 3240 13796
rect 2906 13756 3240 13784
rect 2906 13753 2918 13756
rect 2860 13747 2918 13753
rect 3234 13744 3240 13756
rect 3292 13744 3298 13796
rect 4154 13744 4160 13796
rect 4212 13784 4218 13796
rect 4678 13787 4736 13793
rect 4678 13784 4690 13787
rect 4212 13756 4690 13784
rect 4212 13744 4218 13756
rect 4678 13753 4690 13756
rect 4724 13753 4736 13787
rect 7193 13787 7251 13793
rect 4678 13747 4736 13753
rect 5828 13756 7144 13784
rect 3252 13716 3280 13744
rect 5828 13728 5856 13756
rect 5810 13716 5816 13728
rect 3252 13688 5816 13716
rect 5810 13676 5816 13688
rect 5868 13676 5874 13728
rect 5902 13676 5908 13728
rect 5960 13716 5966 13728
rect 5960 13688 6005 13716
rect 5960 13676 5966 13688
rect 6086 13676 6092 13728
rect 6144 13716 6150 13728
rect 6273 13719 6331 13725
rect 6273 13716 6285 13719
rect 6144 13688 6285 13716
rect 6144 13676 6150 13688
rect 6273 13685 6285 13688
rect 6319 13685 6331 13719
rect 6273 13679 6331 13685
rect 6365 13719 6423 13725
rect 6365 13685 6377 13719
rect 6411 13716 6423 13719
rect 6825 13719 6883 13725
rect 6825 13716 6837 13719
rect 6411 13688 6837 13716
rect 6411 13685 6423 13688
rect 6365 13679 6423 13685
rect 6825 13685 6837 13688
rect 6871 13685 6883 13719
rect 7116 13716 7144 13756
rect 7193 13753 7205 13787
rect 7239 13784 7251 13787
rect 8680 13784 8708 13892
rect 9030 13880 9036 13892
rect 9088 13880 9094 13932
rect 9398 13880 9404 13932
rect 9456 13920 9462 13932
rect 9493 13923 9551 13929
rect 9493 13920 9505 13923
rect 9456 13892 9505 13920
rect 9456 13880 9462 13892
rect 9493 13889 9505 13892
rect 9539 13889 9551 13923
rect 9493 13883 9551 13889
rect 8757 13855 8815 13861
rect 8757 13821 8769 13855
rect 8803 13852 8815 13855
rect 8846 13852 8852 13864
rect 8803 13824 8852 13852
rect 8803 13821 8815 13824
rect 8757 13815 8815 13821
rect 8846 13812 8852 13824
rect 8904 13812 8910 13864
rect 9214 13812 9220 13864
rect 9272 13852 9278 13864
rect 9309 13855 9367 13861
rect 9309 13852 9321 13855
rect 9272 13824 9321 13852
rect 9272 13812 9278 13824
rect 9309 13821 9321 13824
rect 9355 13821 9367 13855
rect 9508 13852 9536 13883
rect 9858 13880 9864 13932
rect 9916 13880 9922 13932
rect 9968 13852 9996 13960
rect 10134 13920 10140 13932
rect 10095 13892 10140 13920
rect 10134 13880 10140 13892
rect 10192 13880 10198 13932
rect 10336 13929 10364 13960
rect 10502 13948 10508 13960
rect 10560 13948 10566 14000
rect 11425 13991 11483 13997
rect 11425 13988 11437 13991
rect 11348 13960 11437 13988
rect 10321 13923 10379 13929
rect 10321 13889 10333 13923
rect 10367 13920 10379 13923
rect 11057 13923 11115 13929
rect 11057 13920 11069 13923
rect 10367 13892 11069 13920
rect 10367 13889 10379 13892
rect 10321 13883 10379 13889
rect 11057 13889 11069 13892
rect 11103 13889 11115 13923
rect 11057 13883 11115 13889
rect 9508 13824 9996 13852
rect 9309 13815 9367 13821
rect 10042 13812 10048 13864
rect 10100 13852 10106 13864
rect 10873 13855 10931 13861
rect 10873 13852 10885 13855
rect 10100 13824 10885 13852
rect 10100 13812 10106 13824
rect 10873 13821 10885 13824
rect 10919 13821 10931 13855
rect 10873 13815 10931 13821
rect 10965 13855 11023 13861
rect 10965 13821 10977 13855
rect 11011 13852 11023 13855
rect 11348 13852 11376 13960
rect 11425 13957 11437 13960
rect 11471 13988 11483 13991
rect 12250 13988 12256 14000
rect 11471 13960 12256 13988
rect 11471 13957 11483 13960
rect 11425 13951 11483 13957
rect 12250 13948 12256 13960
rect 12308 13948 12314 14000
rect 13372 13929 13400 14028
rect 13814 14016 13820 14028
rect 13872 14016 13878 14068
rect 15286 14016 15292 14068
rect 15344 14056 15350 14068
rect 15841 14059 15899 14065
rect 15841 14056 15853 14059
rect 15344 14028 15853 14056
rect 15344 14016 15350 14028
rect 15841 14025 15853 14028
rect 15887 14025 15899 14059
rect 17129 14059 17187 14065
rect 17129 14056 17141 14059
rect 15841 14019 15899 14025
rect 15948 14028 17141 14056
rect 14734 13948 14740 14000
rect 14792 13988 14798 14000
rect 14921 13991 14979 13997
rect 14921 13988 14933 13991
rect 14792 13960 14933 13988
rect 14792 13948 14798 13960
rect 14921 13957 14933 13960
rect 14967 13988 14979 13991
rect 15378 13988 15384 14000
rect 14967 13960 15384 13988
rect 14967 13957 14979 13960
rect 14921 13951 14979 13957
rect 15378 13948 15384 13960
rect 15436 13948 15442 14000
rect 15746 13948 15752 14000
rect 15804 13988 15810 14000
rect 15948 13988 15976 14028
rect 17129 14025 17141 14028
rect 17175 14025 17187 14059
rect 17586 14056 17592 14068
rect 17547 14028 17592 14056
rect 17129 14019 17187 14025
rect 17586 14016 17592 14028
rect 17644 14016 17650 14068
rect 17954 14016 17960 14068
rect 18012 14056 18018 14068
rect 18049 14059 18107 14065
rect 18049 14056 18061 14059
rect 18012 14028 18061 14056
rect 18012 14016 18018 14028
rect 18049 14025 18061 14028
rect 18095 14025 18107 14059
rect 18049 14019 18107 14025
rect 18138 14016 18144 14068
rect 18196 14056 18202 14068
rect 18877 14059 18935 14065
rect 18877 14056 18889 14059
rect 18196 14028 18889 14056
rect 18196 14016 18202 14028
rect 18877 14025 18889 14028
rect 18923 14025 18935 14059
rect 18877 14019 18935 14025
rect 19058 14016 19064 14068
rect 19116 14056 19122 14068
rect 20990 14056 20996 14068
rect 19116 14028 20852 14056
rect 20951 14028 20996 14056
rect 19116 14016 19122 14028
rect 19334 13988 19340 14000
rect 15804 13960 15976 13988
rect 16960 13960 19340 13988
rect 15804 13948 15810 13960
rect 13357 13923 13415 13929
rect 13357 13889 13369 13923
rect 13403 13889 13415 13923
rect 13357 13883 13415 13889
rect 15286 13880 15292 13932
rect 15344 13920 15350 13932
rect 15565 13923 15623 13929
rect 15565 13920 15577 13923
rect 15344 13892 15577 13920
rect 15344 13880 15350 13892
rect 15565 13889 15577 13892
rect 15611 13920 15623 13923
rect 16390 13920 16396 13932
rect 15611 13892 16396 13920
rect 15611 13889 15623 13892
rect 15565 13883 15623 13889
rect 16390 13880 16396 13892
rect 16448 13880 16454 13932
rect 11011 13824 11376 13852
rect 11011 13821 11023 13824
rect 10965 13815 11023 13821
rect 11072 13796 11100 13824
rect 11790 13812 11796 13864
rect 11848 13852 11854 13864
rect 13541 13855 13599 13861
rect 13541 13852 13553 13855
rect 11848 13824 13553 13852
rect 11848 13812 11854 13824
rect 13541 13821 13553 13824
rect 13587 13821 13599 13855
rect 14090 13852 14096 13864
rect 13541 13815 13599 13821
rect 13740 13824 14096 13852
rect 7239 13756 8708 13784
rect 7239 13753 7251 13756
rect 7193 13747 7251 13753
rect 8938 13744 8944 13796
rect 8996 13784 9002 13796
rect 10318 13784 10324 13796
rect 8996 13756 10324 13784
rect 8996 13744 9002 13756
rect 10318 13744 10324 13756
rect 10376 13744 10382 13796
rect 11054 13744 11060 13796
rect 11112 13744 11118 13796
rect 11606 13784 11612 13796
rect 11567 13756 11612 13784
rect 11606 13744 11612 13756
rect 11664 13744 11670 13796
rect 11882 13744 11888 13796
rect 11940 13784 11946 13796
rect 12250 13784 12256 13796
rect 11940 13756 12256 13784
rect 11940 13744 11946 13756
rect 12250 13744 12256 13756
rect 12308 13744 12314 13796
rect 13081 13787 13139 13793
rect 13081 13753 13093 13787
rect 13127 13784 13139 13787
rect 13740 13784 13768 13824
rect 14090 13812 14096 13824
rect 14148 13812 14154 13864
rect 15470 13812 15476 13864
rect 15528 13852 15534 13864
rect 15838 13852 15844 13864
rect 15528 13824 15844 13852
rect 15528 13812 15534 13824
rect 15838 13812 15844 13824
rect 15896 13812 15902 13864
rect 15930 13812 15936 13864
rect 15988 13852 15994 13864
rect 16960 13861 16988 13960
rect 19334 13948 19340 13960
rect 19392 13948 19398 14000
rect 20824 13988 20852 14028
rect 20990 14016 20996 14028
rect 21048 14016 21054 14068
rect 21361 13991 21419 13997
rect 21361 13988 21373 13991
rect 20824 13960 21373 13988
rect 18598 13920 18604 13932
rect 18559 13892 18604 13920
rect 18598 13880 18604 13892
rect 18656 13880 18662 13932
rect 18874 13880 18880 13932
rect 18932 13920 18938 13932
rect 19429 13923 19487 13929
rect 19429 13920 19441 13923
rect 18932 13892 19441 13920
rect 18932 13880 18938 13892
rect 19429 13889 19441 13892
rect 19475 13889 19487 13923
rect 19429 13883 19487 13889
rect 16209 13855 16267 13861
rect 16209 13852 16221 13855
rect 15988 13824 16221 13852
rect 15988 13812 15994 13824
rect 16209 13821 16221 13824
rect 16255 13852 16267 13855
rect 16945 13855 17003 13861
rect 16945 13852 16957 13855
rect 16255 13824 16957 13852
rect 16255 13821 16267 13824
rect 16209 13815 16267 13821
rect 16945 13821 16957 13824
rect 16991 13821 17003 13855
rect 18417 13855 18475 13861
rect 18417 13852 18429 13855
rect 16945 13815 17003 13821
rect 17788 13824 18429 13852
rect 13127 13756 13768 13784
rect 13808 13787 13866 13793
rect 13127 13753 13139 13756
rect 13081 13747 13139 13753
rect 13808 13753 13820 13787
rect 13854 13784 13866 13787
rect 13906 13784 13912 13796
rect 13854 13756 13912 13784
rect 13854 13753 13866 13756
rect 13808 13747 13866 13753
rect 13906 13744 13912 13756
rect 13964 13744 13970 13796
rect 17788 13793 17816 13824
rect 18417 13821 18429 13824
rect 18463 13852 18475 13855
rect 18690 13852 18696 13864
rect 18463 13824 18696 13852
rect 18463 13821 18475 13824
rect 18417 13815 18475 13821
rect 18690 13812 18696 13824
rect 18748 13812 18754 13864
rect 18966 13812 18972 13864
rect 19024 13852 19030 13864
rect 19245 13855 19303 13861
rect 19245 13852 19257 13855
rect 19024 13824 19257 13852
rect 19024 13812 19030 13824
rect 19245 13821 19257 13824
rect 19291 13821 19303 13855
rect 19245 13815 19303 13821
rect 20257 13855 20315 13861
rect 20257 13821 20269 13855
rect 20303 13852 20315 13855
rect 20530 13852 20536 13864
rect 20303 13824 20392 13852
rect 20491 13824 20536 13852
rect 20303 13821 20315 13824
rect 20257 13815 20315 13821
rect 17773 13787 17831 13793
rect 17773 13784 17785 13787
rect 14016 13756 17785 13784
rect 7374 13716 7380 13728
rect 7116 13688 7380 13716
rect 6825 13679 6883 13685
rect 7374 13676 7380 13688
rect 7432 13676 7438 13728
rect 8021 13719 8079 13725
rect 8021 13685 8033 13719
rect 8067 13716 8079 13719
rect 8573 13719 8631 13725
rect 8573 13716 8585 13719
rect 8067 13688 8585 13716
rect 8067 13685 8079 13688
rect 8021 13679 8079 13685
rect 8573 13685 8585 13688
rect 8619 13716 8631 13719
rect 8754 13716 8760 13728
rect 8619 13688 8760 13716
rect 8619 13685 8631 13688
rect 8573 13679 8631 13685
rect 8754 13676 8760 13688
rect 8812 13676 8818 13728
rect 8846 13676 8852 13728
rect 8904 13716 8910 13728
rect 9217 13719 9275 13725
rect 9217 13716 9229 13719
rect 8904 13688 9229 13716
rect 8904 13676 8910 13688
rect 9217 13685 9229 13688
rect 9263 13685 9275 13719
rect 9217 13679 9275 13685
rect 10045 13719 10103 13725
rect 10045 13685 10057 13719
rect 10091 13716 10103 13719
rect 11624 13716 11652 13744
rect 12434 13716 12440 13728
rect 10091 13688 11652 13716
rect 12395 13688 12440 13716
rect 10091 13685 10103 13688
rect 10045 13679 10103 13685
rect 12434 13676 12440 13688
rect 12492 13676 12498 13728
rect 13170 13676 13176 13728
rect 13228 13716 13234 13728
rect 13228 13688 13273 13716
rect 13228 13676 13234 13688
rect 13722 13676 13728 13728
rect 13780 13716 13786 13728
rect 14016 13716 14044 13756
rect 17773 13753 17785 13756
rect 17819 13753 17831 13787
rect 17773 13747 17831 13753
rect 17954 13744 17960 13796
rect 18012 13784 18018 13796
rect 19337 13787 19395 13793
rect 19337 13784 19349 13787
rect 18012 13756 19349 13784
rect 18012 13744 18018 13756
rect 19337 13753 19349 13756
rect 19383 13753 19395 13787
rect 20364 13784 20392 13824
rect 20530 13812 20536 13824
rect 20588 13812 20594 13864
rect 20824 13861 20852 13960
rect 21361 13957 21373 13960
rect 21407 13957 21419 13991
rect 21361 13951 21419 13957
rect 20809 13855 20867 13861
rect 20809 13821 20821 13855
rect 20855 13821 20867 13855
rect 21266 13852 21272 13864
rect 20809 13815 20867 13821
rect 20916 13824 21272 13852
rect 20916 13784 20944 13824
rect 21266 13812 21272 13824
rect 21324 13812 21330 13864
rect 20364 13756 20944 13784
rect 19337 13747 19395 13753
rect 13780 13688 14044 13716
rect 13780 13676 13786 13688
rect 14090 13676 14096 13728
rect 14148 13716 14154 13728
rect 15013 13719 15071 13725
rect 15013 13716 15025 13719
rect 14148 13688 15025 13716
rect 14148 13676 14154 13688
rect 15013 13685 15025 13688
rect 15059 13685 15071 13719
rect 15378 13716 15384 13728
rect 15339 13688 15384 13716
rect 15013 13679 15071 13685
rect 15378 13676 15384 13688
rect 15436 13676 15442 13728
rect 15470 13676 15476 13728
rect 15528 13716 15534 13728
rect 15528 13688 15573 13716
rect 15528 13676 15534 13688
rect 15746 13676 15752 13728
rect 15804 13716 15810 13728
rect 16301 13719 16359 13725
rect 16301 13716 16313 13719
rect 15804 13688 16313 13716
rect 15804 13676 15810 13688
rect 16301 13685 16313 13688
rect 16347 13685 16359 13719
rect 16301 13679 16359 13685
rect 16482 13676 16488 13728
rect 16540 13716 16546 13728
rect 16669 13719 16727 13725
rect 16669 13716 16681 13719
rect 16540 13688 16681 13716
rect 16540 13676 16546 13688
rect 16669 13685 16681 13688
rect 16715 13685 16727 13719
rect 16669 13679 16727 13685
rect 17586 13676 17592 13728
rect 17644 13716 17650 13728
rect 18509 13719 18567 13725
rect 18509 13716 18521 13719
rect 17644 13688 18521 13716
rect 17644 13676 17650 13688
rect 18509 13685 18521 13688
rect 18555 13685 18567 13719
rect 18509 13679 18567 13685
rect 1104 13626 21896 13648
rect 1104 13574 7912 13626
rect 7964 13574 7976 13626
rect 8028 13574 8040 13626
rect 8092 13574 8104 13626
rect 8156 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 15035 13626
rect 15087 13574 21896 13626
rect 1104 13552 21896 13574
rect 2406 13512 2412 13524
rect 2367 13484 2412 13512
rect 2406 13472 2412 13484
rect 2464 13472 2470 13524
rect 2774 13472 2780 13524
rect 2832 13512 2838 13524
rect 3145 13515 3203 13521
rect 2832 13484 2877 13512
rect 2832 13472 2838 13484
rect 3145 13481 3157 13515
rect 3191 13512 3203 13515
rect 3786 13512 3792 13524
rect 3191 13484 3792 13512
rect 3191 13481 3203 13484
rect 3145 13475 3203 13481
rect 3786 13472 3792 13484
rect 3844 13472 3850 13524
rect 4154 13472 4160 13524
rect 4212 13512 4218 13524
rect 5350 13512 5356 13524
rect 4212 13484 5356 13512
rect 4212 13472 4218 13484
rect 5350 13472 5356 13484
rect 5408 13512 5414 13524
rect 5445 13515 5503 13521
rect 5445 13512 5457 13515
rect 5408 13484 5457 13512
rect 5408 13472 5414 13484
rect 5445 13481 5457 13484
rect 5491 13481 5503 13515
rect 6086 13512 6092 13524
rect 6047 13484 6092 13512
rect 5445 13475 5503 13481
rect 6086 13472 6092 13484
rect 6144 13472 6150 13524
rect 6178 13472 6184 13524
rect 6236 13512 6242 13524
rect 6457 13515 6515 13521
rect 6457 13512 6469 13515
rect 6236 13484 6469 13512
rect 6236 13472 6242 13484
rect 6457 13481 6469 13484
rect 6503 13512 6515 13515
rect 6546 13512 6552 13524
rect 6503 13484 6552 13512
rect 6503 13481 6515 13484
rect 6457 13475 6515 13481
rect 6546 13472 6552 13484
rect 6604 13472 6610 13524
rect 7006 13472 7012 13524
rect 7064 13512 7070 13524
rect 7064 13484 7205 13512
rect 7064 13472 7070 13484
rect 4522 13404 4528 13456
rect 4580 13404 4586 13456
rect 5810 13404 5816 13456
rect 5868 13444 5874 13456
rect 7177 13453 7205 13484
rect 8294 13472 8300 13524
rect 8352 13512 8358 13524
rect 8389 13515 8447 13521
rect 8389 13512 8401 13515
rect 8352 13484 8401 13512
rect 8352 13472 8358 13484
rect 8389 13481 8401 13484
rect 8435 13481 8447 13515
rect 9490 13512 9496 13524
rect 9451 13484 9496 13512
rect 8389 13475 8447 13481
rect 9490 13472 9496 13484
rect 9548 13472 9554 13524
rect 9674 13512 9680 13524
rect 9635 13484 9680 13512
rect 9674 13472 9680 13484
rect 9732 13472 9738 13524
rect 10045 13515 10103 13521
rect 10045 13481 10057 13515
rect 10091 13512 10103 13515
rect 10502 13512 10508 13524
rect 10091 13484 10508 13512
rect 10091 13481 10103 13484
rect 10045 13475 10103 13481
rect 10502 13472 10508 13484
rect 10560 13472 10566 13524
rect 13170 13472 13176 13524
rect 13228 13512 13234 13524
rect 13541 13515 13599 13521
rect 13541 13512 13553 13515
rect 13228 13484 13553 13512
rect 13228 13472 13234 13484
rect 13541 13481 13553 13484
rect 13587 13481 13599 13515
rect 13541 13475 13599 13481
rect 13909 13515 13967 13521
rect 13909 13481 13921 13515
rect 13955 13512 13967 13515
rect 14369 13515 14427 13521
rect 14369 13512 14381 13515
rect 13955 13484 14381 13512
rect 13955 13481 13967 13484
rect 13909 13475 13967 13481
rect 14369 13481 14381 13484
rect 14415 13481 14427 13515
rect 14369 13475 14427 13481
rect 14550 13472 14556 13524
rect 14608 13512 14614 13524
rect 14737 13515 14795 13521
rect 14737 13512 14749 13515
rect 14608 13484 14749 13512
rect 14608 13472 14614 13484
rect 14737 13481 14749 13484
rect 14783 13481 14795 13515
rect 14737 13475 14795 13481
rect 15289 13515 15347 13521
rect 15289 13481 15301 13515
rect 15335 13512 15347 13515
rect 15470 13512 15476 13524
rect 15335 13484 15476 13512
rect 15335 13481 15347 13484
rect 15289 13475 15347 13481
rect 15470 13472 15476 13484
rect 15528 13472 15534 13524
rect 16114 13512 16120 13524
rect 16075 13484 16120 13512
rect 16114 13472 16120 13484
rect 16172 13472 16178 13524
rect 16482 13512 16488 13524
rect 16443 13484 16488 13512
rect 16482 13472 16488 13484
rect 16540 13472 16546 13524
rect 17034 13512 17040 13524
rect 16995 13484 17040 13512
rect 17034 13472 17040 13484
rect 17092 13472 17098 13524
rect 17497 13515 17555 13521
rect 17497 13481 17509 13515
rect 17543 13512 17555 13515
rect 17865 13515 17923 13521
rect 17865 13512 17877 13515
rect 17543 13484 17877 13512
rect 17543 13481 17555 13484
rect 17497 13475 17555 13481
rect 17865 13481 17877 13484
rect 17911 13481 17923 13515
rect 21082 13512 21088 13524
rect 21043 13484 21088 13512
rect 17865 13475 17923 13481
rect 21082 13472 21088 13484
rect 21140 13472 21146 13524
rect 7162 13447 7220 13453
rect 5868 13416 6776 13444
rect 5868 13404 5874 13416
rect 1673 13379 1731 13385
rect 1673 13345 1685 13379
rect 1719 13376 1731 13379
rect 1762 13376 1768 13388
rect 1719 13348 1768 13376
rect 1719 13345 1731 13348
rect 1673 13339 1731 13345
rect 1762 13336 1768 13348
rect 1820 13336 1826 13388
rect 2225 13379 2283 13385
rect 2225 13345 2237 13379
rect 2271 13345 2283 13379
rect 2225 13339 2283 13345
rect 1486 13268 1492 13320
rect 1544 13308 1550 13320
rect 1857 13311 1915 13317
rect 1857 13308 1869 13311
rect 1544 13280 1869 13308
rect 1544 13268 1550 13280
rect 1857 13277 1869 13280
rect 1903 13277 1915 13311
rect 2240 13308 2268 13339
rect 2314 13336 2320 13388
rect 2372 13376 2378 13388
rect 2593 13379 2651 13385
rect 2593 13376 2605 13379
rect 2372 13348 2605 13376
rect 2372 13336 2378 13348
rect 2593 13345 2605 13348
rect 2639 13345 2651 13379
rect 2593 13339 2651 13345
rect 3513 13379 3571 13385
rect 3513 13345 3525 13379
rect 3559 13376 3571 13379
rect 3786 13376 3792 13388
rect 3559 13348 3792 13376
rect 3559 13345 3571 13348
rect 3513 13339 3571 13345
rect 3786 13336 3792 13348
rect 3844 13336 3850 13388
rect 4154 13376 4160 13388
rect 3896 13348 4160 13376
rect 3605 13311 3663 13317
rect 2240 13280 3096 13308
rect 1857 13271 1915 13277
rect 3068 13252 3096 13280
rect 3605 13277 3617 13311
rect 3651 13277 3663 13311
rect 3605 13271 3663 13277
rect 3697 13311 3755 13317
rect 3697 13277 3709 13311
rect 3743 13308 3755 13311
rect 3896 13308 3924 13348
rect 4154 13336 4160 13348
rect 4212 13336 4218 13388
rect 4338 13385 4344 13388
rect 4332 13376 4344 13385
rect 4251 13348 4344 13376
rect 4332 13339 4344 13348
rect 4396 13376 4402 13388
rect 4540 13376 4568 13404
rect 4396 13348 4568 13376
rect 5721 13379 5779 13385
rect 4338 13336 4344 13339
rect 4396 13336 4402 13348
rect 5721 13345 5733 13379
rect 5767 13345 5779 13379
rect 5721 13339 5779 13345
rect 5997 13379 6055 13385
rect 5997 13345 6009 13379
rect 6043 13376 6055 13379
rect 6178 13376 6184 13388
rect 6043 13348 6184 13376
rect 6043 13345 6055 13348
rect 5997 13339 6055 13345
rect 3743 13280 3924 13308
rect 3743 13277 3755 13280
rect 3697 13271 3755 13277
rect 3050 13240 3056 13252
rect 3011 13212 3056 13240
rect 3050 13200 3056 13212
rect 3108 13200 3114 13252
rect 3620 13172 3648 13271
rect 3970 13268 3976 13320
rect 4028 13308 4034 13320
rect 4065 13311 4123 13317
rect 4065 13308 4077 13311
rect 4028 13280 4077 13308
rect 4028 13268 4034 13280
rect 4065 13277 4077 13280
rect 4111 13277 4123 13311
rect 5736 13308 5764 13339
rect 6178 13336 6184 13348
rect 6236 13336 6242 13388
rect 5736 13280 6500 13308
rect 4065 13271 4123 13277
rect 4338 13172 4344 13184
rect 3620 13144 4344 13172
rect 4338 13132 4344 13144
rect 4396 13132 4402 13184
rect 5537 13175 5595 13181
rect 5537 13141 5549 13175
rect 5583 13172 5595 13175
rect 6178 13172 6184 13184
rect 5583 13144 6184 13172
rect 5583 13141 5595 13144
rect 5537 13135 5595 13141
rect 6178 13132 6184 13144
rect 6236 13132 6242 13184
rect 6472 13172 6500 13280
rect 6546 13268 6552 13320
rect 6604 13308 6610 13320
rect 6748 13317 6776 13416
rect 7162 13413 7174 13447
rect 7208 13413 7220 13447
rect 7162 13407 7220 13413
rect 7742 13404 7748 13456
rect 7800 13444 7806 13456
rect 8478 13444 8484 13456
rect 7800 13416 8484 13444
rect 7800 13404 7806 13416
rect 8478 13404 8484 13416
rect 8536 13444 8542 13456
rect 8536 13416 8984 13444
rect 8536 13404 8542 13416
rect 6917 13379 6975 13385
rect 6917 13345 6929 13379
rect 6963 13376 6975 13379
rect 8202 13376 8208 13388
rect 6963 13348 8208 13376
rect 6963 13345 6975 13348
rect 6917 13339 6975 13345
rect 8202 13336 8208 13348
rect 8260 13336 8266 13388
rect 8757 13379 8815 13385
rect 8757 13345 8769 13379
rect 8803 13345 8815 13379
rect 8757 13339 8815 13345
rect 6733 13311 6791 13317
rect 6604 13280 6649 13308
rect 6604 13268 6610 13280
rect 6733 13277 6745 13311
rect 6779 13277 6791 13311
rect 6733 13271 6791 13277
rect 7558 13172 7564 13184
rect 6472 13144 7564 13172
rect 7558 13132 7564 13144
rect 7616 13132 7622 13184
rect 8294 13132 8300 13184
rect 8352 13172 8358 13184
rect 8772 13172 8800 13339
rect 8956 13317 8984 13416
rect 9508 13376 9536 13472
rect 9858 13404 9864 13456
rect 9916 13444 9922 13456
rect 10137 13447 10195 13453
rect 10137 13444 10149 13447
rect 9916 13416 10149 13444
rect 9916 13404 9922 13416
rect 10137 13413 10149 13416
rect 10183 13413 10195 13447
rect 10137 13407 10195 13413
rect 10318 13404 10324 13456
rect 10376 13444 10382 13456
rect 10597 13447 10655 13453
rect 10597 13444 10609 13447
rect 10376 13416 10609 13444
rect 10376 13404 10382 13416
rect 10597 13413 10609 13416
rect 10643 13444 10655 13447
rect 11057 13447 11115 13453
rect 11057 13444 11069 13447
rect 10643 13416 11069 13444
rect 10643 13413 10655 13416
rect 10597 13407 10655 13413
rect 11057 13413 11069 13416
rect 11103 13413 11115 13447
rect 13722 13444 13728 13456
rect 11057 13407 11115 13413
rect 11164 13416 13728 13444
rect 11164 13385 11192 13416
rect 13722 13404 13728 13416
rect 13780 13404 13786 13456
rect 13998 13444 14004 13456
rect 13959 13416 14004 13444
rect 13998 13404 14004 13416
rect 14056 13404 14062 13456
rect 14090 13404 14096 13456
rect 14148 13444 14154 13456
rect 14274 13444 14280 13456
rect 14148 13416 14280 13444
rect 14148 13404 14154 13416
rect 14274 13404 14280 13416
rect 14332 13404 14338 13456
rect 14826 13444 14832 13456
rect 14568 13416 14832 13444
rect 11149 13379 11207 13385
rect 11149 13376 11161 13379
rect 9508 13348 11161 13376
rect 11149 13345 11161 13348
rect 11195 13345 11207 13379
rect 11149 13339 11207 13345
rect 11517 13379 11575 13385
rect 11517 13345 11529 13379
rect 11563 13376 11575 13379
rect 11606 13376 11612 13388
rect 11563 13348 11612 13376
rect 11563 13345 11575 13348
rect 11517 13339 11575 13345
rect 11606 13336 11612 13348
rect 11664 13336 11670 13388
rect 11790 13385 11796 13388
rect 11784 13376 11796 13385
rect 11751 13348 11796 13376
rect 11784 13339 11796 13348
rect 11790 13336 11796 13339
rect 11848 13336 11854 13388
rect 8849 13311 8907 13317
rect 8849 13277 8861 13311
rect 8895 13277 8907 13311
rect 8849 13271 8907 13277
rect 8941 13311 8999 13317
rect 8941 13277 8953 13311
rect 8987 13277 8999 13311
rect 8941 13271 8999 13277
rect 8864 13240 8892 13271
rect 9030 13268 9036 13320
rect 9088 13308 9094 13320
rect 10134 13308 10140 13320
rect 9088 13280 10140 13308
rect 9088 13268 9094 13280
rect 10134 13268 10140 13280
rect 10192 13268 10198 13320
rect 10321 13311 10379 13317
rect 10321 13277 10333 13311
rect 10367 13308 10379 13311
rect 10594 13308 10600 13320
rect 10367 13280 10600 13308
rect 10367 13277 10379 13280
rect 10321 13271 10379 13277
rect 10594 13268 10600 13280
rect 10652 13268 10658 13320
rect 11241 13311 11299 13317
rect 11241 13277 11253 13311
rect 11287 13277 11299 13311
rect 11241 13271 11299 13277
rect 14185 13311 14243 13317
rect 14185 13277 14197 13311
rect 14231 13308 14243 13311
rect 14568 13308 14596 13416
rect 14826 13404 14832 13416
rect 14884 13404 14890 13456
rect 15657 13447 15715 13453
rect 15657 13444 15669 13447
rect 14936 13416 15669 13444
rect 14642 13336 14648 13388
rect 14700 13376 14706 13388
rect 14936 13376 14964 13416
rect 15657 13413 15669 13416
rect 15703 13413 15715 13447
rect 15657 13407 15715 13413
rect 15930 13404 15936 13456
rect 15988 13444 15994 13456
rect 16577 13447 16635 13453
rect 16577 13444 16589 13447
rect 15988 13416 16589 13444
rect 15988 13404 15994 13416
rect 16577 13413 16589 13416
rect 16623 13413 16635 13447
rect 16577 13407 16635 13413
rect 17328 13416 20944 13444
rect 14700 13348 14964 13376
rect 14700 13336 14706 13348
rect 15102 13336 15108 13388
rect 15160 13376 15166 13388
rect 17328 13376 17356 13416
rect 15160 13348 17356 13376
rect 17405 13379 17463 13385
rect 15160 13336 15166 13348
rect 17405 13345 17417 13379
rect 17451 13376 17463 13379
rect 18046 13376 18052 13388
rect 17451 13348 18052 13376
rect 17451 13345 17463 13348
rect 17405 13339 17463 13345
rect 18046 13336 18052 13348
rect 18104 13336 18110 13388
rect 18233 13379 18291 13385
rect 18233 13345 18245 13379
rect 18279 13376 18291 13379
rect 18782 13376 18788 13388
rect 18279 13348 18788 13376
rect 18279 13345 18291 13348
rect 18233 13339 18291 13345
rect 18782 13336 18788 13348
rect 18840 13336 18846 13388
rect 20916 13385 20944 13416
rect 20901 13379 20959 13385
rect 20901 13345 20913 13379
rect 20947 13376 20959 13379
rect 21269 13379 21327 13385
rect 21269 13376 21281 13379
rect 20947 13348 21281 13376
rect 20947 13345 20959 13348
rect 20901 13339 20959 13345
rect 21269 13345 21281 13348
rect 21315 13345 21327 13379
rect 21269 13339 21327 13345
rect 14826 13308 14832 13320
rect 14231 13280 14596 13308
rect 14787 13280 14832 13308
rect 14231 13277 14243 13280
rect 14185 13271 14243 13277
rect 8864 13212 9352 13240
rect 9324 13184 9352 13212
rect 9858 13200 9864 13252
rect 9916 13240 9922 13252
rect 10410 13240 10416 13252
rect 9916 13212 10416 13240
rect 9916 13200 9922 13212
rect 10410 13200 10416 13212
rect 10468 13200 10474 13252
rect 10870 13200 10876 13252
rect 10928 13240 10934 13252
rect 11256 13240 11284 13271
rect 14826 13268 14832 13280
rect 14884 13268 14890 13320
rect 14918 13268 14924 13320
rect 14976 13308 14982 13320
rect 15286 13308 15292 13320
rect 14976 13280 15292 13308
rect 14976 13268 14982 13280
rect 15286 13268 15292 13280
rect 15344 13268 15350 13320
rect 15749 13311 15807 13317
rect 15749 13277 15761 13311
rect 15795 13277 15807 13311
rect 15749 13271 15807 13277
rect 15933 13311 15991 13317
rect 15933 13277 15945 13311
rect 15979 13308 15991 13311
rect 16022 13308 16028 13320
rect 15979 13280 16028 13308
rect 15979 13277 15991 13280
rect 15933 13271 15991 13277
rect 10928 13212 11284 13240
rect 10928 13200 10934 13212
rect 12710 13200 12716 13252
rect 12768 13240 12774 13252
rect 15764 13240 15792 13271
rect 16022 13268 16028 13280
rect 16080 13268 16086 13320
rect 16390 13268 16396 13320
rect 16448 13308 16454 13320
rect 16669 13311 16727 13317
rect 16669 13308 16681 13311
rect 16448 13280 16681 13308
rect 16448 13268 16454 13280
rect 16669 13277 16681 13280
rect 16715 13277 16727 13311
rect 16669 13271 16727 13277
rect 17589 13311 17647 13317
rect 17589 13277 17601 13311
rect 17635 13277 17647 13311
rect 17589 13271 17647 13277
rect 16206 13240 16212 13252
rect 12768 13212 12940 13240
rect 15764 13212 16212 13240
rect 12768 13200 12774 13212
rect 9030 13172 9036 13184
rect 8352 13144 8397 13172
rect 8772 13144 9036 13172
rect 8352 13132 8358 13144
rect 9030 13132 9036 13144
rect 9088 13132 9094 13184
rect 9306 13172 9312 13184
rect 9267 13144 9312 13172
rect 9306 13132 9312 13144
rect 9364 13132 9370 13184
rect 10689 13175 10747 13181
rect 10689 13141 10701 13175
rect 10735 13172 10747 13175
rect 12802 13172 12808 13184
rect 10735 13144 12808 13172
rect 10735 13141 10747 13144
rect 10689 13135 10747 13141
rect 12802 13132 12808 13144
rect 12860 13132 12866 13184
rect 12912 13181 12940 13212
rect 16206 13200 16212 13212
rect 16264 13200 16270 13252
rect 17604 13240 17632 13271
rect 17678 13268 17684 13320
rect 17736 13308 17742 13320
rect 18325 13311 18383 13317
rect 18325 13308 18337 13311
rect 17736 13280 18337 13308
rect 17736 13268 17742 13280
rect 18325 13277 18337 13280
rect 18371 13277 18383 13311
rect 18325 13271 18383 13277
rect 18509 13311 18567 13317
rect 18509 13277 18521 13311
rect 18555 13308 18567 13311
rect 18598 13308 18604 13320
rect 18555 13280 18604 13308
rect 18555 13277 18567 13280
rect 18509 13271 18567 13277
rect 18598 13268 18604 13280
rect 18656 13308 18662 13320
rect 19426 13308 19432 13320
rect 18656 13280 19432 13308
rect 18656 13268 18662 13280
rect 19426 13268 19432 13280
rect 19484 13268 19490 13320
rect 18874 13240 18880 13252
rect 17604 13212 18880 13240
rect 18874 13200 18880 13212
rect 18932 13200 18938 13252
rect 12897 13175 12955 13181
rect 12897 13141 12909 13175
rect 12943 13172 12955 13175
rect 13630 13172 13636 13184
rect 12943 13144 13636 13172
rect 12943 13141 12955 13144
rect 12897 13135 12955 13141
rect 13630 13132 13636 13144
rect 13688 13132 13694 13184
rect 13722 13132 13728 13184
rect 13780 13172 13786 13184
rect 14182 13172 14188 13184
rect 13780 13144 14188 13172
rect 13780 13132 13786 13144
rect 14182 13132 14188 13144
rect 14240 13172 14246 13184
rect 19429 13175 19487 13181
rect 19429 13172 19441 13175
rect 14240 13144 19441 13172
rect 14240 13132 14246 13144
rect 19429 13141 19441 13144
rect 19475 13172 19487 13175
rect 19886 13172 19892 13184
rect 19475 13144 19892 13172
rect 19475 13141 19487 13144
rect 19429 13135 19487 13141
rect 19886 13132 19892 13144
rect 19944 13132 19950 13184
rect 1104 13082 21896 13104
rect 1104 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 4575 13082
rect 4627 13030 4639 13082
rect 4691 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 18308 13082
rect 18360 13030 18372 13082
rect 18424 13030 18436 13082
rect 18488 13030 18500 13082
rect 18552 13030 21896 13082
rect 1104 13008 21896 13030
rect 3234 12968 3240 12980
rect 3195 12940 3240 12968
rect 3234 12928 3240 12940
rect 3292 12928 3298 12980
rect 3786 12968 3792 12980
rect 3747 12940 3792 12968
rect 3786 12928 3792 12940
rect 3844 12928 3850 12980
rect 4798 12968 4804 12980
rect 4759 12940 4804 12968
rect 4798 12928 4804 12940
rect 4856 12928 4862 12980
rect 5626 12928 5632 12980
rect 5684 12968 5690 12980
rect 5905 12971 5963 12977
rect 5905 12968 5917 12971
rect 5684 12940 5917 12968
rect 5684 12928 5690 12940
rect 5905 12937 5917 12940
rect 5951 12937 5963 12971
rect 5905 12931 5963 12937
rect 5994 12928 6000 12980
rect 6052 12968 6058 12980
rect 6825 12971 6883 12977
rect 6825 12968 6837 12971
rect 6052 12940 6837 12968
rect 6052 12928 6058 12940
rect 6825 12937 6837 12940
rect 6871 12937 6883 12971
rect 6825 12931 6883 12937
rect 7098 12928 7104 12980
rect 7156 12968 7162 12980
rect 8570 12968 8576 12980
rect 7156 12940 8576 12968
rect 7156 12928 7162 12940
rect 8570 12928 8576 12940
rect 8628 12928 8634 12980
rect 9122 12928 9128 12980
rect 9180 12928 9186 12980
rect 11790 12968 11796 12980
rect 10244 12940 11796 12968
rect 4614 12860 4620 12912
rect 4672 12900 4678 12912
rect 5074 12900 5080 12912
rect 4672 12872 5080 12900
rect 4672 12860 4678 12872
rect 5074 12860 5080 12872
rect 5132 12860 5138 12912
rect 9140 12900 9168 12928
rect 10134 12900 10140 12912
rect 9048 12872 10140 12900
rect 3510 12792 3516 12844
rect 3568 12792 3574 12844
rect 4246 12792 4252 12844
rect 4304 12832 4310 12844
rect 4341 12835 4399 12841
rect 4341 12832 4353 12835
rect 4304 12804 4353 12832
rect 4304 12792 4310 12804
rect 4341 12801 4353 12804
rect 4387 12832 4399 12835
rect 5350 12832 5356 12844
rect 4387 12804 5120 12832
rect 5311 12804 5356 12832
rect 4387 12801 4399 12804
rect 4341 12795 4399 12801
rect 1854 12764 1860 12776
rect 1767 12736 1860 12764
rect 1854 12724 1860 12736
rect 1912 12764 1918 12776
rect 2590 12764 2596 12776
rect 1912 12736 2596 12764
rect 1912 12724 1918 12736
rect 2590 12724 2596 12736
rect 2648 12724 2654 12776
rect 3528 12764 3556 12792
rect 5092 12776 5120 12804
rect 5350 12792 5356 12804
rect 5408 12792 5414 12844
rect 5626 12792 5632 12844
rect 5684 12832 5690 12844
rect 6362 12832 6368 12844
rect 5684 12804 6368 12832
rect 5684 12792 5690 12804
rect 6362 12792 6368 12804
rect 6420 12792 6426 12844
rect 6546 12832 6552 12844
rect 6507 12804 6552 12832
rect 6546 12792 6552 12804
rect 6604 12792 6610 12844
rect 7374 12832 7380 12844
rect 7335 12804 7380 12832
rect 7374 12792 7380 12804
rect 7432 12792 7438 12844
rect 8389 12835 8447 12841
rect 8389 12801 8401 12835
rect 8435 12832 8447 12835
rect 8662 12832 8668 12844
rect 8435 12804 8668 12832
rect 8435 12801 8447 12804
rect 8389 12795 8447 12801
rect 8662 12792 8668 12804
rect 8720 12792 8726 12844
rect 9048 12841 9076 12872
rect 10134 12860 10140 12872
rect 10192 12860 10198 12912
rect 9033 12835 9091 12841
rect 9033 12801 9045 12835
rect 9079 12801 9091 12835
rect 9033 12795 9091 12801
rect 9122 12792 9128 12844
rect 9180 12832 9186 12844
rect 9490 12832 9496 12844
rect 9180 12804 9496 12832
rect 9180 12792 9186 12804
rect 9490 12792 9496 12804
rect 9548 12792 9554 12844
rect 10244 12841 10272 12940
rect 11790 12928 11796 12940
rect 11848 12928 11854 12980
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 14369 12971 14427 12977
rect 14369 12968 14381 12971
rect 12492 12940 14381 12968
rect 12492 12928 12498 12940
rect 14369 12937 14381 12940
rect 14415 12937 14427 12971
rect 14642 12968 14648 12980
rect 14603 12940 14648 12968
rect 14369 12931 14427 12937
rect 10229 12835 10287 12841
rect 10229 12801 10241 12835
rect 10275 12801 10287 12835
rect 11808 12832 11836 12928
rect 13265 12903 13323 12909
rect 13265 12869 13277 12903
rect 13311 12900 13323 12903
rect 13906 12900 13912 12912
rect 13311 12872 13912 12900
rect 13311 12869 13323 12872
rect 13265 12863 13323 12869
rect 13906 12860 13912 12872
rect 13964 12860 13970 12912
rect 14093 12903 14151 12909
rect 14093 12869 14105 12903
rect 14139 12869 14151 12903
rect 14384 12900 14412 12931
rect 14642 12928 14648 12940
rect 14700 12928 14706 12980
rect 14826 12928 14832 12980
rect 14884 12968 14890 12980
rect 14921 12971 14979 12977
rect 14921 12968 14933 12971
rect 14884 12940 14933 12968
rect 14884 12928 14890 12940
rect 14921 12937 14933 12940
rect 14967 12937 14979 12971
rect 14921 12931 14979 12937
rect 15378 12928 15384 12980
rect 15436 12968 15442 12980
rect 16025 12971 16083 12977
rect 16025 12968 16037 12971
rect 15436 12940 16037 12968
rect 15436 12928 15442 12940
rect 16025 12937 16037 12940
rect 16071 12937 16083 12971
rect 16025 12931 16083 12937
rect 17129 12971 17187 12977
rect 17129 12937 17141 12971
rect 17175 12968 17187 12971
rect 17678 12968 17684 12980
rect 17175 12940 17684 12968
rect 17175 12937 17187 12940
rect 17129 12931 17187 12937
rect 17678 12928 17684 12940
rect 17736 12928 17742 12980
rect 18046 12928 18052 12980
rect 18104 12968 18110 12980
rect 19521 12971 19579 12977
rect 19521 12968 19533 12971
rect 18104 12940 19533 12968
rect 18104 12928 18110 12940
rect 19521 12937 19533 12940
rect 19567 12937 19579 12971
rect 20990 12968 20996 12980
rect 20951 12940 20996 12968
rect 19521 12931 19579 12937
rect 20990 12928 20996 12940
rect 21048 12928 21054 12980
rect 14550 12900 14556 12912
rect 14384 12872 14556 12900
rect 14093 12863 14151 12869
rect 12989 12835 13047 12841
rect 12989 12832 13001 12835
rect 11808 12804 13001 12832
rect 10229 12795 10287 12801
rect 12989 12801 13001 12804
rect 13035 12801 13047 12835
rect 12989 12795 13047 12801
rect 13630 12792 13636 12844
rect 13688 12832 13694 12844
rect 13817 12835 13875 12841
rect 13817 12832 13829 12835
rect 13688 12804 13829 12832
rect 13688 12792 13694 12804
rect 13817 12801 13829 12804
rect 13863 12801 13875 12835
rect 13817 12795 13875 12801
rect 13998 12792 14004 12844
rect 14056 12832 14062 12844
rect 14108 12832 14136 12863
rect 14550 12860 14556 12872
rect 14608 12860 14614 12912
rect 19426 12900 19432 12912
rect 19387 12872 19432 12900
rect 19426 12860 19432 12872
rect 19484 12900 19490 12912
rect 19484 12872 20116 12900
rect 19484 12860 19490 12872
rect 14056 12804 14136 12832
rect 15565 12835 15623 12841
rect 14056 12792 14062 12804
rect 15565 12801 15577 12835
rect 15611 12832 15623 12835
rect 16022 12832 16028 12844
rect 15611 12804 16028 12832
rect 15611 12801 15623 12804
rect 15565 12795 15623 12801
rect 16022 12792 16028 12804
rect 16080 12832 16086 12844
rect 20088 12841 20116 12872
rect 16577 12835 16635 12841
rect 16577 12832 16589 12835
rect 16080 12804 16589 12832
rect 16080 12792 16086 12804
rect 16577 12801 16589 12804
rect 16623 12801 16635 12835
rect 16577 12795 16635 12801
rect 17773 12835 17831 12841
rect 17773 12801 17785 12835
rect 17819 12832 17831 12835
rect 20073 12835 20131 12841
rect 17819 12804 18184 12832
rect 17819 12801 17831 12804
rect 17773 12795 17831 12801
rect 3528 12736 4752 12764
rect 2124 12699 2182 12705
rect 2124 12665 2136 12699
rect 2170 12696 2182 12699
rect 2498 12696 2504 12708
rect 2170 12668 2504 12696
rect 2170 12665 2182 12668
rect 2124 12659 2182 12665
rect 2498 12656 2504 12668
rect 2556 12656 2562 12708
rect 3510 12656 3516 12708
rect 3568 12696 3574 12708
rect 3697 12699 3755 12705
rect 3697 12696 3709 12699
rect 3568 12668 3709 12696
rect 3568 12656 3574 12668
rect 3697 12665 3709 12668
rect 3743 12696 3755 12699
rect 4249 12699 4307 12705
rect 4249 12696 4261 12699
rect 3743 12668 4261 12696
rect 3743 12665 3755 12668
rect 3697 12659 3755 12665
rect 4249 12665 4261 12668
rect 4295 12665 4307 12699
rect 4249 12659 4307 12665
rect 4154 12628 4160 12640
rect 4115 12600 4160 12628
rect 4154 12588 4160 12600
rect 4212 12588 4218 12640
rect 4724 12628 4752 12736
rect 4798 12724 4804 12776
rect 4856 12764 4862 12776
rect 4982 12764 4988 12776
rect 4856 12736 4988 12764
rect 4856 12724 4862 12736
rect 4982 12724 4988 12736
rect 5040 12724 5046 12776
rect 5074 12724 5080 12776
rect 5132 12724 5138 12776
rect 5902 12724 5908 12776
rect 5960 12724 5966 12776
rect 7193 12767 7251 12773
rect 7193 12764 7205 12767
rect 6104 12736 7205 12764
rect 5261 12699 5319 12705
rect 5261 12665 5273 12699
rect 5307 12696 5319 12699
rect 5920 12696 5948 12724
rect 5307 12668 5948 12696
rect 5307 12665 5319 12668
rect 5261 12659 5319 12665
rect 4982 12628 4988 12640
rect 4724 12600 4988 12628
rect 4982 12588 4988 12600
rect 5040 12588 5046 12640
rect 5169 12631 5227 12637
rect 5169 12597 5181 12631
rect 5215 12628 5227 12631
rect 5534 12628 5540 12640
rect 5215 12600 5540 12628
rect 5215 12597 5227 12600
rect 5169 12591 5227 12597
rect 5534 12588 5540 12600
rect 5592 12588 5598 12640
rect 5718 12628 5724 12640
rect 5679 12600 5724 12628
rect 5718 12588 5724 12600
rect 5776 12628 5782 12640
rect 6104 12628 6132 12736
rect 7193 12733 7205 12736
rect 7239 12733 7251 12767
rect 7193 12727 7251 12733
rect 8478 12724 8484 12776
rect 8536 12764 8542 12776
rect 8941 12767 8999 12773
rect 8941 12764 8953 12767
rect 8536 12736 8953 12764
rect 8536 12724 8542 12736
rect 8941 12733 8953 12736
rect 8987 12764 8999 12767
rect 9306 12764 9312 12776
rect 8987 12736 9312 12764
rect 8987 12733 8999 12736
rect 8941 12727 8999 12733
rect 9306 12724 9312 12736
rect 9364 12724 9370 12776
rect 9953 12767 10011 12773
rect 9953 12733 9965 12767
rect 9999 12764 10011 12767
rect 10042 12764 10048 12776
rect 9999 12736 10048 12764
rect 9999 12733 10011 12736
rect 9953 12727 10011 12733
rect 10042 12724 10048 12736
rect 10100 12724 10106 12776
rect 10413 12767 10471 12773
rect 10413 12733 10425 12767
rect 10459 12764 10471 12767
rect 10502 12764 10508 12776
rect 10459 12736 10508 12764
rect 10459 12733 10471 12736
rect 10413 12727 10471 12733
rect 10502 12724 10508 12736
rect 10560 12724 10566 12776
rect 13725 12767 13783 12773
rect 13725 12764 13737 12767
rect 10612 12736 13737 12764
rect 6365 12699 6423 12705
rect 6365 12665 6377 12699
rect 6411 12696 6423 12699
rect 7374 12696 7380 12708
rect 6411 12668 7380 12696
rect 6411 12665 6423 12668
rect 6365 12659 6423 12665
rect 7374 12656 7380 12668
rect 7432 12656 7438 12708
rect 8113 12699 8171 12705
rect 8113 12665 8125 12699
rect 8159 12696 8171 12699
rect 10612 12696 10640 12736
rect 13725 12733 13737 12736
rect 13771 12733 13783 12767
rect 13725 12727 13783 12733
rect 14090 12724 14096 12776
rect 14148 12764 14154 12776
rect 14277 12767 14335 12773
rect 14277 12764 14289 12767
rect 14148 12736 14289 12764
rect 14148 12724 14154 12736
rect 14277 12733 14289 12736
rect 14323 12733 14335 12767
rect 14277 12727 14335 12733
rect 14550 12724 14556 12776
rect 14608 12764 14614 12776
rect 16485 12767 16543 12773
rect 16485 12764 16497 12767
rect 14608 12736 16497 12764
rect 14608 12724 14614 12736
rect 16485 12733 16497 12736
rect 16531 12764 16543 12767
rect 16853 12767 16911 12773
rect 16853 12764 16865 12767
rect 16531 12736 16865 12764
rect 16531 12733 16543 12736
rect 16485 12727 16543 12733
rect 16853 12733 16865 12736
rect 16899 12733 16911 12767
rect 16853 12727 16911 12733
rect 17310 12724 17316 12776
rect 17368 12764 17374 12776
rect 18049 12767 18107 12773
rect 18049 12764 18061 12767
rect 17368 12736 18061 12764
rect 17368 12724 17374 12736
rect 18049 12733 18061 12736
rect 18095 12733 18107 12767
rect 18049 12727 18107 12733
rect 8159 12668 8800 12696
rect 8159 12665 8171 12668
rect 8113 12659 8171 12665
rect 8772 12640 8800 12668
rect 9600 12668 10640 12696
rect 10680 12699 10738 12705
rect 6270 12628 6276 12640
rect 5776 12600 6132 12628
rect 6231 12600 6276 12628
rect 5776 12588 5782 12600
rect 6270 12588 6276 12600
rect 6328 12588 6334 12640
rect 6546 12588 6552 12640
rect 6604 12628 6610 12640
rect 6822 12628 6828 12640
rect 6604 12600 6828 12628
rect 6604 12588 6610 12600
rect 6822 12588 6828 12600
rect 6880 12588 6886 12640
rect 6914 12588 6920 12640
rect 6972 12628 6978 12640
rect 7282 12628 7288 12640
rect 6972 12600 7288 12628
rect 6972 12588 6978 12600
rect 7282 12588 7288 12600
rect 7340 12588 7346 12640
rect 7558 12588 7564 12640
rect 7616 12628 7622 12640
rect 7745 12631 7803 12637
rect 7745 12628 7757 12631
rect 7616 12600 7757 12628
rect 7616 12588 7622 12600
rect 7745 12597 7757 12600
rect 7791 12597 7803 12631
rect 7745 12591 7803 12597
rect 8205 12631 8263 12637
rect 8205 12597 8217 12631
rect 8251 12628 8263 12631
rect 8573 12631 8631 12637
rect 8573 12628 8585 12631
rect 8251 12600 8585 12628
rect 8251 12597 8263 12600
rect 8205 12591 8263 12597
rect 8573 12597 8585 12600
rect 8619 12597 8631 12631
rect 8573 12591 8631 12597
rect 8754 12588 8760 12640
rect 8812 12588 8818 12640
rect 9122 12588 9128 12640
rect 9180 12628 9186 12640
rect 9600 12637 9628 12668
rect 10680 12665 10692 12699
rect 10726 12696 10738 12699
rect 10870 12696 10876 12708
rect 10726 12668 10876 12696
rect 10726 12665 10738 12668
rect 10680 12659 10738 12665
rect 10870 12656 10876 12668
rect 10928 12656 10934 12708
rect 11422 12656 11428 12708
rect 11480 12696 11486 12708
rect 12161 12699 12219 12705
rect 12161 12696 12173 12699
rect 11480 12668 12173 12696
rect 11480 12656 11486 12668
rect 12161 12665 12173 12668
rect 12207 12665 12219 12699
rect 13633 12699 13691 12705
rect 13633 12696 13645 12699
rect 12161 12659 12219 12665
rect 12452 12668 13645 12696
rect 9401 12631 9459 12637
rect 9401 12628 9413 12631
rect 9180 12600 9413 12628
rect 9180 12588 9186 12600
rect 9401 12597 9413 12600
rect 9447 12597 9459 12631
rect 9401 12591 9459 12597
rect 9585 12631 9643 12637
rect 9585 12597 9597 12631
rect 9631 12597 9643 12631
rect 9585 12591 9643 12597
rect 10045 12631 10103 12637
rect 10045 12597 10057 12631
rect 10091 12628 10103 12631
rect 11238 12628 11244 12640
rect 10091 12600 11244 12628
rect 10091 12597 10103 12600
rect 10045 12591 10103 12597
rect 11238 12588 11244 12600
rect 11296 12588 11302 12640
rect 11882 12588 11888 12640
rect 11940 12628 11946 12640
rect 12452 12637 12480 12668
rect 13633 12665 13645 12668
rect 13679 12665 13691 12699
rect 13633 12659 13691 12665
rect 13906 12656 13912 12708
rect 13964 12696 13970 12708
rect 14737 12699 14795 12705
rect 14737 12696 14749 12699
rect 13964 12668 14749 12696
rect 13964 12656 13970 12668
rect 14737 12665 14749 12668
rect 14783 12696 14795 12699
rect 15289 12699 15347 12705
rect 15289 12696 15301 12699
rect 14783 12668 15301 12696
rect 14783 12665 14795 12668
rect 14737 12659 14795 12665
rect 15289 12665 15301 12668
rect 15335 12665 15347 12699
rect 15289 12659 15347 12665
rect 15381 12699 15439 12705
rect 15381 12665 15393 12699
rect 15427 12696 15439 12699
rect 15470 12696 15476 12708
rect 15427 12668 15476 12696
rect 15427 12665 15439 12668
rect 15381 12659 15439 12665
rect 15470 12656 15476 12668
rect 15528 12656 15534 12708
rect 16393 12699 16451 12705
rect 16393 12665 16405 12699
rect 16439 12696 16451 12699
rect 16666 12696 16672 12708
rect 16439 12668 16672 12696
rect 16439 12665 16451 12668
rect 16393 12659 16451 12665
rect 16666 12656 16672 12668
rect 16724 12656 16730 12708
rect 16942 12656 16948 12708
rect 17000 12696 17006 12708
rect 17589 12699 17647 12705
rect 17589 12696 17601 12699
rect 17000 12668 17601 12696
rect 17000 12656 17006 12668
rect 17589 12665 17601 12668
rect 17635 12665 17647 12699
rect 18156 12696 18184 12804
rect 20073 12801 20085 12835
rect 20119 12801 20131 12835
rect 20073 12795 20131 12801
rect 19886 12764 19892 12776
rect 19847 12736 19892 12764
rect 19886 12724 19892 12736
rect 19944 12724 19950 12776
rect 20254 12724 20260 12776
rect 20312 12764 20318 12776
rect 20809 12767 20867 12773
rect 20809 12764 20821 12767
rect 20312 12736 20821 12764
rect 20312 12724 20318 12736
rect 20809 12733 20821 12736
rect 20855 12733 20867 12767
rect 20809 12727 20867 12733
rect 18316 12699 18374 12705
rect 18316 12696 18328 12699
rect 18156 12668 18328 12696
rect 17589 12659 17647 12665
rect 18316 12665 18328 12668
rect 18362 12696 18374 12699
rect 18690 12696 18696 12708
rect 18362 12668 18696 12696
rect 18362 12665 18374 12668
rect 18316 12659 18374 12665
rect 18690 12656 18696 12668
rect 18748 12656 18754 12708
rect 19334 12656 19340 12708
rect 19392 12696 19398 12708
rect 19981 12699 20039 12705
rect 19981 12696 19993 12699
rect 19392 12668 19993 12696
rect 19392 12656 19398 12668
rect 19981 12665 19993 12668
rect 20027 12665 20039 12699
rect 19981 12659 20039 12665
rect 12437 12631 12495 12637
rect 11940 12600 11985 12628
rect 11940 12588 11946 12600
rect 12437 12597 12449 12631
rect 12483 12597 12495 12631
rect 12437 12591 12495 12597
rect 12526 12588 12532 12640
rect 12584 12628 12590 12640
rect 12805 12631 12863 12637
rect 12805 12628 12817 12631
rect 12584 12600 12817 12628
rect 12584 12588 12590 12600
rect 12805 12597 12817 12600
rect 12851 12597 12863 12631
rect 12805 12591 12863 12597
rect 12894 12588 12900 12640
rect 12952 12628 12958 12640
rect 12952 12600 12997 12628
rect 12952 12588 12958 12600
rect 13814 12588 13820 12640
rect 13872 12628 13878 12640
rect 13998 12628 14004 12640
rect 13872 12600 14004 12628
rect 13872 12588 13878 12600
rect 13998 12588 14004 12600
rect 14056 12628 14062 12640
rect 15841 12631 15899 12637
rect 15841 12628 15853 12631
rect 14056 12600 15853 12628
rect 14056 12588 14062 12600
rect 15841 12597 15853 12600
rect 15887 12628 15899 12631
rect 15930 12628 15936 12640
rect 15887 12600 15936 12628
rect 15887 12597 15899 12600
rect 15841 12591 15899 12597
rect 15930 12588 15936 12600
rect 15988 12588 15994 12640
rect 16758 12588 16764 12640
rect 16816 12628 16822 12640
rect 17497 12631 17555 12637
rect 17497 12628 17509 12631
rect 16816 12600 17509 12628
rect 16816 12588 16822 12600
rect 17497 12597 17509 12600
rect 17543 12597 17555 12631
rect 17497 12591 17555 12597
rect 1104 12538 21896 12560
rect 1104 12486 7912 12538
rect 7964 12486 7976 12538
rect 8028 12486 8040 12538
rect 8092 12486 8104 12538
rect 8156 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 15035 12538
rect 15087 12486 21896 12538
rect 1104 12464 21896 12486
rect 1670 12424 1676 12436
rect 1631 12396 1676 12424
rect 1670 12384 1676 12396
rect 1728 12384 1734 12436
rect 1762 12384 1768 12436
rect 1820 12424 1826 12436
rect 1857 12427 1915 12433
rect 1857 12424 1869 12427
rect 1820 12396 1869 12424
rect 1820 12384 1826 12396
rect 1857 12393 1869 12396
rect 1903 12393 1915 12427
rect 1857 12387 1915 12393
rect 2317 12427 2375 12433
rect 2317 12393 2329 12427
rect 2363 12424 2375 12427
rect 2777 12427 2835 12433
rect 2777 12424 2789 12427
rect 2363 12396 2789 12424
rect 2363 12393 2375 12396
rect 2317 12387 2375 12393
rect 2777 12393 2789 12396
rect 2823 12393 2835 12427
rect 2777 12387 2835 12393
rect 4065 12427 4123 12433
rect 4065 12393 4077 12427
rect 4111 12424 4123 12427
rect 4154 12424 4160 12436
rect 4111 12396 4160 12424
rect 4111 12393 4123 12396
rect 4065 12387 4123 12393
rect 4154 12384 4160 12396
rect 4212 12384 4218 12436
rect 4338 12384 4344 12436
rect 4396 12424 4402 12436
rect 4525 12427 4583 12433
rect 4525 12424 4537 12427
rect 4396 12396 4537 12424
rect 4396 12384 4402 12396
rect 4525 12393 4537 12396
rect 4571 12393 4583 12427
rect 4525 12387 4583 12393
rect 4985 12427 5043 12433
rect 4985 12393 4997 12427
rect 5031 12424 5043 12427
rect 5445 12427 5503 12433
rect 5445 12424 5457 12427
rect 5031 12396 5457 12424
rect 5031 12393 5043 12396
rect 4985 12387 5043 12393
rect 5445 12393 5457 12396
rect 5491 12424 5503 12427
rect 7285 12427 7343 12433
rect 5491 12396 6684 12424
rect 5491 12393 5503 12396
rect 5445 12387 5503 12393
rect 3970 12316 3976 12368
rect 4028 12356 4034 12368
rect 6178 12356 6184 12368
rect 4028 12328 6184 12356
rect 4028 12316 4034 12328
rect 1486 12288 1492 12300
rect 1447 12260 1492 12288
rect 1486 12248 1492 12260
rect 1544 12248 1550 12300
rect 2222 12288 2228 12300
rect 2183 12260 2228 12288
rect 2222 12248 2228 12260
rect 2280 12248 2286 12300
rect 3145 12291 3203 12297
rect 3145 12257 3157 12291
rect 3191 12288 3203 12291
rect 4246 12288 4252 12300
rect 3191 12260 4252 12288
rect 3191 12257 3203 12260
rect 3145 12251 3203 12257
rect 4246 12248 4252 12260
rect 4304 12248 4310 12300
rect 4893 12291 4951 12297
rect 4893 12288 4905 12291
rect 4356 12260 4905 12288
rect 2498 12220 2504 12232
rect 2459 12192 2504 12220
rect 2498 12180 2504 12192
rect 2556 12180 2562 12232
rect 3234 12220 3240 12232
rect 3195 12192 3240 12220
rect 3234 12180 3240 12192
rect 3292 12180 3298 12232
rect 3329 12223 3387 12229
rect 3329 12189 3341 12223
rect 3375 12189 3387 12223
rect 3329 12183 3387 12189
rect 2682 12112 2688 12164
rect 2740 12152 2746 12164
rect 3344 12152 3372 12183
rect 2740 12124 3372 12152
rect 2740 12112 2746 12124
rect 3970 12044 3976 12096
rect 4028 12084 4034 12096
rect 4356 12093 4384 12260
rect 4893 12257 4905 12260
rect 4939 12257 4951 12291
rect 4893 12251 4951 12257
rect 5828 12232 5856 12328
rect 6178 12316 6184 12328
rect 6236 12316 6242 12368
rect 6656 12356 6684 12396
rect 7285 12393 7297 12427
rect 7331 12424 7343 12427
rect 7466 12424 7472 12436
rect 7331 12396 7472 12424
rect 7331 12393 7343 12396
rect 7285 12387 7343 12393
rect 7466 12384 7472 12396
rect 7524 12384 7530 12436
rect 8478 12424 8484 12436
rect 7567 12396 8484 12424
rect 7567 12356 7595 12396
rect 8478 12384 8484 12396
rect 8536 12384 8542 12436
rect 8662 12384 8668 12436
rect 8720 12424 8726 12436
rect 9401 12427 9459 12433
rect 9401 12424 9413 12427
rect 8720 12396 9413 12424
rect 8720 12384 8726 12396
rect 9401 12393 9413 12396
rect 9447 12393 9459 12427
rect 9401 12387 9459 12393
rect 10042 12384 10048 12436
rect 10100 12424 10106 12436
rect 10137 12427 10195 12433
rect 10137 12424 10149 12427
rect 10100 12396 10149 12424
rect 10100 12384 10106 12396
rect 10137 12393 10149 12396
rect 10183 12393 10195 12427
rect 11422 12424 11428 12436
rect 11383 12396 11428 12424
rect 10137 12387 10195 12393
rect 11422 12384 11428 12396
rect 11480 12384 11486 12436
rect 11793 12427 11851 12433
rect 11793 12393 11805 12427
rect 11839 12393 11851 12427
rect 11793 12387 11851 12393
rect 8294 12365 8300 12368
rect 6656 12328 7595 12356
rect 8288 12319 8300 12365
rect 8352 12356 8358 12368
rect 8352 12328 8388 12356
rect 8294 12316 8300 12319
rect 8352 12316 8358 12328
rect 8938 12316 8944 12368
rect 8996 12316 9002 12368
rect 9766 12316 9772 12368
rect 9824 12356 9830 12368
rect 9861 12359 9919 12365
rect 9861 12356 9873 12359
rect 9824 12328 9873 12356
rect 9824 12316 9830 12328
rect 9861 12325 9873 12328
rect 9907 12356 9919 12359
rect 11808 12356 11836 12387
rect 11882 12384 11888 12436
rect 11940 12424 11946 12436
rect 12161 12427 12219 12433
rect 12161 12424 12173 12427
rect 11940 12396 12173 12424
rect 11940 12384 11946 12396
rect 12161 12393 12173 12396
rect 12207 12393 12219 12427
rect 12161 12387 12219 12393
rect 12434 12384 12440 12436
rect 12492 12424 12498 12436
rect 16758 12424 16764 12436
rect 12492 12396 16764 12424
rect 12492 12384 12498 12396
rect 16758 12384 16764 12396
rect 16816 12384 16822 12436
rect 16942 12424 16948 12436
rect 16903 12396 16948 12424
rect 16942 12384 16948 12396
rect 17000 12384 17006 12436
rect 17126 12384 17132 12436
rect 17184 12424 17190 12436
rect 17221 12427 17279 12433
rect 17221 12424 17233 12427
rect 17184 12396 17233 12424
rect 17184 12384 17190 12396
rect 17221 12393 17233 12396
rect 17267 12424 17279 12427
rect 17678 12424 17684 12436
rect 17267 12396 17684 12424
rect 17267 12393 17279 12396
rect 17221 12387 17279 12393
rect 17678 12384 17684 12396
rect 17736 12384 17742 12436
rect 18782 12424 18788 12436
rect 18743 12396 18788 12424
rect 18782 12384 18788 12396
rect 18840 12384 18846 12436
rect 19245 12427 19303 12433
rect 19245 12393 19257 12427
rect 19291 12424 19303 12427
rect 19426 12424 19432 12436
rect 19291 12396 19432 12424
rect 19291 12393 19303 12396
rect 19245 12387 19303 12393
rect 19426 12384 19432 12396
rect 19484 12384 19490 12436
rect 12526 12356 12532 12368
rect 9907 12328 11376 12356
rect 11808 12328 12532 12356
rect 9907 12325 9919 12328
rect 9861 12319 9919 12325
rect 6086 12297 6092 12300
rect 6080 12288 6092 12297
rect 6047 12260 6092 12288
rect 6080 12251 6092 12260
rect 6086 12248 6092 12251
rect 6144 12248 6150 12300
rect 7466 12288 7472 12300
rect 7427 12260 7472 12288
rect 7466 12248 7472 12260
rect 7524 12248 7530 12300
rect 7929 12291 7987 12297
rect 7929 12257 7941 12291
rect 7975 12288 7987 12291
rect 8956 12288 8984 12316
rect 9122 12288 9128 12300
rect 7975 12260 9128 12288
rect 7975 12257 7987 12260
rect 7929 12251 7987 12257
rect 9122 12248 9128 12260
rect 9180 12248 9186 12300
rect 11348 12297 11376 12328
rect 12526 12316 12532 12328
rect 12584 12316 12590 12368
rect 12802 12316 12808 12368
rect 12860 12356 12866 12368
rect 12958 12359 13016 12365
rect 12958 12356 12970 12359
rect 12860 12328 12970 12356
rect 12860 12316 12866 12328
rect 12958 12325 12970 12328
rect 13004 12325 13016 12359
rect 12958 12319 13016 12325
rect 14182 12316 14188 12368
rect 14240 12356 14246 12368
rect 15534 12359 15592 12365
rect 15534 12356 15546 12359
rect 14240 12328 15546 12356
rect 14240 12316 14246 12328
rect 15534 12325 15546 12328
rect 15580 12325 15592 12359
rect 15534 12319 15592 12325
rect 15654 12316 15660 12368
rect 15712 12356 15718 12368
rect 20254 12356 20260 12368
rect 15712 12328 20024 12356
rect 20215 12328 20260 12356
rect 15712 12316 15718 12328
rect 9677 12291 9735 12297
rect 9677 12257 9689 12291
rect 9723 12288 9735 12291
rect 10505 12291 10563 12297
rect 10505 12288 10517 12291
rect 9723 12260 10517 12288
rect 9723 12257 9735 12260
rect 9677 12251 9735 12257
rect 10505 12257 10517 12260
rect 10551 12257 10563 12291
rect 10505 12251 10563 12257
rect 11333 12291 11391 12297
rect 11333 12257 11345 12291
rect 11379 12288 11391 12291
rect 11422 12288 11428 12300
rect 11379 12260 11428 12288
rect 11379 12257 11391 12260
rect 11333 12251 11391 12257
rect 11422 12248 11428 12260
rect 11480 12248 11486 12300
rect 11698 12248 11704 12300
rect 11756 12288 11762 12300
rect 12713 12291 12771 12297
rect 12713 12288 12725 12291
rect 11756 12260 12725 12288
rect 11756 12248 11762 12260
rect 12713 12257 12725 12260
rect 12759 12257 12771 12291
rect 12713 12251 12771 12257
rect 13906 12248 13912 12300
rect 13964 12288 13970 12300
rect 14274 12288 14280 12300
rect 13964 12260 14280 12288
rect 13964 12248 13970 12260
rect 14274 12248 14280 12260
rect 14332 12248 14338 12300
rect 17310 12288 17316 12300
rect 15304 12260 17316 12288
rect 15304 12232 15332 12260
rect 17310 12248 17316 12260
rect 17368 12248 17374 12300
rect 17586 12297 17592 12300
rect 17580 12288 17592 12297
rect 17547 12260 17592 12288
rect 17580 12251 17592 12260
rect 17586 12248 17592 12251
rect 17644 12248 17650 12300
rect 19996 12297 20024 12328
rect 20254 12316 20260 12328
rect 20312 12316 20318 12368
rect 19153 12291 19211 12297
rect 19153 12257 19165 12291
rect 19199 12288 19211 12291
rect 19981 12291 20039 12297
rect 19199 12260 19748 12288
rect 19199 12257 19211 12260
rect 19153 12251 19211 12257
rect 5074 12180 5080 12232
rect 5132 12220 5138 12232
rect 5810 12220 5816 12232
rect 5132 12192 5177 12220
rect 5771 12192 5816 12220
rect 5132 12180 5138 12192
rect 5810 12180 5816 12192
rect 5868 12180 5874 12232
rect 8018 12220 8024 12232
rect 7979 12192 8024 12220
rect 8018 12180 8024 12192
rect 8076 12180 8082 12232
rect 9398 12180 9404 12232
rect 9456 12180 9462 12232
rect 9858 12180 9864 12232
rect 9916 12220 9922 12232
rect 10226 12220 10232 12232
rect 9916 12192 10232 12220
rect 9916 12180 9922 12192
rect 10226 12180 10232 12192
rect 10284 12180 10290 12232
rect 10594 12220 10600 12232
rect 10555 12192 10600 12220
rect 10594 12180 10600 12192
rect 10652 12180 10658 12232
rect 10781 12223 10839 12229
rect 10781 12189 10793 12223
rect 10827 12220 10839 12223
rect 10870 12220 10876 12232
rect 10827 12192 10876 12220
rect 10827 12189 10839 12192
rect 10781 12183 10839 12189
rect 10870 12180 10876 12192
rect 10928 12180 10934 12232
rect 11146 12180 11152 12232
rect 11204 12220 11210 12232
rect 11517 12223 11575 12229
rect 11517 12220 11529 12223
rect 11204 12192 11529 12220
rect 11204 12180 11210 12192
rect 11517 12189 11529 12192
rect 11563 12189 11575 12223
rect 11517 12183 11575 12189
rect 11882 12180 11888 12232
rect 11940 12220 11946 12232
rect 12253 12223 12311 12229
rect 12253 12220 12265 12223
rect 11940 12192 12265 12220
rect 11940 12180 11946 12192
rect 12253 12189 12265 12192
rect 12299 12189 12311 12223
rect 12253 12183 12311 12189
rect 12437 12223 12495 12229
rect 12437 12189 12449 12223
rect 12483 12220 12495 12223
rect 12526 12220 12532 12232
rect 12483 12192 12532 12220
rect 12483 12189 12495 12192
rect 12437 12183 12495 12189
rect 12526 12180 12532 12192
rect 12584 12180 12590 12232
rect 14185 12223 14243 12229
rect 14185 12189 14197 12223
rect 14231 12220 14243 12223
rect 14734 12220 14740 12232
rect 14231 12192 14740 12220
rect 14231 12189 14243 12192
rect 14185 12183 14243 12189
rect 14734 12180 14740 12192
rect 14792 12180 14798 12232
rect 15286 12220 15292 12232
rect 15247 12192 15292 12220
rect 15286 12180 15292 12192
rect 15344 12180 15350 12232
rect 16666 12180 16672 12232
rect 16724 12220 16730 12232
rect 17126 12220 17132 12232
rect 16724 12192 17132 12220
rect 16724 12180 16730 12192
rect 17126 12180 17132 12192
rect 17184 12180 17190 12232
rect 19337 12223 19395 12229
rect 19337 12189 19349 12223
rect 19383 12189 19395 12223
rect 19337 12183 19395 12189
rect 9416 12152 9444 12180
rect 14642 12152 14648 12164
rect 9416 12124 12756 12152
rect 4341 12087 4399 12093
rect 4341 12084 4353 12087
rect 4028 12056 4353 12084
rect 4028 12044 4034 12056
rect 4341 12053 4353 12056
rect 4387 12053 4399 12087
rect 4341 12047 4399 12053
rect 4890 12044 4896 12096
rect 4948 12084 4954 12096
rect 5350 12084 5356 12096
rect 4948 12056 5356 12084
rect 4948 12044 4954 12056
rect 5350 12044 5356 12056
rect 5408 12044 5414 12096
rect 5534 12044 5540 12096
rect 5592 12084 5598 12096
rect 5629 12087 5687 12093
rect 5629 12084 5641 12087
rect 5592 12056 5641 12084
rect 5592 12044 5598 12056
rect 5629 12053 5641 12056
rect 5675 12053 5687 12087
rect 7190 12084 7196 12096
rect 7151 12056 7196 12084
rect 5629 12047 5687 12053
rect 7190 12044 7196 12056
rect 7248 12044 7254 12096
rect 7282 12044 7288 12096
rect 7340 12084 7346 12096
rect 7745 12087 7803 12093
rect 7745 12084 7757 12087
rect 7340 12056 7757 12084
rect 7340 12044 7346 12056
rect 7745 12053 7757 12056
rect 7791 12084 7803 12087
rect 7834 12084 7840 12096
rect 7791 12056 7840 12084
rect 7791 12053 7803 12056
rect 7745 12047 7803 12053
rect 7834 12044 7840 12056
rect 7892 12044 7898 12096
rect 8938 12044 8944 12096
rect 8996 12084 9002 12096
rect 9677 12087 9735 12093
rect 9677 12084 9689 12087
rect 8996 12056 9689 12084
rect 8996 12044 9002 12056
rect 9677 12053 9689 12056
rect 9723 12084 9735 12087
rect 9953 12087 10011 12093
rect 9953 12084 9965 12087
rect 9723 12056 9965 12084
rect 9723 12053 9735 12056
rect 9677 12047 9735 12053
rect 9953 12053 9965 12056
rect 9999 12053 10011 12087
rect 9953 12047 10011 12053
rect 10965 12087 11023 12093
rect 10965 12053 10977 12087
rect 11011 12084 11023 12087
rect 12434 12084 12440 12096
rect 11011 12056 12440 12084
rect 11011 12053 11023 12056
rect 10965 12047 11023 12053
rect 12434 12044 12440 12056
rect 12492 12044 12498 12096
rect 12728 12084 12756 12124
rect 13832 12124 14648 12152
rect 13832 12084 13860 12124
rect 14642 12112 14648 12124
rect 14700 12112 14706 12164
rect 18690 12152 18696 12164
rect 18651 12124 18696 12152
rect 18690 12112 18696 12124
rect 18748 12152 18754 12164
rect 19352 12152 19380 12183
rect 18748 12124 19380 12152
rect 18748 12112 18754 12124
rect 12728 12056 13860 12084
rect 13906 12044 13912 12096
rect 13964 12084 13970 12096
rect 14093 12087 14151 12093
rect 14093 12084 14105 12087
rect 13964 12056 14105 12084
rect 13964 12044 13970 12056
rect 14093 12053 14105 12056
rect 14139 12053 14151 12087
rect 14826 12084 14832 12096
rect 14787 12056 14832 12084
rect 14093 12047 14151 12053
rect 14826 12044 14832 12056
rect 14884 12044 14890 12096
rect 15013 12087 15071 12093
rect 15013 12053 15025 12087
rect 15059 12084 15071 12087
rect 16022 12084 16028 12096
rect 15059 12056 16028 12084
rect 15059 12053 15071 12056
rect 15013 12047 15071 12053
rect 16022 12044 16028 12056
rect 16080 12084 16086 12096
rect 16206 12084 16212 12096
rect 16080 12056 16212 12084
rect 16080 12044 16086 12056
rect 16206 12044 16212 12056
rect 16264 12044 16270 12096
rect 16574 12044 16580 12096
rect 16632 12084 16638 12096
rect 16669 12087 16727 12093
rect 16669 12084 16681 12087
rect 16632 12056 16681 12084
rect 16632 12044 16638 12056
rect 16669 12053 16681 12056
rect 16715 12053 16727 12087
rect 16669 12047 16727 12053
rect 16758 12044 16764 12096
rect 16816 12084 16822 12096
rect 17034 12084 17040 12096
rect 16816 12056 17040 12084
rect 16816 12044 16822 12056
rect 17034 12044 17040 12056
rect 17092 12044 17098 12096
rect 19720 12093 19748 12260
rect 19981 12257 19993 12291
rect 20027 12257 20039 12291
rect 19981 12251 20039 12257
rect 19705 12087 19763 12093
rect 19705 12053 19717 12087
rect 19751 12084 19763 12087
rect 20070 12084 20076 12096
rect 19751 12056 20076 12084
rect 19751 12053 19763 12056
rect 19705 12047 19763 12053
rect 20070 12044 20076 12056
rect 20128 12044 20134 12096
rect 22002 12016 22008 12028
rect 1104 11994 21896 12016
rect 1104 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 4575 11994
rect 4627 11942 4639 11994
rect 4691 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 18308 11994
rect 18360 11942 18372 11994
rect 18424 11942 18436 11994
rect 18488 11942 18500 11994
rect 18552 11942 21896 11994
rect 21963 11988 22008 12016
rect 22002 11976 22008 11988
rect 22060 11976 22066 12028
rect 1104 11920 21896 11942
rect 1854 11880 1860 11892
rect 1504 11852 1860 11880
rect 1504 11753 1532 11852
rect 1854 11840 1860 11852
rect 1912 11840 1918 11892
rect 2498 11840 2504 11892
rect 2556 11880 2562 11892
rect 2869 11883 2927 11889
rect 2869 11880 2881 11883
rect 2556 11852 2881 11880
rect 2556 11840 2562 11852
rect 2869 11849 2881 11852
rect 2915 11849 2927 11883
rect 3142 11880 3148 11892
rect 3103 11852 3148 11880
rect 2869 11843 2927 11849
rect 3142 11840 3148 11852
rect 3200 11840 3206 11892
rect 3234 11840 3240 11892
rect 3292 11880 3298 11892
rect 3421 11883 3479 11889
rect 3421 11880 3433 11883
rect 3292 11852 3433 11880
rect 3292 11840 3298 11852
rect 3421 11849 3433 11852
rect 3467 11849 3479 11883
rect 4246 11880 4252 11892
rect 4207 11852 4252 11880
rect 3421 11843 3479 11849
rect 4246 11840 4252 11852
rect 4304 11840 4310 11892
rect 6362 11880 6368 11892
rect 4356 11852 6368 11880
rect 3878 11772 3884 11824
rect 3936 11812 3942 11824
rect 4356 11812 4384 11852
rect 6362 11840 6368 11852
rect 6420 11840 6426 11892
rect 6914 11880 6920 11892
rect 6875 11852 6920 11880
rect 6914 11840 6920 11852
rect 6972 11840 6978 11892
rect 7101 11883 7159 11889
rect 7101 11849 7113 11883
rect 7147 11880 7159 11883
rect 7374 11880 7380 11892
rect 7147 11852 7380 11880
rect 7147 11849 7159 11852
rect 7101 11843 7159 11849
rect 7374 11840 7380 11852
rect 7432 11840 7438 11892
rect 8754 11880 8760 11892
rect 8715 11852 8760 11880
rect 8754 11840 8760 11852
rect 8812 11840 8818 11892
rect 10134 11880 10140 11892
rect 10095 11852 10140 11880
rect 10134 11840 10140 11852
rect 10192 11840 10198 11892
rect 10502 11880 10508 11892
rect 10336 11852 10508 11880
rect 3936 11784 4384 11812
rect 3936 11772 3942 11784
rect 6454 11772 6460 11824
rect 6512 11812 6518 11824
rect 6512 11784 6960 11812
rect 6512 11772 6518 11784
rect 6932 11756 6960 11784
rect 7190 11772 7196 11824
rect 7248 11812 7254 11824
rect 10042 11812 10048 11824
rect 7248 11784 7696 11812
rect 7248 11772 7254 11784
rect 1489 11747 1547 11753
rect 1489 11713 1501 11747
rect 1535 11713 1547 11747
rect 1489 11707 1547 11713
rect 3694 11704 3700 11756
rect 3752 11744 3758 11756
rect 4065 11747 4123 11753
rect 4065 11744 4077 11747
rect 3752 11716 4077 11744
rect 3752 11704 3758 11716
rect 4065 11713 4077 11716
rect 4111 11744 4123 11747
rect 4801 11747 4859 11753
rect 4801 11744 4813 11747
rect 4111 11716 4813 11744
rect 4111 11713 4123 11716
rect 4065 11707 4123 11713
rect 4801 11713 4813 11716
rect 4847 11713 4859 11747
rect 4801 11707 4859 11713
rect 6914 11704 6920 11756
rect 6972 11704 6978 11756
rect 2774 11636 2780 11688
rect 2832 11676 2838 11688
rect 2961 11679 3019 11685
rect 2961 11676 2973 11679
rect 2832 11648 2973 11676
rect 2832 11636 2838 11648
rect 2961 11645 2973 11648
rect 3007 11645 3019 11679
rect 2961 11639 3019 11645
rect 4338 11636 4344 11688
rect 4396 11676 4402 11688
rect 4982 11676 4988 11688
rect 4396 11648 4988 11676
rect 4396 11636 4402 11648
rect 4982 11636 4988 11648
rect 5040 11636 5046 11688
rect 5261 11679 5319 11685
rect 5261 11645 5273 11679
rect 5307 11645 5319 11679
rect 5261 11639 5319 11645
rect 5528 11679 5586 11685
rect 5528 11645 5540 11679
rect 5574 11676 5586 11679
rect 6362 11676 6368 11688
rect 5574 11648 6368 11676
rect 5574 11645 5586 11648
rect 5528 11639 5586 11645
rect 1756 11611 1814 11617
rect 1756 11577 1768 11611
rect 1802 11608 1814 11611
rect 2130 11608 2136 11620
rect 1802 11580 2136 11608
rect 1802 11577 1814 11580
rect 1756 11571 1814 11577
rect 2130 11568 2136 11580
rect 2188 11608 2194 11620
rect 2682 11608 2688 11620
rect 2188 11580 2688 11608
rect 2188 11568 2194 11580
rect 2682 11568 2688 11580
rect 2740 11568 2746 11620
rect 5276 11608 5304 11639
rect 6362 11636 6368 11648
rect 6420 11676 6426 11688
rect 7208 11676 7236 11772
rect 7558 11744 7564 11756
rect 7519 11716 7564 11744
rect 7558 11704 7564 11716
rect 7616 11704 7622 11756
rect 7668 11753 7696 11784
rect 7760 11784 9076 11812
rect 7653 11747 7711 11753
rect 7653 11713 7665 11747
rect 7699 11713 7711 11747
rect 7653 11707 7711 11713
rect 6420 11648 7236 11676
rect 6420 11636 6426 11648
rect 7282 11636 7288 11688
rect 7340 11676 7346 11688
rect 7760 11676 7788 11784
rect 8294 11704 8300 11756
rect 8352 11744 8358 11756
rect 8481 11747 8539 11753
rect 8481 11744 8493 11747
rect 8352 11716 8493 11744
rect 8352 11704 8358 11716
rect 8481 11713 8493 11716
rect 8527 11713 8539 11747
rect 8481 11707 8539 11713
rect 7340 11648 7788 11676
rect 8389 11679 8447 11685
rect 7340 11636 7346 11648
rect 8389 11645 8401 11679
rect 8435 11676 8447 11679
rect 8435 11648 8984 11676
rect 8435 11645 8447 11648
rect 8389 11639 8447 11645
rect 5810 11608 5816 11620
rect 5276 11580 5816 11608
rect 5810 11568 5816 11580
rect 5868 11568 5874 11620
rect 7834 11568 7840 11620
rect 7892 11608 7898 11620
rect 8754 11608 8760 11620
rect 7892 11580 8760 11608
rect 7892 11568 7898 11580
rect 8754 11568 8760 11580
rect 8812 11568 8818 11620
rect 3786 11540 3792 11552
rect 3747 11512 3792 11540
rect 3786 11500 3792 11512
rect 3844 11500 3850 11552
rect 3881 11543 3939 11549
rect 3881 11509 3893 11543
rect 3927 11540 3939 11543
rect 4154 11540 4160 11552
rect 3927 11512 4160 11540
rect 3927 11509 3939 11512
rect 3881 11503 3939 11509
rect 4154 11500 4160 11512
rect 4212 11500 4218 11552
rect 4614 11540 4620 11552
rect 4575 11512 4620 11540
rect 4614 11500 4620 11512
rect 4672 11500 4678 11552
rect 4709 11543 4767 11549
rect 4709 11509 4721 11543
rect 4755 11540 4767 11543
rect 4798 11540 4804 11552
rect 4755 11512 4804 11540
rect 4755 11509 4767 11512
rect 4709 11503 4767 11509
rect 4798 11500 4804 11512
rect 4856 11500 4862 11552
rect 5074 11540 5080 11552
rect 5035 11512 5080 11540
rect 5074 11500 5080 11512
rect 5132 11500 5138 11552
rect 6178 11500 6184 11552
rect 6236 11540 6242 11552
rect 6638 11540 6644 11552
rect 6236 11512 6644 11540
rect 6236 11500 6242 11512
rect 6638 11500 6644 11512
rect 6696 11500 6702 11552
rect 7466 11540 7472 11552
rect 7427 11512 7472 11540
rect 7466 11500 7472 11512
rect 7524 11500 7530 11552
rect 7929 11543 7987 11549
rect 7929 11509 7941 11543
rect 7975 11540 7987 11543
rect 8202 11540 8208 11552
rect 7975 11512 8208 11540
rect 7975 11509 7987 11512
rect 7929 11503 7987 11509
rect 8202 11500 8208 11512
rect 8260 11500 8266 11552
rect 8294 11500 8300 11552
rect 8352 11540 8358 11552
rect 8956 11540 8984 11648
rect 9048 11608 9076 11784
rect 9232 11784 10048 11812
rect 9232 11744 9260 11784
rect 10042 11772 10048 11784
rect 10100 11772 10106 11824
rect 9140 11716 9260 11744
rect 9401 11747 9459 11753
rect 9140 11685 9168 11716
rect 9401 11713 9413 11747
rect 9447 11744 9459 11747
rect 9490 11744 9496 11756
rect 9447 11716 9496 11744
rect 9447 11713 9459 11716
rect 9401 11707 9459 11713
rect 9490 11704 9496 11716
rect 9548 11704 9554 11756
rect 9766 11704 9772 11756
rect 9824 11744 9830 11756
rect 10336 11753 10364 11852
rect 10502 11840 10508 11852
rect 10560 11840 10566 11892
rect 10686 11840 10692 11892
rect 10744 11880 10750 11892
rect 11054 11880 11060 11892
rect 10744 11852 11060 11880
rect 10744 11840 10750 11852
rect 11054 11840 11060 11852
rect 11112 11840 11118 11892
rect 11238 11840 11244 11892
rect 11296 11880 11302 11892
rect 12437 11883 12495 11889
rect 12437 11880 12449 11883
rect 11296 11852 12449 11880
rect 11296 11840 11302 11852
rect 12437 11849 12449 11852
rect 12483 11849 12495 11883
rect 12437 11843 12495 11849
rect 13630 11840 13636 11892
rect 13688 11880 13694 11892
rect 15194 11880 15200 11892
rect 13688 11852 15200 11880
rect 13688 11840 13694 11852
rect 15194 11840 15200 11852
rect 15252 11840 15258 11892
rect 15381 11883 15439 11889
rect 15381 11849 15393 11883
rect 15427 11880 15439 11883
rect 15654 11880 15660 11892
rect 15427 11852 15660 11880
rect 15427 11849 15439 11852
rect 15381 11843 15439 11849
rect 15654 11840 15660 11852
rect 15712 11840 15718 11892
rect 17586 11880 17592 11892
rect 16040 11852 17592 11880
rect 11422 11772 11428 11824
rect 11480 11812 11486 11824
rect 11701 11815 11759 11821
rect 11701 11812 11713 11815
rect 11480 11784 11713 11812
rect 11480 11772 11486 11784
rect 11701 11781 11713 11784
rect 11747 11812 11759 11815
rect 12526 11812 12532 11824
rect 11747 11784 12532 11812
rect 11747 11781 11759 11784
rect 11701 11775 11759 11781
rect 12526 11772 12532 11784
rect 12584 11812 12590 11824
rect 12584 11784 13032 11812
rect 12584 11772 12590 11784
rect 9953 11747 10011 11753
rect 9953 11744 9965 11747
rect 9824 11716 9965 11744
rect 9824 11704 9830 11716
rect 9953 11713 9965 11716
rect 9999 11713 10011 11747
rect 9953 11707 10011 11713
rect 10321 11747 10379 11753
rect 10321 11713 10333 11747
rect 10367 11713 10379 11747
rect 10321 11707 10379 11713
rect 12434 11704 12440 11756
rect 12492 11744 12498 11756
rect 13004 11753 13032 11784
rect 12897 11747 12955 11753
rect 12897 11744 12909 11747
rect 12492 11716 12909 11744
rect 12492 11704 12498 11716
rect 12897 11713 12909 11716
rect 12943 11713 12955 11747
rect 12897 11707 12955 11713
rect 12989 11747 13047 11753
rect 12989 11713 13001 11747
rect 13035 11713 13047 11747
rect 12989 11707 13047 11713
rect 14826 11704 14832 11756
rect 14884 11744 14890 11756
rect 15470 11744 15476 11756
rect 14884 11716 15476 11744
rect 14884 11704 14890 11716
rect 15470 11704 15476 11716
rect 15528 11744 15534 11756
rect 15654 11744 15660 11756
rect 15528 11716 15660 11744
rect 15528 11704 15534 11716
rect 15654 11704 15660 11716
rect 15712 11704 15718 11756
rect 16040 11753 16068 11852
rect 17586 11840 17592 11852
rect 17644 11840 17650 11892
rect 18141 11883 18199 11889
rect 18141 11849 18153 11883
rect 18187 11880 18199 11883
rect 19334 11880 19340 11892
rect 18187 11852 19340 11880
rect 18187 11849 18199 11852
rect 18141 11843 18199 11849
rect 19334 11840 19340 11852
rect 19392 11840 19398 11892
rect 20990 11880 20996 11892
rect 20951 11852 20996 11880
rect 20990 11840 20996 11852
rect 21048 11840 21054 11892
rect 21358 11880 21364 11892
rect 21319 11852 21364 11880
rect 21358 11840 21364 11852
rect 21416 11840 21422 11892
rect 18966 11812 18972 11824
rect 18927 11784 18972 11812
rect 18966 11772 18972 11784
rect 19024 11812 19030 11824
rect 19426 11812 19432 11824
rect 19024 11784 19432 11812
rect 19024 11772 19030 11784
rect 19426 11772 19432 11784
rect 19484 11772 19490 11824
rect 16025 11747 16083 11753
rect 16025 11713 16037 11747
rect 16071 11713 16083 11747
rect 18690 11744 18696 11756
rect 18651 11716 18696 11744
rect 16025 11707 16083 11713
rect 18690 11704 18696 11716
rect 18748 11704 18754 11756
rect 9125 11679 9183 11685
rect 9125 11645 9137 11679
rect 9171 11645 9183 11679
rect 9125 11639 9183 11645
rect 9217 11679 9275 11685
rect 9217 11645 9229 11679
rect 9263 11676 9275 11679
rect 9784 11676 9812 11704
rect 9263 11648 9812 11676
rect 10520 11648 11928 11676
rect 9263 11645 9275 11648
rect 9217 11639 9275 11645
rect 10520 11608 10548 11648
rect 9048 11580 10548 11608
rect 10588 11611 10646 11617
rect 10588 11577 10600 11611
rect 10634 11608 10646 11611
rect 11146 11608 11152 11620
rect 10634 11580 11152 11608
rect 10634 11577 10646 11580
rect 10588 11571 10646 11577
rect 11146 11568 11152 11580
rect 11204 11568 11210 11620
rect 11790 11608 11796 11620
rect 11751 11580 11796 11608
rect 11790 11568 11796 11580
rect 11848 11568 11854 11620
rect 9674 11540 9680 11552
rect 8352 11512 8397 11540
rect 8956 11512 9680 11540
rect 8352 11500 8358 11512
rect 9674 11500 9680 11512
rect 9732 11500 9738 11552
rect 9769 11543 9827 11549
rect 9769 11509 9781 11543
rect 9815 11540 9827 11543
rect 10042 11540 10048 11552
rect 9815 11512 10048 11540
rect 9815 11509 9827 11512
rect 9769 11503 9827 11509
rect 10042 11500 10048 11512
rect 10100 11540 10106 11552
rect 10318 11540 10324 11552
rect 10100 11512 10324 11540
rect 10100 11500 10106 11512
rect 10318 11500 10324 11512
rect 10376 11500 10382 11552
rect 10870 11500 10876 11552
rect 10928 11540 10934 11552
rect 11422 11540 11428 11552
rect 10928 11512 11428 11540
rect 10928 11500 10934 11512
rect 11422 11500 11428 11512
rect 11480 11500 11486 11552
rect 11900 11540 11928 11648
rect 11974 11636 11980 11688
rect 12032 11676 12038 11688
rect 13265 11679 13323 11685
rect 13265 11676 13277 11679
rect 12032 11648 13277 11676
rect 12032 11636 12038 11648
rect 13265 11645 13277 11648
rect 13311 11676 13323 11679
rect 13354 11676 13360 11688
rect 13311 11648 13360 11676
rect 13311 11645 13323 11648
rect 13265 11639 13323 11645
rect 13354 11636 13360 11648
rect 13412 11636 13418 11688
rect 13449 11679 13507 11685
rect 13449 11645 13461 11679
rect 13495 11676 13507 11679
rect 15286 11676 15292 11688
rect 13495 11648 15292 11676
rect 13495 11645 13507 11648
rect 13449 11639 13507 11645
rect 15286 11636 15292 11648
rect 15344 11676 15350 11688
rect 16209 11679 16267 11685
rect 16209 11676 16221 11679
rect 15344 11648 16221 11676
rect 15344 11636 15350 11648
rect 16209 11645 16221 11648
rect 16255 11645 16267 11679
rect 16209 11639 16267 11645
rect 20530 11636 20536 11688
rect 20588 11676 20594 11688
rect 20809 11679 20867 11685
rect 20809 11676 20821 11679
rect 20588 11648 20821 11676
rect 20588 11636 20594 11648
rect 20809 11645 20821 11648
rect 20855 11645 20867 11679
rect 21174 11676 21180 11688
rect 21135 11648 21180 11676
rect 20809 11639 20867 11645
rect 21174 11636 21180 11648
rect 21232 11636 21238 11688
rect 12161 11611 12219 11617
rect 12161 11577 12173 11611
rect 12207 11608 12219 11611
rect 12434 11608 12440 11620
rect 12207 11580 12440 11608
rect 12207 11577 12219 11580
rect 12161 11571 12219 11577
rect 12434 11568 12440 11580
rect 12492 11568 12498 11620
rect 13538 11608 13544 11620
rect 12697 11580 13544 11608
rect 12697 11540 12725 11580
rect 13538 11568 13544 11580
rect 13596 11568 13602 11620
rect 13716 11611 13774 11617
rect 13716 11577 13728 11611
rect 13762 11608 13774 11611
rect 13906 11608 13912 11620
rect 13762 11580 13912 11608
rect 13762 11577 13774 11580
rect 13716 11571 13774 11577
rect 13906 11568 13912 11580
rect 13964 11568 13970 11620
rect 16476 11611 16534 11617
rect 16476 11577 16488 11611
rect 16522 11608 16534 11611
rect 17494 11608 17500 11620
rect 16522 11580 17500 11608
rect 16522 11577 16534 11580
rect 16476 11571 16534 11577
rect 17494 11568 17500 11580
rect 17552 11568 17558 11620
rect 18601 11611 18659 11617
rect 18601 11577 18613 11611
rect 18647 11608 18659 11611
rect 19153 11611 19211 11617
rect 19153 11608 19165 11611
rect 18647 11580 19165 11608
rect 18647 11577 18659 11580
rect 18601 11571 18659 11577
rect 19153 11577 19165 11580
rect 19199 11608 19211 11611
rect 20254 11608 20260 11620
rect 19199 11580 20260 11608
rect 19199 11577 19211 11580
rect 19153 11571 19211 11577
rect 20254 11568 20260 11580
rect 20312 11568 20318 11620
rect 12802 11540 12808 11552
rect 11900 11512 12725 11540
rect 12763 11512 12808 11540
rect 12802 11500 12808 11512
rect 12860 11500 12866 11552
rect 14182 11500 14188 11552
rect 14240 11540 14246 11552
rect 14829 11543 14887 11549
rect 14829 11540 14841 11543
rect 14240 11512 14841 11540
rect 14240 11500 14246 11512
rect 14829 11509 14841 11512
rect 14875 11509 14887 11543
rect 14829 11503 14887 11509
rect 15013 11543 15071 11549
rect 15013 11509 15025 11543
rect 15059 11540 15071 11543
rect 15194 11540 15200 11552
rect 15059 11512 15200 11540
rect 15059 11509 15071 11512
rect 15013 11503 15071 11509
rect 15194 11500 15200 11512
rect 15252 11500 15258 11552
rect 15746 11540 15752 11552
rect 15707 11512 15752 11540
rect 15746 11500 15752 11512
rect 15804 11500 15810 11552
rect 15841 11543 15899 11549
rect 15841 11509 15853 11543
rect 15887 11540 15899 11543
rect 16942 11540 16948 11552
rect 15887 11512 16948 11540
rect 15887 11509 15899 11512
rect 15841 11503 15899 11509
rect 16942 11500 16948 11512
rect 17000 11500 17006 11552
rect 17770 11540 17776 11552
rect 17731 11512 17776 11540
rect 17770 11500 17776 11512
rect 17828 11540 17834 11552
rect 18509 11543 18567 11549
rect 18509 11540 18521 11543
rect 17828 11512 18521 11540
rect 17828 11500 17834 11512
rect 18509 11509 18521 11512
rect 18555 11509 18567 11543
rect 18509 11503 18567 11509
rect 1104 11450 21896 11472
rect 1104 11398 7912 11450
rect 7964 11398 7976 11450
rect 8028 11398 8040 11450
rect 8092 11398 8104 11450
rect 8156 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 15035 11450
rect 15087 11398 21896 11450
rect 1104 11376 21896 11398
rect 1578 11336 1584 11348
rect 1539 11308 1584 11336
rect 1578 11296 1584 11308
rect 1636 11296 1642 11348
rect 2682 11296 2688 11348
rect 2740 11336 2746 11348
rect 3145 11339 3203 11345
rect 3145 11336 3157 11339
rect 2740 11308 3157 11336
rect 2740 11296 2746 11308
rect 3145 11305 3157 11308
rect 3191 11305 3203 11339
rect 3145 11299 3203 11305
rect 4157 11339 4215 11345
rect 4157 11305 4169 11339
rect 4203 11336 4215 11339
rect 4614 11336 4620 11348
rect 4203 11308 4620 11336
rect 4203 11305 4215 11308
rect 4157 11299 4215 11305
rect 4614 11296 4620 11308
rect 4672 11296 4678 11348
rect 4982 11336 4988 11348
rect 4943 11308 4988 11336
rect 4982 11296 4988 11308
rect 5040 11296 5046 11348
rect 6454 11296 6460 11348
rect 6512 11336 6518 11348
rect 6549 11339 6607 11345
rect 6549 11336 6561 11339
rect 6512 11308 6561 11336
rect 6512 11296 6518 11308
rect 6549 11305 6561 11308
rect 6595 11305 6607 11339
rect 6549 11299 6607 11305
rect 6638 11296 6644 11348
rect 6696 11336 6702 11348
rect 7377 11339 7435 11345
rect 7377 11336 7389 11339
rect 6696 11308 7389 11336
rect 6696 11296 6702 11308
rect 3418 11228 3424 11280
rect 3476 11268 3482 11280
rect 5629 11271 5687 11277
rect 3476 11240 4844 11268
rect 3476 11228 3482 11240
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11200 1455 11203
rect 1670 11200 1676 11212
rect 1443 11172 1676 11200
rect 1443 11169 1455 11172
rect 1397 11163 1455 11169
rect 1670 11160 1676 11172
rect 1728 11160 1734 11212
rect 1765 11203 1823 11209
rect 1765 11169 1777 11203
rect 1811 11200 1823 11203
rect 1854 11200 1860 11212
rect 1811 11172 1860 11200
rect 1811 11169 1823 11172
rect 1765 11163 1823 11169
rect 1854 11160 1860 11172
rect 1912 11160 1918 11212
rect 2032 11203 2090 11209
rect 2032 11169 2044 11203
rect 2078 11200 2090 11203
rect 2866 11200 2872 11212
rect 2078 11172 2872 11200
rect 2078 11169 2090 11172
rect 2032 11163 2090 11169
rect 2866 11160 2872 11172
rect 2924 11200 2930 11212
rect 3694 11200 3700 11212
rect 2924 11172 3700 11200
rect 2924 11160 2930 11172
rect 3694 11160 3700 11172
rect 3752 11160 3758 11212
rect 4525 11203 4583 11209
rect 4525 11169 4537 11203
rect 4571 11169 4583 11203
rect 4525 11163 4583 11169
rect 4617 11203 4675 11209
rect 4617 11169 4629 11203
rect 4663 11200 4675 11203
rect 4706 11200 4712 11212
rect 4663 11172 4712 11200
rect 4663 11169 4675 11172
rect 4617 11163 4675 11169
rect 3234 11092 3240 11144
rect 3292 11132 3298 11144
rect 3789 11135 3847 11141
rect 3789 11132 3801 11135
rect 3292 11104 3801 11132
rect 3292 11092 3298 11104
rect 3789 11101 3801 11104
rect 3835 11132 3847 11135
rect 3970 11132 3976 11144
rect 3835 11104 3976 11132
rect 3835 11101 3847 11104
rect 3789 11095 3847 11101
rect 3970 11092 3976 11104
rect 4028 11132 4034 11144
rect 4540 11132 4568 11163
rect 4706 11160 4712 11172
rect 4764 11160 4770 11212
rect 4816 11200 4844 11240
rect 5629 11237 5641 11271
rect 5675 11268 5687 11271
rect 6917 11271 6975 11277
rect 6917 11268 6929 11271
rect 5675 11240 6929 11268
rect 5675 11237 5687 11240
rect 5629 11231 5687 11237
rect 6917 11237 6929 11240
rect 6963 11237 6975 11271
rect 6917 11231 6975 11237
rect 5534 11200 5540 11212
rect 4816 11172 5540 11200
rect 5534 11160 5540 11172
rect 5592 11200 5598 11212
rect 6457 11203 6515 11209
rect 6457 11200 6469 11203
rect 5592 11172 6469 11200
rect 5592 11160 5598 11172
rect 6457 11169 6469 11172
rect 6503 11169 6515 11203
rect 6457 11163 6515 11169
rect 4028 11104 4568 11132
rect 4801 11135 4859 11141
rect 4028 11092 4034 11104
rect 4801 11101 4813 11135
rect 4847 11132 4859 11135
rect 4982 11132 4988 11144
rect 4847 11104 4988 11132
rect 4847 11101 4859 11104
rect 4801 11095 4859 11101
rect 4982 11092 4988 11104
rect 5040 11092 5046 11144
rect 5721 11135 5779 11141
rect 5721 11132 5733 11135
rect 5092 11104 5733 11132
rect 3142 11024 3148 11076
rect 3200 11064 3206 11076
rect 3697 11067 3755 11073
rect 3697 11064 3709 11067
rect 3200 11036 3709 11064
rect 3200 11024 3206 11036
rect 3697 11033 3709 11036
rect 3743 11064 3755 11067
rect 5092 11064 5120 11104
rect 5721 11101 5733 11104
rect 5767 11101 5779 11135
rect 5721 11095 5779 11101
rect 5905 11135 5963 11141
rect 5905 11101 5917 11135
rect 5951 11132 5963 11135
rect 6086 11132 6092 11144
rect 5951 11104 6092 11132
rect 5951 11101 5963 11104
rect 5905 11095 5963 11101
rect 6086 11092 6092 11104
rect 6144 11092 6150 11144
rect 6641 11135 6699 11141
rect 6641 11101 6653 11135
rect 6687 11101 6699 11135
rect 6641 11095 6699 11101
rect 3743 11036 5120 11064
rect 5261 11067 5319 11073
rect 3743 11033 3755 11036
rect 3697 11027 3755 11033
rect 5261 11033 5273 11067
rect 5307 11064 5319 11067
rect 5994 11064 6000 11076
rect 5307 11036 6000 11064
rect 5307 11033 5319 11036
rect 5261 11027 5319 11033
rect 5994 11024 6000 11036
rect 6052 11024 6058 11076
rect 6104 11064 6132 11092
rect 6656 11064 6684 11095
rect 6104 11036 6684 11064
rect 6086 10996 6092 11008
rect 6047 10968 6092 10996
rect 6086 10956 6092 10968
rect 6144 10956 6150 11008
rect 7116 10996 7144 11308
rect 7377 11305 7389 11308
rect 7423 11305 7435 11339
rect 7377 11299 7435 11305
rect 7466 11296 7472 11348
rect 7524 11336 7530 11348
rect 7929 11339 7987 11345
rect 7929 11336 7941 11339
rect 7524 11308 7941 11336
rect 7524 11296 7530 11308
rect 7929 11305 7941 11308
rect 7975 11305 7987 11339
rect 7929 11299 7987 11305
rect 8202 11296 8208 11348
rect 8260 11336 8266 11348
rect 8389 11339 8447 11345
rect 8389 11336 8401 11339
rect 8260 11308 8401 11336
rect 8260 11296 8266 11308
rect 8389 11305 8401 11308
rect 8435 11305 8447 11339
rect 8389 11299 8447 11305
rect 8938 11296 8944 11348
rect 8996 11336 9002 11348
rect 9950 11336 9956 11348
rect 8996 11308 9956 11336
rect 8996 11296 9002 11308
rect 9950 11296 9956 11308
rect 10008 11296 10014 11348
rect 10594 11296 10600 11348
rect 10652 11336 10658 11348
rect 12253 11339 12311 11345
rect 12253 11336 12265 11339
rect 10652 11308 12265 11336
rect 10652 11296 10658 11308
rect 12253 11305 12265 11308
rect 12299 11305 12311 11339
rect 12253 11299 12311 11305
rect 12526 11296 12532 11348
rect 12584 11336 12590 11348
rect 12802 11336 12808 11348
rect 12584 11308 12808 11336
rect 12584 11296 12590 11308
rect 12802 11296 12808 11308
rect 12860 11296 12866 11348
rect 13081 11339 13139 11345
rect 13081 11305 13093 11339
rect 13127 11336 13139 11339
rect 14090 11336 14096 11348
rect 13127 11308 14096 11336
rect 13127 11305 13139 11308
rect 13081 11299 13139 11305
rect 14090 11296 14096 11308
rect 14148 11296 14154 11348
rect 14369 11339 14427 11345
rect 14369 11305 14381 11339
rect 14415 11336 14427 11339
rect 15657 11339 15715 11345
rect 15657 11336 15669 11339
rect 14415 11308 15669 11336
rect 14415 11305 14427 11308
rect 14369 11299 14427 11305
rect 15657 11305 15669 11308
rect 15703 11305 15715 11339
rect 15657 11299 15715 11305
rect 16117 11339 16175 11345
rect 16117 11305 16129 11339
rect 16163 11336 16175 11339
rect 17405 11339 17463 11345
rect 17405 11336 17417 11339
rect 16163 11308 17417 11336
rect 16163 11305 16175 11308
rect 16117 11299 16175 11305
rect 17405 11305 17417 11308
rect 17451 11305 17463 11339
rect 17405 11299 17463 11305
rect 17865 11339 17923 11345
rect 17865 11305 17877 11339
rect 17911 11336 17923 11339
rect 19061 11339 19119 11345
rect 19061 11336 19073 11339
rect 17911 11308 19073 11336
rect 17911 11305 17923 11308
rect 17865 11299 17923 11305
rect 19061 11305 19073 11308
rect 19107 11305 19119 11339
rect 19061 11299 19119 11305
rect 21085 11339 21143 11345
rect 21085 11305 21097 11339
rect 21131 11336 21143 11339
rect 22005 11339 22063 11345
rect 22005 11336 22017 11339
rect 21131 11308 22017 11336
rect 21131 11305 21143 11308
rect 21085 11299 21143 11305
rect 22005 11305 22017 11308
rect 22051 11305 22063 11339
rect 22005 11299 22063 11305
rect 10134 11268 10140 11280
rect 8312 11240 10140 11268
rect 7285 11203 7343 11209
rect 7285 11169 7297 11203
rect 7331 11200 7343 11203
rect 7466 11200 7472 11212
rect 7331 11172 7472 11200
rect 7331 11169 7343 11172
rect 7285 11163 7343 11169
rect 7466 11160 7472 11172
rect 7524 11160 7530 11212
rect 8312 11209 8340 11240
rect 10134 11228 10140 11240
rect 10192 11228 10198 11280
rect 10413 11271 10471 11277
rect 10413 11237 10425 11271
rect 10459 11268 10471 11271
rect 10502 11268 10508 11280
rect 10459 11240 10508 11268
rect 10459 11237 10471 11240
rect 10413 11231 10471 11237
rect 10502 11228 10508 11240
rect 10560 11228 10566 11280
rect 12713 11271 12771 11277
rect 12713 11268 12725 11271
rect 10603 11240 12725 11268
rect 8297 11203 8355 11209
rect 8297 11200 8309 11203
rect 7576 11172 8309 11200
rect 7576 11144 7604 11172
rect 8297 11169 8309 11172
rect 8343 11169 8355 11203
rect 8297 11163 8355 11169
rect 8941 11203 8999 11209
rect 8941 11169 8953 11203
rect 8987 11169 8999 11203
rect 9766 11200 9772 11212
rect 9727 11172 9772 11200
rect 8941 11163 8999 11169
rect 7558 11132 7564 11144
rect 7519 11104 7564 11132
rect 7558 11092 7564 11104
rect 7616 11092 7622 11144
rect 8573 11135 8631 11141
rect 8573 11101 8585 11135
rect 8619 11132 8631 11135
rect 8662 11132 8668 11144
rect 8619 11104 8668 11132
rect 8619 11101 8631 11104
rect 8573 11095 8631 11101
rect 8662 11092 8668 11104
rect 8720 11092 8726 11144
rect 7374 11024 7380 11076
rect 7432 11064 7438 11076
rect 8757 11067 8815 11073
rect 8757 11064 8769 11067
rect 7432 11036 8769 11064
rect 7432 11024 7438 11036
rect 8757 11033 8769 11036
rect 8803 11033 8815 11067
rect 8956 11064 8984 11163
rect 9766 11160 9772 11172
rect 9824 11160 9830 11212
rect 9490 11132 9496 11144
rect 9451 11104 9496 11132
rect 9490 11092 9496 11104
rect 9548 11092 9554 11144
rect 9674 11092 9680 11144
rect 9732 11132 9738 11144
rect 10603 11132 10631 11240
rect 12268 11212 12296 11240
rect 12713 11237 12725 11240
rect 12759 11268 12771 11271
rect 13449 11271 13507 11277
rect 12759 11240 13400 11268
rect 12759 11237 12771 11240
rect 12713 11231 12771 11237
rect 12250 11160 12256 11212
rect 12308 11160 12314 11212
rect 12434 11160 12440 11212
rect 12492 11200 12498 11212
rect 12621 11203 12679 11209
rect 12621 11200 12633 11203
rect 12492 11172 12633 11200
rect 12492 11160 12498 11172
rect 12621 11169 12633 11172
rect 12667 11169 12679 11203
rect 12621 11163 12679 11169
rect 13265 11203 13323 11209
rect 13265 11169 13277 11203
rect 13311 11169 13323 11203
rect 13372 11200 13400 11240
rect 13449 11237 13461 11271
rect 13495 11268 13507 11271
rect 13538 11268 13544 11280
rect 13495 11240 13544 11268
rect 13495 11237 13507 11240
rect 13449 11231 13507 11237
rect 13538 11228 13544 11240
rect 13596 11268 13602 11280
rect 13909 11271 13967 11277
rect 13909 11268 13921 11271
rect 13596 11240 13921 11268
rect 13596 11228 13602 11240
rect 13909 11237 13921 11240
rect 13955 11268 13967 11271
rect 13998 11268 14004 11280
rect 13955 11240 14004 11268
rect 13955 11237 13967 11240
rect 13909 11231 13967 11237
rect 13998 11228 14004 11240
rect 14056 11228 14062 11280
rect 14642 11228 14648 11280
rect 14700 11268 14706 11280
rect 14829 11271 14887 11277
rect 14829 11268 14841 11271
rect 14700 11240 14841 11268
rect 14700 11228 14706 11240
rect 14829 11237 14841 11240
rect 14875 11237 14887 11271
rect 14829 11231 14887 11237
rect 15746 11228 15752 11280
rect 15804 11268 15810 11280
rect 17773 11271 17831 11277
rect 17773 11268 17785 11271
rect 15804 11240 17785 11268
rect 15804 11228 15810 11240
rect 17773 11237 17785 11240
rect 17819 11237 17831 11271
rect 17773 11231 17831 11237
rect 18138 11228 18144 11280
rect 18196 11268 18202 11280
rect 18325 11271 18383 11277
rect 18325 11268 18337 11271
rect 18196 11240 18337 11268
rect 18196 11228 18202 11240
rect 18325 11237 18337 11240
rect 18371 11237 18383 11271
rect 18325 11231 18383 11237
rect 18432 11240 19288 11268
rect 13814 11200 13820 11212
rect 13372 11172 13820 11200
rect 13265 11163 13323 11169
rect 9732 11104 10631 11132
rect 9732 11092 9738 11104
rect 11146 11092 11152 11144
rect 11204 11132 11210 11144
rect 12805 11135 12863 11141
rect 12805 11132 12817 11135
rect 11204 11104 12817 11132
rect 11204 11092 11210 11104
rect 12805 11101 12817 11104
rect 12851 11101 12863 11135
rect 12805 11095 12863 11101
rect 11701 11067 11759 11073
rect 11701 11064 11713 11067
rect 8956 11036 11713 11064
rect 8757 11027 8815 11033
rect 11701 11033 11713 11036
rect 11747 11064 11759 11067
rect 13280 11064 13308 11163
rect 13814 11160 13820 11172
rect 13872 11160 13878 11212
rect 14734 11200 14740 11212
rect 14695 11172 14740 11200
rect 14734 11160 14740 11172
rect 14792 11160 14798 11212
rect 15102 11160 15108 11212
rect 15160 11200 15166 11212
rect 16485 11203 16543 11209
rect 15160 11172 15792 11200
rect 15160 11160 15166 11172
rect 13354 11092 13360 11144
rect 13412 11132 13418 11144
rect 14001 11135 14059 11141
rect 14001 11132 14013 11135
rect 13412 11104 14013 11132
rect 13412 11092 13418 11104
rect 14001 11101 14013 11104
rect 14047 11101 14059 11135
rect 14182 11132 14188 11144
rect 14143 11104 14188 11132
rect 14001 11095 14059 11101
rect 14182 11092 14188 11104
rect 14240 11132 14246 11144
rect 15764 11141 15792 11172
rect 16485 11169 16497 11203
rect 16531 11200 16543 11203
rect 17126 11200 17132 11212
rect 16531 11172 17132 11200
rect 16531 11169 16543 11172
rect 16485 11163 16543 11169
rect 17126 11160 17132 11172
rect 17184 11160 17190 11212
rect 17310 11200 17316 11212
rect 17271 11172 17316 11200
rect 17310 11160 17316 11172
rect 17368 11160 17374 11212
rect 18230 11200 18236 11212
rect 18191 11172 18236 11200
rect 18230 11160 18236 11172
rect 18288 11160 18294 11212
rect 14921 11135 14979 11141
rect 14921 11132 14933 11135
rect 14240 11104 14933 11132
rect 14240 11092 14246 11104
rect 14921 11101 14933 11104
rect 14967 11101 14979 11135
rect 14921 11095 14979 11101
rect 15749 11135 15807 11141
rect 15749 11101 15761 11135
rect 15795 11101 15807 11135
rect 15930 11132 15936 11144
rect 15891 11104 15936 11132
rect 15749 11095 15807 11101
rect 15930 11092 15936 11104
rect 15988 11092 15994 11144
rect 16114 11092 16120 11144
rect 16172 11132 16178 11144
rect 16577 11135 16635 11141
rect 16577 11132 16589 11135
rect 16172 11104 16589 11132
rect 16172 11092 16178 11104
rect 16577 11101 16589 11104
rect 16623 11101 16635 11135
rect 16577 11095 16635 11101
rect 16761 11135 16819 11141
rect 16761 11101 16773 11135
rect 16807 11132 16819 11135
rect 17589 11135 17647 11141
rect 17589 11132 17601 11135
rect 16807 11104 17448 11132
rect 16807 11101 16819 11104
rect 16761 11095 16819 11101
rect 11747 11036 13308 11064
rect 13541 11067 13599 11073
rect 11747 11033 11759 11036
rect 11701 11027 11759 11033
rect 13541 11033 13553 11067
rect 13587 11064 13599 11067
rect 15102 11064 15108 11076
rect 13587 11036 15108 11064
rect 13587 11033 13599 11036
rect 13541 11027 13599 11033
rect 15102 11024 15108 11036
rect 15160 11024 15166 11076
rect 15286 11064 15292 11076
rect 15247 11036 15292 11064
rect 15286 11024 15292 11036
rect 15344 11024 15350 11076
rect 16206 11024 16212 11076
rect 16264 11064 16270 11076
rect 16776 11064 16804 11095
rect 16942 11064 16948 11076
rect 16264 11036 16804 11064
rect 16903 11036 16948 11064
rect 16264 11024 16270 11036
rect 16942 11024 16948 11036
rect 17000 11024 17006 11076
rect 7650 10996 7656 11008
rect 7116 10968 7656 10996
rect 7650 10956 7656 10968
rect 7708 10956 7714 11008
rect 7837 10999 7895 11005
rect 7837 10965 7849 10999
rect 7883 10996 7895 10999
rect 7926 10996 7932 11008
rect 7883 10968 7932 10996
rect 7883 10965 7895 10968
rect 7837 10959 7895 10965
rect 7926 10956 7932 10968
rect 7984 10996 7990 11008
rect 8294 10996 8300 11008
rect 7984 10968 8300 10996
rect 7984 10956 7990 10968
rect 8294 10956 8300 10968
rect 8352 10956 8358 11008
rect 8662 10956 8668 11008
rect 8720 10996 8726 11008
rect 9033 10999 9091 11005
rect 9033 10996 9045 10999
rect 8720 10968 9045 10996
rect 8720 10956 8726 10968
rect 9033 10965 9045 10968
rect 9079 10965 9091 10999
rect 9214 10996 9220 11008
rect 9175 10968 9220 10996
rect 9033 10959 9091 10965
rect 9214 10956 9220 10968
rect 9272 10996 9278 11008
rect 16758 10996 16764 11008
rect 9272 10968 16764 10996
rect 9272 10956 9278 10968
rect 16758 10956 16764 10968
rect 16816 10956 16822 11008
rect 17420 10996 17448 11104
rect 17512 11104 17601 11132
rect 17512 11076 17540 11104
rect 17589 11101 17601 11104
rect 17635 11132 17647 11135
rect 18432 11132 18460 11240
rect 17635 11104 18460 11132
rect 18509 11135 18567 11141
rect 17635 11101 17647 11104
rect 17589 11095 17647 11101
rect 18509 11101 18521 11135
rect 18555 11132 18567 11135
rect 18598 11132 18604 11144
rect 18555 11104 18604 11132
rect 18555 11101 18567 11104
rect 18509 11095 18567 11101
rect 18598 11092 18604 11104
rect 18656 11092 18662 11144
rect 19150 11132 19156 11144
rect 19111 11104 19156 11132
rect 19150 11092 19156 11104
rect 19208 11092 19214 11144
rect 19260 11141 19288 11240
rect 20438 11160 20444 11212
rect 20496 11200 20502 11212
rect 20901 11203 20959 11209
rect 20901 11200 20913 11203
rect 20496 11172 20913 11200
rect 20496 11160 20502 11172
rect 20901 11169 20913 11172
rect 20947 11169 20959 11203
rect 20901 11163 20959 11169
rect 19245 11135 19303 11141
rect 19245 11101 19257 11135
rect 19291 11101 19303 11135
rect 19245 11095 19303 11101
rect 17494 11024 17500 11076
rect 17552 11024 17558 11076
rect 17773 11067 17831 11073
rect 17773 11033 17785 11067
rect 17819 11064 17831 11067
rect 18693 11067 18751 11073
rect 18693 11064 18705 11067
rect 17819 11036 18705 11064
rect 17819 11033 17831 11036
rect 17773 11027 17831 11033
rect 18693 11033 18705 11036
rect 18739 11033 18751 11067
rect 18693 11027 18751 11033
rect 18598 10996 18604 11008
rect 17420 10968 18604 10996
rect 18598 10956 18604 10968
rect 18656 10956 18662 11008
rect 1104 10906 21896 10928
rect 1104 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 4575 10906
rect 4627 10854 4639 10906
rect 4691 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 18308 10906
rect 18360 10854 18372 10906
rect 18424 10854 18436 10906
rect 18488 10854 18500 10906
rect 18552 10854 21896 10906
rect 1104 10832 21896 10854
rect 1489 10795 1547 10801
rect 1489 10761 1501 10795
rect 1535 10792 1547 10795
rect 2222 10792 2228 10804
rect 1535 10764 2228 10792
rect 1535 10761 1547 10764
rect 1489 10755 1547 10761
rect 2222 10752 2228 10764
rect 2280 10752 2286 10804
rect 3694 10792 3700 10804
rect 3655 10764 3700 10792
rect 3694 10752 3700 10764
rect 3752 10752 3758 10804
rect 3786 10752 3792 10804
rect 3844 10792 3850 10804
rect 3881 10795 3939 10801
rect 3881 10792 3893 10795
rect 3844 10764 3893 10792
rect 3844 10752 3850 10764
rect 3881 10761 3893 10764
rect 3927 10761 3939 10795
rect 3881 10755 3939 10761
rect 4709 10795 4767 10801
rect 4709 10761 4721 10795
rect 4755 10792 4767 10795
rect 4798 10792 4804 10804
rect 4755 10764 4804 10792
rect 4755 10761 4767 10764
rect 4709 10755 4767 10761
rect 4798 10752 4804 10764
rect 4856 10752 4862 10804
rect 5074 10752 5080 10804
rect 5132 10792 5138 10804
rect 5626 10792 5632 10804
rect 5132 10764 5632 10792
rect 5132 10752 5138 10764
rect 5626 10752 5632 10764
rect 5684 10752 5690 10804
rect 5721 10795 5779 10801
rect 5721 10761 5733 10795
rect 5767 10792 5779 10795
rect 6270 10792 6276 10804
rect 5767 10764 6276 10792
rect 5767 10761 5779 10764
rect 5721 10755 5779 10761
rect 6270 10752 6276 10764
rect 6328 10752 6334 10804
rect 7006 10752 7012 10804
rect 7064 10792 7070 10804
rect 8297 10795 8355 10801
rect 8297 10792 8309 10795
rect 7064 10764 8309 10792
rect 7064 10752 7070 10764
rect 8297 10761 8309 10764
rect 8343 10761 8355 10795
rect 8297 10755 8355 10761
rect 8662 10752 8668 10804
rect 8720 10792 8726 10804
rect 9674 10792 9680 10804
rect 8720 10764 9680 10792
rect 8720 10752 8726 10764
rect 9674 10752 9680 10764
rect 9732 10792 9738 10804
rect 10962 10792 10968 10804
rect 9732 10764 10968 10792
rect 9732 10752 9738 10764
rect 10962 10752 10968 10764
rect 11020 10752 11026 10804
rect 11146 10752 11152 10804
rect 11204 10792 11210 10804
rect 11333 10795 11391 10801
rect 11333 10792 11345 10795
rect 11204 10764 11345 10792
rect 11204 10752 11210 10764
rect 11333 10761 11345 10764
rect 11379 10761 11391 10795
rect 11333 10755 11391 10761
rect 11425 10795 11483 10801
rect 11425 10761 11437 10795
rect 11471 10792 11483 10795
rect 12526 10792 12532 10804
rect 11471 10764 12532 10792
rect 11471 10761 11483 10764
rect 11425 10755 11483 10761
rect 8205 10727 8263 10733
rect 8205 10693 8217 10727
rect 8251 10724 8263 10727
rect 8251 10696 8285 10724
rect 8251 10693 8263 10696
rect 8205 10687 8263 10693
rect 2130 10656 2136 10668
rect 2091 10628 2136 10656
rect 2130 10616 2136 10628
rect 2188 10616 2194 10668
rect 4338 10656 4344 10668
rect 4299 10628 4344 10656
rect 4338 10616 4344 10628
rect 4396 10616 4402 10668
rect 4525 10659 4583 10665
rect 4525 10625 4537 10659
rect 4571 10656 4583 10659
rect 4982 10656 4988 10668
rect 4571 10628 4988 10656
rect 4571 10625 4583 10628
rect 4525 10619 4583 10625
rect 4982 10616 4988 10628
rect 5040 10656 5046 10668
rect 5353 10659 5411 10665
rect 5353 10656 5365 10659
rect 5040 10628 5365 10656
rect 5040 10616 5046 10628
rect 5353 10625 5365 10628
rect 5399 10656 5411 10659
rect 5442 10656 5448 10668
rect 5399 10628 5448 10656
rect 5399 10625 5411 10628
rect 5353 10619 5411 10625
rect 5442 10616 5448 10628
rect 5500 10616 5506 10668
rect 5629 10659 5687 10665
rect 5629 10625 5641 10659
rect 5675 10656 5687 10659
rect 5718 10656 5724 10668
rect 5675 10628 5724 10656
rect 5675 10625 5687 10628
rect 5629 10619 5687 10625
rect 2317 10591 2375 10597
rect 2317 10557 2329 10591
rect 2363 10588 2375 10591
rect 3878 10588 3884 10600
rect 2363 10560 3884 10588
rect 2363 10557 2375 10560
rect 2317 10551 2375 10557
rect 3878 10548 3884 10560
rect 3936 10548 3942 10600
rect 4249 10591 4307 10597
rect 4249 10557 4261 10591
rect 4295 10588 4307 10591
rect 5644 10588 5672 10619
rect 5718 10616 5724 10628
rect 5776 10616 5782 10668
rect 6086 10616 6092 10668
rect 6144 10656 6150 10668
rect 6181 10659 6239 10665
rect 6181 10656 6193 10659
rect 6144 10628 6193 10656
rect 6144 10616 6150 10628
rect 6181 10625 6193 10628
rect 6227 10625 6239 10659
rect 6362 10656 6368 10668
rect 6323 10628 6368 10656
rect 6181 10619 6239 10625
rect 6362 10616 6368 10628
rect 6420 10616 6426 10668
rect 8220 10656 8248 10687
rect 9306 10684 9312 10736
rect 9364 10724 9370 10736
rect 9364 10696 9996 10724
rect 9364 10684 9370 10696
rect 8849 10659 8907 10665
rect 8849 10656 8861 10659
rect 8220 10628 8861 10656
rect 8220 10600 8248 10628
rect 8849 10625 8861 10628
rect 8895 10625 8907 10659
rect 8849 10619 8907 10625
rect 8938 10616 8944 10668
rect 8996 10656 9002 10668
rect 9490 10656 9496 10668
rect 8996 10628 9496 10656
rect 8996 10616 9002 10628
rect 9490 10616 9496 10628
rect 9548 10616 9554 10668
rect 9582 10616 9588 10668
rect 9640 10656 9646 10668
rect 9968 10665 9996 10696
rect 9677 10659 9735 10665
rect 9677 10656 9689 10659
rect 9640 10628 9689 10656
rect 9640 10616 9646 10628
rect 9677 10625 9689 10628
rect 9723 10625 9735 10659
rect 9677 10619 9735 10625
rect 9953 10659 10011 10665
rect 9953 10625 9965 10659
rect 9999 10625 10011 10659
rect 11348 10656 11376 10755
rect 12526 10752 12532 10764
rect 12584 10752 12590 10804
rect 13170 10752 13176 10804
rect 13228 10792 13234 10804
rect 13909 10795 13967 10801
rect 13909 10792 13921 10795
rect 13228 10764 13921 10792
rect 13228 10752 13234 10764
rect 13909 10761 13921 10764
rect 13955 10792 13967 10795
rect 15105 10795 15163 10801
rect 13955 10764 14964 10792
rect 13955 10761 13967 10764
rect 13909 10755 13967 10761
rect 11790 10684 11796 10736
rect 11848 10724 11854 10736
rect 12434 10724 12440 10736
rect 11848 10696 12440 10724
rect 11848 10684 11854 10696
rect 12434 10684 12440 10696
rect 12492 10684 12498 10736
rect 14642 10684 14648 10736
rect 14700 10724 14706 10736
rect 14829 10727 14887 10733
rect 14829 10724 14841 10727
rect 14700 10696 14841 10724
rect 14700 10684 14706 10696
rect 14829 10693 14841 10696
rect 14875 10693 14887 10727
rect 14936 10724 14964 10764
rect 15105 10761 15117 10795
rect 15151 10792 15163 10795
rect 17310 10792 17316 10804
rect 15151 10764 17316 10792
rect 15151 10761 15163 10764
rect 15105 10755 15163 10761
rect 17310 10752 17316 10764
rect 17368 10752 17374 10804
rect 17773 10795 17831 10801
rect 17773 10761 17785 10795
rect 17819 10792 17831 10795
rect 18138 10792 18144 10804
rect 17819 10764 18144 10792
rect 17819 10761 17831 10764
rect 17773 10755 17831 10761
rect 18138 10752 18144 10764
rect 18196 10752 18202 10804
rect 15930 10724 15936 10736
rect 14936 10696 15936 10724
rect 14829 10687 14887 10693
rect 15930 10684 15936 10696
rect 15988 10684 15994 10736
rect 18049 10727 18107 10733
rect 18049 10693 18061 10727
rect 18095 10724 18107 10727
rect 19150 10724 19156 10736
rect 18095 10696 19156 10724
rect 18095 10693 18107 10696
rect 18049 10687 18107 10693
rect 19150 10684 19156 10696
rect 19208 10684 19214 10736
rect 19337 10727 19395 10733
rect 19337 10693 19349 10727
rect 19383 10724 19395 10727
rect 19383 10696 20760 10724
rect 19383 10693 19395 10696
rect 19337 10687 19395 10693
rect 11977 10659 12035 10665
rect 11977 10656 11989 10659
rect 11348 10628 11989 10656
rect 9953 10619 10011 10625
rect 11977 10625 11989 10628
rect 12023 10625 12035 10659
rect 11977 10619 12035 10625
rect 12360 10628 12664 10656
rect 4295 10560 5672 10588
rect 4295 10557 4307 10560
rect 4249 10551 4307 10557
rect 5810 10548 5816 10600
rect 5868 10588 5874 10600
rect 6825 10591 6883 10597
rect 6825 10588 6837 10591
rect 5868 10560 6837 10588
rect 5868 10548 5874 10560
rect 6825 10557 6837 10560
rect 6871 10557 6883 10591
rect 6825 10551 6883 10557
rect 7466 10548 7472 10600
rect 7524 10588 7530 10600
rect 7926 10588 7932 10600
rect 7524 10560 7932 10588
rect 7524 10548 7530 10560
rect 7926 10548 7932 10560
rect 7984 10548 7990 10600
rect 8202 10548 8208 10600
rect 8260 10548 8266 10600
rect 8757 10591 8815 10597
rect 8757 10557 8769 10591
rect 8803 10588 8815 10591
rect 9766 10588 9772 10600
rect 8803 10560 9772 10588
rect 8803 10557 8815 10560
rect 8757 10551 8815 10557
rect 9766 10548 9772 10560
rect 9824 10548 9830 10600
rect 9858 10548 9864 10600
rect 9916 10588 9922 10600
rect 10209 10591 10267 10597
rect 10209 10588 10221 10591
rect 9916 10560 10221 10588
rect 9916 10548 9922 10560
rect 10209 10557 10221 10560
rect 10255 10557 10267 10591
rect 10209 10551 10267 10557
rect 11054 10548 11060 10600
rect 11112 10588 11118 10600
rect 11330 10588 11336 10600
rect 11112 10560 11336 10588
rect 11112 10548 11118 10560
rect 11330 10548 11336 10560
rect 11388 10588 11394 10600
rect 11885 10591 11943 10597
rect 11885 10588 11897 10591
rect 11388 10560 11897 10588
rect 11388 10548 11394 10560
rect 11885 10557 11897 10560
rect 11931 10588 11943 10591
rect 12360 10588 12388 10628
rect 11931 10560 12388 10588
rect 11931 10557 11943 10560
rect 11885 10551 11943 10557
rect 12434 10548 12440 10600
rect 12492 10588 12498 10600
rect 12529 10591 12587 10597
rect 12529 10588 12541 10591
rect 12492 10560 12541 10588
rect 12492 10548 12498 10560
rect 12529 10557 12541 10560
rect 12575 10557 12587 10591
rect 12636 10588 12664 10628
rect 13538 10616 13544 10668
rect 13596 10656 13602 10668
rect 14182 10656 14188 10668
rect 13596 10628 14188 10656
rect 13596 10616 13602 10628
rect 14182 10616 14188 10628
rect 14240 10656 14246 10668
rect 14553 10659 14611 10665
rect 14553 10656 14565 10659
rect 14240 10628 14565 10656
rect 14240 10616 14246 10628
rect 14553 10625 14565 10628
rect 14599 10625 14611 10659
rect 15749 10659 15807 10665
rect 14553 10619 14611 10625
rect 14660 10628 15599 10656
rect 14660 10588 14688 10628
rect 12636 10560 14688 10588
rect 12529 10551 12587 10557
rect 15194 10548 15200 10600
rect 15252 10588 15258 10600
rect 15473 10591 15531 10597
rect 15473 10588 15485 10591
rect 15252 10560 15485 10588
rect 15252 10548 15258 10560
rect 15473 10557 15485 10560
rect 15519 10557 15531 10591
rect 15473 10551 15531 10557
rect 2584 10523 2642 10529
rect 2584 10489 2596 10523
rect 2630 10520 2642 10523
rect 2682 10520 2688 10532
rect 2630 10492 2688 10520
rect 2630 10489 2642 10492
rect 2584 10483 2642 10489
rect 2682 10480 2688 10492
rect 2740 10480 2746 10532
rect 4982 10480 4988 10532
rect 5040 10520 5046 10532
rect 5169 10523 5227 10529
rect 5169 10520 5181 10523
rect 5040 10492 5181 10520
rect 5040 10480 5046 10492
rect 5169 10489 5181 10492
rect 5215 10489 5227 10523
rect 5169 10483 5227 10489
rect 1854 10452 1860 10464
rect 1815 10424 1860 10452
rect 1854 10412 1860 10424
rect 1912 10412 1918 10464
rect 1949 10455 2007 10461
rect 1949 10421 1961 10455
rect 1995 10452 2007 10455
rect 2038 10452 2044 10464
rect 1995 10424 2044 10452
rect 1995 10421 2007 10424
rect 1949 10415 2007 10421
rect 2038 10412 2044 10424
rect 2096 10412 2102 10464
rect 5074 10452 5080 10464
rect 5035 10424 5080 10452
rect 5074 10412 5080 10424
rect 5132 10412 5138 10464
rect 5184 10452 5212 10483
rect 5994 10480 6000 10532
rect 6052 10520 6058 10532
rect 6089 10523 6147 10529
rect 6089 10520 6101 10523
rect 6052 10492 6101 10520
rect 6052 10480 6058 10492
rect 6089 10489 6101 10492
rect 6135 10489 6147 10523
rect 6089 10483 6147 10489
rect 6178 10480 6184 10532
rect 6236 10520 6242 10532
rect 7070 10523 7128 10529
rect 7070 10520 7082 10523
rect 6236 10492 7082 10520
rect 6236 10480 6242 10492
rect 7070 10489 7082 10492
rect 7116 10489 7128 10523
rect 7070 10483 7128 10489
rect 8665 10523 8723 10529
rect 8665 10489 8677 10523
rect 8711 10520 8723 10523
rect 8938 10520 8944 10532
rect 8711 10492 8944 10520
rect 8711 10489 8723 10492
rect 8665 10483 8723 10489
rect 8938 10480 8944 10492
rect 8996 10480 9002 10532
rect 9493 10523 9551 10529
rect 9493 10489 9505 10523
rect 9539 10520 9551 10523
rect 10042 10520 10048 10532
rect 9539 10492 10048 10520
rect 9539 10489 9551 10492
rect 9493 10483 9551 10489
rect 10042 10480 10048 10492
rect 10100 10480 10106 10532
rect 10318 10480 10324 10532
rect 10376 10520 10382 10532
rect 11793 10523 11851 10529
rect 11793 10520 11805 10523
rect 10376 10492 11805 10520
rect 10376 10480 10382 10492
rect 11793 10489 11805 10492
rect 11839 10520 11851 10523
rect 12796 10523 12854 10529
rect 11839 10492 12664 10520
rect 11839 10489 11851 10492
rect 11793 10483 11851 10489
rect 6549 10455 6607 10461
rect 6549 10452 6561 10455
rect 5184 10424 6561 10452
rect 6549 10421 6561 10424
rect 6595 10452 6607 10455
rect 6822 10452 6828 10464
rect 6595 10424 6828 10452
rect 6595 10421 6607 10424
rect 6549 10415 6607 10421
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 7190 10412 7196 10464
rect 7248 10452 7254 10464
rect 9125 10455 9183 10461
rect 9125 10452 9137 10455
rect 7248 10424 9137 10452
rect 7248 10412 7254 10424
rect 9125 10421 9137 10424
rect 9171 10421 9183 10455
rect 9125 10415 9183 10421
rect 9585 10455 9643 10461
rect 9585 10421 9597 10455
rect 9631 10452 9643 10455
rect 9674 10452 9680 10464
rect 9631 10424 9680 10452
rect 9631 10421 9643 10424
rect 9585 10415 9643 10421
rect 9674 10412 9680 10424
rect 9732 10412 9738 10464
rect 11054 10412 11060 10464
rect 11112 10452 11118 10464
rect 11882 10452 11888 10464
rect 11112 10424 11888 10452
rect 11112 10412 11118 10424
rect 11882 10412 11888 10424
rect 11940 10412 11946 10464
rect 11974 10412 11980 10464
rect 12032 10452 12038 10464
rect 12526 10452 12532 10464
rect 12032 10424 12532 10452
rect 12032 10412 12038 10424
rect 12526 10412 12532 10424
rect 12584 10412 12590 10464
rect 12636 10452 12664 10492
rect 12796 10489 12808 10523
rect 12842 10520 12854 10523
rect 13446 10520 13452 10532
rect 12842 10492 13452 10520
rect 12842 10489 12854 10492
rect 12796 10483 12854 10489
rect 13446 10480 13452 10492
rect 13504 10480 13510 10532
rect 14369 10523 14427 10529
rect 14369 10489 14381 10523
rect 14415 10520 14427 10523
rect 15286 10520 15292 10532
rect 14415 10492 15292 10520
rect 14415 10489 14427 10492
rect 14369 10483 14427 10489
rect 15286 10480 15292 10492
rect 15344 10480 15350 10532
rect 15571 10520 15599 10628
rect 15749 10625 15761 10659
rect 15795 10656 15807 10659
rect 15795 10628 16068 10656
rect 15795 10625 15807 10628
rect 15749 10619 15807 10625
rect 15930 10588 15936 10600
rect 15891 10560 15936 10588
rect 15930 10548 15936 10560
rect 15988 10548 15994 10600
rect 16040 10588 16068 10628
rect 17862 10616 17868 10668
rect 17920 10656 17926 10668
rect 18509 10659 18567 10665
rect 18509 10656 18521 10659
rect 17920 10628 18521 10656
rect 17920 10616 17926 10628
rect 18509 10625 18521 10628
rect 18555 10625 18567 10659
rect 18690 10656 18696 10668
rect 18651 10628 18696 10656
rect 18509 10619 18567 10625
rect 16206 10597 16212 10600
rect 16200 10588 16212 10597
rect 16040 10560 16212 10588
rect 16200 10551 16212 10560
rect 16206 10548 16212 10551
rect 16264 10548 16270 10600
rect 16758 10548 16764 10600
rect 16816 10588 16822 10600
rect 17497 10591 17555 10597
rect 17497 10588 17509 10591
rect 16816 10560 17509 10588
rect 16816 10548 16822 10560
rect 17497 10557 17509 10560
rect 17543 10588 17555 10591
rect 18417 10591 18475 10597
rect 18417 10588 18429 10591
rect 17543 10560 18429 10588
rect 17543 10557 17555 10560
rect 17497 10551 17555 10557
rect 18417 10557 18429 10560
rect 18463 10557 18475 10591
rect 18524 10588 18552 10619
rect 18690 10616 18696 10628
rect 18748 10616 18754 10668
rect 18782 10616 18788 10668
rect 18840 10656 18846 10668
rect 18877 10659 18935 10665
rect 18877 10656 18889 10659
rect 18840 10628 18889 10656
rect 18840 10616 18846 10628
rect 18877 10625 18889 10628
rect 18923 10625 18935 10659
rect 19886 10656 19892 10668
rect 19847 10628 19892 10656
rect 18877 10619 18935 10625
rect 19886 10616 19892 10628
rect 19944 10616 19950 10668
rect 20438 10656 20444 10668
rect 20399 10628 20444 10656
rect 20438 10616 20444 10628
rect 20496 10616 20502 10668
rect 19153 10591 19211 10597
rect 19153 10588 19165 10591
rect 18524 10560 19165 10588
rect 18417 10551 18475 10557
rect 19153 10557 19165 10560
rect 19199 10557 19211 10591
rect 19153 10551 19211 10557
rect 18138 10520 18144 10532
rect 15571 10492 18144 10520
rect 18138 10480 18144 10492
rect 18196 10480 18202 10532
rect 18432 10520 18460 10551
rect 19426 10548 19432 10600
rect 19484 10588 19490 10600
rect 20732 10597 20760 10696
rect 20993 10659 21051 10665
rect 20993 10625 21005 10659
rect 21039 10656 21051 10659
rect 21174 10656 21180 10668
rect 21039 10628 21180 10656
rect 21039 10625 21051 10628
rect 20993 10619 21051 10625
rect 21174 10616 21180 10628
rect 21232 10616 21238 10668
rect 20165 10591 20223 10597
rect 20165 10588 20177 10591
rect 19484 10560 20177 10588
rect 19484 10548 19490 10560
rect 20165 10557 20177 10560
rect 20211 10557 20223 10591
rect 20165 10551 20223 10557
rect 20717 10591 20775 10597
rect 20717 10557 20729 10591
rect 20763 10557 20775 10591
rect 20717 10551 20775 10557
rect 20346 10520 20352 10532
rect 18432 10492 20352 10520
rect 20346 10480 20352 10492
rect 20404 10480 20410 10532
rect 13630 10452 13636 10464
rect 12636 10424 13636 10452
rect 13630 10412 13636 10424
rect 13688 10412 13694 10464
rect 13998 10452 14004 10464
rect 13959 10424 14004 10452
rect 13998 10412 14004 10424
rect 14056 10412 14062 10464
rect 14182 10412 14188 10464
rect 14240 10452 14246 10464
rect 14461 10455 14519 10461
rect 14461 10452 14473 10455
rect 14240 10424 14473 10452
rect 14240 10412 14246 10424
rect 14461 10421 14473 10424
rect 14507 10421 14519 10455
rect 14461 10415 14519 10421
rect 14734 10412 14740 10464
rect 14792 10452 14798 10464
rect 15565 10455 15623 10461
rect 15565 10452 15577 10455
rect 14792 10424 15577 10452
rect 14792 10412 14798 10424
rect 15565 10421 15577 10424
rect 15611 10421 15623 10455
rect 15565 10415 15623 10421
rect 15746 10412 15752 10464
rect 15804 10452 15810 10464
rect 16850 10452 16856 10464
rect 15804 10424 16856 10452
rect 15804 10412 15810 10424
rect 16850 10412 16856 10424
rect 16908 10412 16914 10464
rect 17313 10455 17371 10461
rect 17313 10421 17325 10455
rect 17359 10452 17371 10455
rect 17494 10452 17500 10464
rect 17359 10424 17500 10452
rect 17359 10421 17371 10424
rect 17313 10415 17371 10421
rect 17494 10412 17500 10424
rect 17552 10412 17558 10464
rect 19702 10452 19708 10464
rect 19663 10424 19708 10452
rect 19702 10412 19708 10424
rect 19760 10412 19766 10464
rect 19797 10455 19855 10461
rect 19797 10421 19809 10455
rect 19843 10452 19855 10455
rect 20438 10452 20444 10464
rect 19843 10424 20444 10452
rect 19843 10421 19855 10424
rect 19797 10415 19855 10421
rect 20438 10412 20444 10424
rect 20496 10412 20502 10464
rect 1104 10362 21896 10384
rect 1104 10310 7912 10362
rect 7964 10310 7976 10362
rect 8028 10310 8040 10362
rect 8092 10310 8104 10362
rect 8156 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 15035 10362
rect 15087 10310 21896 10362
rect 1104 10288 21896 10310
rect 2038 10248 2044 10260
rect 1999 10220 2044 10248
rect 2038 10208 2044 10220
rect 2096 10208 2102 10260
rect 3142 10248 3148 10260
rect 3103 10220 3148 10248
rect 3142 10208 3148 10220
rect 3200 10208 3206 10260
rect 4154 10208 4160 10260
rect 4212 10248 4218 10260
rect 4341 10251 4399 10257
rect 4341 10248 4353 10251
rect 4212 10220 4353 10248
rect 4212 10208 4218 10220
rect 4341 10217 4353 10220
rect 4387 10217 4399 10251
rect 4341 10211 4399 10217
rect 4890 10208 4896 10260
rect 4948 10248 4954 10260
rect 5261 10251 5319 10257
rect 5261 10248 5273 10251
rect 4948 10220 5273 10248
rect 4948 10208 4954 10220
rect 5261 10217 5273 10220
rect 5307 10217 5319 10251
rect 5261 10211 5319 10217
rect 5626 10208 5632 10260
rect 5684 10248 5690 10260
rect 6086 10248 6092 10260
rect 5684 10220 6092 10248
rect 5684 10208 5690 10220
rect 6086 10208 6092 10220
rect 6144 10208 6150 10260
rect 6733 10251 6791 10257
rect 6733 10217 6745 10251
rect 6779 10248 6791 10251
rect 7101 10251 7159 10257
rect 7101 10248 7113 10251
rect 6779 10220 7113 10248
rect 6779 10217 6791 10220
rect 6733 10211 6791 10217
rect 7101 10217 7113 10220
rect 7147 10217 7159 10251
rect 7101 10211 7159 10217
rect 8294 10208 8300 10260
rect 8352 10208 8358 10260
rect 8478 10208 8484 10260
rect 8536 10248 8542 10260
rect 11330 10248 11336 10260
rect 8536 10220 11192 10248
rect 11291 10220 11336 10248
rect 8536 10208 8542 10220
rect 4249 10183 4307 10189
rect 4249 10149 4261 10183
rect 4295 10180 4307 10183
rect 4709 10183 4767 10189
rect 4709 10180 4721 10183
rect 4295 10152 4721 10180
rect 4295 10149 4307 10152
rect 4249 10143 4307 10149
rect 4709 10149 4721 10152
rect 4755 10180 4767 10183
rect 6454 10180 6460 10192
rect 4755 10152 6460 10180
rect 4755 10149 4767 10152
rect 4709 10143 4767 10149
rect 6454 10140 6460 10152
rect 6512 10140 6518 10192
rect 6641 10183 6699 10189
rect 6641 10149 6653 10183
rect 6687 10180 6699 10183
rect 7006 10180 7012 10192
rect 6687 10152 7012 10180
rect 6687 10149 6699 10152
rect 6641 10143 6699 10149
rect 7006 10140 7012 10152
rect 7064 10140 7070 10192
rect 7190 10140 7196 10192
rect 7248 10180 7254 10192
rect 8312 10180 8340 10208
rect 8846 10180 8852 10192
rect 7248 10152 8248 10180
rect 8312 10152 8852 10180
rect 7248 10140 7254 10152
rect 2406 10112 2412 10124
rect 2367 10084 2412 10112
rect 2406 10072 2412 10084
rect 2464 10072 2470 10124
rect 3326 10072 3332 10124
rect 3384 10112 3390 10124
rect 3786 10112 3792 10124
rect 3384 10084 3792 10112
rect 3384 10072 3390 10084
rect 3786 10072 3792 10084
rect 3844 10072 3850 10124
rect 5534 10072 5540 10124
rect 5592 10112 5598 10124
rect 5629 10115 5687 10121
rect 5629 10112 5641 10115
rect 5592 10084 5641 10112
rect 5592 10072 5598 10084
rect 5629 10081 5641 10084
rect 5675 10081 5687 10115
rect 5629 10075 5687 10081
rect 5721 10115 5779 10121
rect 5721 10081 5733 10115
rect 5767 10112 5779 10115
rect 6730 10112 6736 10124
rect 5767 10084 6736 10112
rect 5767 10081 5779 10084
rect 5721 10075 5779 10081
rect 6730 10072 6736 10084
rect 6788 10072 6794 10124
rect 6914 10072 6920 10124
rect 6972 10112 6978 10124
rect 7466 10112 7472 10124
rect 6972 10084 7472 10112
rect 6972 10072 6978 10084
rect 7466 10072 7472 10084
rect 7524 10072 7530 10124
rect 7561 10115 7619 10121
rect 7561 10081 7573 10115
rect 7607 10112 7619 10115
rect 7650 10112 7656 10124
rect 7607 10084 7656 10112
rect 7607 10081 7619 10084
rect 7561 10075 7619 10081
rect 7650 10072 7656 10084
rect 7708 10072 7714 10124
rect 8220 10112 8248 10152
rect 8846 10140 8852 10152
rect 8904 10140 8910 10192
rect 9125 10183 9183 10189
rect 9125 10180 9137 10183
rect 8956 10152 9137 10180
rect 8297 10115 8355 10121
rect 8297 10112 8309 10115
rect 8220 10084 8309 10112
rect 8297 10081 8309 10084
rect 8343 10081 8355 10115
rect 8297 10075 8355 10081
rect 8754 10072 8760 10124
rect 8812 10112 8818 10124
rect 8956 10112 8984 10152
rect 9125 10149 9137 10152
rect 9171 10149 9183 10183
rect 9922 10183 9980 10189
rect 9922 10180 9934 10183
rect 9125 10143 9183 10149
rect 9416 10152 9934 10180
rect 9416 10112 9444 10152
rect 9922 10149 9934 10152
rect 9968 10180 9980 10183
rect 10134 10180 10140 10192
rect 9968 10152 10140 10180
rect 9968 10149 9980 10152
rect 9922 10143 9980 10149
rect 10134 10140 10140 10152
rect 10192 10140 10198 10192
rect 11164 10180 11192 10220
rect 11330 10208 11336 10220
rect 11388 10208 11394 10260
rect 11514 10208 11520 10260
rect 11572 10248 11578 10260
rect 11793 10251 11851 10257
rect 11793 10248 11805 10251
rect 11572 10220 11805 10248
rect 11572 10208 11578 10220
rect 11793 10217 11805 10220
rect 11839 10217 11851 10251
rect 11793 10211 11851 10217
rect 11885 10251 11943 10257
rect 11885 10217 11897 10251
rect 11931 10248 11943 10251
rect 11974 10248 11980 10260
rect 11931 10220 11980 10248
rect 11931 10217 11943 10220
rect 11885 10211 11943 10217
rect 11974 10208 11980 10220
rect 12032 10208 12038 10260
rect 12066 10208 12072 10260
rect 12124 10248 12130 10260
rect 12342 10248 12348 10260
rect 12124 10220 12348 10248
rect 12124 10208 12130 10220
rect 12342 10208 12348 10220
rect 12400 10208 12406 10260
rect 13633 10251 13691 10257
rect 13633 10217 13645 10251
rect 13679 10217 13691 10251
rect 13633 10211 13691 10217
rect 11698 10180 11704 10192
rect 11164 10152 11704 10180
rect 11698 10140 11704 10152
rect 11756 10140 11762 10192
rect 13648 10180 13676 10211
rect 13814 10208 13820 10260
rect 13872 10248 13878 10260
rect 13909 10251 13967 10257
rect 13909 10248 13921 10251
rect 13872 10220 13921 10248
rect 13872 10208 13878 10220
rect 13909 10217 13921 10220
rect 13955 10217 13967 10251
rect 13909 10211 13967 10217
rect 14182 10208 14188 10260
rect 14240 10248 14246 10260
rect 14277 10251 14335 10257
rect 14277 10248 14289 10251
rect 14240 10220 14289 10248
rect 14240 10208 14246 10220
rect 14277 10217 14289 10220
rect 14323 10217 14335 10251
rect 14642 10248 14648 10260
rect 14603 10220 14648 10248
rect 14277 10211 14335 10217
rect 14642 10208 14648 10220
rect 14700 10208 14706 10260
rect 15286 10248 15292 10260
rect 15247 10220 15292 10248
rect 15286 10208 15292 10220
rect 15344 10208 15350 10260
rect 16114 10248 16120 10260
rect 15396 10220 15884 10248
rect 16075 10220 16120 10248
rect 14737 10183 14795 10189
rect 14737 10180 14749 10183
rect 12084 10152 13676 10180
rect 14200 10152 14749 10180
rect 8812 10084 8984 10112
rect 9140 10084 9444 10112
rect 8812 10072 8818 10084
rect 2498 10044 2504 10056
rect 2459 10016 2504 10044
rect 2498 10004 2504 10016
rect 2556 10004 2562 10056
rect 2685 10047 2743 10053
rect 2685 10013 2697 10047
rect 2731 10044 2743 10047
rect 2866 10044 2872 10056
rect 2731 10016 2872 10044
rect 2731 10013 2743 10016
rect 2685 10007 2743 10013
rect 2866 10004 2872 10016
rect 2924 10004 2930 10056
rect 4798 10044 4804 10056
rect 4759 10016 4804 10044
rect 4798 10004 4804 10016
rect 4856 10004 4862 10056
rect 4985 10047 5043 10053
rect 4985 10013 4997 10047
rect 5031 10044 5043 10047
rect 5442 10044 5448 10056
rect 5031 10016 5448 10044
rect 5031 10013 5043 10016
rect 4985 10007 5043 10013
rect 5442 10004 5448 10016
rect 5500 10004 5506 10056
rect 5902 10044 5908 10056
rect 5863 10016 5908 10044
rect 5902 10004 5908 10016
rect 5960 10004 5966 10056
rect 6822 10044 6828 10056
rect 6783 10016 6828 10044
rect 6822 10004 6828 10016
rect 6880 10004 6886 10056
rect 2961 9979 3019 9985
rect 2961 9945 2973 9979
rect 3007 9976 3019 9979
rect 3326 9976 3332 9988
rect 3007 9948 3332 9976
rect 3007 9945 3019 9948
rect 2961 9939 3019 9945
rect 3326 9936 3332 9948
rect 3384 9976 3390 9988
rect 3510 9976 3516 9988
rect 3384 9948 3516 9976
rect 3384 9936 3390 9948
rect 3510 9936 3516 9948
rect 3568 9936 3574 9988
rect 7668 9976 7696 10072
rect 7742 10004 7748 10056
rect 7800 10044 7806 10056
rect 8202 10044 8208 10056
rect 7800 10016 8208 10044
rect 7800 10004 7806 10016
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 8389 10047 8447 10053
rect 8389 10013 8401 10047
rect 8435 10013 8447 10047
rect 8389 10007 8447 10013
rect 8573 10047 8631 10053
rect 8573 10013 8585 10047
rect 8619 10044 8631 10047
rect 9140 10044 9168 10084
rect 9490 10072 9496 10124
rect 9548 10112 9554 10124
rect 11882 10112 11888 10124
rect 9548 10084 11888 10112
rect 9548 10072 9554 10084
rect 11882 10072 11888 10084
rect 11940 10072 11946 10124
rect 8619 10016 9168 10044
rect 8619 10013 8631 10016
rect 8573 10007 8631 10013
rect 8294 9976 8300 9988
rect 7668 9948 8300 9976
rect 8294 9936 8300 9948
rect 8352 9936 8358 9988
rect 8404 9976 8432 10007
rect 9214 10004 9220 10056
rect 9272 10044 9278 10056
rect 9401 10047 9459 10053
rect 9272 10016 9317 10044
rect 9272 10004 9278 10016
rect 9401 10013 9413 10047
rect 9447 10044 9459 10047
rect 9582 10044 9588 10056
rect 9447 10016 9588 10044
rect 9447 10013 9459 10016
rect 9401 10007 9459 10013
rect 9582 10004 9588 10016
rect 9640 10004 9646 10056
rect 9677 10047 9735 10053
rect 9677 10013 9689 10047
rect 9723 10013 9735 10047
rect 9677 10007 9735 10013
rect 8757 9979 8815 9985
rect 8757 9976 8769 9979
rect 8404 9948 8769 9976
rect 8757 9945 8769 9948
rect 8803 9945 8815 9979
rect 8757 9939 8815 9945
rect 9306 9936 9312 9988
rect 9364 9976 9370 9988
rect 9692 9976 9720 10007
rect 11974 10004 11980 10056
rect 12032 10044 12038 10056
rect 12084 10053 12112 10152
rect 14200 10124 14228 10152
rect 14737 10149 14749 10152
rect 14783 10180 14795 10183
rect 15396 10180 15424 10220
rect 15746 10180 15752 10192
rect 14783 10152 15424 10180
rect 15707 10152 15752 10180
rect 14783 10149 14795 10152
rect 14737 10143 14795 10149
rect 15746 10140 15752 10152
rect 15804 10140 15810 10192
rect 15856 10180 15884 10220
rect 16114 10208 16120 10220
rect 16172 10208 16178 10260
rect 16482 10248 16488 10260
rect 16395 10220 16488 10248
rect 16482 10208 16488 10220
rect 16540 10248 16546 10260
rect 18414 10248 18420 10260
rect 16540 10220 18420 10248
rect 16540 10208 16546 10220
rect 18414 10208 18420 10220
rect 18472 10208 18478 10260
rect 18690 10208 18696 10260
rect 18748 10248 18754 10260
rect 18785 10251 18843 10257
rect 18785 10248 18797 10251
rect 18748 10220 18797 10248
rect 18748 10208 18754 10220
rect 18785 10217 18797 10220
rect 18831 10217 18843 10251
rect 18785 10211 18843 10217
rect 20625 10251 20683 10257
rect 20625 10217 20637 10251
rect 20671 10217 20683 10251
rect 20625 10211 20683 10217
rect 16022 10180 16028 10192
rect 15856 10152 16028 10180
rect 16022 10140 16028 10152
rect 16080 10140 16086 10192
rect 17678 10189 17684 10192
rect 17129 10183 17187 10189
rect 17129 10180 17141 10183
rect 16132 10152 17141 10180
rect 12253 10115 12311 10121
rect 12253 10081 12265 10115
rect 12299 10112 12311 10115
rect 12342 10112 12348 10124
rect 12299 10084 12348 10112
rect 12299 10081 12311 10084
rect 12253 10075 12311 10081
rect 12342 10072 12348 10084
rect 12400 10072 12406 10124
rect 12520 10115 12578 10121
rect 12520 10081 12532 10115
rect 12566 10112 12578 10115
rect 13262 10112 13268 10124
rect 12566 10084 13268 10112
rect 12566 10081 12578 10084
rect 12520 10075 12578 10081
rect 13262 10072 13268 10084
rect 13320 10072 13326 10124
rect 14182 10072 14188 10124
rect 14240 10072 14246 10124
rect 15470 10072 15476 10124
rect 15528 10112 15534 10124
rect 15657 10115 15715 10121
rect 15657 10112 15669 10115
rect 15528 10084 15669 10112
rect 15528 10072 15534 10084
rect 15657 10081 15669 10084
rect 15703 10112 15715 10115
rect 16132 10112 16160 10152
rect 17129 10149 17141 10152
rect 17175 10149 17187 10183
rect 17129 10143 17187 10149
rect 17313 10183 17371 10189
rect 17313 10149 17325 10183
rect 17359 10180 17371 10183
rect 17650 10183 17684 10189
rect 17650 10180 17662 10183
rect 17359 10152 17662 10180
rect 17359 10149 17371 10152
rect 17313 10143 17371 10149
rect 17650 10149 17662 10152
rect 17736 10180 17742 10192
rect 20640 10180 20668 10211
rect 17736 10152 20668 10180
rect 17650 10143 17684 10149
rect 15703 10084 16160 10112
rect 15703 10081 15715 10084
rect 15657 10075 15715 10081
rect 16390 10072 16396 10124
rect 16448 10112 16454 10124
rect 16577 10115 16635 10121
rect 16577 10112 16589 10115
rect 16448 10084 16589 10112
rect 16448 10072 16454 10084
rect 16577 10081 16589 10084
rect 16623 10081 16635 10115
rect 17144 10112 17172 10143
rect 17678 10140 17684 10143
rect 17736 10140 17742 10152
rect 18782 10112 18788 10124
rect 17144 10084 18788 10112
rect 16577 10075 16635 10081
rect 18782 10072 18788 10084
rect 18840 10072 18846 10124
rect 19512 10115 19570 10121
rect 19512 10081 19524 10115
rect 19558 10112 19570 10115
rect 19886 10112 19892 10124
rect 19558 10084 19892 10112
rect 19558 10081 19570 10084
rect 19512 10075 19570 10081
rect 19886 10072 19892 10084
rect 19944 10112 19950 10124
rect 20346 10112 20352 10124
rect 19944 10084 20352 10112
rect 19944 10072 19950 10084
rect 20346 10072 20352 10084
rect 20404 10072 20410 10124
rect 12069 10047 12127 10053
rect 12069 10044 12081 10047
rect 12032 10016 12081 10044
rect 12032 10004 12038 10016
rect 12069 10013 12081 10016
rect 12115 10013 12127 10047
rect 12069 10007 12127 10013
rect 13538 10004 13544 10056
rect 13596 10044 13602 10056
rect 13725 10047 13783 10053
rect 13725 10044 13737 10047
rect 13596 10016 13737 10044
rect 13596 10004 13602 10016
rect 13725 10013 13737 10016
rect 13771 10013 13783 10047
rect 13725 10007 13783 10013
rect 14921 10047 14979 10053
rect 14921 10013 14933 10047
rect 14967 10044 14979 10047
rect 15841 10047 15899 10053
rect 15841 10044 15853 10047
rect 14967 10016 15853 10044
rect 14967 10013 14979 10016
rect 14921 10007 14979 10013
rect 15028 9988 15056 10016
rect 15841 10013 15853 10016
rect 15887 10013 15899 10047
rect 15841 10007 15899 10013
rect 16761 10047 16819 10053
rect 16761 10013 16773 10047
rect 16807 10013 16819 10047
rect 16761 10007 16819 10013
rect 9364 9948 9720 9976
rect 9364 9936 9370 9948
rect 13630 9936 13636 9988
rect 13688 9976 13694 9988
rect 14185 9979 14243 9985
rect 14185 9976 14197 9979
rect 13688 9948 14197 9976
rect 13688 9936 13694 9948
rect 14185 9945 14197 9948
rect 14231 9976 14243 9979
rect 14826 9976 14832 9988
rect 14231 9948 14832 9976
rect 14231 9945 14243 9948
rect 14185 9939 14243 9945
rect 14826 9936 14832 9948
rect 14884 9936 14890 9988
rect 15010 9936 15016 9988
rect 15068 9936 15074 9988
rect 15470 9936 15476 9988
rect 15528 9976 15534 9988
rect 16776 9976 16804 10007
rect 16850 10004 16856 10056
rect 16908 10044 16914 10056
rect 17405 10047 17463 10053
rect 17405 10044 17417 10047
rect 16908 10016 17417 10044
rect 16908 10004 16914 10016
rect 17405 10013 17417 10016
rect 17451 10013 17463 10047
rect 17405 10007 17463 10013
rect 17313 9979 17371 9985
rect 17313 9976 17325 9979
rect 15528 9948 17325 9976
rect 15528 9936 15534 9948
rect 17313 9945 17325 9948
rect 17359 9945 17371 9979
rect 17313 9939 17371 9945
rect 3237 9911 3295 9917
rect 3237 9877 3249 9911
rect 3283 9908 3295 9911
rect 3694 9908 3700 9920
rect 3283 9880 3700 9908
rect 3283 9877 3295 9880
rect 3237 9871 3295 9877
rect 3694 9868 3700 9880
rect 3752 9868 3758 9920
rect 6273 9911 6331 9917
rect 6273 9877 6285 9911
rect 6319 9908 6331 9911
rect 7190 9908 7196 9920
rect 6319 9880 7196 9908
rect 6319 9877 6331 9880
rect 6273 9871 6331 9877
rect 7190 9868 7196 9880
rect 7248 9868 7254 9920
rect 7929 9911 7987 9917
rect 7929 9877 7941 9911
rect 7975 9908 7987 9911
rect 8202 9908 8208 9920
rect 7975 9880 8208 9908
rect 7975 9877 7987 9880
rect 7929 9871 7987 9877
rect 8202 9868 8208 9880
rect 8260 9868 8266 9920
rect 9858 9868 9864 9920
rect 9916 9908 9922 9920
rect 11057 9911 11115 9917
rect 11057 9908 11069 9911
rect 9916 9880 11069 9908
rect 9916 9868 9922 9880
rect 11057 9877 11069 9880
rect 11103 9877 11115 9911
rect 11057 9871 11115 9877
rect 11425 9911 11483 9917
rect 11425 9877 11437 9911
rect 11471 9908 11483 9911
rect 11882 9908 11888 9920
rect 11471 9880 11888 9908
rect 11471 9877 11483 9880
rect 11425 9871 11483 9877
rect 11882 9868 11888 9880
rect 11940 9868 11946 9920
rect 12066 9868 12072 9920
rect 12124 9908 12130 9920
rect 15746 9908 15752 9920
rect 12124 9880 15752 9908
rect 12124 9868 12130 9880
rect 15746 9868 15752 9880
rect 15804 9868 15810 9920
rect 15930 9868 15936 9920
rect 15988 9908 15994 9920
rect 16206 9908 16212 9920
rect 15988 9880 16212 9908
rect 15988 9868 15994 9880
rect 16206 9868 16212 9880
rect 16264 9908 16270 9920
rect 16758 9908 16764 9920
rect 16264 9880 16764 9908
rect 16264 9868 16270 9880
rect 16758 9868 16764 9880
rect 16816 9868 16822 9920
rect 16942 9908 16948 9920
rect 16903 9880 16948 9908
rect 16942 9868 16948 9880
rect 17000 9868 17006 9920
rect 17420 9908 17448 10007
rect 18414 10004 18420 10056
rect 18472 10044 18478 10056
rect 18877 10047 18935 10053
rect 18877 10044 18889 10047
rect 18472 10016 18889 10044
rect 18472 10004 18478 10016
rect 18877 10013 18889 10016
rect 18923 10013 18935 10047
rect 18877 10007 18935 10013
rect 18966 10004 18972 10056
rect 19024 10044 19030 10056
rect 19245 10047 19303 10053
rect 19245 10044 19257 10047
rect 19024 10016 19257 10044
rect 19024 10004 19030 10016
rect 19245 10013 19257 10016
rect 19291 10013 19303 10047
rect 19245 10007 19303 10013
rect 18598 9908 18604 9920
rect 17420 9880 18604 9908
rect 18598 9868 18604 9880
rect 18656 9868 18662 9920
rect 19150 9908 19156 9920
rect 19111 9880 19156 9908
rect 19150 9868 19156 9880
rect 19208 9868 19214 9920
rect 1104 9818 21896 9840
rect 1104 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 4575 9818
rect 4627 9766 4639 9818
rect 4691 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 18308 9818
rect 18360 9766 18372 9818
rect 18424 9766 18436 9818
rect 18488 9766 18500 9818
rect 18552 9766 21896 9818
rect 1104 9744 21896 9766
rect 1581 9707 1639 9713
rect 1581 9673 1593 9707
rect 1627 9704 1639 9707
rect 1854 9704 1860 9716
rect 1627 9676 1860 9704
rect 1627 9673 1639 9676
rect 1581 9667 1639 9673
rect 1854 9664 1860 9676
rect 1912 9664 1918 9716
rect 2406 9704 2412 9716
rect 2367 9676 2412 9704
rect 2406 9664 2412 9676
rect 2464 9664 2470 9716
rect 2608 9676 2912 9704
rect 2608 9636 2636 9676
rect 2056 9608 2636 9636
rect 2884 9636 2912 9676
rect 2958 9664 2964 9716
rect 3016 9704 3022 9716
rect 3510 9704 3516 9716
rect 3016 9676 3516 9704
rect 3016 9664 3022 9676
rect 3510 9664 3516 9676
rect 3568 9664 3574 9716
rect 4249 9707 4307 9713
rect 4249 9673 4261 9707
rect 4295 9704 4307 9707
rect 4798 9704 4804 9716
rect 4295 9676 4804 9704
rect 4295 9673 4307 9676
rect 4249 9667 4307 9673
rect 4798 9664 4804 9676
rect 4856 9664 4862 9716
rect 8570 9664 8576 9716
rect 8628 9704 8634 9716
rect 8754 9704 8760 9716
rect 8628 9676 8760 9704
rect 8628 9664 8634 9676
rect 8754 9664 8760 9676
rect 8812 9664 8818 9716
rect 9490 9664 9496 9716
rect 9548 9704 9554 9716
rect 10134 9704 10140 9716
rect 9548 9676 9996 9704
rect 10095 9676 10140 9704
rect 9548 9664 9554 9676
rect 3237 9639 3295 9645
rect 3237 9636 3249 9639
rect 2884 9608 3249 9636
rect 2056 9577 2084 9608
rect 3237 9605 3249 9608
rect 3283 9605 3295 9639
rect 3237 9599 3295 9605
rect 4157 9639 4215 9645
rect 4157 9605 4169 9639
rect 4203 9636 4215 9639
rect 4706 9636 4712 9648
rect 4203 9608 4712 9636
rect 4203 9605 4215 9608
rect 4157 9599 4215 9605
rect 4264 9580 4292 9608
rect 4706 9596 4712 9608
rect 4764 9596 4770 9648
rect 5077 9639 5135 9645
rect 5077 9605 5089 9639
rect 5123 9636 5135 9639
rect 5534 9636 5540 9648
rect 5123 9608 5540 9636
rect 5123 9605 5135 9608
rect 5077 9599 5135 9605
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 9968 9636 9996 9676
rect 10134 9664 10140 9676
rect 10192 9664 10198 9716
rect 10428 9676 12112 9704
rect 10428 9636 10456 9676
rect 9968 9608 10456 9636
rect 12084 9636 12112 9676
rect 12158 9664 12164 9716
rect 12216 9704 12222 9716
rect 12253 9707 12311 9713
rect 12253 9704 12265 9707
rect 12216 9676 12265 9704
rect 12216 9664 12222 9676
rect 12253 9673 12265 9676
rect 12299 9673 12311 9707
rect 12526 9704 12532 9716
rect 12487 9676 12532 9704
rect 12253 9667 12311 9673
rect 12526 9664 12532 9676
rect 12584 9664 12590 9716
rect 13354 9664 13360 9716
rect 13412 9704 13418 9716
rect 14645 9707 14703 9713
rect 14645 9704 14657 9707
rect 13412 9676 14657 9704
rect 13412 9664 13418 9676
rect 14645 9673 14657 9676
rect 14691 9704 14703 9707
rect 14691 9676 15148 9704
rect 14691 9673 14703 9676
rect 14645 9667 14703 9673
rect 12342 9636 12348 9648
rect 12084 9608 12348 9636
rect 12342 9596 12348 9608
rect 12400 9596 12406 9648
rect 13722 9636 13728 9648
rect 13004 9608 13728 9636
rect 2041 9571 2099 9577
rect 2041 9537 2053 9571
rect 2087 9537 2099 9571
rect 2041 9531 2099 9537
rect 2225 9571 2283 9577
rect 2225 9537 2237 9571
rect 2271 9568 2283 9571
rect 2866 9568 2872 9580
rect 2271 9540 2872 9568
rect 2271 9537 2283 9540
rect 2225 9531 2283 9537
rect 2866 9528 2872 9540
rect 2924 9528 2930 9580
rect 3050 9568 3056 9580
rect 2963 9540 3056 9568
rect 3050 9528 3056 9540
rect 3108 9568 3114 9580
rect 3881 9571 3939 9577
rect 3881 9568 3893 9571
rect 3108 9540 3893 9568
rect 3108 9528 3114 9540
rect 3881 9537 3893 9540
rect 3927 9537 3939 9571
rect 3881 9531 3939 9537
rect 2682 9460 2688 9512
rect 2740 9500 2746 9512
rect 3068 9500 3096 9528
rect 2740 9472 3096 9500
rect 2740 9460 2746 9472
rect 3142 9460 3148 9512
rect 3200 9500 3206 9512
rect 3697 9503 3755 9509
rect 3697 9500 3709 9503
rect 3200 9472 3709 9500
rect 3200 9460 3206 9472
rect 3697 9469 3709 9472
rect 3743 9469 3755 9503
rect 3896 9500 3924 9531
rect 4246 9528 4252 9580
rect 4304 9528 4310 9580
rect 4798 9568 4804 9580
rect 4759 9540 4804 9568
rect 4798 9528 4804 9540
rect 4856 9528 4862 9580
rect 5629 9571 5687 9577
rect 5629 9537 5641 9571
rect 5675 9537 5687 9571
rect 5629 9531 5687 9537
rect 6549 9571 6607 9577
rect 6549 9537 6561 9571
rect 6595 9568 6607 9571
rect 8754 9568 8760 9580
rect 6595 9540 7144 9568
rect 8715 9540 8760 9568
rect 6595 9537 6607 9540
rect 6549 9531 6607 9537
rect 5442 9500 5448 9512
rect 3896 9472 5448 9500
rect 3697 9463 3755 9469
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 5534 9460 5540 9512
rect 5592 9500 5598 9512
rect 5644 9500 5672 9531
rect 5592 9472 5672 9500
rect 5592 9460 5598 9472
rect 6454 9460 6460 9512
rect 6512 9500 6518 9512
rect 7009 9503 7067 9509
rect 7009 9500 7021 9503
rect 6512 9472 7021 9500
rect 6512 9460 6518 9472
rect 7009 9469 7021 9472
rect 7055 9469 7067 9503
rect 7116 9500 7144 9540
rect 8754 9528 8760 9540
rect 8812 9528 8818 9580
rect 10042 9528 10048 9580
rect 10100 9568 10106 9580
rect 10229 9571 10287 9577
rect 10229 9568 10241 9571
rect 10100 9540 10241 9568
rect 10100 9528 10106 9540
rect 10229 9537 10241 9540
rect 10275 9537 10287 9571
rect 10229 9531 10287 9537
rect 12618 9528 12624 9580
rect 12676 9568 12682 9580
rect 13004 9568 13032 9608
rect 13722 9596 13728 9608
rect 13780 9636 13786 9648
rect 14185 9639 14243 9645
rect 14185 9636 14197 9639
rect 13780 9608 14197 9636
rect 13780 9596 13786 9608
rect 14185 9605 14197 9608
rect 14231 9605 14243 9639
rect 14185 9599 14243 9605
rect 14734 9596 14740 9648
rect 14792 9636 14798 9648
rect 14829 9639 14887 9645
rect 14829 9636 14841 9639
rect 14792 9608 14841 9636
rect 14792 9596 14798 9608
rect 14829 9605 14841 9608
rect 14875 9605 14887 9639
rect 14829 9599 14887 9605
rect 13170 9568 13176 9580
rect 12676 9540 13032 9568
rect 13131 9540 13176 9568
rect 12676 9528 12682 9540
rect 13170 9528 13176 9540
rect 13228 9528 13234 9580
rect 13538 9528 13544 9580
rect 13596 9568 13602 9580
rect 13596 9540 13768 9568
rect 13596 9528 13602 9540
rect 7265 9503 7323 9509
rect 7265 9500 7277 9503
rect 7116 9472 7277 9500
rect 7009 9463 7067 9469
rect 7265 9469 7277 9472
rect 7311 9500 7323 9503
rect 7742 9500 7748 9512
rect 7311 9472 7748 9500
rect 7311 9469 7323 9472
rect 7265 9463 7323 9469
rect 7742 9460 7748 9472
rect 7800 9460 7806 9512
rect 9024 9503 9082 9509
rect 9024 9469 9036 9503
rect 9070 9500 9082 9503
rect 9582 9500 9588 9512
rect 9070 9472 9588 9500
rect 9070 9469 9082 9472
rect 9024 9463 9082 9469
rect 9582 9460 9588 9472
rect 9640 9460 9646 9512
rect 10873 9503 10931 9509
rect 10873 9469 10885 9503
rect 10919 9469 10931 9503
rect 10873 9463 10931 9469
rect 11140 9503 11198 9509
rect 11140 9469 11152 9503
rect 11186 9500 11198 9503
rect 11974 9500 11980 9512
rect 11186 9472 11980 9500
rect 11186 9469 11198 9472
rect 11140 9463 11198 9469
rect 2869 9435 2927 9441
rect 2869 9432 2881 9435
rect 1412 9404 2881 9432
rect 1302 9324 1308 9376
rect 1360 9364 1366 9376
rect 1412 9373 1440 9404
rect 2869 9401 2881 9404
rect 2915 9401 2927 9435
rect 2869 9395 2927 9401
rect 6638 9392 6644 9444
rect 6696 9432 6702 9444
rect 7926 9432 7932 9444
rect 6696 9404 7932 9432
rect 6696 9392 6702 9404
rect 7926 9392 7932 9404
rect 7984 9392 7990 9444
rect 8312 9404 9067 9432
rect 1397 9367 1455 9373
rect 1397 9364 1409 9367
rect 1360 9336 1409 9364
rect 1360 9324 1366 9336
rect 1397 9333 1409 9336
rect 1443 9333 1455 9367
rect 1397 9327 1455 9333
rect 1578 9324 1584 9376
rect 1636 9364 1642 9376
rect 1949 9367 2007 9373
rect 1949 9364 1961 9367
rect 1636 9336 1961 9364
rect 1636 9324 1642 9336
rect 1949 9333 1961 9336
rect 1995 9333 2007 9367
rect 1949 9327 2007 9333
rect 2130 9324 2136 9376
rect 2188 9364 2194 9376
rect 2777 9367 2835 9373
rect 2777 9364 2789 9367
rect 2188 9336 2789 9364
rect 2188 9324 2194 9336
rect 2777 9333 2789 9336
rect 2823 9364 2835 9367
rect 3326 9364 3332 9376
rect 2823 9336 3332 9364
rect 2823 9333 2835 9336
rect 2777 9327 2835 9333
rect 3326 9324 3332 9336
rect 3384 9324 3390 9376
rect 3605 9367 3663 9373
rect 3605 9333 3617 9367
rect 3651 9364 3663 9367
rect 3694 9364 3700 9376
rect 3651 9336 3700 9364
rect 3651 9333 3663 9336
rect 3605 9327 3663 9333
rect 3694 9324 3700 9336
rect 3752 9324 3758 9376
rect 4614 9364 4620 9376
rect 4575 9336 4620 9364
rect 4614 9324 4620 9336
rect 4672 9324 4678 9376
rect 4706 9324 4712 9376
rect 4764 9364 4770 9376
rect 5074 9364 5080 9376
rect 4764 9336 5080 9364
rect 4764 9324 4770 9336
rect 5074 9324 5080 9336
rect 5132 9324 5138 9376
rect 5166 9324 5172 9376
rect 5224 9364 5230 9376
rect 5445 9367 5503 9373
rect 5445 9364 5457 9367
rect 5224 9336 5457 9364
rect 5224 9324 5230 9336
rect 5445 9333 5457 9336
rect 5491 9333 5503 9367
rect 5445 9327 5503 9333
rect 5537 9367 5595 9373
rect 5537 9333 5549 9367
rect 5583 9364 5595 9367
rect 5810 9364 5816 9376
rect 5583 9336 5816 9364
rect 5583 9333 5595 9336
rect 5537 9327 5595 9333
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 5905 9367 5963 9373
rect 5905 9333 5917 9367
rect 5951 9364 5963 9367
rect 6086 9364 6092 9376
rect 5951 9336 6092 9364
rect 5951 9333 5963 9336
rect 5905 9327 5963 9333
rect 6086 9324 6092 9336
rect 6144 9324 6150 9376
rect 6270 9364 6276 9376
rect 6231 9336 6276 9364
rect 6270 9324 6276 9336
rect 6328 9324 6334 9376
rect 6365 9367 6423 9373
rect 6365 9333 6377 9367
rect 6411 9364 6423 9367
rect 6917 9367 6975 9373
rect 6917 9364 6929 9367
rect 6411 9336 6929 9364
rect 6411 9333 6423 9336
rect 6365 9327 6423 9333
rect 6917 9333 6929 9336
rect 6963 9364 6975 9367
rect 8312 9364 8340 9404
rect 6963 9336 8340 9364
rect 6963 9333 6975 9336
rect 6917 9327 6975 9333
rect 8386 9324 8392 9376
rect 8444 9364 8450 9376
rect 8570 9364 8576 9376
rect 8444 9336 8489 9364
rect 8531 9336 8576 9364
rect 8444 9324 8450 9336
rect 8570 9324 8576 9336
rect 8628 9324 8634 9376
rect 8754 9324 8760 9376
rect 8812 9364 8818 9376
rect 8938 9364 8944 9376
rect 8812 9336 8944 9364
rect 8812 9324 8818 9336
rect 8938 9324 8944 9336
rect 8996 9324 9002 9376
rect 9039 9364 9067 9404
rect 10042 9392 10048 9444
rect 10100 9432 10106 9444
rect 10502 9432 10508 9444
rect 10100 9404 10508 9432
rect 10100 9392 10106 9404
rect 10502 9392 10508 9404
rect 10560 9392 10566 9444
rect 10888 9432 10916 9463
rect 11974 9460 11980 9472
rect 12032 9460 12038 9512
rect 12158 9500 12164 9512
rect 12084 9472 12164 9500
rect 11330 9432 11336 9444
rect 10888 9404 11336 9432
rect 11330 9392 11336 9404
rect 11388 9392 11394 9444
rect 11698 9392 11704 9444
rect 11756 9432 11762 9444
rect 12084 9432 12112 9472
rect 12158 9460 12164 9472
rect 12216 9460 12222 9512
rect 12989 9503 13047 9509
rect 12989 9469 13001 9503
rect 13035 9500 13047 9503
rect 13630 9500 13636 9512
rect 13035 9472 13636 9500
rect 13035 9469 13047 9472
rect 12989 9463 13047 9469
rect 13630 9460 13636 9472
rect 13688 9460 13694 9512
rect 13740 9509 13768 9540
rect 13906 9528 13912 9580
rect 13964 9568 13970 9580
rect 14001 9571 14059 9577
rect 14001 9568 14013 9571
rect 13964 9540 14013 9568
rect 13964 9528 13970 9540
rect 14001 9537 14013 9540
rect 14047 9568 14059 9571
rect 15010 9568 15016 9580
rect 14047 9540 15016 9568
rect 14047 9537 14059 9540
rect 14001 9531 14059 9537
rect 15010 9528 15016 9540
rect 15068 9528 15074 9580
rect 13725 9503 13783 9509
rect 13725 9469 13737 9503
rect 13771 9469 13783 9503
rect 13725 9463 13783 9469
rect 14090 9460 14096 9512
rect 14148 9500 14154 9512
rect 14369 9503 14427 9509
rect 14369 9500 14381 9503
rect 14148 9472 14381 9500
rect 14148 9460 14154 9472
rect 14369 9469 14381 9472
rect 14415 9469 14427 9503
rect 14369 9463 14427 9469
rect 13817 9435 13875 9441
rect 13817 9432 13829 9435
rect 11756 9404 12112 9432
rect 12176 9404 13829 9432
rect 11756 9392 11762 9404
rect 12176 9364 12204 9404
rect 12728 9376 12756 9404
rect 13817 9401 13829 9404
rect 13863 9432 13875 9435
rect 14461 9435 14519 9441
rect 14461 9432 14473 9435
rect 13863 9404 14473 9432
rect 13863 9401 13875 9404
rect 13817 9395 13875 9401
rect 14461 9401 14473 9404
rect 14507 9401 14519 9435
rect 15120 9432 15148 9676
rect 16390 9664 16396 9716
rect 16448 9704 16454 9716
rect 17497 9707 17555 9713
rect 17497 9704 17509 9707
rect 16448 9676 17509 9704
rect 16448 9664 16454 9676
rect 17497 9673 17509 9676
rect 17543 9673 17555 9707
rect 19610 9704 19616 9716
rect 17497 9667 17555 9673
rect 18984 9676 19616 9704
rect 15657 9639 15715 9645
rect 15657 9605 15669 9639
rect 15703 9636 15715 9639
rect 16666 9636 16672 9648
rect 15703 9608 16672 9636
rect 15703 9605 15715 9608
rect 15657 9599 15715 9605
rect 16666 9596 16672 9608
rect 16724 9596 16730 9648
rect 18984 9636 19012 9676
rect 19610 9664 19616 9676
rect 19668 9664 19674 9716
rect 20438 9704 20444 9716
rect 20399 9676 20444 9704
rect 20438 9664 20444 9676
rect 20496 9664 20502 9716
rect 20806 9664 20812 9716
rect 20864 9704 20870 9716
rect 21450 9704 21456 9716
rect 20864 9676 21456 9704
rect 20864 9664 20870 9676
rect 21450 9664 21456 9676
rect 21508 9664 21514 9716
rect 20346 9636 20352 9648
rect 18064 9608 19012 9636
rect 20307 9608 20352 9636
rect 15194 9528 15200 9580
rect 15252 9568 15258 9580
rect 15289 9571 15347 9577
rect 15289 9568 15301 9571
rect 15252 9540 15301 9568
rect 15252 9528 15258 9540
rect 15289 9537 15301 9540
rect 15335 9537 15347 9571
rect 15470 9568 15476 9580
rect 15431 9540 15476 9568
rect 15289 9531 15347 9537
rect 15470 9528 15476 9540
rect 15528 9528 15534 9580
rect 15746 9528 15752 9580
rect 15804 9568 15810 9580
rect 16206 9568 16212 9580
rect 15804 9540 16212 9568
rect 15804 9528 15810 9540
rect 16206 9528 16212 9540
rect 16264 9528 16270 9580
rect 16301 9571 16359 9577
rect 16301 9537 16313 9571
rect 16347 9568 16359 9571
rect 16574 9568 16580 9580
rect 16347 9540 16580 9568
rect 16347 9537 16359 9540
rect 16301 9531 16359 9537
rect 16574 9528 16580 9540
rect 16632 9568 16638 9580
rect 16758 9568 16764 9580
rect 16632 9540 16764 9568
rect 16632 9528 16638 9540
rect 16758 9528 16764 9540
rect 16816 9528 16822 9580
rect 16850 9528 16856 9580
rect 16908 9568 16914 9580
rect 17037 9571 17095 9577
rect 17037 9568 17049 9571
rect 16908 9540 17049 9568
rect 16908 9528 16914 9540
rect 17037 9537 17049 9540
rect 17083 9537 17095 9571
rect 17037 9531 17095 9537
rect 18064 9500 18092 9608
rect 20346 9596 20352 9608
rect 20404 9596 20410 9648
rect 21634 9596 21640 9648
rect 21692 9636 21698 9648
rect 21818 9636 21824 9648
rect 21692 9608 21824 9636
rect 21692 9596 21698 9608
rect 21818 9596 21824 9608
rect 21876 9596 21882 9648
rect 18785 9571 18843 9577
rect 18785 9537 18797 9571
rect 18831 9568 18843 9571
rect 18831 9540 19104 9568
rect 18831 9537 18843 9540
rect 18785 9531 18843 9537
rect 16316 9472 18092 9500
rect 15197 9435 15255 9441
rect 15197 9432 15209 9435
rect 15120 9404 15209 9432
rect 14461 9395 14519 9401
rect 15197 9401 15209 9404
rect 15243 9401 15255 9435
rect 15197 9395 15255 9401
rect 9039 9336 12204 9364
rect 12710 9324 12716 9376
rect 12768 9324 12774 9376
rect 12894 9364 12900 9376
rect 12855 9336 12900 9364
rect 12894 9324 12900 9336
rect 12952 9324 12958 9376
rect 13357 9367 13415 9373
rect 13357 9333 13369 9367
rect 13403 9364 13415 9367
rect 13630 9364 13636 9376
rect 13403 9336 13636 9364
rect 13403 9333 13415 9336
rect 13357 9327 13415 9333
rect 13630 9324 13636 9336
rect 13688 9324 13694 9376
rect 15838 9324 15844 9376
rect 15896 9364 15902 9376
rect 16025 9367 16083 9373
rect 16025 9364 16037 9367
rect 15896 9336 16037 9364
rect 15896 9324 15902 9336
rect 16025 9333 16037 9336
rect 16071 9333 16083 9367
rect 16025 9327 16083 9333
rect 16117 9367 16175 9373
rect 16117 9333 16129 9367
rect 16163 9364 16175 9367
rect 16206 9364 16212 9376
rect 16163 9336 16212 9364
rect 16163 9333 16175 9336
rect 16117 9327 16175 9333
rect 16206 9324 16212 9336
rect 16264 9324 16270 9376
rect 16316 9364 16344 9472
rect 18598 9460 18604 9512
rect 18656 9500 18662 9512
rect 18966 9500 18972 9512
rect 18656 9472 18972 9500
rect 18656 9460 18662 9472
rect 18966 9460 18972 9472
rect 19024 9460 19030 9512
rect 19076 9500 19104 9540
rect 20162 9528 20168 9580
rect 20220 9568 20226 9580
rect 20993 9571 21051 9577
rect 20993 9568 21005 9571
rect 20220 9540 21005 9568
rect 20220 9528 20226 9540
rect 20993 9537 21005 9540
rect 21039 9537 21051 9571
rect 20993 9531 21051 9537
rect 19236 9503 19294 9509
rect 19236 9500 19248 9503
rect 19076 9472 19248 9500
rect 19236 9469 19248 9472
rect 19282 9500 19294 9503
rect 20180 9500 20208 9528
rect 19282 9472 20208 9500
rect 19282 9469 19294 9472
rect 19236 9463 19294 9469
rect 20898 9460 20904 9512
rect 20956 9500 20962 9512
rect 21910 9500 21916 9512
rect 20956 9472 21916 9500
rect 20956 9460 20962 9472
rect 21910 9460 21916 9472
rect 21968 9460 21974 9512
rect 16390 9392 16396 9444
rect 16448 9432 16454 9444
rect 17681 9435 17739 9441
rect 17681 9432 17693 9435
rect 16448 9404 17693 9432
rect 16448 9392 16454 9404
rect 17681 9401 17693 9404
rect 17727 9401 17739 9435
rect 19702 9432 19708 9444
rect 17681 9395 17739 9401
rect 18156 9404 19708 9432
rect 16485 9367 16543 9373
rect 16485 9364 16497 9367
rect 16316 9336 16497 9364
rect 16485 9333 16497 9336
rect 16531 9333 16543 9367
rect 16485 9327 16543 9333
rect 16574 9324 16580 9376
rect 16632 9364 16638 9376
rect 16853 9367 16911 9373
rect 16853 9364 16865 9367
rect 16632 9336 16865 9364
rect 16632 9324 16638 9336
rect 16853 9333 16865 9336
rect 16899 9333 16911 9367
rect 16853 9327 16911 9333
rect 16942 9324 16948 9376
rect 17000 9364 17006 9376
rect 17402 9364 17408 9376
rect 17000 9336 17045 9364
rect 17363 9336 17408 9364
rect 17000 9324 17006 9336
rect 17402 9324 17408 9336
rect 17460 9324 17466 9376
rect 18156 9373 18184 9404
rect 19702 9392 19708 9404
rect 19760 9392 19766 9444
rect 18141 9367 18199 9373
rect 18141 9333 18153 9367
rect 18187 9333 18199 9367
rect 18506 9364 18512 9376
rect 18467 9336 18512 9364
rect 18141 9327 18199 9333
rect 18506 9324 18512 9336
rect 18564 9324 18570 9376
rect 18601 9367 18659 9373
rect 18601 9333 18613 9367
rect 18647 9364 18659 9367
rect 18874 9364 18880 9376
rect 18647 9336 18880 9364
rect 18647 9333 18659 9336
rect 18601 9327 18659 9333
rect 18874 9324 18880 9336
rect 18932 9324 18938 9376
rect 18966 9324 18972 9376
rect 19024 9364 19030 9376
rect 20809 9367 20867 9373
rect 20809 9364 20821 9367
rect 19024 9336 20821 9364
rect 19024 9324 19030 9336
rect 20809 9333 20821 9336
rect 20855 9333 20867 9367
rect 20809 9327 20867 9333
rect 20898 9324 20904 9376
rect 20956 9364 20962 9376
rect 20956 9336 21001 9364
rect 20956 9324 20962 9336
rect 1104 9274 21896 9296
rect 1104 9222 7912 9274
rect 7964 9222 7976 9274
rect 8028 9222 8040 9274
rect 8092 9222 8104 9274
rect 8156 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 15035 9274
rect 15087 9222 21896 9274
rect 1104 9200 21896 9222
rect 1578 9160 1584 9172
rect 1539 9132 1584 9160
rect 1578 9120 1584 9132
rect 1636 9120 1642 9172
rect 2409 9163 2467 9169
rect 2409 9129 2421 9163
rect 2455 9160 2467 9163
rect 2498 9160 2504 9172
rect 2455 9132 2504 9160
rect 2455 9129 2467 9132
rect 2409 9123 2467 9129
rect 2498 9120 2504 9132
rect 2556 9120 2562 9172
rect 2866 9160 2872 9172
rect 2779 9132 2872 9160
rect 2866 9120 2872 9132
rect 2924 9160 2930 9172
rect 3418 9160 3424 9172
rect 2924 9132 3424 9160
rect 2924 9120 2930 9132
rect 3418 9120 3424 9132
rect 3476 9120 3482 9172
rect 4614 9120 4620 9172
rect 4672 9160 4678 9172
rect 5442 9160 5448 9172
rect 4672 9132 4936 9160
rect 5403 9132 5448 9160
rect 4672 9120 4678 9132
rect 1949 9095 2007 9101
rect 1949 9061 1961 9095
rect 1995 9092 2007 9095
rect 3237 9095 3295 9101
rect 3237 9092 3249 9095
rect 1995 9064 3249 9092
rect 1995 9061 2007 9064
rect 1949 9055 2007 9061
rect 3237 9061 3249 9064
rect 3283 9061 3295 9095
rect 3237 9055 3295 9061
rect 4321 9095 4379 9101
rect 4321 9061 4333 9095
rect 4367 9092 4379 9095
rect 4798 9092 4804 9104
rect 4367 9064 4804 9092
rect 4367 9061 4379 9064
rect 4321 9055 4379 9061
rect 4798 9052 4804 9064
rect 4856 9052 4862 9104
rect 4908 9092 4936 9132
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 6270 9120 6276 9172
rect 6328 9160 6334 9172
rect 7837 9163 7895 9169
rect 7837 9160 7849 9163
rect 6328 9132 7849 9160
rect 6328 9120 6334 9132
rect 7837 9129 7849 9132
rect 7883 9129 7895 9163
rect 7837 9123 7895 9129
rect 8202 9120 8208 9172
rect 8260 9160 8266 9172
rect 8297 9163 8355 9169
rect 8297 9160 8309 9163
rect 8260 9132 8309 9160
rect 8260 9120 8266 9132
rect 8297 9129 8309 9132
rect 8343 9129 8355 9163
rect 8297 9123 8355 9129
rect 8389 9163 8447 9169
rect 8389 9129 8401 9163
rect 8435 9160 8447 9163
rect 8757 9163 8815 9169
rect 8757 9160 8769 9163
rect 8435 9132 8769 9160
rect 8435 9129 8447 9132
rect 8389 9123 8447 9129
rect 8757 9129 8769 9132
rect 8803 9129 8815 9163
rect 8757 9123 8815 9129
rect 9125 9163 9183 9169
rect 9125 9129 9137 9163
rect 9171 9160 9183 9163
rect 9677 9163 9735 9169
rect 9677 9160 9689 9163
rect 9171 9132 9689 9160
rect 9171 9129 9183 9132
rect 9125 9123 9183 9129
rect 9677 9129 9689 9132
rect 9723 9129 9735 9163
rect 10134 9160 10140 9172
rect 9677 9123 9735 9129
rect 9784 9132 10140 9160
rect 5626 9092 5632 9104
rect 4908 9064 5632 9092
rect 5626 9052 5632 9064
rect 5684 9052 5690 9104
rect 6454 9092 6460 9104
rect 5736 9064 6460 9092
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 2777 9027 2835 9033
rect 1443 8996 2452 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 2424 8968 2452 8996
rect 2777 8993 2789 9027
rect 2823 9024 2835 9027
rect 2823 8996 3648 9024
rect 2823 8993 2835 8996
rect 2777 8987 2835 8993
rect 1486 8916 1492 8968
rect 1544 8956 1550 8968
rect 2041 8959 2099 8965
rect 2041 8956 2053 8959
rect 1544 8928 2053 8956
rect 1544 8916 1550 8928
rect 2041 8925 2053 8928
rect 2087 8925 2099 8959
rect 2041 8919 2099 8925
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8925 2283 8959
rect 2406 8956 2412 8968
rect 2319 8928 2412 8956
rect 2225 8919 2283 8925
rect 2240 8888 2268 8919
rect 2406 8916 2412 8928
rect 2464 8956 2470 8968
rect 2866 8956 2872 8968
rect 2464 8928 2872 8956
rect 2464 8916 2470 8928
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 3050 8956 3056 8968
rect 3011 8928 3056 8956
rect 3050 8916 3056 8928
rect 3108 8916 3114 8968
rect 3068 8888 3096 8916
rect 2240 8860 3096 8888
rect 2498 8780 2504 8832
rect 2556 8820 2562 8832
rect 3142 8820 3148 8832
rect 2556 8792 3148 8820
rect 2556 8780 2562 8792
rect 3142 8780 3148 8792
rect 3200 8780 3206 8832
rect 3620 8829 3648 8996
rect 3878 8984 3884 9036
rect 3936 9024 3942 9036
rect 5736 9033 5764 9064
rect 6454 9052 6460 9064
rect 6512 9052 6518 9104
rect 7282 9052 7288 9104
rect 7340 9092 7346 9104
rect 8018 9092 8024 9104
rect 7340 9064 8024 9092
rect 7340 9052 7346 9064
rect 8018 9052 8024 9064
rect 8076 9052 8082 9104
rect 8478 9052 8484 9104
rect 8536 9092 8542 9104
rect 9030 9092 9036 9104
rect 8536 9064 9036 9092
rect 8536 9052 8542 9064
rect 9030 9052 9036 9064
rect 9088 9052 9094 9104
rect 9784 9092 9812 9132
rect 10134 9120 10140 9132
rect 10192 9120 10198 9172
rect 10594 9120 10600 9172
rect 10652 9160 10658 9172
rect 10652 9132 10824 9160
rect 10652 9120 10658 9132
rect 9508 9064 9812 9092
rect 4065 9027 4123 9033
rect 4065 9024 4077 9027
rect 3936 8996 4077 9024
rect 3936 8984 3942 8996
rect 4065 8993 4077 8996
rect 4111 9024 4123 9027
rect 5721 9027 5779 9033
rect 5721 9024 5733 9027
rect 4111 8996 5733 9024
rect 4111 8993 4123 8996
rect 4065 8987 4123 8993
rect 5721 8993 5733 8996
rect 5767 8993 5779 9027
rect 5721 8987 5779 8993
rect 5988 9027 6046 9033
rect 5988 8993 6000 9027
rect 6034 9024 6046 9027
rect 6822 9024 6828 9036
rect 6034 8996 6828 9024
rect 6034 8993 6046 8996
rect 5988 8987 6046 8993
rect 6822 8984 6828 8996
rect 6880 8984 6886 9036
rect 7374 9024 7380 9036
rect 7335 8996 7380 9024
rect 7374 8984 7380 8996
rect 7432 8984 7438 9036
rect 7466 8984 7472 9036
rect 7524 9024 7530 9036
rect 7745 9027 7803 9033
rect 7745 9024 7757 9027
rect 7524 8996 7757 9024
rect 7524 8984 7530 8996
rect 7745 8993 7757 8996
rect 7791 9024 7803 9027
rect 8202 9024 8208 9036
rect 7791 8996 8208 9024
rect 7791 8993 7803 8996
rect 7745 8987 7803 8993
rect 8202 8984 8208 8996
rect 8260 8984 8266 9036
rect 8294 8984 8300 9036
rect 8352 9024 8358 9036
rect 9217 9027 9275 9033
rect 9217 9024 9229 9027
rect 8352 8996 9229 9024
rect 8352 8984 8358 8996
rect 9217 8993 9229 8996
rect 9263 8993 9275 9027
rect 9217 8987 9275 8993
rect 5074 8916 5080 8968
rect 5132 8956 5138 8968
rect 5534 8956 5540 8968
rect 5132 8928 5540 8956
rect 5132 8916 5138 8928
rect 5534 8916 5540 8928
rect 5592 8916 5598 8968
rect 8573 8959 8631 8965
rect 6748 8928 8524 8956
rect 3605 8823 3663 8829
rect 3605 8789 3617 8823
rect 3651 8820 3663 8823
rect 5074 8820 5080 8832
rect 3651 8792 5080 8820
rect 3651 8789 3663 8792
rect 3605 8783 3663 8789
rect 5074 8780 5080 8792
rect 5132 8780 5138 8832
rect 5626 8820 5632 8832
rect 5587 8792 5632 8820
rect 5626 8780 5632 8792
rect 5684 8780 5690 8832
rect 5718 8780 5724 8832
rect 5776 8820 5782 8832
rect 6748 8820 6776 8928
rect 7006 8848 7012 8900
rect 7064 8888 7070 8900
rect 7193 8891 7251 8897
rect 7193 8888 7205 8891
rect 7064 8860 7205 8888
rect 7064 8848 7070 8860
rect 7193 8857 7205 8860
rect 7239 8857 7251 8891
rect 7193 8851 7251 8857
rect 7561 8891 7619 8897
rect 7561 8857 7573 8891
rect 7607 8888 7619 8891
rect 7837 8891 7895 8897
rect 7837 8888 7849 8891
rect 7607 8860 7849 8888
rect 7607 8857 7619 8860
rect 7561 8851 7619 8857
rect 7837 8857 7849 8860
rect 7883 8888 7895 8891
rect 8202 8888 8208 8900
rect 7883 8860 8208 8888
rect 7883 8857 7895 8860
rect 7837 8851 7895 8857
rect 8202 8848 8208 8860
rect 8260 8848 8266 8900
rect 5776 8792 6776 8820
rect 7101 8823 7159 8829
rect 5776 8780 5782 8792
rect 7101 8789 7113 8823
rect 7147 8820 7159 8823
rect 7282 8820 7288 8832
rect 7147 8792 7288 8820
rect 7147 8789 7159 8792
rect 7101 8783 7159 8789
rect 7282 8780 7288 8792
rect 7340 8780 7346 8832
rect 7926 8820 7932 8832
rect 7887 8792 7932 8820
rect 7926 8780 7932 8792
rect 7984 8780 7990 8832
rect 8496 8820 8524 8928
rect 8573 8925 8585 8959
rect 8619 8925 8631 8959
rect 8573 8919 8631 8925
rect 9401 8959 9459 8965
rect 9401 8925 9413 8959
rect 9447 8956 9459 8959
rect 9508 8956 9536 9064
rect 9858 9052 9864 9104
rect 9916 9052 9922 9104
rect 10318 9092 10324 9104
rect 10060 9064 10324 9092
rect 9867 9024 9895 9052
rect 10060 9033 10088 9064
rect 10318 9052 10324 9064
rect 10376 9052 10382 9104
rect 10502 9052 10508 9104
rect 10560 9092 10566 9104
rect 10689 9095 10747 9101
rect 10689 9092 10701 9095
rect 10560 9064 10701 9092
rect 10560 9052 10566 9064
rect 10689 9061 10701 9064
rect 10735 9061 10747 9095
rect 10796 9092 10824 9132
rect 10962 9120 10968 9172
rect 11020 9160 11026 9172
rect 11330 9160 11336 9172
rect 11020 9132 11336 9160
rect 11020 9120 11026 9132
rect 11330 9120 11336 9132
rect 11388 9120 11394 9172
rect 12894 9120 12900 9172
rect 12952 9160 12958 9172
rect 13173 9163 13231 9169
rect 13173 9160 13185 9163
rect 12952 9132 13185 9160
rect 12952 9120 12958 9132
rect 13173 9129 13185 9132
rect 13219 9129 13231 9163
rect 13541 9163 13599 9169
rect 13541 9160 13553 9163
rect 13173 9123 13231 9129
rect 13280 9132 13553 9160
rect 11241 9095 11299 9101
rect 11241 9092 11253 9095
rect 10796 9064 11253 9092
rect 10689 9055 10747 9061
rect 11241 9061 11253 9064
rect 11287 9061 11299 9095
rect 13078 9092 13084 9104
rect 12991 9064 13084 9092
rect 11241 9055 11299 9061
rect 13078 9052 13084 9064
rect 13136 9092 13142 9104
rect 13280 9092 13308 9132
rect 13541 9129 13553 9132
rect 13587 9129 13599 9163
rect 14734 9160 14740 9172
rect 13541 9123 13599 9129
rect 13648 9132 14740 9160
rect 13648 9092 13676 9132
rect 14734 9120 14740 9132
rect 14792 9120 14798 9172
rect 15194 9120 15200 9172
rect 15252 9160 15258 9172
rect 15289 9163 15347 9169
rect 15289 9160 15301 9163
rect 15252 9132 15301 9160
rect 15252 9120 15258 9132
rect 15289 9129 15301 9132
rect 15335 9160 15347 9163
rect 15746 9160 15752 9172
rect 15335 9132 15752 9160
rect 15335 9129 15347 9132
rect 15289 9123 15347 9129
rect 15746 9120 15752 9132
rect 15804 9120 15810 9172
rect 17126 9160 17132 9172
rect 17087 9132 17132 9160
rect 17126 9120 17132 9132
rect 17184 9120 17190 9172
rect 17402 9120 17408 9172
rect 17460 9160 17466 9172
rect 17589 9163 17647 9169
rect 17589 9160 17601 9163
rect 17460 9132 17601 9160
rect 17460 9120 17466 9132
rect 17589 9129 17601 9132
rect 17635 9129 17647 9163
rect 17589 9123 17647 9129
rect 17957 9163 18015 9169
rect 17957 9129 17969 9163
rect 18003 9160 18015 9163
rect 18506 9160 18512 9172
rect 18003 9132 18512 9160
rect 18003 9129 18015 9132
rect 17957 9123 18015 9129
rect 18506 9120 18512 9132
rect 18564 9120 18570 9172
rect 20162 9160 20168 9172
rect 20123 9132 20168 9160
rect 20162 9120 20168 9132
rect 20220 9120 20226 9172
rect 13136 9064 13308 9092
rect 13372 9064 13676 9092
rect 13136 9052 13142 9064
rect 10045 9027 10103 9033
rect 10045 9024 10057 9027
rect 9447 8928 9536 8956
rect 9784 8996 9895 9024
rect 9959 8996 10057 9024
rect 9447 8925 9459 8928
rect 9401 8919 9459 8925
rect 8588 8888 8616 8919
rect 9784 8888 9812 8996
rect 9858 8916 9864 8968
rect 9916 8956 9922 8968
rect 9959 8956 9987 8996
rect 10045 8993 10057 8996
rect 10091 8993 10103 9027
rect 10045 8987 10103 8993
rect 10244 8996 10364 9024
rect 10134 8956 10140 8968
rect 9916 8928 9987 8956
rect 10095 8928 10140 8956
rect 9916 8916 9922 8928
rect 10134 8916 10140 8928
rect 10192 8916 10198 8968
rect 10244 8965 10272 8996
rect 10229 8959 10287 8965
rect 10229 8925 10241 8959
rect 10275 8925 10287 8959
rect 10229 8919 10287 8925
rect 8588 8860 9812 8888
rect 9490 8820 9496 8832
rect 8496 8792 9496 8820
rect 9490 8780 9496 8792
rect 9548 8780 9554 8832
rect 9582 8780 9588 8832
rect 9640 8820 9646 8832
rect 10336 8820 10364 8996
rect 10410 8984 10416 9036
rect 10468 9024 10474 9036
rect 11422 9024 11428 9036
rect 10468 8996 11428 9024
rect 10468 8984 10474 8996
rect 11422 8984 11428 8996
rect 11480 8984 11486 9036
rect 11882 8984 11888 9036
rect 11940 9024 11946 9036
rect 13372 9024 13400 9064
rect 13722 9052 13728 9104
rect 13780 9052 13786 9104
rect 14182 9052 14188 9104
rect 14240 9092 14246 9104
rect 14277 9095 14335 9101
rect 14277 9092 14289 9095
rect 14240 9064 14289 9092
rect 14240 9052 14246 9064
rect 14277 9061 14289 9064
rect 14323 9061 14335 9095
rect 14277 9055 14335 9061
rect 14550 9052 14556 9104
rect 14608 9092 14614 9104
rect 14645 9095 14703 9101
rect 14645 9092 14657 9095
rect 14608 9064 14657 9092
rect 14608 9052 14614 9064
rect 14645 9061 14657 9064
rect 14691 9092 14703 9095
rect 15838 9092 15844 9104
rect 14691 9064 15844 9092
rect 14691 9061 14703 9064
rect 14645 9055 14703 9061
rect 15838 9052 15844 9064
rect 15896 9052 15902 9104
rect 17497 9095 17555 9101
rect 17497 9061 17509 9095
rect 17543 9061 17555 9095
rect 17497 9055 17555 9061
rect 18325 9095 18383 9101
rect 18325 9061 18337 9095
rect 18371 9092 18383 9095
rect 19242 9092 19248 9104
rect 18371 9064 19248 9092
rect 18371 9061 18383 9064
rect 18325 9055 18383 9061
rect 13630 9024 13636 9036
rect 11940 8996 13400 9024
rect 13591 8996 13636 9024
rect 11940 8984 11946 8996
rect 13630 8984 13636 8996
rect 13688 8984 13694 9036
rect 13740 9024 13768 9052
rect 15473 9027 15531 9033
rect 15473 9024 15485 9027
rect 13740 8996 15485 9024
rect 15473 8993 15485 8996
rect 15519 8993 15531 9027
rect 15473 8987 15531 8993
rect 15657 9027 15715 9033
rect 15657 8993 15669 9027
rect 15703 9024 15715 9027
rect 15746 9024 15752 9036
rect 15703 8996 15752 9024
rect 15703 8993 15715 8996
rect 15657 8987 15715 8993
rect 15746 8984 15752 8996
rect 15804 8984 15810 9036
rect 15924 9027 15982 9033
rect 15924 8993 15936 9027
rect 15970 9024 15982 9027
rect 16482 9024 16488 9036
rect 15970 8996 16488 9024
rect 15970 8993 15982 8996
rect 15924 8987 15982 8993
rect 16482 8984 16488 8996
rect 16540 8984 16546 9036
rect 17512 8968 17540 9055
rect 19242 9052 19248 9064
rect 19300 9052 19306 9104
rect 19052 9027 19110 9033
rect 19052 9024 19064 9027
rect 18616 8996 19064 9024
rect 10870 8916 10876 8968
rect 10928 8956 10934 8968
rect 11333 8959 11391 8965
rect 11333 8956 11345 8959
rect 10928 8928 11345 8956
rect 10928 8916 10934 8928
rect 11333 8925 11345 8928
rect 11379 8925 11391 8959
rect 11333 8919 11391 8925
rect 11517 8959 11575 8965
rect 11517 8925 11529 8959
rect 11563 8956 11575 8959
rect 12250 8956 12256 8968
rect 11563 8928 12256 8956
rect 11563 8925 11575 8928
rect 11517 8919 11575 8925
rect 12250 8916 12256 8928
rect 12308 8916 12314 8968
rect 12526 8916 12532 8968
rect 12584 8956 12590 8968
rect 12802 8956 12808 8968
rect 12584 8928 12808 8956
rect 12584 8916 12590 8928
rect 12802 8916 12808 8928
rect 12860 8916 12866 8968
rect 13446 8916 13452 8968
rect 13504 8956 13510 8968
rect 13725 8959 13783 8965
rect 13725 8956 13737 8959
rect 13504 8928 13737 8956
rect 13504 8916 13510 8928
rect 13725 8925 13737 8928
rect 13771 8925 13783 8959
rect 13725 8919 13783 8925
rect 14182 8916 14188 8968
rect 14240 8956 14246 8968
rect 14921 8959 14979 8965
rect 14921 8956 14933 8959
rect 14240 8928 14933 8956
rect 14240 8916 14246 8928
rect 14921 8925 14933 8928
rect 14967 8925 14979 8959
rect 14921 8919 14979 8925
rect 17494 8916 17500 8968
rect 17552 8916 17558 8968
rect 17678 8956 17684 8968
rect 17639 8928 17684 8956
rect 17678 8916 17684 8928
rect 17736 8916 17742 8968
rect 18046 8916 18052 8968
rect 18104 8956 18110 8968
rect 18616 8965 18644 8996
rect 19052 8993 19064 8996
rect 19098 9024 19110 9027
rect 19334 9024 19340 9036
rect 19098 8996 19340 9024
rect 19098 8993 19110 8996
rect 19052 8987 19110 8993
rect 19334 8984 19340 8996
rect 19392 8984 19398 9036
rect 18417 8959 18475 8965
rect 18417 8956 18429 8959
rect 18104 8928 18429 8956
rect 18104 8916 18110 8928
rect 18417 8925 18429 8928
rect 18463 8925 18475 8959
rect 18417 8919 18475 8925
rect 18601 8959 18659 8965
rect 18601 8925 18613 8959
rect 18647 8925 18659 8959
rect 18601 8919 18659 8925
rect 18785 8959 18843 8965
rect 18785 8925 18797 8959
rect 18831 8925 18843 8959
rect 18785 8919 18843 8925
rect 10410 8848 10416 8900
rect 10468 8888 10474 8900
rect 10505 8891 10563 8897
rect 10505 8888 10517 8891
rect 10468 8860 10517 8888
rect 10468 8848 10474 8860
rect 10505 8857 10517 8860
rect 10551 8857 10563 8891
rect 10505 8851 10563 8857
rect 10686 8848 10692 8900
rect 10744 8888 10750 8900
rect 10744 8860 14780 8888
rect 10744 8848 10750 8860
rect 9640 8792 10364 8820
rect 10873 8823 10931 8829
rect 9640 8780 9646 8792
rect 10873 8789 10885 8823
rect 10919 8820 10931 8823
rect 12802 8820 12808 8832
rect 10919 8792 12808 8820
rect 10919 8789 10931 8792
rect 10873 8783 10931 8789
rect 12802 8780 12808 8792
rect 12860 8780 12866 8832
rect 13446 8780 13452 8832
rect 13504 8820 13510 8832
rect 14185 8823 14243 8829
rect 14185 8820 14197 8823
rect 13504 8792 14197 8820
rect 13504 8780 13510 8792
rect 14185 8789 14197 8792
rect 14231 8820 14243 8823
rect 14642 8820 14648 8832
rect 14231 8792 14648 8820
rect 14231 8789 14243 8792
rect 14185 8783 14243 8789
rect 14642 8780 14648 8792
rect 14700 8780 14706 8832
rect 14752 8820 14780 8860
rect 14826 8848 14832 8900
rect 14884 8888 14890 8900
rect 14884 8860 14929 8888
rect 14884 8848 14890 8860
rect 15930 8820 15936 8832
rect 14752 8792 15936 8820
rect 15930 8780 15936 8792
rect 15988 8780 15994 8832
rect 16850 8780 16856 8832
rect 16908 8820 16914 8832
rect 17037 8823 17095 8829
rect 17037 8820 17049 8823
rect 16908 8792 17049 8820
rect 16908 8780 16914 8792
rect 17037 8789 17049 8792
rect 17083 8789 17095 8823
rect 17037 8783 17095 8789
rect 17954 8780 17960 8832
rect 18012 8820 18018 8832
rect 18598 8820 18604 8832
rect 18012 8792 18604 8820
rect 18012 8780 18018 8792
rect 18598 8780 18604 8792
rect 18656 8820 18662 8832
rect 18800 8820 18828 8919
rect 18656 8792 18828 8820
rect 18656 8780 18662 8792
rect 19518 8780 19524 8832
rect 19576 8820 19582 8832
rect 20349 8823 20407 8829
rect 20349 8820 20361 8823
rect 19576 8792 20361 8820
rect 19576 8780 19582 8792
rect 20349 8789 20361 8792
rect 20395 8820 20407 8823
rect 20438 8820 20444 8832
rect 20395 8792 20444 8820
rect 20395 8789 20407 8792
rect 20349 8783 20407 8789
rect 20438 8780 20444 8792
rect 20496 8780 20502 8832
rect 1104 8730 21896 8752
rect 1104 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 4575 8730
rect 4627 8678 4639 8730
rect 4691 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 18308 8730
rect 18360 8678 18372 8730
rect 18424 8678 18436 8730
rect 18488 8678 18500 8730
rect 18552 8678 21896 8730
rect 1104 8656 21896 8678
rect 3142 8616 3148 8628
rect 1412 8588 3148 8616
rect 1412 8421 1440 8588
rect 3142 8576 3148 8588
rect 3200 8576 3206 8628
rect 4249 8619 4307 8625
rect 4249 8585 4261 8619
rect 4295 8616 4307 8619
rect 4798 8616 4804 8628
rect 4295 8588 4804 8616
rect 4295 8585 4307 8588
rect 4249 8579 4307 8585
rect 4798 8576 4804 8588
rect 4856 8576 4862 8628
rect 5902 8576 5908 8628
rect 5960 8616 5966 8628
rect 6181 8619 6239 8625
rect 6181 8616 6193 8619
rect 5960 8588 6193 8616
rect 5960 8576 5966 8588
rect 6181 8585 6193 8588
rect 6227 8585 6239 8619
rect 6181 8579 6239 8585
rect 6914 8576 6920 8628
rect 6972 8616 6978 8628
rect 7193 8619 7251 8625
rect 7193 8616 7205 8619
rect 6972 8588 7205 8616
rect 6972 8576 6978 8588
rect 7193 8585 7205 8588
rect 7239 8616 7251 8619
rect 7466 8616 7472 8628
rect 7239 8588 7472 8616
rect 7239 8585 7251 8588
rect 7193 8579 7251 8585
rect 7466 8576 7472 8588
rect 7524 8576 7530 8628
rect 8754 8616 8760 8628
rect 8496 8588 8760 8616
rect 1949 8551 2007 8557
rect 1949 8517 1961 8551
rect 1995 8548 2007 8551
rect 2866 8548 2872 8560
rect 1995 8520 2872 8548
rect 1995 8517 2007 8520
rect 1949 8511 2007 8517
rect 2866 8508 2872 8520
rect 2924 8508 2930 8560
rect 6822 8508 6828 8560
rect 6880 8548 6886 8560
rect 6880 8520 8064 8548
rect 6880 8508 6886 8520
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8480 1731 8483
rect 2593 8483 2651 8489
rect 1719 8452 2544 8480
rect 1719 8449 1731 8452
rect 1673 8443 1731 8449
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8381 1455 8415
rect 1397 8375 1455 8381
rect 1946 8372 1952 8424
rect 2004 8412 2010 8424
rect 2409 8415 2467 8421
rect 2409 8412 2421 8415
rect 2004 8384 2421 8412
rect 2004 8372 2010 8384
rect 2409 8381 2421 8384
rect 2455 8381 2467 8415
rect 2516 8412 2544 8452
rect 2593 8449 2605 8483
rect 2639 8480 2651 8483
rect 2682 8480 2688 8492
rect 2639 8452 2688 8480
rect 2639 8449 2651 8452
rect 2593 8443 2651 8449
rect 2682 8440 2688 8452
rect 2740 8440 2746 8492
rect 6178 8440 6184 8492
rect 6236 8480 6242 8492
rect 8036 8489 8064 8520
rect 8496 8492 8524 8588
rect 8754 8576 8760 8588
rect 8812 8576 8818 8628
rect 9953 8619 10011 8625
rect 9953 8585 9965 8619
rect 9999 8616 10011 8619
rect 10134 8616 10140 8628
rect 9999 8588 10140 8616
rect 9999 8585 10011 8588
rect 9953 8579 10011 8585
rect 10134 8576 10140 8588
rect 10192 8576 10198 8628
rect 12437 8619 12495 8625
rect 12437 8585 12449 8619
rect 12483 8616 12495 8619
rect 12710 8616 12716 8628
rect 12483 8588 12716 8616
rect 12483 8585 12495 8588
rect 12437 8579 12495 8585
rect 12710 8576 12716 8588
rect 12768 8576 12774 8628
rect 13262 8616 13268 8628
rect 13223 8588 13268 8616
rect 13262 8576 13268 8588
rect 13320 8576 13326 8628
rect 16390 8616 16396 8628
rect 13740 8588 16396 8616
rect 9582 8508 9588 8560
rect 9640 8548 9646 8560
rect 9861 8551 9919 8557
rect 9861 8548 9873 8551
rect 9640 8520 9873 8548
rect 9640 8508 9646 8520
rect 9861 8517 9873 8520
rect 9907 8517 9919 8551
rect 9861 8511 9919 8517
rect 11882 8508 11888 8560
rect 11940 8548 11946 8560
rect 13740 8548 13768 8588
rect 16390 8576 16396 8588
rect 16448 8576 16454 8628
rect 16482 8576 16488 8628
rect 16540 8616 16546 8628
rect 16577 8619 16635 8625
rect 16577 8616 16589 8619
rect 16540 8588 16589 8616
rect 16540 8576 16546 8588
rect 16577 8585 16589 8588
rect 16623 8585 16635 8619
rect 16577 8579 16635 8585
rect 17494 8576 17500 8628
rect 17552 8616 17558 8628
rect 18877 8619 18935 8625
rect 17552 8588 18000 8616
rect 17552 8576 17558 8588
rect 11940 8520 13768 8548
rect 16408 8548 16436 8576
rect 17972 8548 18000 8588
rect 18877 8585 18889 8619
rect 18923 8616 18935 8619
rect 18966 8616 18972 8628
rect 18923 8588 18972 8616
rect 18923 8585 18935 8588
rect 18877 8579 18935 8585
rect 18966 8576 18972 8588
rect 19024 8576 19030 8628
rect 19150 8576 19156 8628
rect 19208 8616 19214 8628
rect 19334 8616 19340 8628
rect 19208 8588 19340 8616
rect 19208 8576 19214 8588
rect 19334 8576 19340 8588
rect 19392 8576 19398 8628
rect 19705 8619 19763 8625
rect 19705 8585 19717 8619
rect 19751 8616 19763 8619
rect 20898 8616 20904 8628
rect 19751 8588 20904 8616
rect 19751 8585 19763 8588
rect 19705 8579 19763 8585
rect 20898 8576 20904 8588
rect 20956 8576 20962 8628
rect 19518 8548 19524 8560
rect 16408 8520 17908 8548
rect 17972 8520 19524 8548
rect 11940 8508 11946 8520
rect 7837 8483 7895 8489
rect 7837 8480 7849 8483
rect 6236 8452 7849 8480
rect 6236 8440 6242 8452
rect 7837 8449 7849 8452
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 8021 8483 8079 8489
rect 8021 8449 8033 8483
rect 8067 8480 8079 8483
rect 8386 8480 8392 8492
rect 8067 8452 8392 8480
rect 8067 8449 8079 8452
rect 8021 8443 8079 8449
rect 8386 8440 8392 8452
rect 8444 8440 8450 8492
rect 8478 8440 8484 8492
rect 8536 8480 8542 8492
rect 8536 8452 8629 8480
rect 8536 8440 8542 8452
rect 10042 8440 10048 8492
rect 10100 8480 10106 8492
rect 10502 8480 10508 8492
rect 10100 8452 10364 8480
rect 10463 8452 10508 8480
rect 10100 8440 10106 8452
rect 2774 8412 2780 8424
rect 2516 8384 2780 8412
rect 2409 8375 2467 8381
rect 2774 8372 2780 8384
rect 2832 8372 2838 8424
rect 2869 8415 2927 8421
rect 2869 8381 2881 8415
rect 2915 8412 2927 8415
rect 3878 8412 3884 8424
rect 2915 8384 3884 8412
rect 2915 8381 2927 8384
rect 2869 8375 2927 8381
rect 3878 8372 3884 8384
rect 3936 8412 3942 8424
rect 4801 8415 4859 8421
rect 4801 8412 4813 8415
rect 3936 8384 4813 8412
rect 3936 8372 3942 8384
rect 4801 8381 4813 8384
rect 4847 8412 4859 8415
rect 6454 8412 6460 8424
rect 4847 8384 6460 8412
rect 4847 8381 4859 8384
rect 4801 8375 4859 8381
rect 6454 8372 6460 8384
rect 6512 8372 6518 8424
rect 7006 8412 7012 8424
rect 6967 8384 7012 8412
rect 7006 8372 7012 8384
rect 7064 8372 7070 8424
rect 7374 8372 7380 8424
rect 7432 8412 7438 8424
rect 7432 8384 7512 8412
rect 7432 8372 7438 8384
rect 7484 8356 7512 8384
rect 9766 8372 9772 8424
rect 9824 8412 9830 8424
rect 10336 8412 10364 8452
rect 10502 8440 10508 8452
rect 10560 8440 10566 8492
rect 10781 8483 10839 8489
rect 10781 8449 10793 8483
rect 10827 8480 10839 8483
rect 10873 8483 10931 8489
rect 10873 8480 10885 8483
rect 10827 8452 10885 8480
rect 10827 8449 10839 8452
rect 10781 8443 10839 8449
rect 10873 8449 10885 8452
rect 10919 8449 10931 8483
rect 10873 8443 10931 8449
rect 12434 8440 12440 8492
rect 12492 8480 12498 8492
rect 13078 8480 13084 8492
rect 12492 8452 12940 8480
rect 13039 8452 13084 8480
rect 12492 8440 12498 8452
rect 10413 8415 10471 8421
rect 10413 8412 10425 8415
rect 9824 8384 10272 8412
rect 10336 8384 10425 8412
rect 9824 8372 9830 8384
rect 2038 8304 2044 8356
rect 2096 8344 2102 8356
rect 2317 8347 2375 8353
rect 2317 8344 2329 8347
rect 2096 8316 2329 8344
rect 2096 8304 2102 8316
rect 2317 8313 2329 8316
rect 2363 8313 2375 8347
rect 2317 8307 2375 8313
rect 3050 8304 3056 8356
rect 3108 8353 3114 8356
rect 3108 8347 3172 8353
rect 3108 8313 3126 8347
rect 3160 8313 3172 8347
rect 3108 8307 3172 8313
rect 5068 8347 5126 8353
rect 5068 8313 5080 8347
rect 5114 8344 5126 8347
rect 5442 8344 5448 8356
rect 5114 8316 5448 8344
rect 5114 8313 5126 8316
rect 5068 8307 5126 8313
rect 3108 8304 3114 8307
rect 5442 8304 5448 8316
rect 5500 8344 5506 8356
rect 7282 8344 7288 8356
rect 5500 8316 7288 8344
rect 5500 8304 5506 8316
rect 7282 8304 7288 8316
rect 7340 8304 7346 8356
rect 7466 8304 7472 8356
rect 7524 8304 7530 8356
rect 7650 8304 7656 8356
rect 7708 8344 7714 8356
rect 8018 8344 8024 8356
rect 7708 8316 8024 8344
rect 7708 8304 7714 8316
rect 8018 8304 8024 8316
rect 8076 8304 8082 8356
rect 8748 8347 8806 8353
rect 8748 8313 8760 8347
rect 8794 8344 8806 8347
rect 9490 8344 9496 8356
rect 8794 8316 9496 8344
rect 8794 8313 8806 8316
rect 8748 8307 8806 8313
rect 9490 8304 9496 8316
rect 9548 8304 9554 8356
rect 10244 8344 10272 8384
rect 10413 8381 10425 8384
rect 10459 8381 10471 8415
rect 11129 8415 11187 8421
rect 11129 8412 11141 8415
rect 10413 8375 10471 8381
rect 10704 8384 11141 8412
rect 10704 8356 10732 8384
rect 11129 8381 11141 8384
rect 11175 8381 11187 8415
rect 12342 8412 12348 8424
rect 11129 8375 11187 8381
rect 11808 8384 12348 8412
rect 10321 8347 10379 8353
rect 10321 8344 10333 8347
rect 10244 8316 10333 8344
rect 10321 8313 10333 8316
rect 10367 8313 10379 8347
rect 10321 8307 10379 8313
rect 10686 8304 10692 8356
rect 10744 8304 10750 8356
rect 10781 8347 10839 8353
rect 10781 8313 10793 8347
rect 10827 8344 10839 8347
rect 10962 8344 10968 8356
rect 10827 8316 10968 8344
rect 10827 8313 10839 8316
rect 10781 8307 10839 8313
rect 10962 8304 10968 8316
rect 11020 8304 11026 8356
rect 3970 8236 3976 8288
rect 4028 8276 4034 8288
rect 6086 8276 6092 8288
rect 4028 8248 6092 8276
rect 4028 8236 4034 8248
rect 6086 8236 6092 8248
rect 6144 8236 6150 8288
rect 6270 8276 6276 8288
rect 6231 8248 6276 8276
rect 6270 8236 6276 8248
rect 6328 8236 6334 8288
rect 6454 8236 6460 8288
rect 6512 8276 6518 8288
rect 6825 8279 6883 8285
rect 6825 8276 6837 8279
rect 6512 8248 6837 8276
rect 6512 8236 6518 8248
rect 6825 8245 6837 8248
rect 6871 8245 6883 8279
rect 7374 8276 7380 8288
rect 7335 8248 7380 8276
rect 6825 8239 6883 8245
rect 7374 8236 7380 8248
rect 7432 8236 7438 8288
rect 7745 8279 7803 8285
rect 7745 8245 7757 8279
rect 7791 8276 7803 8279
rect 8297 8279 8355 8285
rect 8297 8276 8309 8279
rect 7791 8248 8309 8276
rect 7791 8245 7803 8248
rect 7745 8239 7803 8245
rect 8297 8245 8309 8248
rect 8343 8276 8355 8279
rect 8846 8276 8852 8288
rect 8343 8248 8852 8276
rect 8343 8245 8355 8248
rect 8297 8239 8355 8245
rect 8846 8236 8852 8248
rect 8904 8236 8910 8288
rect 9030 8236 9036 8288
rect 9088 8276 9094 8288
rect 11808 8276 11836 8384
rect 12342 8372 12348 8384
rect 12400 8372 12406 8424
rect 12802 8412 12808 8424
rect 12763 8384 12808 8412
rect 12802 8372 12808 8384
rect 12860 8372 12866 8424
rect 12912 8412 12940 8452
rect 13078 8440 13084 8452
rect 13136 8440 13142 8492
rect 13262 8440 13268 8492
rect 13320 8480 13326 8492
rect 13541 8483 13599 8489
rect 13541 8480 13553 8483
rect 13320 8452 13553 8480
rect 13320 8440 13326 8452
rect 13541 8449 13553 8452
rect 13587 8449 13599 8483
rect 15194 8480 15200 8492
rect 15155 8452 15200 8480
rect 13541 8443 13599 8449
rect 15194 8440 15200 8452
rect 15252 8440 15258 8492
rect 16758 8440 16764 8492
rect 16816 8480 16822 8492
rect 17221 8483 17279 8489
rect 17221 8480 17233 8483
rect 16816 8452 17233 8480
rect 16816 8440 16822 8452
rect 13725 8415 13783 8421
rect 13725 8412 13737 8415
rect 12912 8384 13737 8412
rect 13725 8381 13737 8384
rect 13771 8381 13783 8415
rect 13725 8375 13783 8381
rect 13992 8415 14050 8421
rect 13992 8381 14004 8415
rect 14038 8412 14050 8415
rect 16850 8412 16856 8424
rect 14038 8384 16856 8412
rect 14038 8381 14050 8384
rect 13992 8375 14050 8381
rect 16850 8372 16856 8384
rect 16908 8372 16914 8424
rect 11882 8304 11888 8356
rect 11940 8344 11946 8356
rect 14642 8344 14648 8356
rect 11940 8316 14648 8344
rect 11940 8304 11946 8316
rect 14642 8304 14648 8316
rect 14700 8304 14706 8356
rect 15464 8347 15522 8353
rect 15464 8313 15476 8347
rect 15510 8344 15522 8347
rect 15930 8344 15936 8356
rect 15510 8316 15936 8344
rect 15510 8313 15522 8316
rect 15464 8307 15522 8313
rect 15930 8304 15936 8316
rect 15988 8344 15994 8356
rect 16960 8344 16988 8452
rect 17221 8449 17233 8452
rect 17267 8480 17279 8483
rect 17678 8480 17684 8492
rect 17267 8452 17684 8480
rect 17267 8449 17279 8452
rect 17221 8443 17279 8449
rect 17678 8440 17684 8452
rect 17736 8440 17742 8492
rect 17126 8412 17132 8424
rect 17087 8384 17132 8412
rect 17126 8372 17132 8384
rect 17184 8412 17190 8424
rect 17773 8415 17831 8421
rect 17773 8412 17785 8415
rect 17184 8384 17785 8412
rect 17184 8372 17190 8384
rect 17773 8381 17785 8384
rect 17819 8381 17831 8415
rect 17773 8375 17831 8381
rect 15988 8316 16988 8344
rect 17037 8347 17095 8353
rect 15988 8304 15994 8316
rect 17037 8313 17049 8347
rect 17083 8344 17095 8347
rect 17497 8347 17555 8353
rect 17497 8344 17509 8347
rect 17083 8316 17509 8344
rect 17083 8313 17095 8316
rect 17037 8307 17095 8313
rect 17497 8313 17509 8316
rect 17543 8313 17555 8347
rect 17880 8344 17908 8520
rect 19518 8508 19524 8520
rect 19576 8508 19582 8560
rect 19610 8508 19616 8560
rect 19668 8548 19674 8560
rect 20533 8551 20591 8557
rect 20533 8548 20545 8551
rect 19668 8520 20545 8548
rect 19668 8508 19674 8520
rect 20533 8517 20545 8520
rect 20579 8517 20591 8551
rect 20533 8511 20591 8517
rect 18598 8480 18604 8492
rect 18559 8452 18604 8480
rect 18598 8440 18604 8452
rect 18656 8440 18662 8492
rect 19150 8440 19156 8492
rect 19208 8480 19214 8492
rect 19429 8483 19487 8489
rect 19429 8480 19441 8483
rect 19208 8452 19441 8480
rect 19208 8440 19214 8452
rect 19429 8449 19441 8452
rect 19475 8480 19487 8483
rect 20257 8483 20315 8489
rect 20257 8480 20269 8483
rect 19475 8452 20269 8480
rect 19475 8449 19487 8452
rect 19429 8443 19487 8449
rect 20257 8449 20269 8452
rect 20303 8449 20315 8483
rect 21082 8480 21088 8492
rect 21043 8452 21088 8480
rect 20257 8443 20315 8449
rect 21082 8440 21088 8452
rect 21140 8440 21146 8492
rect 18506 8412 18512 8424
rect 18467 8384 18512 8412
rect 18506 8372 18512 8384
rect 18564 8372 18570 8424
rect 18690 8372 18696 8424
rect 18748 8412 18754 8424
rect 20165 8415 20223 8421
rect 20165 8412 20177 8415
rect 18748 8384 20177 8412
rect 18748 8372 18754 8384
rect 20165 8381 20177 8384
rect 20211 8381 20223 8415
rect 20165 8375 20223 8381
rect 18417 8347 18475 8353
rect 18417 8344 18429 8347
rect 17880 8316 18429 8344
rect 17497 8307 17555 8313
rect 18417 8313 18429 8316
rect 18463 8313 18475 8347
rect 18417 8307 18475 8313
rect 19245 8347 19303 8353
rect 19245 8313 19257 8347
rect 19291 8344 19303 8347
rect 19978 8344 19984 8356
rect 19291 8316 19984 8344
rect 19291 8313 19303 8316
rect 19245 8307 19303 8313
rect 19978 8304 19984 8316
rect 20036 8304 20042 8356
rect 9088 8248 11836 8276
rect 9088 8236 9094 8248
rect 12250 8236 12256 8288
rect 12308 8276 12314 8288
rect 12308 8248 12353 8276
rect 12308 8236 12314 8248
rect 12802 8236 12808 8288
rect 12860 8276 12866 8288
rect 12897 8279 12955 8285
rect 12897 8276 12909 8279
rect 12860 8248 12909 8276
rect 12860 8236 12866 8248
rect 12897 8245 12909 8248
rect 12943 8245 12955 8279
rect 12897 8239 12955 8245
rect 13265 8279 13323 8285
rect 13265 8245 13277 8279
rect 13311 8276 13323 8279
rect 13449 8279 13507 8285
rect 13449 8276 13461 8279
rect 13311 8248 13461 8276
rect 13311 8245 13323 8248
rect 13265 8239 13323 8245
rect 13449 8245 13461 8248
rect 13495 8276 13507 8279
rect 13906 8276 13912 8288
rect 13495 8248 13912 8276
rect 13495 8245 13507 8248
rect 13449 8239 13507 8245
rect 13906 8236 13912 8248
rect 13964 8236 13970 8288
rect 14734 8236 14740 8288
rect 14792 8276 14798 8288
rect 15105 8279 15163 8285
rect 15105 8276 15117 8279
rect 14792 8248 15117 8276
rect 14792 8236 14798 8248
rect 15105 8245 15117 8248
rect 15151 8245 15163 8279
rect 15105 8239 15163 8245
rect 16669 8279 16727 8285
rect 16669 8245 16681 8279
rect 16715 8276 16727 8279
rect 16758 8276 16764 8288
rect 16715 8248 16764 8276
rect 16715 8245 16727 8248
rect 16669 8239 16727 8245
rect 16758 8236 16764 8248
rect 16816 8236 16822 8288
rect 16850 8236 16856 8288
rect 16908 8276 16914 8288
rect 17402 8276 17408 8288
rect 16908 8248 17408 8276
rect 16908 8236 16914 8248
rect 17402 8236 17408 8248
rect 17460 8236 17466 8288
rect 18049 8279 18107 8285
rect 18049 8245 18061 8279
rect 18095 8276 18107 8279
rect 18138 8276 18144 8288
rect 18095 8248 18144 8276
rect 18095 8245 18107 8248
rect 18049 8239 18107 8245
rect 18138 8236 18144 8248
rect 18196 8236 18202 8288
rect 19337 8279 19395 8285
rect 19337 8245 19349 8279
rect 19383 8276 19395 8279
rect 19610 8276 19616 8288
rect 19383 8248 19616 8276
rect 19383 8245 19395 8248
rect 19337 8239 19395 8245
rect 19610 8236 19616 8248
rect 19668 8236 19674 8288
rect 20070 8276 20076 8288
rect 20031 8248 20076 8276
rect 20070 8236 20076 8248
rect 20128 8236 20134 8288
rect 20714 8236 20720 8288
rect 20772 8276 20778 8288
rect 20901 8279 20959 8285
rect 20901 8276 20913 8279
rect 20772 8248 20913 8276
rect 20772 8236 20778 8248
rect 20901 8245 20913 8248
rect 20947 8245 20959 8279
rect 20901 8239 20959 8245
rect 20993 8279 21051 8285
rect 20993 8245 21005 8279
rect 21039 8276 21051 8279
rect 21450 8276 21456 8288
rect 21039 8248 21456 8276
rect 21039 8245 21051 8248
rect 20993 8239 21051 8245
rect 21450 8236 21456 8248
rect 21508 8236 21514 8288
rect 1104 8186 21896 8208
rect 1104 8134 7912 8186
rect 7964 8134 7976 8186
rect 8028 8134 8040 8186
rect 8092 8134 8104 8186
rect 8156 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 15035 8186
rect 15087 8134 21896 8186
rect 1104 8112 21896 8134
rect 1486 8072 1492 8084
rect 1447 8044 1492 8072
rect 1486 8032 1492 8044
rect 1544 8032 1550 8084
rect 2866 8032 2872 8084
rect 2924 8072 2930 8084
rect 3513 8075 3571 8081
rect 3513 8072 3525 8075
rect 2924 8044 3525 8072
rect 2924 8032 2930 8044
rect 3513 8041 3525 8044
rect 3559 8041 3571 8075
rect 3513 8035 3571 8041
rect 5077 8075 5135 8081
rect 5077 8041 5089 8075
rect 5123 8072 5135 8075
rect 5166 8072 5172 8084
rect 5123 8044 5172 8072
rect 5123 8041 5135 8044
rect 5077 8035 5135 8041
rect 5166 8032 5172 8044
rect 5224 8032 5230 8084
rect 5445 8075 5503 8081
rect 5445 8041 5457 8075
rect 5491 8072 5503 8075
rect 6270 8072 6276 8084
rect 5491 8044 6276 8072
rect 5491 8041 5503 8044
rect 5445 8035 5503 8041
rect 6270 8032 6276 8044
rect 6328 8032 6334 8084
rect 6730 8072 6736 8084
rect 6691 8044 6736 8072
rect 6730 8032 6736 8044
rect 6788 8032 6794 8084
rect 7101 8075 7159 8081
rect 7101 8041 7113 8075
rect 7147 8072 7159 8075
rect 7374 8072 7380 8084
rect 7147 8044 7380 8072
rect 7147 8041 7159 8044
rect 7101 8035 7159 8041
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 7929 8075 7987 8081
rect 7929 8041 7941 8075
rect 7975 8072 7987 8075
rect 8294 8072 8300 8084
rect 7975 8044 8300 8072
rect 7975 8041 7987 8044
rect 7929 8035 7987 8041
rect 8294 8032 8300 8044
rect 8352 8032 8358 8084
rect 8389 8075 8447 8081
rect 8389 8041 8401 8075
rect 8435 8072 8447 8075
rect 8757 8075 8815 8081
rect 8757 8072 8769 8075
rect 8435 8044 8769 8072
rect 8435 8041 8447 8044
rect 8389 8035 8447 8041
rect 8757 8041 8769 8044
rect 8803 8041 8815 8075
rect 8938 8072 8944 8084
rect 8757 8035 8815 8041
rect 8864 8044 8944 8072
rect 3602 7964 3608 8016
rect 3660 8004 3666 8016
rect 6638 8004 6644 8016
rect 3660 7976 6644 8004
rect 3660 7964 3666 7976
rect 6638 7964 6644 7976
rect 6696 7964 6702 8016
rect 7190 8004 7196 8016
rect 7151 7976 7196 8004
rect 7190 7964 7196 7976
rect 7248 7964 7254 8016
rect 8662 7964 8668 8016
rect 8720 8004 8726 8016
rect 8864 8004 8892 8044
rect 8938 8032 8944 8044
rect 8996 8072 9002 8084
rect 9217 8075 9275 8081
rect 9217 8072 9229 8075
rect 8996 8044 9229 8072
rect 8996 8032 9002 8044
rect 9217 8041 9229 8044
rect 9263 8041 9275 8075
rect 9217 8035 9275 8041
rect 10137 8075 10195 8081
rect 10137 8041 10149 8075
rect 10183 8072 10195 8075
rect 10318 8072 10324 8084
rect 10183 8044 10324 8072
rect 10183 8041 10195 8044
rect 10137 8035 10195 8041
rect 10318 8032 10324 8044
rect 10376 8032 10382 8084
rect 11238 8072 11244 8084
rect 10428 8044 11244 8072
rect 9122 8004 9128 8016
rect 8720 7976 8892 8004
rect 9035 7976 9128 8004
rect 8720 7964 8726 7976
rect 9122 7964 9128 7976
rect 9180 8004 9186 8016
rect 10428 8004 10456 8044
rect 11238 8032 11244 8044
rect 11296 8032 11302 8084
rect 11330 8032 11336 8084
rect 11388 8072 11394 8084
rect 11974 8072 11980 8084
rect 11388 8044 11980 8072
rect 11388 8032 11394 8044
rect 11974 8032 11980 8044
rect 12032 8032 12038 8084
rect 12434 8072 12440 8084
rect 12395 8044 12440 8072
rect 12434 8032 12440 8044
rect 12492 8032 12498 8084
rect 12713 8075 12771 8081
rect 12713 8041 12725 8075
rect 12759 8072 12771 8075
rect 12802 8072 12808 8084
rect 12759 8044 12808 8072
rect 12759 8041 12771 8044
rect 12713 8035 12771 8041
rect 12802 8032 12808 8044
rect 12860 8032 12866 8084
rect 13173 8075 13231 8081
rect 13173 8041 13185 8075
rect 13219 8072 13231 8075
rect 13541 8075 13599 8081
rect 13541 8072 13553 8075
rect 13219 8044 13553 8072
rect 13219 8041 13231 8044
rect 13173 8035 13231 8041
rect 13541 8041 13553 8044
rect 13587 8041 13599 8075
rect 13541 8035 13599 8041
rect 14369 8075 14427 8081
rect 14369 8041 14381 8075
rect 14415 8041 14427 8075
rect 14369 8035 14427 8041
rect 9180 7976 10456 8004
rect 10597 8007 10655 8013
rect 9180 7964 9186 7976
rect 10597 7973 10609 8007
rect 10643 8004 10655 8007
rect 13081 8007 13139 8013
rect 10643 7976 12747 8004
rect 10643 7973 10655 7976
rect 10597 7967 10655 7973
rect 1940 7939 1998 7945
rect 1940 7905 1952 7939
rect 1986 7936 1998 7939
rect 2682 7936 2688 7948
rect 1986 7908 2688 7936
rect 1986 7905 1998 7908
rect 1940 7899 1998 7905
rect 2682 7896 2688 7908
rect 2740 7896 2746 7948
rect 5074 7896 5080 7948
rect 5132 7936 5138 7948
rect 6273 7939 6331 7945
rect 6273 7936 6285 7939
rect 5132 7908 6285 7936
rect 5132 7896 5138 7908
rect 6273 7905 6285 7908
rect 6319 7905 6331 7939
rect 6273 7899 6331 7905
rect 6365 7939 6423 7945
rect 6365 7905 6377 7939
rect 6411 7936 6423 7939
rect 6914 7936 6920 7948
rect 6411 7908 6920 7936
rect 6411 7905 6423 7908
rect 6365 7899 6423 7905
rect 6914 7896 6920 7908
rect 6972 7896 6978 7948
rect 7742 7936 7748 7948
rect 7116 7908 7748 7936
rect 1670 7868 1676 7880
rect 1631 7840 1676 7868
rect 1670 7828 1676 7840
rect 1728 7828 1734 7880
rect 3602 7868 3608 7880
rect 3563 7840 3608 7868
rect 3602 7828 3608 7840
rect 3660 7828 3666 7880
rect 3697 7871 3755 7877
rect 3697 7837 3709 7871
rect 3743 7837 3755 7871
rect 5537 7871 5595 7877
rect 5537 7868 5549 7871
rect 3697 7831 3755 7837
rect 4724 7840 5549 7868
rect 3050 7800 3056 7812
rect 2963 7772 3056 7800
rect 3050 7760 3056 7772
rect 3108 7800 3114 7812
rect 3712 7800 3740 7831
rect 3108 7772 3740 7800
rect 3108 7760 3114 7772
rect 3142 7732 3148 7744
rect 3103 7704 3148 7732
rect 3142 7692 3148 7704
rect 3200 7692 3206 7744
rect 3694 7692 3700 7744
rect 3752 7732 3758 7744
rect 4724 7741 4752 7840
rect 5537 7837 5549 7840
rect 5583 7837 5595 7871
rect 5537 7831 5595 7837
rect 5721 7871 5779 7877
rect 5721 7837 5733 7871
rect 5767 7868 5779 7871
rect 6549 7871 6607 7877
rect 5767 7840 6316 7868
rect 5767 7837 5779 7840
rect 5721 7831 5779 7837
rect 5810 7760 5816 7812
rect 5868 7800 5874 7812
rect 5905 7803 5963 7809
rect 5905 7800 5917 7803
rect 5868 7772 5917 7800
rect 5868 7760 5874 7772
rect 5905 7769 5917 7772
rect 5951 7769 5963 7803
rect 6288 7800 6316 7840
rect 6549 7837 6561 7871
rect 6595 7868 6607 7871
rect 6822 7868 6828 7880
rect 6595 7840 6828 7868
rect 6595 7837 6607 7840
rect 6549 7831 6607 7837
rect 6564 7800 6592 7831
rect 6822 7828 6828 7840
rect 6880 7828 6886 7880
rect 7116 7868 7144 7908
rect 7742 7896 7748 7908
rect 7800 7896 7806 7948
rect 7837 7939 7895 7945
rect 7837 7905 7849 7939
rect 7883 7905 7895 7939
rect 8294 7936 8300 7948
rect 8255 7908 8300 7936
rect 7837 7899 7895 7905
rect 7282 7868 7288 7880
rect 6932 7840 7144 7868
rect 7243 7840 7288 7868
rect 6288 7772 6592 7800
rect 5905 7763 5963 7769
rect 6730 7760 6736 7812
rect 6788 7800 6794 7812
rect 6932 7800 6960 7840
rect 7282 7828 7288 7840
rect 7340 7828 7346 7880
rect 7852 7868 7880 7899
rect 8294 7896 8300 7908
rect 8352 7896 8358 7948
rect 9582 7936 9588 7948
rect 8588 7908 9588 7936
rect 8588 7877 8616 7908
rect 9582 7896 9588 7908
rect 9640 7896 9646 7948
rect 9950 7896 9956 7948
rect 10008 7936 10014 7948
rect 10505 7939 10563 7945
rect 10505 7936 10517 7939
rect 10008 7908 10517 7936
rect 10008 7896 10014 7908
rect 10505 7905 10517 7908
rect 10551 7905 10563 7939
rect 10505 7899 10563 7905
rect 7392 7840 7880 7868
rect 8573 7871 8631 7877
rect 6788 7772 6960 7800
rect 6788 7760 6794 7772
rect 7006 7760 7012 7812
rect 7064 7800 7070 7812
rect 7392 7800 7420 7840
rect 8573 7837 8585 7871
rect 8619 7837 8631 7871
rect 8573 7831 8631 7837
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7868 9459 7871
rect 9490 7868 9496 7880
rect 9447 7840 9496 7868
rect 9447 7837 9459 7840
rect 9401 7831 9459 7837
rect 9490 7828 9496 7840
rect 9548 7828 9554 7880
rect 10612 7868 10640 7967
rect 10686 7896 10692 7948
rect 10744 7936 10750 7948
rect 11054 7936 11060 7948
rect 10744 7908 11060 7936
rect 10744 7896 10750 7908
rect 10796 7877 10824 7908
rect 11054 7896 11060 7908
rect 11112 7896 11118 7948
rect 11232 7939 11290 7945
rect 11232 7905 11244 7939
rect 11278 7936 11290 7939
rect 12618 7936 12624 7948
rect 11278 7908 12388 7936
rect 12579 7908 12624 7936
rect 11278 7905 11290 7908
rect 11232 7899 11290 7905
rect 12360 7880 12388 7908
rect 12618 7896 12624 7908
rect 12676 7896 12682 7948
rect 12719 7936 12747 7976
rect 13081 7973 13093 8007
rect 13127 8004 13139 8007
rect 14384 8004 14412 8035
rect 14642 8032 14648 8084
rect 14700 8072 14706 8084
rect 14737 8075 14795 8081
rect 14737 8072 14749 8075
rect 14700 8044 14749 8072
rect 14700 8032 14706 8044
rect 14737 8041 14749 8044
rect 14783 8041 14795 8075
rect 14737 8035 14795 8041
rect 16577 8075 16635 8081
rect 16577 8041 16589 8075
rect 16623 8072 16635 8075
rect 17129 8075 17187 8081
rect 17129 8072 17141 8075
rect 16623 8044 17141 8072
rect 16623 8041 16635 8044
rect 16577 8035 16635 8041
rect 17129 8041 17141 8044
rect 17175 8041 17187 8075
rect 17129 8035 17187 8041
rect 18230 8032 18236 8084
rect 18288 8072 18294 8084
rect 18966 8072 18972 8084
rect 18288 8044 18972 8072
rect 18288 8032 18294 8044
rect 18966 8032 18972 8044
rect 19024 8032 19030 8084
rect 19334 8032 19340 8084
rect 19392 8072 19398 8084
rect 19429 8075 19487 8081
rect 19429 8072 19441 8075
rect 19392 8044 19441 8072
rect 19392 8032 19398 8044
rect 19429 8041 19441 8044
rect 19475 8041 19487 8075
rect 19978 8072 19984 8084
rect 19939 8044 19984 8072
rect 19429 8035 19487 8041
rect 19978 8032 19984 8044
rect 20036 8032 20042 8084
rect 20254 8032 20260 8084
rect 20312 8072 20318 8084
rect 20349 8075 20407 8081
rect 20349 8072 20361 8075
rect 20312 8044 20361 8072
rect 20312 8032 20318 8044
rect 20349 8041 20361 8044
rect 20395 8072 20407 8075
rect 21085 8075 21143 8081
rect 21085 8072 21097 8075
rect 20395 8044 21097 8072
rect 20395 8041 20407 8044
rect 20349 8035 20407 8041
rect 21085 8041 21097 8044
rect 21131 8041 21143 8075
rect 21085 8035 21143 8041
rect 13127 7976 14412 8004
rect 13127 7973 13139 7976
rect 13081 7967 13139 7973
rect 14550 7964 14556 8016
rect 14608 8004 14614 8016
rect 14829 8007 14887 8013
rect 14829 8004 14841 8007
rect 14608 7976 14841 8004
rect 14608 7964 14614 7976
rect 14829 7973 14841 7976
rect 14875 8004 14887 8007
rect 15194 8004 15200 8016
rect 14875 7976 15200 8004
rect 14875 7973 14887 7976
rect 14829 7967 14887 7973
rect 15194 7964 15200 7976
rect 15252 7964 15258 8016
rect 16666 8004 16672 8016
rect 16627 7976 16672 8004
rect 16666 7964 16672 7976
rect 16724 7964 16730 8016
rect 17497 8007 17555 8013
rect 17497 7973 17509 8007
rect 17543 8004 17555 8007
rect 17543 7976 19380 8004
rect 17543 7973 17555 7976
rect 17497 7967 17555 7973
rect 19352 7948 19380 7976
rect 13538 7936 13544 7948
rect 12719 7908 13544 7936
rect 13538 7896 13544 7908
rect 13596 7896 13602 7948
rect 13906 7936 13912 7948
rect 13867 7908 13912 7936
rect 13906 7896 13912 7908
rect 13964 7896 13970 7948
rect 14182 7896 14188 7948
rect 14240 7936 14246 7948
rect 15657 7939 15715 7945
rect 15657 7936 15669 7939
rect 14240 7908 15669 7936
rect 14240 7896 14246 7908
rect 15657 7905 15669 7908
rect 15703 7905 15715 7939
rect 15657 7899 15715 7905
rect 16482 7896 16488 7948
rect 16540 7936 16546 7948
rect 17954 7936 17960 7948
rect 16540 7908 16804 7936
rect 17915 7908 17960 7936
rect 16540 7896 16546 7908
rect 9968 7840 10640 7868
rect 10781 7871 10839 7877
rect 7064 7772 7420 7800
rect 7653 7803 7711 7809
rect 7064 7760 7070 7772
rect 7653 7769 7665 7803
rect 7699 7800 7711 7803
rect 7742 7800 7748 7812
rect 7699 7772 7748 7800
rect 7699 7769 7711 7772
rect 7653 7763 7711 7769
rect 7742 7760 7748 7772
rect 7800 7800 7806 7812
rect 8478 7800 8484 7812
rect 7800 7772 8484 7800
rect 7800 7760 7806 7772
rect 8478 7760 8484 7772
rect 8536 7760 8542 7812
rect 8938 7760 8944 7812
rect 8996 7800 9002 7812
rect 9306 7800 9312 7812
rect 8996 7772 9312 7800
rect 8996 7760 9002 7772
rect 9306 7760 9312 7772
rect 9364 7760 9370 7812
rect 9858 7760 9864 7812
rect 9916 7800 9922 7812
rect 9968 7809 9996 7840
rect 10781 7837 10793 7871
rect 10827 7837 10839 7871
rect 10962 7868 10968 7880
rect 10923 7840 10968 7868
rect 10781 7831 10839 7837
rect 10962 7828 10968 7840
rect 11020 7828 11026 7880
rect 12342 7828 12348 7880
rect 12400 7868 12406 7880
rect 13357 7871 13415 7877
rect 13357 7868 13369 7871
rect 12400 7840 13369 7868
rect 12400 7828 12406 7840
rect 13357 7837 13369 7840
rect 13403 7868 13415 7871
rect 13630 7868 13636 7880
rect 13403 7840 13636 7868
rect 13403 7837 13415 7840
rect 13357 7831 13415 7837
rect 13630 7828 13636 7840
rect 13688 7828 13694 7880
rect 13998 7868 14004 7880
rect 13959 7840 14004 7868
rect 13998 7828 14004 7840
rect 14056 7828 14062 7880
rect 14090 7828 14096 7880
rect 14148 7868 14154 7880
rect 14734 7868 14740 7880
rect 14148 7840 14740 7868
rect 14148 7828 14154 7840
rect 14734 7828 14740 7840
rect 14792 7868 14798 7880
rect 14921 7871 14979 7877
rect 14921 7868 14933 7871
rect 14792 7840 14933 7868
rect 14792 7828 14798 7840
rect 14921 7837 14933 7840
rect 14967 7837 14979 7871
rect 14921 7831 14979 7837
rect 15470 7828 15476 7880
rect 15528 7868 15534 7880
rect 15749 7871 15807 7877
rect 15749 7868 15761 7871
rect 15528 7840 15761 7868
rect 15528 7828 15534 7840
rect 15749 7837 15761 7840
rect 15795 7837 15807 7871
rect 15930 7868 15936 7880
rect 15891 7840 15936 7868
rect 15749 7831 15807 7837
rect 15930 7828 15936 7840
rect 15988 7828 15994 7880
rect 16298 7868 16304 7880
rect 16040 7840 16304 7868
rect 9953 7803 10011 7809
rect 9953 7800 9965 7803
rect 9916 7772 9965 7800
rect 9916 7760 9922 7772
rect 9953 7769 9965 7772
rect 9999 7769 10011 7803
rect 10686 7800 10692 7812
rect 9953 7763 10011 7769
rect 10244 7772 10692 7800
rect 4709 7735 4767 7741
rect 4709 7732 4721 7735
rect 3752 7704 4721 7732
rect 3752 7692 3758 7704
rect 4709 7701 4721 7704
rect 4755 7701 4767 7735
rect 4709 7695 4767 7701
rect 4985 7735 5043 7741
rect 4985 7701 4997 7735
rect 5031 7732 5043 7735
rect 5074 7732 5080 7744
rect 5031 7704 5080 7732
rect 5031 7701 5043 7704
rect 4985 7695 5043 7701
rect 5074 7692 5080 7704
rect 5132 7692 5138 7744
rect 6454 7692 6460 7744
rect 6512 7732 6518 7744
rect 8754 7732 8760 7744
rect 6512 7704 8760 7732
rect 6512 7692 6518 7704
rect 8754 7692 8760 7704
rect 8812 7692 8818 7744
rect 9766 7732 9772 7744
rect 9727 7704 9772 7732
rect 9766 7692 9772 7704
rect 9824 7732 9830 7744
rect 10244 7732 10272 7772
rect 10686 7760 10692 7772
rect 10744 7760 10750 7812
rect 16040 7800 16068 7840
rect 16298 7828 16304 7840
rect 16356 7828 16362 7880
rect 16776 7877 16804 7908
rect 17954 7896 17960 7908
rect 18012 7896 18018 7948
rect 18224 7939 18282 7945
rect 18224 7905 18236 7939
rect 18270 7936 18282 7939
rect 18598 7936 18604 7948
rect 18270 7908 18604 7936
rect 18270 7905 18282 7908
rect 18224 7899 18282 7905
rect 18598 7896 18604 7908
rect 18656 7896 18662 7948
rect 19334 7896 19340 7948
rect 19392 7896 19398 7948
rect 20993 7939 21051 7945
rect 20993 7936 21005 7939
rect 20456 7908 21005 7936
rect 16761 7871 16819 7877
rect 16761 7837 16773 7871
rect 16807 7837 16819 7871
rect 16761 7831 16819 7837
rect 17589 7871 17647 7877
rect 17589 7837 17601 7871
rect 17635 7837 17647 7871
rect 17589 7831 17647 7837
rect 11891 7772 16068 7800
rect 16209 7803 16267 7809
rect 9824 7704 10272 7732
rect 9824 7692 9830 7704
rect 10318 7692 10324 7744
rect 10376 7732 10382 7744
rect 11891 7732 11919 7772
rect 16209 7769 16221 7803
rect 16255 7800 16267 7803
rect 16942 7800 16948 7812
rect 16255 7772 16948 7800
rect 16255 7769 16267 7772
rect 16209 7763 16267 7769
rect 16942 7760 16948 7772
rect 17000 7760 17006 7812
rect 12342 7732 12348 7744
rect 10376 7704 11919 7732
rect 12255 7704 12348 7732
rect 10376 7692 10382 7704
rect 12342 7692 12348 7704
rect 12400 7732 12406 7744
rect 12986 7732 12992 7744
rect 12400 7704 12992 7732
rect 12400 7692 12406 7704
rect 12986 7692 12992 7704
rect 13044 7692 13050 7744
rect 13906 7692 13912 7744
rect 13964 7732 13970 7744
rect 14550 7732 14556 7744
rect 13964 7704 14556 7732
rect 13964 7692 13970 7704
rect 14550 7692 14556 7704
rect 14608 7692 14614 7744
rect 15289 7735 15347 7741
rect 15289 7701 15301 7735
rect 15335 7732 15347 7735
rect 15562 7732 15568 7744
rect 15335 7704 15568 7732
rect 15335 7701 15347 7704
rect 15289 7695 15347 7701
rect 15562 7692 15568 7704
rect 15620 7692 15626 7744
rect 17604 7732 17632 7831
rect 17678 7828 17684 7880
rect 17736 7868 17742 7880
rect 17736 7840 17781 7868
rect 17736 7828 17742 7840
rect 19058 7828 19064 7880
rect 19116 7868 19122 7880
rect 20456 7877 20484 7908
rect 20993 7905 21005 7908
rect 21039 7905 21051 7939
rect 20993 7899 21051 7905
rect 20441 7871 20499 7877
rect 20441 7868 20453 7871
rect 19116 7840 20453 7868
rect 19116 7828 19122 7840
rect 20441 7837 20453 7840
rect 20487 7837 20499 7871
rect 20441 7831 20499 7837
rect 20625 7871 20683 7877
rect 20625 7837 20637 7871
rect 20671 7868 20683 7871
rect 20898 7868 20904 7880
rect 20671 7840 20904 7868
rect 20671 7837 20683 7840
rect 20625 7831 20683 7837
rect 20898 7828 20904 7840
rect 20956 7868 20962 7880
rect 21082 7868 21088 7880
rect 20956 7840 21088 7868
rect 20956 7828 20962 7840
rect 21082 7828 21088 7840
rect 21140 7828 21146 7880
rect 19610 7800 19616 7812
rect 19076 7772 19616 7800
rect 19076 7732 19104 7772
rect 19610 7760 19616 7772
rect 19668 7800 19674 7812
rect 20714 7800 20720 7812
rect 19668 7772 20720 7800
rect 19668 7760 19674 7772
rect 20714 7760 20720 7772
rect 20772 7800 20778 7812
rect 21453 7803 21511 7809
rect 21453 7800 21465 7803
rect 20772 7772 21465 7800
rect 20772 7760 20778 7772
rect 21453 7769 21465 7772
rect 21499 7769 21511 7803
rect 21453 7763 21511 7769
rect 17604 7704 19104 7732
rect 19150 7692 19156 7744
rect 19208 7732 19214 7744
rect 19337 7735 19395 7741
rect 19337 7732 19349 7735
rect 19208 7704 19349 7732
rect 19208 7692 19214 7704
rect 19337 7701 19349 7704
rect 19383 7701 19395 7735
rect 19337 7695 19395 7701
rect 1104 7642 21896 7664
rect 1104 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 4575 7642
rect 4627 7590 4639 7642
rect 4691 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 18308 7642
rect 18360 7590 18372 7642
rect 18424 7590 18436 7642
rect 18488 7590 18500 7642
rect 18552 7590 21896 7642
rect 1104 7568 21896 7590
rect 3602 7488 3608 7540
rect 3660 7528 3666 7540
rect 3697 7531 3755 7537
rect 3697 7528 3709 7531
rect 3660 7500 3709 7528
rect 3660 7488 3666 7500
rect 3697 7497 3709 7500
rect 3743 7497 3755 7531
rect 5813 7531 5871 7537
rect 5813 7528 5825 7531
rect 3697 7491 3755 7497
rect 5276 7500 5825 7528
rect 5276 7460 5304 7500
rect 5813 7497 5825 7500
rect 5859 7497 5871 7531
rect 8018 7528 8024 7540
rect 5813 7491 5871 7497
rect 7576 7500 8024 7528
rect 4172 7432 5304 7460
rect 3878 7392 3884 7404
rect 3160 7364 3884 7392
rect 1670 7284 1676 7336
rect 1728 7324 1734 7336
rect 1857 7327 1915 7333
rect 1857 7324 1869 7327
rect 1728 7296 1869 7324
rect 1728 7284 1734 7296
rect 1857 7293 1869 7296
rect 1903 7324 1915 7327
rect 3160 7324 3188 7364
rect 3878 7352 3884 7364
rect 3936 7352 3942 7404
rect 4172 7401 4200 7432
rect 5442 7420 5448 7472
rect 5500 7460 5506 7472
rect 6178 7460 6184 7472
rect 5500 7432 6184 7460
rect 5500 7420 5506 7432
rect 6178 7420 6184 7432
rect 6236 7420 6242 7472
rect 6641 7463 6699 7469
rect 6641 7429 6653 7463
rect 6687 7460 6699 7463
rect 6825 7463 6883 7469
rect 6825 7460 6837 7463
rect 6687 7432 6837 7460
rect 6687 7429 6699 7432
rect 6641 7423 6699 7429
rect 6825 7429 6837 7432
rect 6871 7429 6883 7463
rect 6825 7423 6883 7429
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 4249 7395 4307 7401
rect 4249 7361 4261 7395
rect 4295 7361 4307 7395
rect 4249 7355 4307 7361
rect 4264 7324 4292 7355
rect 5166 7352 5172 7404
rect 5224 7392 5230 7404
rect 5537 7395 5595 7401
rect 5537 7392 5549 7395
rect 5224 7364 5549 7392
rect 5224 7352 5230 7364
rect 5537 7361 5549 7364
rect 5583 7361 5595 7395
rect 6365 7395 6423 7401
rect 6365 7392 6377 7395
rect 5537 7355 5595 7361
rect 5644 7364 6377 7392
rect 1903 7296 3188 7324
rect 3252 7296 4292 7324
rect 4709 7327 4767 7333
rect 1903 7293 1915 7296
rect 1857 7287 1915 7293
rect 2124 7259 2182 7265
rect 2124 7225 2136 7259
rect 2170 7256 2182 7259
rect 2590 7256 2596 7268
rect 2170 7228 2596 7256
rect 2170 7225 2182 7228
rect 2124 7219 2182 7225
rect 2590 7216 2596 7228
rect 2648 7216 2654 7268
rect 2682 7148 2688 7200
rect 2740 7188 2746 7200
rect 3252 7197 3280 7296
rect 4709 7293 4721 7327
rect 4755 7324 4767 7327
rect 4798 7324 4804 7336
rect 4755 7296 4804 7324
rect 4755 7293 4767 7296
rect 4709 7287 4767 7293
rect 4798 7284 4804 7296
rect 4856 7324 4862 7336
rect 5350 7324 5356 7336
rect 4856 7296 5356 7324
rect 4856 7284 4862 7296
rect 5350 7284 5356 7296
rect 5408 7284 5414 7336
rect 5442 7284 5448 7336
rect 5500 7324 5506 7336
rect 5644 7324 5672 7364
rect 6365 7361 6377 7364
rect 6411 7361 6423 7395
rect 7374 7392 7380 7404
rect 7335 7364 7380 7392
rect 6365 7355 6423 7361
rect 7374 7352 7380 7364
rect 7432 7352 7438 7404
rect 5500 7296 5672 7324
rect 6273 7327 6331 7333
rect 5500 7284 5506 7296
rect 6273 7293 6285 7327
rect 6319 7324 6331 7327
rect 7006 7324 7012 7336
rect 6319 7296 7012 7324
rect 6319 7293 6331 7296
rect 6273 7287 6331 7293
rect 7006 7284 7012 7296
rect 7064 7284 7070 7336
rect 7098 7284 7104 7336
rect 7156 7324 7162 7336
rect 7193 7327 7251 7333
rect 7193 7324 7205 7327
rect 7156 7296 7205 7324
rect 7156 7284 7162 7296
rect 7193 7293 7205 7296
rect 7239 7293 7251 7327
rect 7576 7324 7604 7500
rect 8018 7488 8024 7500
rect 8076 7488 8082 7540
rect 8294 7488 8300 7540
rect 8352 7528 8358 7540
rect 9125 7531 9183 7537
rect 9125 7528 9137 7531
rect 8352 7500 9137 7528
rect 8352 7488 8358 7500
rect 9125 7497 9137 7500
rect 9171 7497 9183 7531
rect 9125 7491 9183 7497
rect 10042 7488 10048 7540
rect 10100 7528 10106 7540
rect 10502 7528 10508 7540
rect 10100 7500 10508 7528
rect 10100 7488 10106 7500
rect 10502 7488 10508 7500
rect 10560 7488 10566 7540
rect 10686 7528 10692 7540
rect 10647 7500 10692 7528
rect 10686 7488 10692 7500
rect 10744 7488 10750 7540
rect 10870 7528 10876 7540
rect 10831 7500 10876 7528
rect 10870 7488 10876 7500
rect 10928 7488 10934 7540
rect 11701 7531 11759 7537
rect 11701 7497 11713 7531
rect 11747 7528 11759 7531
rect 12066 7528 12072 7540
rect 11747 7500 12072 7528
rect 11747 7497 11759 7500
rect 11701 7491 11759 7497
rect 12066 7488 12072 7500
rect 12124 7488 12130 7540
rect 13078 7528 13084 7540
rect 12176 7500 13084 7528
rect 9033 7463 9091 7469
rect 9033 7429 9045 7463
rect 9079 7429 9091 7463
rect 9033 7423 9091 7429
rect 9048 7392 9076 7423
rect 9306 7420 9312 7472
rect 9364 7460 9370 7472
rect 12176 7469 12204 7500
rect 13078 7488 13084 7500
rect 13136 7528 13142 7540
rect 13722 7528 13728 7540
rect 13136 7500 13728 7528
rect 13136 7488 13142 7500
rect 13722 7488 13728 7500
rect 13780 7488 13786 7540
rect 14642 7488 14648 7540
rect 14700 7528 14706 7540
rect 15013 7531 15071 7537
rect 15013 7528 15025 7531
rect 14700 7500 15025 7528
rect 14700 7488 14706 7500
rect 15013 7497 15025 7500
rect 15059 7497 15071 7531
rect 16574 7528 16580 7540
rect 15013 7491 15071 7497
rect 15948 7500 16580 7528
rect 12161 7463 12219 7469
rect 12161 7460 12173 7463
rect 9364 7432 12173 7460
rect 9364 7420 9370 7432
rect 12161 7429 12173 7432
rect 12207 7429 12219 7463
rect 12161 7423 12219 7429
rect 12437 7463 12495 7469
rect 12437 7429 12449 7463
rect 12483 7429 12495 7463
rect 12437 7423 12495 7429
rect 9490 7392 9496 7404
rect 9048 7364 9496 7392
rect 9490 7352 9496 7364
rect 9548 7392 9554 7404
rect 9677 7395 9735 7401
rect 9677 7392 9689 7395
rect 9548 7364 9689 7392
rect 9548 7352 9554 7364
rect 9677 7361 9689 7364
rect 9723 7361 9735 7395
rect 9677 7355 9735 7361
rect 9766 7352 9772 7404
rect 9824 7392 9830 7404
rect 10042 7392 10048 7404
rect 9824 7364 10048 7392
rect 9824 7352 9830 7364
rect 10042 7352 10048 7364
rect 10100 7352 10106 7404
rect 10226 7352 10232 7404
rect 10284 7392 10290 7404
rect 10686 7392 10692 7404
rect 10284 7364 10692 7392
rect 10284 7352 10290 7364
rect 10686 7352 10692 7364
rect 10744 7352 10750 7404
rect 11054 7352 11060 7404
rect 11112 7392 11118 7404
rect 11517 7395 11575 7401
rect 11517 7392 11529 7395
rect 11112 7364 11529 7392
rect 11112 7352 11118 7364
rect 11517 7361 11529 7364
rect 11563 7361 11575 7395
rect 12452 7392 12480 7423
rect 12986 7420 12992 7472
rect 13044 7460 13050 7472
rect 15197 7463 15255 7469
rect 13044 7432 14688 7460
rect 13044 7420 13050 7432
rect 12618 7392 12624 7404
rect 12452 7364 12624 7392
rect 11517 7355 11575 7361
rect 7193 7287 7251 7293
rect 7484 7296 7604 7324
rect 7653 7327 7711 7333
rect 4065 7259 4123 7265
rect 4065 7225 4077 7259
rect 4111 7256 4123 7259
rect 4338 7256 4344 7268
rect 4111 7228 4344 7256
rect 4111 7225 4123 7228
rect 4065 7219 4123 7225
rect 4338 7216 4344 7228
rect 4396 7216 4402 7268
rect 4893 7259 4951 7265
rect 4893 7225 4905 7259
rect 4939 7256 4951 7259
rect 4939 7228 5488 7256
rect 4939 7225 4951 7228
rect 4893 7219 4951 7225
rect 3237 7191 3295 7197
rect 3237 7188 3249 7191
rect 2740 7160 3249 7188
rect 2740 7148 2746 7160
rect 3237 7157 3249 7160
rect 3283 7157 3295 7191
rect 4982 7188 4988 7200
rect 4943 7160 4988 7188
rect 3237 7151 3295 7157
rect 4982 7148 4988 7160
rect 5040 7148 5046 7200
rect 5460 7197 5488 7228
rect 5626 7216 5632 7268
rect 5684 7256 5690 7268
rect 6086 7256 6092 7268
rect 5684 7228 6092 7256
rect 5684 7216 5690 7228
rect 6086 7216 6092 7228
rect 6144 7216 6150 7268
rect 6181 7259 6239 7265
rect 6181 7225 6193 7259
rect 6227 7256 6239 7259
rect 6641 7259 6699 7265
rect 6641 7256 6653 7259
rect 6227 7228 6653 7256
rect 6227 7225 6239 7228
rect 6181 7219 6239 7225
rect 6641 7225 6653 7228
rect 6687 7225 6699 7259
rect 7484 7256 7512 7296
rect 7653 7293 7665 7327
rect 7699 7324 7711 7327
rect 7742 7324 7748 7336
rect 7699 7296 7748 7324
rect 7699 7293 7711 7296
rect 7653 7287 7711 7293
rect 7742 7284 7748 7296
rect 7800 7284 7806 7336
rect 9585 7327 9643 7333
rect 9585 7293 9597 7327
rect 9631 7324 9643 7327
rect 10244 7324 10272 7352
rect 9631 7296 10272 7324
rect 10597 7327 10655 7333
rect 9631 7293 9643 7296
rect 9585 7287 9643 7293
rect 10597 7293 10609 7327
rect 10643 7324 10655 7327
rect 11238 7324 11244 7336
rect 10643 7296 11244 7324
rect 10643 7293 10655 7296
rect 10597 7287 10655 7293
rect 11238 7284 11244 7296
rect 11296 7284 11302 7336
rect 11532 7324 11560 7355
rect 12618 7352 12624 7364
rect 12676 7352 12682 7404
rect 13081 7395 13139 7401
rect 13081 7361 13093 7395
rect 13127 7392 13139 7395
rect 13630 7392 13636 7404
rect 13127 7364 13636 7392
rect 13127 7361 13139 7364
rect 13081 7355 13139 7361
rect 13630 7352 13636 7364
rect 13688 7352 13694 7404
rect 13722 7352 13728 7404
rect 13780 7392 13786 7404
rect 13909 7395 13967 7401
rect 13780 7364 13825 7392
rect 13780 7352 13786 7364
rect 13909 7361 13921 7395
rect 13955 7392 13967 7395
rect 14090 7392 14096 7404
rect 13955 7364 14096 7392
rect 13955 7361 13967 7364
rect 13909 7355 13967 7361
rect 13924 7324 13952 7355
rect 14090 7352 14096 7364
rect 14148 7352 14154 7404
rect 14660 7401 14688 7432
rect 15197 7429 15209 7463
rect 15243 7460 15255 7463
rect 15948 7460 15976 7500
rect 16574 7488 16580 7500
rect 16632 7488 16638 7540
rect 16666 7488 16672 7540
rect 16724 7528 16730 7540
rect 16850 7528 16856 7540
rect 16724 7500 16856 7528
rect 16724 7488 16730 7500
rect 16850 7488 16856 7500
rect 16908 7488 16914 7540
rect 17126 7528 17132 7540
rect 17039 7500 17132 7528
rect 17126 7488 17132 7500
rect 17184 7528 17190 7540
rect 17494 7528 17500 7540
rect 17184 7500 17500 7528
rect 17184 7488 17190 7500
rect 17494 7488 17500 7500
rect 17552 7488 17558 7540
rect 17681 7531 17739 7537
rect 17681 7497 17693 7531
rect 17727 7528 17739 7531
rect 17770 7528 17776 7540
rect 17727 7500 17776 7528
rect 17727 7497 17739 7500
rect 17681 7491 17739 7497
rect 17770 7488 17776 7500
rect 17828 7488 17834 7540
rect 18046 7528 18052 7540
rect 18007 7500 18052 7528
rect 18046 7488 18052 7500
rect 18104 7488 18110 7540
rect 18598 7488 18604 7540
rect 18656 7528 18662 7540
rect 19794 7528 19800 7540
rect 18656 7500 19800 7528
rect 18656 7488 18662 7500
rect 19794 7488 19800 7500
rect 19852 7488 19858 7540
rect 20070 7488 20076 7540
rect 20128 7528 20134 7540
rect 20349 7531 20407 7537
rect 20349 7528 20361 7531
rect 20128 7500 20361 7528
rect 20128 7488 20134 7500
rect 20349 7497 20361 7500
rect 20395 7497 20407 7531
rect 20349 7491 20407 7497
rect 15243 7432 15976 7460
rect 16025 7463 16083 7469
rect 15243 7429 15255 7432
rect 15197 7423 15255 7429
rect 16025 7429 16037 7463
rect 16071 7460 16083 7463
rect 19426 7460 19432 7472
rect 16071 7432 19432 7460
rect 16071 7429 16083 7432
rect 16025 7423 16083 7429
rect 19426 7420 19432 7432
rect 19484 7420 19490 7472
rect 20806 7460 20812 7472
rect 19720 7432 20812 7460
rect 14645 7395 14703 7401
rect 14645 7361 14657 7395
rect 14691 7361 14703 7395
rect 14645 7355 14703 7361
rect 15562 7352 15568 7404
rect 15620 7392 15626 7404
rect 15657 7395 15715 7401
rect 15657 7392 15669 7395
rect 15620 7364 15669 7392
rect 15620 7352 15626 7364
rect 15657 7361 15669 7364
rect 15703 7361 15715 7395
rect 15657 7355 15715 7361
rect 15841 7395 15899 7401
rect 15841 7361 15853 7395
rect 15887 7392 15899 7395
rect 16482 7392 16488 7404
rect 15887 7364 16488 7392
rect 15887 7361 15899 7364
rect 15841 7355 15899 7361
rect 16482 7352 16488 7364
rect 16540 7352 16546 7404
rect 16577 7395 16635 7401
rect 16577 7361 16589 7395
rect 16623 7361 16635 7395
rect 16850 7392 16856 7404
rect 16811 7364 16856 7392
rect 16577 7355 16635 7361
rect 11532 7296 13952 7324
rect 16390 7284 16396 7336
rect 16448 7324 16454 7336
rect 16592 7324 16620 7355
rect 16850 7352 16856 7364
rect 16908 7392 16914 7404
rect 17034 7392 17040 7404
rect 16908 7364 17040 7392
rect 16908 7352 16914 7364
rect 17034 7352 17040 7364
rect 17092 7352 17098 7404
rect 18598 7392 18604 7404
rect 18559 7364 18604 7392
rect 18598 7352 18604 7364
rect 18656 7352 18662 7404
rect 19720 7392 19748 7432
rect 20806 7420 20812 7432
rect 20864 7420 20870 7472
rect 18708 7364 19748 7392
rect 16448 7296 16620 7324
rect 16448 7284 16454 7296
rect 17770 7284 17776 7336
rect 17828 7324 17834 7336
rect 18509 7327 18567 7333
rect 18509 7324 18521 7327
rect 17828 7296 18521 7324
rect 17828 7284 17834 7296
rect 18509 7293 18521 7296
rect 18555 7293 18567 7327
rect 18509 7287 18567 7293
rect 6641 7219 6699 7225
rect 7208 7228 7512 7256
rect 5445 7191 5503 7197
rect 5445 7157 5457 7191
rect 5491 7188 5503 7191
rect 7208 7188 7236 7228
rect 7558 7216 7564 7268
rect 7616 7256 7622 7268
rect 7898 7259 7956 7265
rect 7898 7256 7910 7259
rect 7616 7228 7910 7256
rect 7616 7216 7622 7228
rect 7898 7225 7910 7228
rect 7944 7225 7956 7259
rect 7898 7219 7956 7225
rect 8018 7216 8024 7268
rect 8076 7256 8082 7268
rect 9030 7256 9036 7268
rect 8076 7228 9036 7256
rect 8076 7216 8082 7228
rect 9030 7216 9036 7228
rect 9088 7216 9094 7268
rect 9493 7259 9551 7265
rect 9493 7225 9505 7259
rect 9539 7256 9551 7259
rect 10410 7256 10416 7268
rect 9539 7228 10416 7256
rect 9539 7225 9551 7228
rect 9493 7219 9551 7225
rect 10410 7216 10416 7228
rect 10468 7256 10474 7268
rect 10778 7256 10784 7268
rect 10468 7228 10784 7256
rect 10468 7216 10474 7228
rect 10778 7216 10784 7228
rect 10836 7216 10842 7268
rect 11333 7259 11391 7265
rect 11333 7225 11345 7259
rect 11379 7256 11391 7259
rect 11514 7256 11520 7268
rect 11379 7228 11520 7256
rect 11379 7225 11391 7228
rect 11333 7219 11391 7225
rect 11514 7216 11520 7228
rect 11572 7256 11578 7268
rect 11701 7259 11759 7265
rect 11701 7256 11713 7259
rect 11572 7228 11713 7256
rect 11572 7216 11578 7228
rect 11701 7225 11713 7228
rect 11747 7225 11759 7259
rect 11701 7219 11759 7225
rect 11808 7228 12572 7256
rect 5491 7160 7236 7188
rect 7285 7191 7343 7197
rect 5491 7157 5503 7160
rect 5445 7151 5503 7157
rect 7285 7157 7297 7191
rect 7331 7188 7343 7191
rect 8294 7188 8300 7200
rect 7331 7160 8300 7188
rect 7331 7157 7343 7160
rect 7285 7151 7343 7157
rect 8294 7148 8300 7160
rect 8352 7148 8358 7200
rect 9950 7188 9956 7200
rect 9911 7160 9956 7188
rect 9950 7148 9956 7160
rect 10008 7148 10014 7200
rect 10042 7148 10048 7200
rect 10100 7188 10106 7200
rect 11241 7191 11299 7197
rect 11241 7188 11253 7191
rect 10100 7160 11253 7188
rect 10100 7148 10106 7160
rect 11241 7157 11253 7160
rect 11287 7157 11299 7191
rect 11241 7151 11299 7157
rect 11422 7148 11428 7200
rect 11480 7188 11486 7200
rect 11808 7197 11836 7228
rect 11793 7191 11851 7197
rect 11793 7188 11805 7191
rect 11480 7160 11805 7188
rect 11480 7148 11486 7160
rect 11793 7157 11805 7160
rect 11839 7157 11851 7191
rect 11793 7151 11851 7157
rect 12066 7148 12072 7200
rect 12124 7188 12130 7200
rect 12544 7188 12572 7228
rect 12618 7216 12624 7268
rect 12676 7256 12682 7268
rect 14553 7259 14611 7265
rect 14553 7256 14565 7259
rect 12676 7228 14565 7256
rect 12676 7216 12682 7228
rect 14553 7225 14565 7228
rect 14599 7225 14611 7259
rect 14553 7219 14611 7225
rect 15565 7259 15623 7265
rect 15565 7225 15577 7259
rect 15611 7256 15623 7259
rect 16758 7256 16764 7268
rect 15611 7228 16764 7256
rect 15611 7225 15623 7228
rect 15565 7219 15623 7225
rect 16758 7216 16764 7228
rect 16816 7216 16822 7268
rect 17402 7216 17408 7268
rect 17460 7256 17466 7268
rect 17865 7259 17923 7265
rect 17865 7256 17877 7259
rect 17460 7228 17877 7256
rect 17460 7216 17466 7228
rect 17865 7225 17877 7228
rect 17911 7256 17923 7259
rect 18417 7259 18475 7265
rect 18417 7256 18429 7259
rect 17911 7228 18429 7256
rect 17911 7225 17923 7228
rect 17865 7219 17923 7225
rect 18417 7225 18429 7228
rect 18463 7256 18475 7259
rect 18708 7256 18736 7364
rect 19794 7352 19800 7404
rect 19852 7392 19858 7404
rect 20165 7395 20223 7401
rect 20165 7392 20177 7395
rect 19852 7364 20177 7392
rect 19852 7352 19858 7364
rect 20165 7361 20177 7364
rect 20211 7392 20223 7395
rect 20898 7392 20904 7404
rect 20211 7364 20904 7392
rect 20211 7361 20223 7364
rect 20165 7355 20223 7361
rect 20898 7352 20904 7364
rect 20956 7352 20962 7404
rect 18969 7327 19027 7333
rect 18969 7293 18981 7327
rect 19015 7324 19027 7327
rect 19334 7324 19340 7336
rect 19015 7296 19340 7324
rect 19015 7293 19027 7296
rect 18969 7287 19027 7293
rect 19334 7284 19340 7296
rect 19392 7324 19398 7336
rect 19889 7327 19947 7333
rect 19889 7324 19901 7327
rect 19392 7296 19901 7324
rect 19392 7284 19398 7296
rect 19889 7293 19901 7296
rect 19935 7324 19947 7327
rect 20346 7324 20352 7336
rect 19935 7296 20352 7324
rect 19935 7293 19947 7296
rect 19889 7287 19947 7293
rect 20346 7284 20352 7296
rect 20404 7284 20410 7336
rect 20438 7284 20444 7336
rect 20496 7324 20502 7336
rect 20806 7324 20812 7336
rect 20496 7296 20812 7324
rect 20496 7284 20502 7296
rect 20806 7284 20812 7296
rect 20864 7284 20870 7336
rect 18463 7228 18736 7256
rect 19245 7259 19303 7265
rect 18463 7225 18475 7228
rect 18417 7219 18475 7225
rect 19245 7225 19257 7259
rect 19291 7256 19303 7259
rect 20070 7256 20076 7268
rect 19291 7228 20076 7256
rect 19291 7225 19303 7228
rect 19245 7219 19303 7225
rect 20070 7216 20076 7228
rect 20128 7216 20134 7268
rect 20162 7216 20168 7268
rect 20220 7256 20226 7268
rect 21361 7259 21419 7265
rect 21361 7256 21373 7259
rect 20220 7228 21373 7256
rect 20220 7216 20226 7228
rect 20732 7200 20760 7228
rect 21361 7225 21373 7228
rect 21407 7225 21419 7259
rect 21361 7219 21419 7225
rect 12802 7188 12808 7200
rect 12124 7160 12169 7188
rect 12544 7160 12808 7188
rect 12124 7148 12130 7160
rect 12802 7148 12808 7160
rect 12860 7148 12866 7200
rect 12897 7191 12955 7197
rect 12897 7157 12909 7191
rect 12943 7188 12955 7191
rect 13265 7191 13323 7197
rect 13265 7188 13277 7191
rect 12943 7160 13277 7188
rect 12943 7157 12955 7160
rect 12897 7151 12955 7157
rect 13265 7157 13277 7160
rect 13311 7157 13323 7191
rect 13265 7151 13323 7157
rect 13633 7191 13691 7197
rect 13633 7157 13645 7191
rect 13679 7188 13691 7191
rect 13722 7188 13728 7200
rect 13679 7160 13728 7188
rect 13679 7157 13691 7160
rect 13633 7151 13691 7157
rect 13722 7148 13728 7160
rect 13780 7148 13786 7200
rect 14090 7188 14096 7200
rect 14051 7160 14096 7188
rect 14090 7148 14096 7160
rect 14148 7148 14154 7200
rect 14458 7188 14464 7200
rect 14419 7160 14464 7188
rect 14458 7148 14464 7160
rect 14516 7148 14522 7200
rect 14642 7148 14648 7200
rect 14700 7188 14706 7200
rect 16022 7188 16028 7200
rect 14700 7160 16028 7188
rect 14700 7148 14706 7160
rect 16022 7148 16028 7160
rect 16080 7148 16086 7200
rect 16298 7148 16304 7200
rect 16356 7188 16362 7200
rect 16393 7191 16451 7197
rect 16393 7188 16405 7191
rect 16356 7160 16405 7188
rect 16356 7148 16362 7160
rect 16393 7157 16405 7160
rect 16439 7157 16451 7191
rect 16393 7151 16451 7157
rect 16485 7191 16543 7197
rect 16485 7157 16497 7191
rect 16531 7188 16543 7191
rect 16574 7188 16580 7200
rect 16531 7160 16580 7188
rect 16531 7157 16543 7160
rect 16485 7151 16543 7157
rect 16574 7148 16580 7160
rect 16632 7148 16638 7200
rect 16666 7148 16672 7200
rect 16724 7188 16730 7200
rect 19334 7188 19340 7200
rect 16724 7160 19340 7188
rect 16724 7148 16730 7160
rect 19334 7148 19340 7160
rect 19392 7148 19398 7200
rect 19518 7188 19524 7200
rect 19479 7160 19524 7188
rect 19518 7148 19524 7160
rect 19576 7148 19582 7200
rect 19978 7188 19984 7200
rect 19939 7160 19984 7188
rect 19978 7148 19984 7160
rect 20036 7148 20042 7200
rect 20714 7188 20720 7200
rect 20675 7160 20720 7188
rect 20714 7148 20720 7160
rect 20772 7148 20778 7200
rect 20806 7148 20812 7200
rect 20864 7188 20870 7200
rect 21177 7191 21235 7197
rect 21177 7188 21189 7191
rect 20864 7160 21189 7188
rect 20864 7148 20870 7160
rect 21177 7157 21189 7160
rect 21223 7157 21235 7191
rect 21177 7151 21235 7157
rect 1104 7098 21896 7120
rect 1104 7046 7912 7098
rect 7964 7046 7976 7098
rect 8028 7046 8040 7098
rect 8092 7046 8104 7098
rect 8156 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 15035 7098
rect 15087 7046 21896 7098
rect 1104 7024 21896 7046
rect 2406 6944 2412 6996
rect 2464 6984 2470 6996
rect 3050 6984 3056 6996
rect 2464 6956 3056 6984
rect 2464 6944 2470 6956
rect 3050 6944 3056 6956
rect 3108 6944 3114 6996
rect 7006 6984 7012 6996
rect 6967 6956 7012 6984
rect 7006 6944 7012 6956
rect 7064 6944 7070 6996
rect 7190 6944 7196 6996
rect 7248 6984 7254 6996
rect 9950 6984 9956 6996
rect 7248 6956 9956 6984
rect 7248 6944 7254 6956
rect 9950 6944 9956 6956
rect 10008 6944 10014 6996
rect 10318 6984 10324 6996
rect 10279 6956 10324 6984
rect 10318 6944 10324 6956
rect 10376 6944 10382 6996
rect 11514 6984 11520 6996
rect 11475 6956 11520 6984
rect 11514 6944 11520 6956
rect 11572 6944 11578 6996
rect 11698 6984 11704 6996
rect 11624 6956 11704 6984
rect 2498 6916 2504 6928
rect 2332 6888 2504 6916
rect 1762 6808 1768 6860
rect 1820 6848 1826 6860
rect 2332 6857 2360 6888
rect 2498 6876 2504 6888
rect 2556 6876 2562 6928
rect 3418 6876 3424 6928
rect 3476 6916 3482 6928
rect 3694 6916 3700 6928
rect 3476 6888 3700 6916
rect 3476 6876 3482 6888
rect 3694 6876 3700 6888
rect 3752 6876 3758 6928
rect 4062 6876 4068 6928
rect 4120 6916 4126 6928
rect 9769 6919 9827 6925
rect 9769 6916 9781 6919
rect 4120 6888 9781 6916
rect 4120 6876 4126 6888
rect 9769 6885 9781 6888
rect 9815 6916 9827 6919
rect 10336 6916 10364 6944
rect 11624 6916 11652 6956
rect 11698 6944 11704 6956
rect 11756 6944 11762 6996
rect 12894 6944 12900 6996
rect 12952 6984 12958 6996
rect 14550 6984 14556 6996
rect 12952 6956 14412 6984
rect 14511 6956 14556 6984
rect 12952 6944 12958 6956
rect 9815 6888 10364 6916
rect 11532 6888 11652 6916
rect 13449 6919 13507 6925
rect 9815 6885 9827 6888
rect 9769 6879 9827 6885
rect 2317 6851 2375 6857
rect 2317 6848 2329 6851
rect 1820 6820 2329 6848
rect 1820 6808 1826 6820
rect 2317 6817 2329 6820
rect 2363 6817 2375 6851
rect 3145 6851 3203 6857
rect 3145 6848 3157 6851
rect 2317 6811 2375 6817
rect 2884 6820 3157 6848
rect 1670 6780 1676 6792
rect 1631 6752 1676 6780
rect 1670 6740 1676 6752
rect 1728 6740 1734 6792
rect 2409 6783 2467 6789
rect 2409 6749 2421 6783
rect 2455 6749 2467 6783
rect 2590 6780 2596 6792
rect 2551 6752 2596 6780
rect 2409 6743 2467 6749
rect 1946 6712 1952 6724
rect 1907 6684 1952 6712
rect 1946 6672 1952 6684
rect 2004 6672 2010 6724
rect 2424 6712 2452 6743
rect 2590 6740 2596 6752
rect 2648 6740 2654 6792
rect 2777 6715 2835 6721
rect 2777 6712 2789 6715
rect 2424 6684 2789 6712
rect 2777 6681 2789 6684
rect 2823 6681 2835 6715
rect 2777 6675 2835 6681
rect 1302 6604 1308 6656
rect 1360 6644 1366 6656
rect 1489 6647 1547 6653
rect 1489 6644 1501 6647
rect 1360 6616 1501 6644
rect 1360 6604 1366 6616
rect 1489 6613 1501 6616
rect 1535 6644 1547 6647
rect 2884 6644 2912 6820
rect 3145 6817 3157 6820
rect 3191 6817 3203 6851
rect 4321 6851 4379 6857
rect 4321 6848 4333 6851
rect 3145 6811 3203 6817
rect 3436 6820 4333 6848
rect 3436 6792 3464 6820
rect 4321 6817 4333 6820
rect 4367 6848 4379 6851
rect 5166 6848 5172 6860
rect 4367 6820 5172 6848
rect 4367 6817 4379 6820
rect 4321 6811 4379 6817
rect 5166 6808 5172 6820
rect 5224 6808 5230 6860
rect 5810 6857 5816 6860
rect 5804 6848 5816 6857
rect 5771 6820 5816 6848
rect 5804 6811 5816 6820
rect 5810 6808 5816 6811
rect 5868 6808 5874 6860
rect 6178 6808 6184 6860
rect 6236 6848 6242 6860
rect 7377 6851 7435 6857
rect 6236 6820 7328 6848
rect 6236 6808 6242 6820
rect 3050 6740 3056 6792
rect 3108 6780 3114 6792
rect 3237 6783 3295 6789
rect 3237 6780 3249 6783
rect 3108 6752 3249 6780
rect 3108 6740 3114 6752
rect 3237 6749 3249 6752
rect 3283 6749 3295 6783
rect 3418 6780 3424 6792
rect 3379 6752 3424 6780
rect 3237 6743 3295 6749
rect 3418 6740 3424 6752
rect 3476 6740 3482 6792
rect 3878 6740 3884 6792
rect 3936 6780 3942 6792
rect 4065 6783 4123 6789
rect 4065 6780 4077 6783
rect 3936 6752 4077 6780
rect 3936 6740 3942 6752
rect 4065 6749 4077 6752
rect 4111 6749 4123 6783
rect 5537 6783 5595 6789
rect 5537 6780 5549 6783
rect 4065 6743 4123 6749
rect 5083 6752 5549 6780
rect 1535 6616 2912 6644
rect 4080 6644 4108 6743
rect 5083 6644 5111 6752
rect 5537 6749 5549 6752
rect 5583 6749 5595 6783
rect 5537 6743 5595 6749
rect 7300 6780 7328 6820
rect 7377 6817 7389 6851
rect 7423 6848 7435 6851
rect 7650 6848 7656 6860
rect 7423 6820 7656 6848
rect 7423 6817 7435 6820
rect 7377 6811 7435 6817
rect 7650 6808 7656 6820
rect 7708 6848 7714 6860
rect 8297 6851 8355 6857
rect 7708 6820 8248 6848
rect 7708 6808 7714 6820
rect 8220 6792 8248 6820
rect 8297 6817 8309 6851
rect 8343 6848 8355 6851
rect 8343 6820 8616 6848
rect 8343 6817 8355 6820
rect 8297 6811 8355 6817
rect 7469 6783 7527 6789
rect 7469 6780 7481 6783
rect 7300 6752 7481 6780
rect 5442 6644 5448 6656
rect 4080 6616 5111 6644
rect 5403 6616 5448 6644
rect 1535 6613 1547 6616
rect 1489 6607 1547 6613
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 6914 6644 6920 6656
rect 6875 6616 6920 6644
rect 6914 6604 6920 6616
rect 6972 6604 6978 6656
rect 7300 6644 7328 6752
rect 7469 6749 7481 6752
rect 7515 6749 7527 6783
rect 7469 6743 7527 6749
rect 7561 6783 7619 6789
rect 7561 6749 7573 6783
rect 7607 6749 7619 6783
rect 7834 6780 7840 6792
rect 7795 6752 7840 6780
rect 7561 6743 7619 6749
rect 7374 6672 7380 6724
rect 7432 6712 7438 6724
rect 7576 6712 7604 6743
rect 7834 6740 7840 6752
rect 7892 6740 7898 6792
rect 8018 6740 8024 6792
rect 8076 6780 8082 6792
rect 8076 6752 8121 6780
rect 8076 6740 8082 6752
rect 8202 6740 8208 6792
rect 8260 6780 8266 6792
rect 8389 6783 8447 6789
rect 8389 6780 8401 6783
rect 8260 6752 8401 6780
rect 8260 6740 8266 6752
rect 8389 6749 8401 6752
rect 8435 6749 8447 6783
rect 8588 6780 8616 6820
rect 8662 6808 8668 6860
rect 8720 6848 8726 6860
rect 8941 6851 8999 6857
rect 8941 6848 8953 6851
rect 8720 6820 8953 6848
rect 8720 6808 8726 6820
rect 8941 6817 8953 6820
rect 8987 6817 8999 6851
rect 8941 6811 8999 6817
rect 10229 6851 10287 6857
rect 10229 6817 10241 6851
rect 10275 6848 10287 6851
rect 10689 6851 10747 6857
rect 10689 6848 10701 6851
rect 10275 6820 10701 6848
rect 10275 6817 10287 6820
rect 10229 6811 10287 6817
rect 10689 6817 10701 6820
rect 10735 6817 10747 6851
rect 10689 6811 10747 6817
rect 9398 6780 9404 6792
rect 8588 6752 9404 6780
rect 8389 6743 8447 6749
rect 9398 6740 9404 6752
rect 9456 6780 9462 6792
rect 10318 6780 10324 6792
rect 9456 6752 10324 6780
rect 9456 6740 9462 6752
rect 10318 6740 10324 6752
rect 10376 6740 10382 6792
rect 10505 6783 10563 6789
rect 10505 6749 10517 6783
rect 10551 6780 10563 6783
rect 11532 6780 11560 6888
rect 13449 6885 13461 6919
rect 13495 6916 13507 6919
rect 14384 6916 14412 6956
rect 14550 6944 14556 6956
rect 14608 6984 14614 6996
rect 15013 6987 15071 6993
rect 15013 6984 15025 6987
rect 14608 6956 15025 6984
rect 14608 6944 14614 6956
rect 15013 6953 15025 6956
rect 15059 6953 15071 6987
rect 15013 6947 15071 6953
rect 15194 6944 15200 6996
rect 15252 6984 15258 6996
rect 15381 6987 15439 6993
rect 15381 6984 15393 6987
rect 15252 6956 15393 6984
rect 15252 6944 15258 6956
rect 15381 6953 15393 6956
rect 15427 6984 15439 6987
rect 16022 6984 16028 6996
rect 15427 6956 16028 6984
rect 15427 6953 15439 6956
rect 15381 6947 15439 6953
rect 16022 6944 16028 6956
rect 16080 6944 16086 6996
rect 16482 6984 16488 6996
rect 16224 6956 16488 6984
rect 16224 6916 16252 6956
rect 16482 6944 16488 6956
rect 16540 6944 16546 6996
rect 16577 6987 16635 6993
rect 16577 6953 16589 6987
rect 16623 6984 16635 6987
rect 17126 6984 17132 6996
rect 16623 6956 17132 6984
rect 16623 6953 16635 6956
rect 16577 6947 16635 6953
rect 17126 6944 17132 6956
rect 17184 6944 17190 6996
rect 18138 6944 18144 6996
rect 18196 6984 18202 6996
rect 19245 6987 19303 6993
rect 19245 6984 19257 6987
rect 18196 6956 19257 6984
rect 18196 6944 18202 6956
rect 19245 6953 19257 6956
rect 19291 6953 19303 6987
rect 19245 6947 19303 6953
rect 19337 6987 19395 6993
rect 19337 6953 19349 6987
rect 19383 6984 19395 6987
rect 19518 6984 19524 6996
rect 19383 6956 19524 6984
rect 19383 6953 19395 6956
rect 19337 6947 19395 6953
rect 19518 6944 19524 6956
rect 19576 6944 19582 6996
rect 19794 6944 19800 6996
rect 19852 6944 19858 6996
rect 20070 6984 20076 6996
rect 20031 6956 20076 6984
rect 20070 6944 20076 6956
rect 20128 6944 20134 6996
rect 13495 6888 13952 6916
rect 14384 6888 16252 6916
rect 13495 6885 13507 6888
rect 13449 6879 13507 6885
rect 11876 6851 11934 6857
rect 11876 6817 11888 6851
rect 11922 6848 11934 6851
rect 12342 6848 12348 6860
rect 11922 6820 12348 6848
rect 11922 6817 11934 6820
rect 11876 6811 11934 6817
rect 12342 6808 12348 6820
rect 12400 6808 12406 6860
rect 13924 6857 13952 6888
rect 16298 6876 16304 6928
rect 16356 6916 16362 6928
rect 17586 6916 17592 6928
rect 16356 6888 17592 6916
rect 16356 6876 16362 6888
rect 17586 6876 17592 6888
rect 17644 6876 17650 6928
rect 18417 6919 18475 6925
rect 18417 6885 18429 6919
rect 18463 6916 18475 6919
rect 18506 6916 18512 6928
rect 18463 6888 18512 6916
rect 18463 6885 18475 6888
rect 18417 6879 18475 6885
rect 18506 6876 18512 6888
rect 18564 6876 18570 6928
rect 19426 6876 19432 6928
rect 19484 6916 19490 6928
rect 19812 6916 19840 6944
rect 19484 6888 19840 6916
rect 19484 6876 19490 6888
rect 13909 6851 13967 6857
rect 12820 6820 13860 6848
rect 10551 6752 11560 6780
rect 11609 6783 11667 6789
rect 10551 6749 10563 6752
rect 10505 6743 10563 6749
rect 11609 6749 11621 6783
rect 11655 6749 11667 6783
rect 11609 6743 11667 6749
rect 7432 6684 7604 6712
rect 7852 6712 7880 6740
rect 8110 6712 8116 6724
rect 7852 6684 8116 6712
rect 7432 6672 7438 6684
rect 8110 6672 8116 6684
rect 8168 6672 8174 6724
rect 8294 6672 8300 6724
rect 8352 6712 8358 6724
rect 8665 6715 8723 6721
rect 8665 6712 8677 6715
rect 8352 6684 8677 6712
rect 8352 6672 8358 6684
rect 8665 6681 8677 6684
rect 8711 6712 8723 6715
rect 10594 6712 10600 6724
rect 8711 6684 10600 6712
rect 8711 6681 8723 6684
rect 8665 6675 8723 6681
rect 10594 6672 10600 6684
rect 10652 6672 10658 6724
rect 10962 6672 10968 6724
rect 11020 6712 11026 6724
rect 11624 6712 11652 6743
rect 11020 6684 11652 6712
rect 11020 6672 11026 6684
rect 8478 6644 8484 6656
rect 7300 6616 8484 6644
rect 8478 6604 8484 6616
rect 8536 6644 8542 6656
rect 8757 6647 8815 6653
rect 8757 6644 8769 6647
rect 8536 6616 8769 6644
rect 8536 6604 8542 6616
rect 8757 6613 8769 6616
rect 8803 6613 8815 6647
rect 8757 6607 8815 6613
rect 9030 6604 9036 6656
rect 9088 6644 9094 6656
rect 9401 6647 9459 6653
rect 9401 6644 9413 6647
rect 9088 6616 9413 6644
rect 9088 6604 9094 6616
rect 9401 6613 9413 6616
rect 9447 6613 9459 6647
rect 9401 6607 9459 6613
rect 9861 6647 9919 6653
rect 9861 6613 9873 6647
rect 9907 6644 9919 6647
rect 10318 6644 10324 6656
rect 9907 6616 10324 6644
rect 9907 6613 9919 6616
rect 9861 6607 9919 6613
rect 10318 6604 10324 6616
rect 10376 6604 10382 6656
rect 10612 6644 10640 6672
rect 12820 6644 12848 6820
rect 13354 6740 13360 6792
rect 13412 6780 13418 6792
rect 13541 6783 13599 6789
rect 13541 6780 13553 6783
rect 13412 6752 13553 6780
rect 13412 6740 13418 6752
rect 13541 6749 13553 6752
rect 13587 6749 13599 6783
rect 13541 6743 13599 6749
rect 13630 6740 13636 6792
rect 13688 6780 13694 6792
rect 13832 6780 13860 6820
rect 13909 6817 13921 6851
rect 13955 6817 13967 6851
rect 13909 6811 13967 6817
rect 13998 6808 14004 6860
rect 14056 6848 14062 6860
rect 14645 6851 14703 6857
rect 14645 6848 14657 6851
rect 14056 6820 14657 6848
rect 14056 6808 14062 6820
rect 14645 6817 14657 6820
rect 14691 6817 14703 6851
rect 17218 6848 17224 6860
rect 14645 6811 14703 6817
rect 14844 6820 17224 6848
rect 14844 6792 14872 6820
rect 14826 6780 14832 6792
rect 13688 6752 13733 6780
rect 13832 6752 14596 6780
rect 14739 6752 14832 6780
rect 13688 6740 13694 6752
rect 13081 6715 13139 6721
rect 13081 6681 13093 6715
rect 13127 6712 13139 6715
rect 14458 6712 14464 6724
rect 13127 6684 14464 6712
rect 13127 6681 13139 6684
rect 13081 6675 13139 6681
rect 14458 6672 14464 6684
rect 14516 6672 14522 6724
rect 14568 6712 14596 6752
rect 14826 6740 14832 6752
rect 14884 6740 14890 6792
rect 15746 6740 15752 6792
rect 15804 6780 15810 6792
rect 16114 6780 16120 6792
rect 15804 6752 16120 6780
rect 15804 6740 15810 6752
rect 16114 6740 16120 6752
rect 16172 6740 16178 6792
rect 16868 6789 16896 6820
rect 17218 6808 17224 6820
rect 17276 6808 17282 6860
rect 17402 6848 17408 6860
rect 17363 6820 17408 6848
rect 17402 6808 17408 6820
rect 17460 6808 17466 6860
rect 16669 6783 16727 6789
rect 16669 6749 16681 6783
rect 16715 6749 16727 6783
rect 16669 6743 16727 6749
rect 16853 6783 16911 6789
rect 16853 6749 16865 6783
rect 16899 6749 16911 6783
rect 16853 6743 16911 6749
rect 16025 6715 16083 6721
rect 16025 6712 16037 6715
rect 14568 6684 16037 6712
rect 16025 6681 16037 6684
rect 16071 6712 16083 6715
rect 16684 6712 16712 6743
rect 17034 6740 17040 6792
rect 17092 6780 17098 6792
rect 17497 6783 17555 6789
rect 17497 6780 17509 6783
rect 17092 6752 17509 6780
rect 17092 6740 17098 6752
rect 17497 6749 17509 6752
rect 17543 6749 17555 6783
rect 17497 6743 17555 6749
rect 17589 6783 17647 6789
rect 17589 6749 17601 6783
rect 17635 6749 17647 6783
rect 17589 6743 17647 6749
rect 16071 6684 16712 6712
rect 16071 6681 16083 6684
rect 16025 6675 16083 6681
rect 17218 6672 17224 6724
rect 17276 6712 17282 6724
rect 17604 6712 17632 6743
rect 18138 6740 18144 6792
rect 18196 6780 18202 6792
rect 18509 6783 18567 6789
rect 18509 6780 18521 6783
rect 18196 6752 18521 6780
rect 18196 6740 18202 6752
rect 18509 6749 18521 6752
rect 18555 6749 18567 6783
rect 18509 6743 18567 6749
rect 18598 6740 18604 6792
rect 18656 6780 18662 6792
rect 18693 6783 18751 6789
rect 18693 6780 18705 6783
rect 18656 6752 18705 6780
rect 18656 6740 18662 6752
rect 18693 6749 18705 6752
rect 18739 6749 18751 6783
rect 18693 6743 18751 6749
rect 19150 6740 19156 6792
rect 19208 6780 19214 6792
rect 19429 6783 19487 6789
rect 19429 6780 19441 6783
rect 19208 6752 19441 6780
rect 19208 6740 19214 6752
rect 19429 6749 19441 6752
rect 19475 6749 19487 6783
rect 19812 6780 19840 6888
rect 20533 6851 20591 6857
rect 20533 6848 20545 6851
rect 20180 6820 20545 6848
rect 20180 6789 20208 6820
rect 20533 6817 20545 6820
rect 20579 6817 20591 6851
rect 20533 6811 20591 6817
rect 20165 6783 20223 6789
rect 20165 6780 20177 6783
rect 19812 6752 20177 6780
rect 19429 6743 19487 6749
rect 20165 6749 20177 6752
rect 20211 6749 20223 6783
rect 20165 6743 20223 6749
rect 20349 6783 20407 6789
rect 20349 6749 20361 6783
rect 20395 6780 20407 6783
rect 20898 6780 20904 6792
rect 20395 6752 20904 6780
rect 20395 6749 20407 6752
rect 20349 6743 20407 6749
rect 20898 6740 20904 6752
rect 20956 6740 20962 6792
rect 17276 6684 17632 6712
rect 18049 6715 18107 6721
rect 17276 6672 17282 6684
rect 18049 6681 18061 6715
rect 18095 6712 18107 6715
rect 18874 6712 18880 6724
rect 18095 6684 18736 6712
rect 18835 6684 18880 6712
rect 18095 6681 18107 6684
rect 18049 6675 18107 6681
rect 18708 6656 18736 6684
rect 18874 6672 18880 6684
rect 18932 6672 18938 6724
rect 19242 6672 19248 6724
rect 19300 6712 19306 6724
rect 19705 6715 19763 6721
rect 19705 6712 19717 6715
rect 19300 6684 19717 6712
rect 19300 6672 19306 6684
rect 19705 6681 19717 6684
rect 19751 6681 19763 6715
rect 21082 6712 21088 6724
rect 21043 6684 21088 6712
rect 19705 6675 19763 6681
rect 21082 6672 21088 6684
rect 21140 6672 21146 6724
rect 12986 6644 12992 6656
rect 10612 6616 12848 6644
rect 12947 6616 12992 6644
rect 12986 6604 12992 6616
rect 13044 6604 13050 6656
rect 13630 6604 13636 6656
rect 13688 6644 13694 6656
rect 13998 6644 14004 6656
rect 13688 6616 14004 6644
rect 13688 6604 13694 6616
rect 13998 6604 14004 6616
rect 14056 6604 14062 6656
rect 14182 6644 14188 6656
rect 14143 6616 14188 6644
rect 14182 6604 14188 6616
rect 14240 6604 14246 6656
rect 15470 6604 15476 6656
rect 15528 6644 15534 6656
rect 15565 6647 15623 6653
rect 15565 6644 15577 6647
rect 15528 6616 15577 6644
rect 15528 6604 15534 6616
rect 15565 6613 15577 6616
rect 15611 6613 15623 6647
rect 15565 6607 15623 6613
rect 16114 6604 16120 6656
rect 16172 6644 16178 6656
rect 16209 6647 16267 6653
rect 16209 6644 16221 6647
rect 16172 6616 16221 6644
rect 16172 6604 16178 6616
rect 16209 6613 16221 6616
rect 16255 6613 16267 6647
rect 16209 6607 16267 6613
rect 17037 6647 17095 6653
rect 17037 6613 17049 6647
rect 17083 6644 17095 6647
rect 17770 6644 17776 6656
rect 17083 6616 17776 6644
rect 17083 6613 17095 6616
rect 17037 6607 17095 6613
rect 17770 6604 17776 6616
rect 17828 6604 17834 6656
rect 17957 6647 18015 6653
rect 17957 6613 17969 6647
rect 18003 6644 18015 6647
rect 18598 6644 18604 6656
rect 18003 6616 18604 6644
rect 18003 6613 18015 6616
rect 17957 6607 18015 6613
rect 18598 6604 18604 6616
rect 18656 6604 18662 6656
rect 18690 6604 18696 6656
rect 18748 6604 18754 6656
rect 19978 6604 19984 6656
rect 20036 6644 20042 6656
rect 20993 6647 21051 6653
rect 20993 6644 21005 6647
rect 20036 6616 21005 6644
rect 20036 6604 20042 6616
rect 20993 6613 21005 6616
rect 21039 6644 21051 6647
rect 22005 6647 22063 6653
rect 22005 6644 22017 6647
rect 21039 6616 22017 6644
rect 21039 6613 21051 6616
rect 20993 6607 21051 6613
rect 22005 6613 22017 6616
rect 22051 6613 22063 6647
rect 22005 6607 22063 6613
rect 1104 6554 21896 6576
rect 1104 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 4575 6554
rect 4627 6502 4639 6554
rect 4691 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 18308 6554
rect 18360 6502 18372 6554
rect 18424 6502 18436 6554
rect 18488 6502 18500 6554
rect 18552 6502 21896 6554
rect 1104 6480 21896 6502
rect 2038 6440 2044 6452
rect 1999 6412 2044 6440
rect 2038 6400 2044 6412
rect 2096 6400 2102 6452
rect 4338 6400 4344 6452
rect 4396 6440 4402 6452
rect 4709 6443 4767 6449
rect 4709 6440 4721 6443
rect 4396 6412 4721 6440
rect 4396 6400 4402 6412
rect 4709 6409 4721 6412
rect 4755 6409 4767 6443
rect 4709 6403 4767 6409
rect 5258 6400 5264 6452
rect 5316 6440 5322 6452
rect 5316 6412 7972 6440
rect 5316 6400 5322 6412
rect 2590 6332 2596 6384
rect 2648 6372 2654 6384
rect 5442 6372 5448 6384
rect 2648 6344 5448 6372
rect 2648 6332 2654 6344
rect 2700 6313 2728 6344
rect 2685 6307 2743 6313
rect 2685 6273 2697 6307
rect 2731 6273 2743 6307
rect 3786 6304 3792 6316
rect 3747 6276 3792 6304
rect 2685 6267 2743 6273
rect 3786 6264 3792 6276
rect 3844 6264 3850 6316
rect 4982 6264 4988 6316
rect 5040 6304 5046 6316
rect 5276 6313 5304 6344
rect 5442 6332 5448 6344
rect 5500 6332 5506 6384
rect 5813 6375 5871 6381
rect 5813 6341 5825 6375
rect 5859 6372 5871 6375
rect 5994 6372 6000 6384
rect 5859 6344 6000 6372
rect 5859 6341 5871 6344
rect 5813 6335 5871 6341
rect 5994 6332 6000 6344
rect 6052 6372 6058 6384
rect 6052 6344 7144 6372
rect 6052 6332 6058 6344
rect 5169 6307 5227 6313
rect 5169 6304 5181 6307
rect 5040 6276 5181 6304
rect 5040 6264 5046 6276
rect 5169 6273 5181 6276
rect 5215 6273 5227 6307
rect 5169 6267 5227 6273
rect 5261 6307 5319 6313
rect 5261 6273 5273 6307
rect 5307 6273 5319 6307
rect 5261 6267 5319 6273
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6304 6607 6307
rect 6914 6304 6920 6316
rect 6595 6276 6920 6304
rect 6595 6273 6607 6276
rect 6549 6267 6607 6273
rect 6914 6264 6920 6276
rect 6972 6264 6978 6316
rect 1670 6196 1676 6248
rect 1728 6236 1734 6248
rect 2409 6239 2467 6245
rect 2409 6236 2421 6239
rect 1728 6208 2421 6236
rect 1728 6196 1734 6208
rect 2409 6205 2421 6208
rect 2455 6205 2467 6239
rect 2409 6199 2467 6205
rect 3510 6196 3516 6248
rect 3568 6236 3574 6248
rect 5537 6239 5595 6245
rect 5537 6236 5549 6239
rect 3568 6208 5549 6236
rect 3568 6196 3574 6208
rect 5537 6205 5549 6208
rect 5583 6236 5595 6239
rect 6362 6236 6368 6248
rect 5583 6208 6368 6236
rect 5583 6205 5595 6208
rect 5537 6199 5595 6205
rect 6362 6196 6368 6208
rect 6420 6196 6426 6248
rect 7116 6236 7144 6344
rect 7374 6304 7380 6316
rect 7335 6276 7380 6304
rect 7374 6264 7380 6276
rect 7432 6264 7438 6316
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 7116 6208 7297 6236
rect 7285 6205 7297 6208
rect 7331 6205 7343 6239
rect 7944 6236 7972 6412
rect 9582 6400 9588 6452
rect 9640 6440 9646 6452
rect 10686 6440 10692 6452
rect 9640 6412 10692 6440
rect 9640 6400 9646 6412
rect 10686 6400 10692 6412
rect 10744 6400 10750 6452
rect 11977 6443 12035 6449
rect 11977 6440 11989 6443
rect 11532 6412 11989 6440
rect 8202 6332 8208 6384
rect 8260 6372 8266 6384
rect 11422 6372 11428 6384
rect 8260 6344 11428 6372
rect 8260 6332 8266 6344
rect 11422 6332 11428 6344
rect 11480 6332 11486 6384
rect 8297 6307 8355 6313
rect 8297 6273 8309 6307
rect 8343 6304 8355 6307
rect 8386 6304 8392 6316
rect 8343 6276 8392 6304
rect 8343 6273 8355 6276
rect 8297 6267 8355 6273
rect 8386 6264 8392 6276
rect 8444 6304 8450 6316
rect 9125 6307 9183 6313
rect 9125 6304 9137 6307
rect 8444 6276 9137 6304
rect 8444 6264 8450 6276
rect 9125 6273 9137 6276
rect 9171 6273 9183 6307
rect 9125 6267 9183 6273
rect 10229 6307 10287 6313
rect 10229 6273 10241 6307
rect 10275 6304 10287 6307
rect 10778 6304 10784 6316
rect 10275 6276 10784 6304
rect 10275 6273 10287 6276
rect 10229 6267 10287 6273
rect 10778 6264 10784 6276
rect 10836 6264 10842 6316
rect 11532 6313 11560 6412
rect 11977 6409 11989 6412
rect 12023 6440 12035 6443
rect 12526 6440 12532 6452
rect 12023 6412 12532 6440
rect 12023 6409 12035 6412
rect 11977 6403 12035 6409
rect 12526 6400 12532 6412
rect 12584 6400 12590 6452
rect 13354 6440 13360 6452
rect 13315 6412 13360 6440
rect 13354 6400 13360 6412
rect 13412 6400 13418 6452
rect 14090 6400 14096 6452
rect 14148 6400 14154 6452
rect 14182 6400 14188 6452
rect 14240 6440 14246 6452
rect 14240 6412 15240 6440
rect 14240 6400 14246 6412
rect 12437 6375 12495 6381
rect 12437 6341 12449 6375
rect 12483 6372 12495 6375
rect 13538 6372 13544 6384
rect 12483 6344 13544 6372
rect 12483 6341 12495 6344
rect 12437 6335 12495 6341
rect 13538 6332 13544 6344
rect 13596 6332 13602 6384
rect 11517 6307 11575 6313
rect 11517 6273 11529 6307
rect 11563 6273 11575 6307
rect 11698 6304 11704 6316
rect 11659 6276 11704 6304
rect 11517 6267 11575 6273
rect 11698 6264 11704 6276
rect 11756 6264 11762 6316
rect 12710 6264 12716 6316
rect 12768 6304 12774 6316
rect 12897 6307 12955 6313
rect 12897 6304 12909 6307
rect 12768 6276 12909 6304
rect 12768 6264 12774 6276
rect 12897 6273 12909 6276
rect 12943 6273 12955 6307
rect 12897 6267 12955 6273
rect 12986 6264 12992 6316
rect 13044 6304 13050 6316
rect 14108 6304 14136 6400
rect 13044 6276 13089 6304
rect 13464 6276 14136 6304
rect 15212 6304 15240 6412
rect 15286 6400 15292 6452
rect 15344 6440 15350 6452
rect 15565 6443 15623 6449
rect 15565 6440 15577 6443
rect 15344 6412 15577 6440
rect 15344 6400 15350 6412
rect 15565 6409 15577 6412
rect 15611 6440 15623 6443
rect 18138 6440 18144 6452
rect 15611 6412 16896 6440
rect 18099 6412 18144 6440
rect 15611 6409 15623 6412
rect 15565 6403 15623 6409
rect 15749 6375 15807 6381
rect 15749 6341 15761 6375
rect 15795 6372 15807 6375
rect 16758 6372 16764 6384
rect 15795 6344 16764 6372
rect 15795 6341 15807 6344
rect 15749 6335 15807 6341
rect 16758 6332 16764 6344
rect 16816 6332 16822 6384
rect 16209 6307 16267 6313
rect 16209 6304 16221 6307
rect 15212 6276 16221 6304
rect 13044 6264 13050 6276
rect 9033 6239 9091 6245
rect 9033 6236 9045 6239
rect 7944 6208 9045 6236
rect 7285 6199 7343 6205
rect 9033 6205 9045 6208
rect 9079 6236 9091 6239
rect 10965 6239 11023 6245
rect 9079 6208 10548 6236
rect 9079 6205 9091 6208
rect 9033 6199 9091 6205
rect 1486 6128 1492 6180
rect 1544 6168 1550 6180
rect 1581 6171 1639 6177
rect 1581 6168 1593 6171
rect 1544 6140 1593 6168
rect 1544 6128 1550 6140
rect 1581 6137 1593 6140
rect 1627 6168 1639 6171
rect 2961 6171 3019 6177
rect 1627 6140 2544 6168
rect 1627 6137 1639 6140
rect 1581 6131 1639 6137
rect 1762 6100 1768 6112
rect 1723 6072 1768 6100
rect 1762 6060 1768 6072
rect 1820 6060 1826 6112
rect 2516 6109 2544 6140
rect 2961 6137 2973 6171
rect 3007 6168 3019 6171
rect 3050 6168 3056 6180
rect 3007 6140 3056 6168
rect 3007 6137 3019 6140
rect 2961 6131 3019 6137
rect 3050 6128 3056 6140
rect 3108 6128 3114 6180
rect 3694 6128 3700 6180
rect 3752 6168 3758 6180
rect 4154 6168 4160 6180
rect 3752 6140 4160 6168
rect 3752 6128 3758 6140
rect 4154 6128 4160 6140
rect 4212 6128 4218 6180
rect 5077 6171 5135 6177
rect 5077 6137 5089 6171
rect 5123 6168 5135 6171
rect 7193 6171 7251 6177
rect 5123 6140 6868 6168
rect 5123 6137 5135 6140
rect 5077 6131 5135 6137
rect 2501 6103 2559 6109
rect 2501 6069 2513 6103
rect 2547 6100 2559 6103
rect 2682 6100 2688 6112
rect 2547 6072 2688 6100
rect 2547 6069 2559 6072
rect 2501 6063 2559 6069
rect 2682 6060 2688 6072
rect 2740 6060 2746 6112
rect 3142 6100 3148 6112
rect 3103 6072 3148 6100
rect 3142 6060 3148 6072
rect 3200 6060 3206 6112
rect 3510 6100 3516 6112
rect 3471 6072 3516 6100
rect 3510 6060 3516 6072
rect 3568 6060 3574 6112
rect 3605 6103 3663 6109
rect 3605 6069 3617 6103
rect 3651 6100 3663 6103
rect 4338 6100 4344 6112
rect 3651 6072 4344 6100
rect 3651 6069 3663 6072
rect 3605 6063 3663 6069
rect 4338 6060 4344 6072
rect 4396 6060 4402 6112
rect 5902 6100 5908 6112
rect 5863 6072 5908 6100
rect 5902 6060 5908 6072
rect 5960 6060 5966 6112
rect 6270 6100 6276 6112
rect 6231 6072 6276 6100
rect 6270 6060 6276 6072
rect 6328 6060 6334 6112
rect 6840 6109 6868 6140
rect 7193 6137 7205 6171
rect 7239 6168 7251 6171
rect 7834 6168 7840 6180
rect 7239 6140 7840 6168
rect 7239 6137 7251 6140
rect 7193 6131 7251 6137
rect 7834 6128 7840 6140
rect 7892 6128 7898 6180
rect 8110 6168 8116 6180
rect 8071 6140 8116 6168
rect 8110 6128 8116 6140
rect 8168 6128 8174 6180
rect 9953 6171 10011 6177
rect 9953 6137 9965 6171
rect 9999 6168 10011 6171
rect 10318 6168 10324 6180
rect 9999 6140 10324 6168
rect 9999 6137 10011 6140
rect 9953 6131 10011 6137
rect 10318 6128 10324 6140
rect 10376 6128 10382 6180
rect 10520 6177 10548 6208
rect 10965 6205 10977 6239
rect 11011 6236 11023 6239
rect 11146 6236 11152 6248
rect 11011 6208 11152 6236
rect 11011 6205 11023 6208
rect 10965 6199 11023 6205
rect 11146 6196 11152 6208
rect 11204 6236 11210 6248
rect 11425 6239 11483 6245
rect 11425 6236 11437 6239
rect 11204 6208 11437 6236
rect 11204 6196 11210 6208
rect 11425 6205 11437 6208
rect 11471 6205 11483 6239
rect 11425 6199 11483 6205
rect 10505 6171 10563 6177
rect 10505 6137 10517 6171
rect 10551 6168 10563 6171
rect 12618 6168 12624 6180
rect 10551 6140 12624 6168
rect 10551 6137 10563 6140
rect 10505 6131 10563 6137
rect 12618 6128 12624 6140
rect 12676 6128 12682 6180
rect 12805 6171 12863 6177
rect 12805 6137 12817 6171
rect 12851 6168 12863 6171
rect 13464 6168 13492 6276
rect 16209 6273 16221 6276
rect 16255 6273 16267 6307
rect 16209 6267 16267 6273
rect 16393 6307 16451 6313
rect 16393 6273 16405 6307
rect 16439 6304 16451 6307
rect 16868 6304 16896 6412
rect 18138 6400 18144 6412
rect 18196 6400 18202 6452
rect 20625 6443 20683 6449
rect 20625 6409 20637 6443
rect 20671 6440 20683 6443
rect 20898 6440 20904 6452
rect 20671 6412 20904 6440
rect 20671 6409 20683 6412
rect 20625 6403 20683 6409
rect 20898 6400 20904 6412
rect 20956 6400 20962 6452
rect 17954 6332 17960 6384
rect 18012 6372 18018 6384
rect 18690 6372 18696 6384
rect 18012 6344 18696 6372
rect 18012 6332 18018 6344
rect 18690 6332 18696 6344
rect 18748 6372 18754 6384
rect 18748 6344 19288 6372
rect 18748 6332 18754 6344
rect 17218 6304 17224 6316
rect 16439 6276 17224 6304
rect 16439 6273 16451 6276
rect 16393 6267 16451 6273
rect 17218 6264 17224 6276
rect 17276 6264 17282 6316
rect 17402 6304 17408 6316
rect 17363 6276 17408 6304
rect 17402 6264 17408 6276
rect 17460 6264 17466 6316
rect 19260 6313 19288 6344
rect 20346 6332 20352 6384
rect 20404 6372 20410 6384
rect 21082 6372 21088 6384
rect 20404 6344 21088 6372
rect 20404 6332 20410 6344
rect 21082 6332 21088 6344
rect 21140 6332 21146 6384
rect 18785 6307 18843 6313
rect 18785 6273 18797 6307
rect 18831 6273 18843 6307
rect 18785 6267 18843 6273
rect 19245 6307 19303 6313
rect 19245 6273 19257 6307
rect 19291 6273 19303 6307
rect 19245 6267 19303 6273
rect 14185 6239 14243 6245
rect 14185 6236 14197 6239
rect 12851 6140 13492 6168
rect 13556 6208 14197 6236
rect 12851 6137 12863 6140
rect 12805 6131 12863 6137
rect 6825 6103 6883 6109
rect 6825 6069 6837 6103
rect 6871 6069 6883 6103
rect 7650 6100 7656 6112
rect 7611 6072 7656 6100
rect 6825 6063 6883 6069
rect 7650 6060 7656 6072
rect 7708 6060 7714 6112
rect 7742 6060 7748 6112
rect 7800 6100 7806 6112
rect 8021 6103 8079 6109
rect 8021 6100 8033 6103
rect 7800 6072 8033 6100
rect 7800 6060 7806 6072
rect 8021 6069 8033 6072
rect 8067 6069 8079 6103
rect 8021 6063 8079 6069
rect 8573 6103 8631 6109
rect 8573 6069 8585 6103
rect 8619 6100 8631 6103
rect 8754 6100 8760 6112
rect 8619 6072 8760 6100
rect 8619 6069 8631 6072
rect 8573 6063 8631 6069
rect 8754 6060 8760 6072
rect 8812 6060 8818 6112
rect 8941 6103 8999 6109
rect 8941 6069 8953 6103
rect 8987 6100 8999 6103
rect 9214 6100 9220 6112
rect 8987 6072 9220 6100
rect 8987 6069 8999 6072
rect 8941 6063 8999 6069
rect 9214 6060 9220 6072
rect 9272 6100 9278 6112
rect 9401 6103 9459 6109
rect 9401 6100 9413 6103
rect 9272 6072 9413 6100
rect 9272 6060 9278 6072
rect 9401 6069 9413 6072
rect 9447 6069 9459 6103
rect 9401 6063 9459 6069
rect 9585 6103 9643 6109
rect 9585 6069 9597 6103
rect 9631 6100 9643 6103
rect 9858 6100 9864 6112
rect 9631 6072 9864 6100
rect 9631 6069 9643 6072
rect 9585 6063 9643 6069
rect 9858 6060 9864 6072
rect 9916 6060 9922 6112
rect 10042 6100 10048 6112
rect 10003 6072 10048 6100
rect 10042 6060 10048 6072
rect 10100 6060 10106 6112
rect 10962 6060 10968 6112
rect 11020 6100 11026 6112
rect 11057 6103 11115 6109
rect 11057 6100 11069 6103
rect 11020 6072 11069 6100
rect 11020 6060 11026 6072
rect 11057 6069 11069 6072
rect 11103 6069 11115 6103
rect 11057 6063 11115 6069
rect 12434 6060 12440 6112
rect 12492 6100 12498 6112
rect 13556 6100 13584 6208
rect 14185 6205 14197 6208
rect 14231 6205 14243 6239
rect 14185 6199 14243 6205
rect 14452 6239 14510 6245
rect 14452 6205 14464 6239
rect 14498 6236 14510 6239
rect 14826 6236 14832 6248
rect 14498 6208 14832 6236
rect 14498 6205 14510 6208
rect 14452 6199 14510 6205
rect 14826 6196 14832 6208
rect 14884 6196 14890 6248
rect 16114 6236 16120 6248
rect 16075 6208 16120 6236
rect 16114 6196 16120 6208
rect 16172 6196 16178 6248
rect 13817 6171 13875 6177
rect 13817 6137 13829 6171
rect 13863 6168 13875 6171
rect 13998 6168 14004 6180
rect 13863 6140 14004 6168
rect 13863 6137 13875 6140
rect 13817 6131 13875 6137
rect 13998 6128 14004 6140
rect 14056 6128 14062 6180
rect 15838 6128 15844 6180
rect 15896 6168 15902 6180
rect 16945 6171 17003 6177
rect 16945 6168 16957 6171
rect 15896 6140 16957 6168
rect 15896 6128 15902 6140
rect 16945 6137 16957 6140
rect 16991 6137 17003 6171
rect 16945 6131 17003 6137
rect 17678 6128 17684 6180
rect 17736 6168 17742 6180
rect 17773 6171 17831 6177
rect 17773 6168 17785 6171
rect 17736 6140 17785 6168
rect 17736 6128 17742 6140
rect 17773 6137 17785 6140
rect 17819 6168 17831 6171
rect 18601 6171 18659 6177
rect 18601 6168 18613 6171
rect 17819 6140 18613 6168
rect 17819 6137 17831 6140
rect 17773 6131 17831 6137
rect 18601 6137 18613 6140
rect 18647 6137 18659 6171
rect 18800 6168 18828 6267
rect 19512 6171 19570 6177
rect 19512 6168 19524 6171
rect 18800 6140 19524 6168
rect 18601 6131 18659 6137
rect 19512 6137 19524 6140
rect 19558 6168 19570 6171
rect 20070 6168 20076 6180
rect 19558 6140 20076 6168
rect 19558 6137 19570 6140
rect 19512 6131 19570 6137
rect 20070 6128 20076 6140
rect 20128 6128 20134 6180
rect 12492 6072 13584 6100
rect 12492 6060 12498 6072
rect 13630 6060 13636 6112
rect 13688 6100 13694 6112
rect 13688 6072 13733 6100
rect 13688 6060 13694 6072
rect 13906 6060 13912 6112
rect 13964 6100 13970 6112
rect 14093 6103 14151 6109
rect 14093 6100 14105 6103
rect 13964 6072 14105 6100
rect 13964 6060 13970 6072
rect 14093 6069 14105 6072
rect 14139 6100 14151 6103
rect 15194 6100 15200 6112
rect 14139 6072 15200 6100
rect 14139 6069 14151 6072
rect 14093 6063 14151 6069
rect 15194 6060 15200 6072
rect 15252 6060 15258 6112
rect 16577 6103 16635 6109
rect 16577 6069 16589 6103
rect 16623 6100 16635 6103
rect 16850 6100 16856 6112
rect 16623 6072 16856 6100
rect 16623 6069 16635 6072
rect 16577 6063 16635 6069
rect 16850 6060 16856 6072
rect 16908 6060 16914 6112
rect 17034 6060 17040 6112
rect 17092 6100 17098 6112
rect 17092 6072 17137 6100
rect 17092 6060 17098 6072
rect 18138 6060 18144 6112
rect 18196 6100 18202 6112
rect 18509 6103 18567 6109
rect 18509 6100 18521 6103
rect 18196 6072 18521 6100
rect 18196 6060 18202 6072
rect 18509 6069 18521 6072
rect 18555 6069 18567 6103
rect 18509 6063 18567 6069
rect 1104 6010 21896 6032
rect 1104 5958 7912 6010
rect 7964 5958 7976 6010
rect 8028 5958 8040 6010
rect 8092 5958 8104 6010
rect 8156 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 15035 6010
rect 15087 5958 21896 6010
rect 1104 5936 21896 5958
rect 2314 5896 2320 5908
rect 2275 5868 2320 5896
rect 2314 5856 2320 5868
rect 2372 5856 2378 5908
rect 2685 5899 2743 5905
rect 2685 5865 2697 5899
rect 2731 5896 2743 5899
rect 3142 5896 3148 5908
rect 2731 5868 3148 5896
rect 2731 5865 2743 5868
rect 2685 5859 2743 5865
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 4062 5856 4068 5908
rect 4120 5896 4126 5908
rect 6181 5899 6239 5905
rect 4120 5868 6132 5896
rect 4120 5856 4126 5868
rect 1854 5788 1860 5840
rect 1912 5828 1918 5840
rect 1949 5831 2007 5837
rect 1949 5828 1961 5831
rect 1912 5800 1961 5828
rect 1912 5788 1918 5800
rect 1949 5797 1961 5800
rect 1995 5797 2007 5831
rect 1949 5791 2007 5797
rect 2777 5831 2835 5837
rect 2777 5797 2789 5831
rect 2823 5828 2835 5831
rect 5534 5828 5540 5840
rect 2823 5800 5540 5828
rect 2823 5797 2835 5800
rect 2777 5791 2835 5797
rect 5534 5788 5540 5800
rect 5592 5788 5598 5840
rect 6104 5828 6132 5868
rect 6181 5865 6193 5899
rect 6227 5896 6239 5899
rect 6270 5896 6276 5908
rect 6227 5868 6276 5896
rect 6227 5865 6239 5868
rect 6181 5859 6239 5865
rect 6270 5856 6276 5868
rect 6328 5856 6334 5908
rect 6733 5899 6791 5905
rect 6733 5865 6745 5899
rect 6779 5896 6791 5899
rect 7006 5896 7012 5908
rect 6779 5868 7012 5896
rect 6779 5865 6791 5868
rect 6733 5859 6791 5865
rect 7006 5856 7012 5868
rect 7064 5856 7070 5908
rect 7469 5899 7527 5905
rect 7469 5865 7481 5899
rect 7515 5896 7527 5899
rect 7742 5896 7748 5908
rect 7515 5868 7748 5896
rect 7515 5865 7527 5868
rect 7469 5859 7527 5865
rect 7742 5856 7748 5868
rect 7800 5856 7806 5908
rect 8570 5896 8576 5908
rect 8531 5868 8576 5896
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 9674 5896 9680 5908
rect 8680 5868 9680 5896
rect 7101 5831 7159 5837
rect 7101 5828 7113 5831
rect 6104 5800 7113 5828
rect 7101 5797 7113 5800
rect 7147 5828 7159 5831
rect 8113 5831 8171 5837
rect 8113 5828 8125 5831
rect 7147 5800 8125 5828
rect 7147 5797 7159 5800
rect 7101 5791 7159 5797
rect 8113 5797 8125 5800
rect 8159 5828 8171 5831
rect 8680 5828 8708 5868
rect 9674 5856 9680 5868
rect 9732 5856 9738 5908
rect 10686 5856 10692 5908
rect 10744 5896 10750 5908
rect 11609 5899 11667 5905
rect 11609 5896 11621 5899
rect 10744 5868 11621 5896
rect 10744 5856 10750 5868
rect 11609 5865 11621 5868
rect 11655 5865 11667 5899
rect 11609 5859 11667 5865
rect 11974 5856 11980 5908
rect 12032 5896 12038 5908
rect 12069 5899 12127 5905
rect 12069 5896 12081 5899
rect 12032 5868 12081 5896
rect 12032 5856 12038 5868
rect 12069 5865 12081 5868
rect 12115 5865 12127 5899
rect 12069 5859 12127 5865
rect 12345 5899 12403 5905
rect 12345 5865 12357 5899
rect 12391 5896 12403 5899
rect 14642 5896 14648 5908
rect 12391 5868 14648 5896
rect 12391 5865 12403 5868
rect 12345 5859 12403 5865
rect 11517 5831 11575 5837
rect 11517 5828 11529 5831
rect 8159 5800 8708 5828
rect 8864 5800 11529 5828
rect 8159 5797 8171 5800
rect 8113 5791 8171 5797
rect 1670 5760 1676 5772
rect 1631 5732 1676 5760
rect 1670 5720 1676 5732
rect 1728 5720 1734 5772
rect 3513 5763 3571 5769
rect 3513 5729 3525 5763
rect 3559 5760 3571 5763
rect 3970 5760 3976 5772
rect 3559 5732 3976 5760
rect 3559 5729 3571 5732
rect 3513 5723 3571 5729
rect 3970 5720 3976 5732
rect 4028 5720 4034 5772
rect 4424 5763 4482 5769
rect 4424 5760 4436 5763
rect 4080 5732 4436 5760
rect 2869 5695 2927 5701
rect 2869 5661 2881 5695
rect 2915 5661 2927 5695
rect 2869 5655 2927 5661
rect 2884 5624 2912 5655
rect 2958 5652 2964 5704
rect 3016 5692 3022 5704
rect 3605 5695 3663 5701
rect 3605 5692 3617 5695
rect 3016 5664 3617 5692
rect 3016 5652 3022 5664
rect 3605 5661 3617 5664
rect 3651 5661 3663 5695
rect 3605 5655 3663 5661
rect 3789 5695 3847 5701
rect 3789 5661 3801 5695
rect 3835 5692 3847 5695
rect 4080 5692 4108 5732
rect 4424 5729 4436 5732
rect 4470 5760 4482 5763
rect 6641 5763 6699 5769
rect 4470 5732 5396 5760
rect 4470 5729 4482 5732
rect 4424 5723 4482 5729
rect 5368 5704 5396 5732
rect 6641 5729 6653 5763
rect 6687 5760 6699 5763
rect 7006 5760 7012 5772
rect 6687 5732 7012 5760
rect 6687 5729 6699 5732
rect 6641 5723 6699 5729
rect 7006 5720 7012 5732
rect 7064 5720 7070 5772
rect 7834 5720 7840 5772
rect 7892 5760 7898 5772
rect 8864 5760 8892 5800
rect 11517 5797 11529 5800
rect 11563 5828 11575 5831
rect 12360 5828 12388 5859
rect 14642 5856 14648 5868
rect 14700 5856 14706 5908
rect 15749 5899 15807 5905
rect 15749 5865 15761 5899
rect 15795 5896 15807 5899
rect 15838 5896 15844 5908
rect 15795 5868 15844 5896
rect 15795 5865 15807 5868
rect 15749 5859 15807 5865
rect 15838 5856 15844 5868
rect 15896 5856 15902 5908
rect 15930 5856 15936 5908
rect 15988 5896 15994 5908
rect 16209 5899 16267 5905
rect 16209 5896 16221 5899
rect 15988 5868 16221 5896
rect 15988 5856 15994 5868
rect 16209 5865 16221 5868
rect 16255 5896 16267 5899
rect 16577 5899 16635 5905
rect 16577 5896 16589 5899
rect 16255 5868 16589 5896
rect 16255 5865 16267 5868
rect 16209 5859 16267 5865
rect 16577 5865 16589 5868
rect 16623 5896 16635 5899
rect 16666 5896 16672 5908
rect 16623 5868 16672 5896
rect 16623 5865 16635 5868
rect 16577 5859 16635 5865
rect 16666 5856 16672 5868
rect 16724 5856 16730 5908
rect 16761 5899 16819 5905
rect 16761 5865 16773 5899
rect 16807 5896 16819 5899
rect 17034 5896 17040 5908
rect 16807 5868 17040 5896
rect 16807 5865 16819 5868
rect 16761 5859 16819 5865
rect 17034 5856 17040 5868
rect 17092 5856 17098 5908
rect 17221 5899 17279 5905
rect 17221 5865 17233 5899
rect 17267 5896 17279 5899
rect 17310 5896 17316 5908
rect 17267 5868 17316 5896
rect 17267 5865 17279 5868
rect 17221 5859 17279 5865
rect 17310 5856 17316 5868
rect 17368 5856 17374 5908
rect 17586 5896 17592 5908
rect 17547 5868 17592 5896
rect 17586 5856 17592 5868
rect 17644 5856 17650 5908
rect 17770 5856 17776 5908
rect 17828 5896 17834 5908
rect 17957 5899 18015 5905
rect 17957 5896 17969 5899
rect 17828 5868 17969 5896
rect 17828 5856 17834 5868
rect 17957 5865 17969 5868
rect 18003 5865 18015 5899
rect 17957 5859 18015 5865
rect 18138 5856 18144 5908
rect 18196 5896 18202 5908
rect 18417 5899 18475 5905
rect 18417 5896 18429 5899
rect 18196 5868 18429 5896
rect 18196 5856 18202 5868
rect 18417 5865 18429 5868
rect 18463 5865 18475 5899
rect 20070 5896 20076 5908
rect 20031 5868 20076 5896
rect 18417 5859 18475 5865
rect 20070 5856 20076 5868
rect 20128 5856 20134 5908
rect 11563 5800 12388 5828
rect 12796 5831 12854 5837
rect 11563 5797 11575 5800
rect 11517 5791 11575 5797
rect 12796 5797 12808 5831
rect 12842 5828 12854 5831
rect 12986 5828 12992 5840
rect 12842 5800 12992 5828
rect 12842 5797 12854 5800
rect 12796 5791 12854 5797
rect 12986 5788 12992 5800
rect 13044 5788 13050 5840
rect 19978 5828 19984 5840
rect 18248 5800 19984 5828
rect 7892 5732 8892 5760
rect 8941 5763 8999 5769
rect 7892 5720 7898 5732
rect 8941 5729 8953 5763
rect 8987 5760 8999 5763
rect 9490 5760 9496 5772
rect 8987 5732 9496 5760
rect 8987 5729 8999 5732
rect 8941 5723 8999 5729
rect 9490 5720 9496 5732
rect 9548 5720 9554 5772
rect 9944 5763 10002 5769
rect 9944 5729 9956 5763
rect 9990 5760 10002 5763
rect 10318 5760 10324 5772
rect 9990 5732 10324 5760
rect 9990 5729 10002 5732
rect 9944 5723 10002 5729
rect 10318 5720 10324 5732
rect 10376 5760 10382 5772
rect 10376 5732 11744 5760
rect 10376 5720 10382 5732
rect 11716 5704 11744 5732
rect 12434 5720 12440 5772
rect 12492 5760 12498 5772
rect 12529 5763 12587 5769
rect 12529 5760 12541 5763
rect 12492 5732 12541 5760
rect 12492 5720 12498 5732
rect 12529 5729 12541 5732
rect 12575 5760 12587 5763
rect 12618 5760 12624 5772
rect 12575 5732 12624 5760
rect 12575 5729 12587 5732
rect 12529 5723 12587 5729
rect 12618 5720 12624 5732
rect 12676 5720 12682 5772
rect 13722 5720 13728 5772
rect 13780 5760 13786 5772
rect 14001 5763 14059 5769
rect 14001 5760 14013 5763
rect 13780 5732 14013 5760
rect 13780 5720 13786 5732
rect 14001 5729 14013 5732
rect 14047 5729 14059 5763
rect 14737 5763 14795 5769
rect 14737 5760 14749 5763
rect 14001 5723 14059 5729
rect 14200 5732 14749 5760
rect 3835 5664 4108 5692
rect 4157 5695 4215 5701
rect 3835 5661 3847 5664
rect 3789 5655 3847 5661
rect 4157 5661 4169 5695
rect 4203 5661 4215 5695
rect 4157 5655 4215 5661
rect 3050 5624 3056 5636
rect 2884 5596 3056 5624
rect 3050 5584 3056 5596
rect 3108 5584 3114 5636
rect 3145 5627 3203 5633
rect 3145 5593 3157 5627
rect 3191 5624 3203 5627
rect 3510 5624 3516 5636
rect 3191 5596 3516 5624
rect 3191 5593 3203 5596
rect 3145 5587 3203 5593
rect 3510 5584 3516 5596
rect 3568 5584 3574 5636
rect 3694 5584 3700 5636
rect 3752 5624 3758 5636
rect 3878 5624 3884 5636
rect 3752 5596 3884 5624
rect 3752 5584 3758 5596
rect 3878 5584 3884 5596
rect 3936 5624 3942 5636
rect 4172 5624 4200 5655
rect 5350 5652 5356 5704
rect 5408 5692 5414 5704
rect 6822 5692 6828 5704
rect 5408 5664 6828 5692
rect 5408 5652 5414 5664
rect 6822 5652 6828 5664
rect 6880 5652 6886 5704
rect 7282 5652 7288 5704
rect 7340 5692 7346 5704
rect 8205 5695 8263 5701
rect 8205 5692 8217 5695
rect 7340 5664 8217 5692
rect 7340 5652 7346 5664
rect 8205 5661 8217 5664
rect 8251 5661 8263 5695
rect 8386 5692 8392 5704
rect 8347 5664 8392 5692
rect 8205 5655 8263 5661
rect 8386 5652 8392 5664
rect 8444 5692 8450 5704
rect 8570 5692 8576 5704
rect 8444 5664 8576 5692
rect 8444 5652 8450 5664
rect 8570 5652 8576 5664
rect 8628 5652 8634 5704
rect 9030 5692 9036 5704
rect 8991 5664 9036 5692
rect 9030 5652 9036 5664
rect 9088 5652 9094 5704
rect 9125 5695 9183 5701
rect 9125 5661 9137 5695
rect 9171 5661 9183 5695
rect 9125 5655 9183 5661
rect 3936 5596 4200 5624
rect 5537 5627 5595 5633
rect 3936 5584 3942 5596
rect 5537 5593 5549 5627
rect 5583 5624 5595 5627
rect 6178 5624 6184 5636
rect 5583 5596 6184 5624
rect 5583 5593 5595 5596
rect 5537 5587 5595 5593
rect 6178 5584 6184 5596
rect 6236 5584 6242 5636
rect 6730 5584 6736 5636
rect 6788 5624 6794 5636
rect 9140 5624 9168 5655
rect 9398 5652 9404 5704
rect 9456 5692 9462 5704
rect 9677 5695 9735 5701
rect 9677 5692 9689 5695
rect 9456 5664 9689 5692
rect 9456 5652 9462 5664
rect 9677 5661 9689 5664
rect 9723 5661 9735 5695
rect 11698 5692 11704 5704
rect 11659 5664 11704 5692
rect 9677 5655 9735 5661
rect 11698 5652 11704 5664
rect 11756 5652 11762 5704
rect 6788 5596 9168 5624
rect 6788 5584 6794 5596
rect 10962 5584 10968 5636
rect 11020 5624 11026 5636
rect 14200 5633 14228 5732
rect 14737 5729 14749 5732
rect 14783 5729 14795 5763
rect 14737 5723 14795 5729
rect 15470 5720 15476 5772
rect 15528 5760 15534 5772
rect 16117 5763 16175 5769
rect 16117 5760 16129 5763
rect 15528 5732 16129 5760
rect 15528 5720 15534 5732
rect 16117 5729 16129 5732
rect 16163 5729 16175 5763
rect 17126 5760 17132 5772
rect 17087 5732 17132 5760
rect 16117 5723 16175 5729
rect 17126 5720 17132 5732
rect 17184 5720 17190 5772
rect 17402 5720 17408 5772
rect 17460 5760 17466 5772
rect 17460 5732 18184 5760
rect 17460 5720 17466 5732
rect 14829 5695 14887 5701
rect 14829 5661 14841 5695
rect 14875 5661 14887 5695
rect 14829 5655 14887 5661
rect 15013 5695 15071 5701
rect 15013 5661 15025 5695
rect 15059 5692 15071 5695
rect 15286 5692 15292 5704
rect 15059 5664 15292 5692
rect 15059 5661 15071 5664
rect 15013 5655 15071 5661
rect 11149 5627 11207 5633
rect 11149 5624 11161 5627
rect 11020 5596 11161 5624
rect 11020 5584 11026 5596
rect 11149 5593 11161 5596
rect 11195 5593 11207 5627
rect 14185 5627 14243 5633
rect 14185 5624 14197 5627
rect 11149 5587 11207 5593
rect 13464 5596 14197 5624
rect 5718 5556 5724 5568
rect 5679 5528 5724 5556
rect 5718 5516 5724 5528
rect 5776 5516 5782 5568
rect 6270 5556 6276 5568
rect 6231 5528 6276 5556
rect 6270 5516 6276 5528
rect 6328 5516 6334 5568
rect 7742 5556 7748 5568
rect 7703 5528 7748 5556
rect 7742 5516 7748 5528
rect 7800 5516 7806 5568
rect 8018 5516 8024 5568
rect 8076 5556 8082 5568
rect 8754 5556 8760 5568
rect 8076 5528 8760 5556
rect 8076 5516 8082 5528
rect 8754 5516 8760 5528
rect 8812 5516 8818 5568
rect 9490 5556 9496 5568
rect 9451 5528 9496 5556
rect 9490 5516 9496 5528
rect 9548 5516 9554 5568
rect 9582 5516 9588 5568
rect 9640 5556 9646 5568
rect 10686 5556 10692 5568
rect 9640 5528 10692 5556
rect 9640 5516 9646 5528
rect 10686 5516 10692 5528
rect 10744 5516 10750 5568
rect 10778 5516 10784 5568
rect 10836 5556 10842 5568
rect 11057 5559 11115 5565
rect 11057 5556 11069 5559
rect 10836 5528 11069 5556
rect 10836 5516 10842 5528
rect 11057 5525 11069 5528
rect 11103 5525 11115 5559
rect 11057 5519 11115 5525
rect 11238 5516 11244 5568
rect 11296 5556 11302 5568
rect 13464 5556 13492 5596
rect 14185 5593 14197 5596
rect 14231 5593 14243 5627
rect 14185 5587 14243 5593
rect 14550 5584 14556 5636
rect 14608 5624 14614 5636
rect 14844 5624 14872 5655
rect 15286 5652 15292 5664
rect 15344 5652 15350 5704
rect 16393 5695 16451 5701
rect 16393 5661 16405 5695
rect 16439 5692 16451 5695
rect 17218 5692 17224 5704
rect 16439 5664 17224 5692
rect 16439 5661 16451 5664
rect 16393 5655 16451 5661
rect 17218 5652 17224 5664
rect 17276 5692 17282 5704
rect 18156 5701 18184 5732
rect 17313 5695 17371 5701
rect 17313 5692 17325 5695
rect 17276 5664 17325 5692
rect 17276 5652 17282 5664
rect 17313 5661 17325 5664
rect 17359 5661 17371 5695
rect 17313 5655 17371 5661
rect 18049 5695 18107 5701
rect 18049 5661 18061 5695
rect 18095 5661 18107 5695
rect 18049 5655 18107 5661
rect 18141 5695 18199 5701
rect 18141 5661 18153 5695
rect 18187 5661 18199 5695
rect 18141 5655 18199 5661
rect 18064 5624 18092 5655
rect 14608 5596 14872 5624
rect 15028 5596 18092 5624
rect 14608 5584 14614 5596
rect 13906 5556 13912 5568
rect 11296 5528 13492 5556
rect 13867 5528 13912 5556
rect 11296 5516 11302 5528
rect 13906 5516 13912 5528
rect 13964 5516 13970 5568
rect 14369 5559 14427 5565
rect 14369 5525 14381 5559
rect 14415 5556 14427 5559
rect 15028 5556 15056 5596
rect 14415 5528 15056 5556
rect 14415 5525 14427 5528
rect 14369 5519 14427 5525
rect 15102 5516 15108 5568
rect 15160 5556 15166 5568
rect 15289 5559 15347 5565
rect 15289 5556 15301 5559
rect 15160 5528 15301 5556
rect 15160 5516 15166 5528
rect 15289 5525 15301 5528
rect 15335 5525 15347 5559
rect 15289 5519 15347 5525
rect 15470 5516 15476 5568
rect 15528 5556 15534 5568
rect 15565 5559 15623 5565
rect 15565 5556 15577 5559
rect 15528 5528 15577 5556
rect 15528 5516 15534 5528
rect 15565 5525 15577 5528
rect 15611 5525 15623 5559
rect 15565 5519 15623 5525
rect 16666 5516 16672 5568
rect 16724 5556 16730 5568
rect 18248 5556 18276 5800
rect 19978 5788 19984 5800
rect 20036 5788 20042 5840
rect 20441 5831 20499 5837
rect 20441 5797 20453 5831
rect 20487 5828 20499 5831
rect 20530 5828 20536 5840
rect 20487 5800 20536 5828
rect 20487 5797 20499 5800
rect 20441 5791 20499 5797
rect 20530 5788 20536 5800
rect 20588 5788 20594 5840
rect 18690 5760 18696 5772
rect 18651 5732 18696 5760
rect 18690 5720 18696 5732
rect 18748 5720 18754 5772
rect 18960 5763 19018 5769
rect 18960 5729 18972 5763
rect 19006 5760 19018 5763
rect 19518 5760 19524 5772
rect 19006 5732 19524 5760
rect 19006 5729 19018 5732
rect 18960 5723 19018 5729
rect 19518 5720 19524 5732
rect 19576 5720 19582 5772
rect 20162 5760 20168 5772
rect 20123 5732 20168 5760
rect 20162 5720 20168 5732
rect 20220 5720 20226 5772
rect 22002 5556 22008 5568
rect 16724 5528 18276 5556
rect 21963 5528 22008 5556
rect 16724 5516 16730 5528
rect 22002 5516 22008 5528
rect 22060 5516 22066 5568
rect 1104 5466 21896 5488
rect 1104 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 4575 5466
rect 4627 5414 4639 5466
rect 4691 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 18308 5466
rect 18360 5414 18372 5466
rect 18424 5414 18436 5466
rect 18488 5414 18500 5466
rect 18552 5414 21896 5466
rect 1104 5392 21896 5414
rect 3050 5312 3056 5364
rect 3108 5352 3114 5364
rect 3878 5352 3884 5364
rect 3108 5324 3884 5352
rect 3108 5312 3114 5324
rect 3878 5312 3884 5324
rect 3936 5352 3942 5364
rect 3936 5324 4200 5352
rect 3936 5312 3942 5324
rect 4172 5284 4200 5324
rect 4338 5312 4344 5364
rect 4396 5352 4402 5364
rect 4709 5355 4767 5361
rect 4709 5352 4721 5355
rect 4396 5324 4721 5352
rect 4396 5312 4402 5324
rect 4709 5321 4721 5324
rect 4755 5321 4767 5355
rect 5534 5352 5540 5364
rect 5495 5324 5540 5352
rect 4709 5315 4767 5321
rect 5534 5312 5540 5324
rect 5592 5312 5598 5364
rect 7006 5352 7012 5364
rect 6967 5324 7012 5352
rect 7006 5312 7012 5324
rect 7064 5312 7070 5364
rect 7098 5312 7104 5364
rect 7156 5352 7162 5364
rect 7193 5355 7251 5361
rect 7193 5352 7205 5355
rect 7156 5324 7205 5352
rect 7156 5312 7162 5324
rect 7193 5321 7205 5324
rect 7239 5352 7251 5355
rect 7834 5352 7840 5364
rect 7239 5324 7840 5352
rect 7239 5321 7251 5324
rect 7193 5315 7251 5321
rect 7834 5312 7840 5324
rect 7892 5312 7898 5364
rect 8297 5355 8355 5361
rect 8297 5321 8309 5355
rect 8343 5352 8355 5355
rect 8386 5352 8392 5364
rect 8343 5324 8392 5352
rect 8343 5321 8355 5324
rect 8297 5315 8355 5321
rect 8386 5312 8392 5324
rect 8444 5312 8450 5364
rect 9398 5352 9404 5364
rect 9140 5324 9404 5352
rect 4617 5287 4675 5293
rect 4617 5284 4629 5287
rect 4172 5256 4629 5284
rect 4617 5253 4629 5256
rect 4663 5253 4675 5287
rect 4617 5247 4675 5253
rect 8662 5244 8668 5296
rect 8720 5284 8726 5296
rect 9140 5284 9168 5324
rect 9398 5312 9404 5324
rect 9456 5312 9462 5364
rect 10778 5352 10784 5364
rect 10152 5324 10784 5352
rect 8720 5256 9168 5284
rect 8720 5244 8726 5256
rect 5350 5216 5356 5228
rect 5311 5188 5356 5216
rect 5350 5176 5356 5188
rect 5408 5176 5414 5228
rect 5902 5176 5908 5228
rect 5960 5216 5966 5228
rect 5997 5219 6055 5225
rect 5997 5216 6009 5219
rect 5960 5188 6009 5216
rect 5960 5176 5966 5188
rect 5997 5185 6009 5188
rect 6043 5185 6055 5219
rect 6178 5216 6184 5228
rect 6139 5188 6184 5216
rect 5997 5179 6055 5185
rect 6178 5176 6184 5188
rect 6236 5176 6242 5228
rect 6457 5219 6515 5225
rect 6457 5185 6469 5219
rect 6503 5216 6515 5219
rect 7098 5216 7104 5228
rect 6503 5188 7104 5216
rect 6503 5185 6515 5188
rect 6457 5179 6515 5185
rect 7098 5176 7104 5188
rect 7156 5216 7162 5228
rect 7374 5216 7380 5228
rect 7156 5188 7380 5216
rect 7156 5176 7162 5188
rect 7374 5176 7380 5188
rect 7432 5176 7438 5228
rect 7742 5176 7748 5228
rect 7800 5216 7806 5228
rect 7837 5219 7895 5225
rect 7837 5216 7849 5219
rect 7800 5188 7849 5216
rect 7800 5176 7806 5188
rect 7837 5185 7849 5188
rect 7883 5185 7895 5219
rect 7837 5179 7895 5185
rect 7926 5176 7932 5228
rect 7984 5216 7990 5228
rect 9140 5225 9168 5256
rect 8849 5219 8907 5225
rect 8849 5216 8861 5219
rect 7984 5188 8616 5216
rect 7984 5176 7990 5188
rect 1394 5108 1400 5160
rect 1452 5148 1458 5160
rect 1765 5151 1823 5157
rect 1765 5148 1777 5151
rect 1452 5120 1777 5148
rect 1452 5108 1458 5120
rect 1765 5117 1777 5120
rect 1811 5148 1823 5151
rect 3237 5151 3295 5157
rect 1811 5120 2912 5148
rect 1811 5117 1823 5120
rect 1765 5111 1823 5117
rect 2884 5092 2912 5120
rect 3237 5117 3249 5151
rect 3283 5117 3295 5151
rect 3237 5111 3295 5117
rect 3504 5151 3562 5157
rect 3504 5117 3516 5151
rect 3550 5148 3562 5151
rect 3786 5148 3792 5160
rect 3550 5120 3792 5148
rect 3550 5117 3562 5120
rect 3504 5111 3562 5117
rect 2032 5083 2090 5089
rect 2032 5049 2044 5083
rect 2078 5080 2090 5083
rect 2774 5080 2780 5092
rect 2078 5052 2780 5080
rect 2078 5049 2090 5052
rect 2032 5043 2090 5049
rect 2774 5040 2780 5052
rect 2832 5040 2838 5092
rect 2866 5040 2872 5092
rect 2924 5080 2930 5092
rect 3252 5080 3280 5111
rect 3786 5108 3792 5120
rect 3844 5148 3850 5160
rect 6196 5148 6224 5176
rect 3844 5120 6224 5148
rect 8588 5148 8616 5188
rect 8763 5188 8861 5216
rect 8763 5148 8791 5188
rect 8849 5185 8861 5188
rect 8895 5185 8907 5219
rect 8849 5179 8907 5185
rect 9125 5219 9183 5225
rect 9125 5185 9137 5219
rect 9171 5185 9183 5219
rect 9125 5179 9183 5185
rect 8588 5120 8791 5148
rect 9392 5151 9450 5157
rect 3844 5108 3850 5120
rect 9392 5117 9404 5151
rect 9438 5148 9450 5151
rect 10152 5148 10180 5324
rect 10778 5312 10784 5324
rect 10836 5312 10842 5364
rect 11698 5312 11704 5364
rect 11756 5352 11762 5364
rect 11974 5352 11980 5364
rect 11756 5324 11980 5352
rect 11756 5312 11762 5324
rect 11974 5312 11980 5324
rect 12032 5352 12038 5364
rect 12710 5352 12716 5364
rect 12032 5324 12716 5352
rect 12032 5312 12038 5324
rect 12710 5312 12716 5324
rect 12768 5312 12774 5364
rect 14185 5355 14243 5361
rect 14185 5321 14197 5355
rect 14231 5352 14243 5355
rect 14550 5352 14556 5364
rect 14231 5324 14556 5352
rect 14231 5321 14243 5324
rect 14185 5315 14243 5321
rect 14550 5312 14556 5324
rect 14608 5312 14614 5364
rect 16574 5352 16580 5364
rect 14936 5324 16160 5352
rect 16535 5324 16580 5352
rect 11330 5244 11336 5296
rect 11388 5284 11394 5296
rect 12250 5284 12256 5296
rect 11388 5256 12256 5284
rect 11388 5244 11394 5256
rect 12250 5244 12256 5256
rect 12308 5244 12314 5296
rect 12894 5244 12900 5296
rect 12952 5284 12958 5296
rect 14936 5284 14964 5324
rect 12952 5256 14964 5284
rect 12952 5244 12958 5256
rect 10778 5176 10784 5228
rect 10836 5176 10842 5228
rect 10962 5176 10968 5228
rect 11020 5216 11026 5228
rect 11057 5219 11115 5225
rect 11057 5216 11069 5219
rect 11020 5188 11069 5216
rect 11020 5176 11026 5188
rect 11057 5185 11069 5188
rect 11103 5185 11115 5219
rect 11057 5179 11115 5185
rect 11149 5219 11207 5225
rect 11149 5185 11161 5219
rect 11195 5185 11207 5219
rect 11974 5216 11980 5228
rect 11935 5188 11980 5216
rect 11149 5179 11207 5185
rect 9438 5120 10180 5148
rect 10796 5148 10824 5176
rect 11164 5148 11192 5179
rect 11974 5176 11980 5188
rect 12032 5176 12038 5228
rect 13078 5216 13084 5228
rect 12991 5188 13084 5216
rect 13078 5176 13084 5188
rect 13136 5216 13142 5228
rect 13906 5216 13912 5228
rect 13136 5188 13912 5216
rect 13136 5176 13142 5188
rect 13906 5176 13912 5188
rect 13964 5216 13970 5228
rect 14001 5219 14059 5225
rect 14001 5216 14013 5219
rect 13964 5188 14013 5216
rect 13964 5176 13970 5188
rect 14001 5185 14013 5188
rect 14047 5216 14059 5219
rect 14734 5216 14740 5228
rect 14047 5188 14740 5216
rect 14047 5185 14059 5188
rect 14001 5179 14059 5185
rect 14734 5176 14740 5188
rect 14792 5176 14798 5228
rect 14826 5176 14832 5228
rect 14884 5216 14890 5228
rect 16132 5216 16160 5324
rect 16574 5312 16580 5324
rect 16632 5312 16638 5364
rect 17126 5312 17132 5364
rect 17184 5352 17190 5364
rect 17865 5355 17923 5361
rect 17865 5352 17877 5355
rect 17184 5324 17877 5352
rect 17184 5312 17190 5324
rect 17865 5321 17877 5324
rect 17911 5352 17923 5355
rect 19058 5352 19064 5364
rect 17911 5324 19064 5352
rect 17911 5321 17923 5324
rect 17865 5315 17923 5321
rect 19058 5312 19064 5324
rect 19116 5312 19122 5364
rect 19518 5352 19524 5364
rect 19479 5324 19524 5352
rect 19518 5312 19524 5324
rect 19576 5312 19582 5364
rect 19613 5355 19671 5361
rect 19613 5321 19625 5355
rect 19659 5352 19671 5355
rect 20162 5352 20168 5364
rect 19659 5324 20168 5352
rect 19659 5321 19671 5324
rect 19613 5315 19671 5321
rect 20162 5312 20168 5324
rect 20220 5312 20226 5364
rect 16485 5287 16543 5293
rect 16485 5253 16497 5287
rect 16531 5284 16543 5287
rect 16666 5284 16672 5296
rect 16531 5256 16672 5284
rect 16531 5253 16543 5256
rect 16485 5247 16543 5253
rect 16666 5244 16672 5256
rect 16724 5284 16730 5296
rect 16724 5256 17264 5284
rect 16724 5244 16730 5256
rect 16574 5216 16580 5228
rect 14884 5188 14929 5216
rect 16132 5188 16580 5216
rect 14884 5176 14890 5188
rect 16574 5176 16580 5188
rect 16632 5176 16638 5228
rect 16758 5176 16764 5228
rect 16816 5216 16822 5228
rect 17236 5225 17264 5256
rect 17586 5244 17592 5296
rect 17644 5284 17650 5296
rect 18138 5284 18144 5296
rect 17644 5256 18144 5284
rect 17644 5244 17650 5256
rect 18138 5244 18144 5256
rect 18196 5244 18202 5296
rect 17037 5219 17095 5225
rect 17037 5216 17049 5219
rect 16816 5188 17049 5216
rect 16816 5176 16822 5188
rect 17037 5185 17049 5188
rect 17083 5185 17095 5219
rect 17037 5179 17095 5185
rect 17221 5219 17279 5225
rect 17221 5185 17233 5219
rect 17267 5216 17279 5219
rect 17402 5216 17408 5228
rect 17267 5188 17408 5216
rect 17267 5185 17279 5188
rect 17221 5179 17279 5185
rect 17402 5176 17408 5188
rect 17460 5176 17466 5228
rect 19536 5216 19564 5312
rect 19702 5244 19708 5296
rect 19760 5284 19766 5296
rect 20070 5284 20076 5296
rect 19760 5256 20076 5284
rect 19760 5244 19766 5256
rect 20070 5244 20076 5256
rect 20128 5244 20134 5296
rect 20165 5219 20223 5225
rect 20165 5216 20177 5219
rect 19536 5188 20177 5216
rect 20165 5185 20177 5188
rect 20211 5185 20223 5219
rect 20165 5179 20223 5185
rect 11790 5148 11796 5160
rect 10796 5120 11192 5148
rect 11751 5120 11796 5148
rect 9438 5117 9450 5120
rect 9392 5111 9450 5117
rect 11790 5108 11796 5120
rect 11848 5108 11854 5160
rect 11885 5151 11943 5157
rect 11885 5117 11897 5151
rect 11931 5148 11943 5151
rect 12434 5148 12440 5160
rect 11931 5120 12440 5148
rect 11931 5117 11943 5120
rect 11885 5111 11943 5117
rect 12434 5108 12440 5120
rect 12492 5148 12498 5160
rect 13170 5148 13176 5160
rect 12492 5120 13176 5148
rect 12492 5108 12498 5120
rect 13170 5108 13176 5120
rect 13228 5108 13234 5160
rect 13722 5108 13728 5160
rect 13780 5148 13786 5160
rect 13817 5151 13875 5157
rect 13817 5148 13829 5151
rect 13780 5120 13829 5148
rect 13780 5108 13786 5120
rect 13817 5117 13829 5120
rect 13863 5117 13875 5151
rect 13817 5111 13875 5117
rect 14645 5151 14703 5157
rect 14645 5117 14657 5151
rect 14691 5148 14703 5151
rect 15105 5151 15163 5157
rect 14691 5120 15056 5148
rect 14691 5117 14703 5120
rect 14645 5111 14703 5117
rect 15028 5092 15056 5120
rect 15105 5117 15117 5151
rect 15151 5148 15163 5151
rect 15194 5148 15200 5160
rect 15151 5120 15200 5148
rect 15151 5117 15163 5120
rect 15105 5111 15163 5117
rect 15194 5108 15200 5120
rect 15252 5108 15258 5160
rect 16850 5108 16856 5160
rect 16908 5148 16914 5160
rect 16945 5151 17003 5157
rect 16945 5148 16957 5151
rect 16908 5120 16957 5148
rect 16908 5108 16914 5120
rect 16945 5117 16957 5120
rect 16991 5117 17003 5151
rect 16945 5111 17003 5117
rect 17310 5108 17316 5160
rect 17368 5148 17374 5160
rect 17681 5151 17739 5157
rect 17681 5148 17693 5151
rect 17368 5120 17693 5148
rect 17368 5108 17374 5120
rect 17681 5117 17693 5120
rect 17727 5148 17739 5151
rect 17862 5148 17868 5160
rect 17727 5120 17868 5148
rect 17727 5117 17739 5120
rect 17681 5111 17739 5117
rect 17862 5108 17868 5120
rect 17920 5108 17926 5160
rect 18046 5108 18052 5160
rect 18104 5148 18110 5160
rect 18141 5151 18199 5157
rect 18141 5148 18153 5151
rect 18104 5120 18153 5148
rect 18104 5108 18110 5120
rect 18141 5117 18153 5120
rect 18187 5148 18199 5151
rect 18690 5148 18696 5160
rect 18187 5120 18696 5148
rect 18187 5117 18199 5120
rect 18141 5111 18199 5117
rect 18690 5108 18696 5120
rect 18748 5108 18754 5160
rect 3694 5080 3700 5092
rect 2924 5052 3700 5080
rect 2924 5040 2930 5052
rect 3694 5040 3700 5052
rect 3752 5040 3758 5092
rect 4246 5040 4252 5092
rect 4304 5080 4310 5092
rect 5077 5083 5135 5089
rect 5077 5080 5089 5083
rect 4304 5052 5089 5080
rect 4304 5040 4310 5052
rect 5077 5049 5089 5052
rect 5123 5049 5135 5083
rect 5077 5043 5135 5049
rect 5905 5083 5963 5089
rect 5905 5049 5917 5083
rect 5951 5080 5963 5083
rect 6270 5080 6276 5092
rect 5951 5052 6276 5080
rect 5951 5049 5963 5052
rect 5905 5043 5963 5049
rect 6270 5040 6276 5052
rect 6328 5040 6334 5092
rect 6638 5080 6644 5092
rect 6551 5052 6644 5080
rect 6638 5040 6644 5052
rect 6696 5080 6702 5092
rect 6696 5052 7604 5080
rect 6696 5040 6702 5052
rect 3145 5015 3203 5021
rect 3145 4981 3157 5015
rect 3191 5012 3203 5015
rect 3418 5012 3424 5024
rect 3191 4984 3424 5012
rect 3191 4981 3203 4984
rect 3145 4975 3203 4981
rect 3418 4972 3424 4984
rect 3476 4972 3482 5024
rect 5169 5015 5227 5021
rect 5169 4981 5181 5015
rect 5215 5012 5227 5015
rect 5718 5012 5724 5024
rect 5215 4984 5724 5012
rect 5215 4981 5227 4984
rect 5169 4975 5227 4981
rect 5718 4972 5724 4984
rect 5776 4972 5782 5024
rect 7374 5012 7380 5024
rect 7335 4984 7380 5012
rect 7374 4972 7380 4984
rect 7432 4972 7438 5024
rect 7576 5012 7604 5052
rect 7650 5040 7656 5092
rect 7708 5080 7714 5092
rect 7745 5083 7803 5089
rect 7745 5080 7757 5083
rect 7708 5052 7757 5080
rect 7708 5040 7714 5052
rect 7745 5049 7757 5052
rect 7791 5049 7803 5083
rect 7745 5043 7803 5049
rect 8018 5040 8024 5092
rect 8076 5080 8082 5092
rect 8665 5083 8723 5089
rect 8665 5080 8677 5083
rect 8076 5052 8677 5080
rect 8076 5040 8082 5052
rect 8665 5049 8677 5052
rect 8711 5049 8723 5083
rect 8665 5043 8723 5049
rect 8754 5040 8760 5092
rect 8812 5080 8818 5092
rect 8812 5052 8857 5080
rect 8812 5040 8818 5052
rect 9214 5040 9220 5092
rect 9272 5080 9278 5092
rect 9272 5052 10824 5080
rect 9272 5040 9278 5052
rect 9674 5012 9680 5024
rect 7576 4984 9680 5012
rect 9674 4972 9680 4984
rect 9732 4972 9738 5024
rect 10502 5012 10508 5024
rect 10463 4984 10508 5012
rect 10502 4972 10508 4984
rect 10560 4972 10566 5024
rect 10594 4972 10600 5024
rect 10652 5012 10658 5024
rect 10796 5012 10824 5052
rect 10870 5040 10876 5092
rect 10928 5080 10934 5092
rect 10965 5083 11023 5089
rect 10965 5080 10977 5083
rect 10928 5052 10977 5080
rect 10928 5040 10934 5052
rect 10965 5049 10977 5052
rect 11011 5049 11023 5083
rect 10965 5043 11023 5049
rect 12250 5040 12256 5092
rect 12308 5080 12314 5092
rect 12308 5052 12664 5080
rect 12308 5040 12314 5052
rect 11238 5012 11244 5024
rect 10652 4984 10697 5012
rect 10796 4984 11244 5012
rect 10652 4972 10658 4984
rect 11238 4972 11244 4984
rect 11296 4972 11302 5024
rect 11425 5015 11483 5021
rect 11425 4981 11437 5015
rect 11471 5012 11483 5015
rect 11698 5012 11704 5024
rect 11471 4984 11704 5012
rect 11471 4981 11483 4984
rect 11425 4975 11483 4981
rect 11698 4972 11704 4984
rect 11756 4972 11762 5024
rect 12437 5015 12495 5021
rect 12437 4981 12449 5015
rect 12483 5012 12495 5015
rect 12526 5012 12532 5024
rect 12483 4984 12532 5012
rect 12483 4981 12495 4984
rect 12437 4975 12495 4981
rect 12526 4972 12532 4984
rect 12584 4972 12590 5024
rect 12636 5012 12664 5052
rect 12710 5040 12716 5092
rect 12768 5080 12774 5092
rect 12805 5083 12863 5089
rect 12805 5080 12817 5083
rect 12768 5052 12817 5080
rect 12768 5040 12774 5052
rect 12805 5049 12817 5052
rect 12851 5049 12863 5083
rect 12805 5043 12863 5049
rect 13906 5040 13912 5092
rect 13964 5080 13970 5092
rect 13964 5052 14964 5080
rect 13964 5040 13970 5052
rect 12897 5015 12955 5021
rect 12897 5012 12909 5015
rect 12636 4984 12909 5012
rect 12897 4981 12909 4984
rect 12943 4981 12955 5015
rect 13354 5012 13360 5024
rect 13315 4984 13360 5012
rect 12897 4975 12955 4981
rect 13354 4972 13360 4984
rect 13412 4972 13418 5024
rect 13722 5012 13728 5024
rect 13683 4984 13728 5012
rect 13722 4972 13728 4984
rect 13780 4972 13786 5024
rect 13998 4972 14004 5024
rect 14056 5012 14062 5024
rect 14553 5015 14611 5021
rect 14553 5012 14565 5015
rect 14056 4984 14565 5012
rect 14056 4972 14062 4984
rect 14553 4981 14565 4984
rect 14599 4981 14611 5015
rect 14936 5012 14964 5052
rect 15010 5040 15016 5092
rect 15068 5040 15074 5092
rect 15286 5040 15292 5092
rect 15344 5089 15350 5092
rect 15344 5083 15408 5089
rect 15344 5049 15362 5083
rect 15396 5049 15408 5083
rect 15344 5043 15408 5049
rect 15344 5040 15350 5043
rect 18322 5040 18328 5092
rect 18380 5089 18386 5092
rect 18380 5083 18444 5089
rect 18380 5049 18398 5083
rect 18432 5049 18444 5083
rect 20073 5083 20131 5089
rect 20073 5080 20085 5083
rect 18380 5043 18444 5049
rect 18524 5052 20085 5080
rect 18380 5040 18386 5043
rect 16114 5012 16120 5024
rect 14936 4984 16120 5012
rect 14553 4975 14611 4981
rect 16114 4972 16120 4984
rect 16172 4972 16178 5024
rect 17862 4972 17868 5024
rect 17920 5012 17926 5024
rect 18524 5012 18552 5052
rect 20073 5049 20085 5052
rect 20119 5049 20131 5083
rect 20073 5043 20131 5049
rect 19978 5012 19984 5024
rect 17920 4984 18552 5012
rect 19939 4984 19984 5012
rect 17920 4972 17926 4984
rect 19978 4972 19984 4984
rect 20036 4972 20042 5024
rect 1104 4922 21896 4944
rect 1104 4870 7912 4922
rect 7964 4870 7976 4922
rect 8028 4870 8040 4922
rect 8092 4870 8104 4922
rect 8156 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 15035 4922
rect 15087 4870 21896 4922
rect 1104 4848 21896 4870
rect 2774 4768 2780 4820
rect 2832 4808 2838 4820
rect 4062 4808 4068 4820
rect 2832 4780 2877 4808
rect 4023 4780 4068 4808
rect 2832 4768 2838 4780
rect 4062 4768 4068 4780
rect 4120 4768 4126 4820
rect 5261 4811 5319 4817
rect 5261 4777 5273 4811
rect 5307 4808 5319 4811
rect 7098 4808 7104 4820
rect 5307 4780 7104 4808
rect 5307 4777 5319 4780
rect 5261 4771 5319 4777
rect 7098 4768 7104 4780
rect 7156 4768 7162 4820
rect 7561 4811 7619 4817
rect 7561 4777 7573 4811
rect 7607 4808 7619 4811
rect 7929 4811 7987 4817
rect 7929 4808 7941 4811
rect 7607 4780 7941 4808
rect 7607 4777 7619 4780
rect 7561 4771 7619 4777
rect 7929 4777 7941 4780
rect 7975 4777 7987 4811
rect 8386 4808 8392 4820
rect 8347 4780 8392 4808
rect 7929 4771 7987 4777
rect 8386 4768 8392 4780
rect 8444 4768 8450 4820
rect 8754 4808 8760 4820
rect 8715 4780 8760 4808
rect 8754 4768 8760 4780
rect 8812 4768 8818 4820
rect 9122 4808 9128 4820
rect 9083 4780 9128 4808
rect 9122 4768 9128 4780
rect 9180 4768 9186 4820
rect 9677 4811 9735 4817
rect 9677 4777 9689 4811
rect 9723 4808 9735 4811
rect 10042 4808 10048 4820
rect 9723 4780 10048 4808
rect 9723 4777 9735 4780
rect 9677 4771 9735 4777
rect 10042 4768 10048 4780
rect 10100 4768 10106 4820
rect 10410 4768 10416 4820
rect 10468 4808 10474 4820
rect 10597 4811 10655 4817
rect 10597 4808 10609 4811
rect 10468 4780 10609 4808
rect 10468 4768 10474 4780
rect 10597 4777 10609 4780
rect 10643 4808 10655 4811
rect 11330 4808 11336 4820
rect 10643 4780 11336 4808
rect 10643 4777 10655 4780
rect 10597 4771 10655 4777
rect 11330 4768 11336 4780
rect 11388 4768 11394 4820
rect 11790 4768 11796 4820
rect 11848 4808 11854 4820
rect 11977 4811 12035 4817
rect 11977 4808 11989 4811
rect 11848 4780 11989 4808
rect 11848 4768 11854 4780
rect 11977 4777 11989 4780
rect 12023 4777 12035 4811
rect 12250 4808 12256 4820
rect 12211 4780 12256 4808
rect 11977 4771 12035 4777
rect 12250 4768 12256 4780
rect 12308 4768 12314 4820
rect 12434 4808 12440 4820
rect 12395 4780 12440 4808
rect 12434 4768 12440 4780
rect 12492 4768 12498 4820
rect 15289 4811 15347 4817
rect 15289 4808 15301 4811
rect 12912 4780 15301 4808
rect 1302 4700 1308 4752
rect 1360 4740 1366 4752
rect 1664 4743 1722 4749
rect 1360 4712 1624 4740
rect 1360 4700 1366 4712
rect 1394 4672 1400 4684
rect 1355 4644 1400 4672
rect 1394 4632 1400 4644
rect 1452 4632 1458 4684
rect 1596 4672 1624 4712
rect 1664 4709 1676 4743
rect 1710 4740 1722 4743
rect 2682 4740 2688 4752
rect 1710 4712 2688 4740
rect 1710 4709 1722 4712
rect 1664 4703 1722 4709
rect 2682 4700 2688 4712
rect 2740 4740 2746 4752
rect 2740 4712 3648 4740
rect 2740 4700 2746 4712
rect 3510 4672 3516 4684
rect 1596 4644 2728 4672
rect 3471 4644 3516 4672
rect 2700 4604 2728 4644
rect 3510 4632 3516 4644
rect 3568 4632 3574 4684
rect 3620 4672 3648 4712
rect 3694 4700 3700 4752
rect 3752 4740 3758 4752
rect 5896 4743 5954 4749
rect 3752 4712 5304 4740
rect 3752 4700 3758 4712
rect 5166 4672 5172 4684
rect 3620 4644 3740 4672
rect 5127 4644 5172 4672
rect 3712 4616 3740 4644
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 5276 4672 5304 4712
rect 5896 4709 5908 4743
rect 5942 4740 5954 4743
rect 10502 4740 10508 4752
rect 5942 4712 10508 4740
rect 5942 4709 5954 4712
rect 5896 4703 5954 4709
rect 10502 4700 10508 4712
rect 10560 4700 10566 4752
rect 12268 4740 12296 4768
rect 10612 4712 12296 4740
rect 7466 4672 7472 4684
rect 5276 4644 5580 4672
rect 7427 4644 7472 4672
rect 3605 4607 3663 4613
rect 2700 4576 3280 4604
rect 2406 4496 2412 4548
rect 2464 4536 2470 4548
rect 3145 4539 3203 4545
rect 3145 4536 3157 4539
rect 2464 4508 3157 4536
rect 2464 4496 2470 4508
rect 3145 4505 3157 4508
rect 3191 4505 3203 4539
rect 3145 4499 3203 4505
rect 2958 4468 2964 4480
rect 2919 4440 2964 4468
rect 2958 4428 2964 4440
rect 3016 4428 3022 4480
rect 3252 4468 3280 4576
rect 3605 4573 3617 4607
rect 3651 4573 3663 4607
rect 3605 4567 3663 4573
rect 3620 4536 3648 4567
rect 3694 4564 3700 4616
rect 3752 4604 3758 4616
rect 3752 4576 3845 4604
rect 3752 4564 3758 4576
rect 5350 4564 5356 4616
rect 5408 4604 5414 4616
rect 5552 4604 5580 4644
rect 7466 4632 7472 4644
rect 7524 4632 7530 4684
rect 8297 4675 8355 4681
rect 8297 4641 8309 4675
rect 8343 4672 8355 4675
rect 8343 4644 8616 4672
rect 8343 4641 8355 4644
rect 8297 4635 8355 4641
rect 5629 4607 5687 4613
rect 5629 4604 5641 4607
rect 5408 4576 5453 4604
rect 5552 4576 5641 4604
rect 5408 4564 5414 4576
rect 5629 4573 5641 4576
rect 5675 4573 5687 4607
rect 5629 4567 5687 4573
rect 7558 4564 7564 4616
rect 7616 4604 7622 4616
rect 7653 4607 7711 4613
rect 7653 4604 7665 4607
rect 7616 4576 7665 4604
rect 7616 4564 7622 4576
rect 7653 4573 7665 4576
rect 7699 4573 7711 4607
rect 7653 4567 7711 4573
rect 8202 4564 8208 4616
rect 8260 4604 8266 4616
rect 8481 4607 8539 4613
rect 8481 4604 8493 4607
rect 8260 4576 8493 4604
rect 8260 4564 8266 4576
rect 8481 4573 8493 4576
rect 8527 4573 8539 4607
rect 8588 4604 8616 4644
rect 8662 4632 8668 4684
rect 8720 4672 8726 4684
rect 8720 4644 8984 4672
rect 8720 4632 8726 4644
rect 8846 4604 8852 4616
rect 8588 4576 8852 4604
rect 8481 4567 8539 4573
rect 8846 4564 8852 4576
rect 8904 4564 8910 4616
rect 8956 4604 8984 4644
rect 9122 4632 9128 4684
rect 9180 4672 9186 4684
rect 9180 4644 9435 4672
rect 9180 4632 9186 4644
rect 9217 4607 9275 4613
rect 9217 4604 9229 4607
rect 8956 4576 9229 4604
rect 9217 4573 9229 4576
rect 9263 4573 9275 4607
rect 9217 4567 9275 4573
rect 9309 4607 9367 4613
rect 9309 4573 9321 4607
rect 9355 4573 9367 4607
rect 9309 4567 9367 4573
rect 4890 4536 4896 4548
rect 3620 4508 4896 4536
rect 4890 4496 4896 4508
rect 4948 4496 4954 4548
rect 8570 4496 8576 4548
rect 8628 4536 8634 4548
rect 9122 4536 9128 4548
rect 8628 4508 9128 4536
rect 8628 4496 8634 4508
rect 9122 4496 9128 4508
rect 9180 4536 9186 4548
rect 9324 4536 9352 4567
rect 9180 4508 9352 4536
rect 9180 4496 9186 4508
rect 4246 4468 4252 4480
rect 3252 4440 4252 4468
rect 4246 4428 4252 4440
rect 4304 4468 4310 4480
rect 4525 4471 4583 4477
rect 4525 4468 4537 4471
rect 4304 4440 4537 4468
rect 4304 4428 4310 4440
rect 4525 4437 4537 4440
rect 4571 4437 4583 4471
rect 4798 4468 4804 4480
rect 4759 4440 4804 4468
rect 4525 4431 4583 4437
rect 4798 4428 4804 4440
rect 4856 4428 4862 4480
rect 5350 4428 5356 4480
rect 5408 4468 5414 4480
rect 7009 4471 7067 4477
rect 7009 4468 7021 4471
rect 5408 4440 7021 4468
rect 5408 4428 5414 4440
rect 7009 4437 7021 4440
rect 7055 4437 7067 4471
rect 7009 4431 7067 4437
rect 7101 4471 7159 4477
rect 7101 4437 7113 4471
rect 7147 4468 7159 4471
rect 8478 4468 8484 4480
rect 7147 4440 8484 4468
rect 7147 4437 7159 4440
rect 7101 4431 7159 4437
rect 8478 4428 8484 4440
rect 8536 4428 8542 4480
rect 9407 4468 9435 4644
rect 9490 4632 9496 4684
rect 9548 4672 9554 4684
rect 10045 4675 10103 4681
rect 10045 4672 10057 4675
rect 9548 4644 10057 4672
rect 9548 4632 9554 4644
rect 10045 4641 10057 4644
rect 10091 4641 10103 4675
rect 10045 4635 10103 4641
rect 10137 4675 10195 4681
rect 10137 4641 10149 4675
rect 10183 4672 10195 4675
rect 10612 4672 10640 4712
rect 12342 4700 12348 4752
rect 12400 4740 12406 4752
rect 12912 4740 12940 4780
rect 15289 4777 15301 4780
rect 15335 4808 15347 4811
rect 15562 4808 15568 4820
rect 15335 4780 15568 4808
rect 15335 4777 15347 4780
rect 15289 4771 15347 4777
rect 15562 4768 15568 4780
rect 15620 4768 15626 4820
rect 16390 4768 16396 4820
rect 16448 4808 16454 4820
rect 16853 4811 16911 4817
rect 16853 4808 16865 4811
rect 16448 4780 16865 4808
rect 16448 4768 16454 4780
rect 16853 4777 16865 4780
rect 16899 4777 16911 4811
rect 16853 4771 16911 4777
rect 17681 4811 17739 4817
rect 17681 4777 17693 4811
rect 17727 4808 17739 4811
rect 17862 4808 17868 4820
rect 17727 4780 17868 4808
rect 17727 4777 17739 4780
rect 17681 4771 17739 4777
rect 17862 4768 17868 4780
rect 17920 4768 17926 4820
rect 18509 4811 18567 4817
rect 18509 4777 18521 4811
rect 18555 4808 18567 4811
rect 19797 4811 19855 4817
rect 19797 4808 19809 4811
rect 18555 4780 19809 4808
rect 18555 4777 18567 4780
rect 18509 4771 18567 4777
rect 19797 4777 19809 4780
rect 19843 4777 19855 4811
rect 19797 4771 19855 4777
rect 12400 4712 12940 4740
rect 12980 4743 13038 4749
rect 12400 4700 12406 4712
rect 12980 4709 12992 4743
rect 13026 4740 13038 4743
rect 13078 4740 13084 4752
rect 13026 4712 13084 4740
rect 13026 4709 13038 4712
rect 12980 4703 13038 4709
rect 13078 4700 13084 4712
rect 13136 4700 13142 4752
rect 14090 4700 14096 4752
rect 14148 4740 14154 4752
rect 14642 4740 14648 4752
rect 14148 4712 14648 4740
rect 14148 4700 14154 4712
rect 14642 4700 14648 4712
rect 14700 4700 14706 4752
rect 15013 4743 15071 4749
rect 15013 4709 15025 4743
rect 15059 4740 15071 4743
rect 15470 4740 15476 4752
rect 15059 4712 15476 4740
rect 15059 4709 15071 4712
rect 15013 4703 15071 4709
rect 10183 4644 10640 4672
rect 10183 4641 10195 4644
rect 10137 4635 10195 4641
rect 9674 4564 9680 4616
rect 9732 4604 9738 4616
rect 10152 4604 10180 4635
rect 10686 4632 10692 4684
rect 10744 4672 10750 4684
rect 10870 4672 10876 4684
rect 10744 4644 10876 4672
rect 10744 4632 10750 4644
rect 10870 4632 10876 4644
rect 10928 4672 10934 4684
rect 11517 4675 11575 4681
rect 11517 4672 11529 4675
rect 10928 4644 11529 4672
rect 10928 4632 10934 4644
rect 11517 4641 11529 4644
rect 11563 4641 11575 4675
rect 13998 4672 14004 4684
rect 11517 4635 11575 4641
rect 12544 4644 14004 4672
rect 10318 4604 10324 4616
rect 9732 4576 10180 4604
rect 10279 4576 10324 4604
rect 9732 4564 9738 4576
rect 10318 4564 10324 4576
rect 10376 4564 10382 4616
rect 10778 4564 10784 4616
rect 10836 4604 10842 4616
rect 11146 4604 11152 4616
rect 10836 4576 11152 4604
rect 10836 4564 10842 4576
rect 11146 4564 11152 4576
rect 11204 4604 11210 4616
rect 11609 4607 11667 4613
rect 11609 4604 11621 4607
rect 11204 4576 11621 4604
rect 11204 4564 11210 4576
rect 11609 4573 11621 4576
rect 11655 4573 11667 4607
rect 11609 4567 11667 4573
rect 11793 4607 11851 4613
rect 11793 4573 11805 4607
rect 11839 4604 11851 4607
rect 11974 4604 11980 4616
rect 11839 4576 11980 4604
rect 11839 4573 11851 4576
rect 11793 4567 11851 4573
rect 11974 4564 11980 4576
rect 12032 4564 12038 4616
rect 9582 4496 9588 4548
rect 9640 4536 9646 4548
rect 12544 4536 12572 4644
rect 13998 4632 14004 4644
rect 14056 4632 14062 4684
rect 14553 4675 14611 4681
rect 14553 4641 14565 4675
rect 14599 4641 14611 4675
rect 14553 4635 14611 4641
rect 12618 4564 12624 4616
rect 12676 4604 12682 4616
rect 12713 4607 12771 4613
rect 12713 4604 12725 4607
rect 12676 4576 12725 4604
rect 12676 4564 12682 4576
rect 12713 4573 12725 4576
rect 12759 4573 12771 4607
rect 14568 4604 14596 4635
rect 14734 4604 14740 4616
rect 12713 4567 12771 4573
rect 13740 4576 14596 4604
rect 14695 4576 14740 4604
rect 9640 4508 12572 4536
rect 9640 4496 9646 4508
rect 10704 4480 10732 4508
rect 13740 4480 13768 4576
rect 14734 4564 14740 4576
rect 14792 4564 14798 4616
rect 13906 4496 13912 4548
rect 13964 4536 13970 4548
rect 15028 4536 15056 4703
rect 15470 4700 15476 4712
rect 15528 4700 15534 4752
rect 15740 4743 15798 4749
rect 15740 4709 15752 4743
rect 15786 4740 15798 4743
rect 16666 4740 16672 4752
rect 15786 4712 16672 4740
rect 15786 4709 15798 4712
rect 15740 4703 15798 4709
rect 16666 4700 16672 4712
rect 16724 4700 16730 4752
rect 18969 4743 19027 4749
rect 18969 4740 18981 4743
rect 16776 4712 18981 4740
rect 15102 4632 15108 4684
rect 15160 4672 15166 4684
rect 16776 4672 16804 4712
rect 18969 4709 18981 4712
rect 19015 4709 19027 4743
rect 19150 4740 19156 4752
rect 18969 4703 19027 4709
rect 19076 4712 19156 4740
rect 15160 4644 16804 4672
rect 15160 4632 15166 4644
rect 17126 4632 17132 4684
rect 17184 4672 17190 4684
rect 18049 4675 18107 4681
rect 18049 4672 18061 4675
rect 17184 4644 18061 4672
rect 17184 4632 17190 4644
rect 18049 4641 18061 4644
rect 18095 4641 18107 4675
rect 18049 4635 18107 4641
rect 18230 4632 18236 4684
rect 18288 4672 18294 4684
rect 18877 4675 18935 4681
rect 18877 4672 18889 4675
rect 18288 4644 18889 4672
rect 18288 4632 18294 4644
rect 18877 4641 18889 4644
rect 18923 4672 18935 4675
rect 19076 4672 19104 4712
rect 19150 4700 19156 4712
rect 19208 4700 19214 4752
rect 19518 4672 19524 4684
rect 18923 4644 19104 4672
rect 19168 4644 19524 4672
rect 18923 4641 18935 4644
rect 18877 4635 18935 4641
rect 15194 4564 15200 4616
rect 15252 4604 15258 4616
rect 15470 4604 15476 4616
rect 15252 4576 15476 4604
rect 15252 4564 15258 4576
rect 15470 4564 15476 4576
rect 15528 4564 15534 4616
rect 18138 4604 18144 4616
rect 18099 4576 18144 4604
rect 18138 4564 18144 4576
rect 18196 4564 18202 4616
rect 18322 4604 18328 4616
rect 18283 4576 18328 4604
rect 18322 4564 18328 4576
rect 18380 4564 18386 4616
rect 19168 4613 19196 4644
rect 19518 4632 19524 4644
rect 19576 4632 19582 4684
rect 19702 4672 19708 4684
rect 19663 4644 19708 4672
rect 19702 4632 19708 4644
rect 19760 4632 19766 4684
rect 19153 4607 19211 4613
rect 19153 4573 19165 4607
rect 19199 4573 19211 4607
rect 19153 4567 19211 4573
rect 19426 4564 19432 4616
rect 19484 4604 19490 4616
rect 19889 4607 19947 4613
rect 19889 4604 19901 4607
rect 19484 4576 19901 4604
rect 19484 4564 19490 4576
rect 19889 4573 19901 4576
rect 19935 4573 19947 4607
rect 19889 4567 19947 4573
rect 13964 4508 15056 4536
rect 13964 4496 13970 4508
rect 16574 4496 16580 4548
rect 16632 4536 16638 4548
rect 17589 4539 17647 4545
rect 17589 4536 17601 4539
rect 16632 4508 17601 4536
rect 16632 4496 16638 4508
rect 17589 4505 17601 4508
rect 17635 4536 17647 4539
rect 18230 4536 18236 4548
rect 17635 4508 18236 4536
rect 17635 4505 17647 4508
rect 17589 4499 17647 4505
rect 18230 4496 18236 4508
rect 18288 4496 18294 4548
rect 10410 4468 10416 4480
rect 9407 4440 10416 4468
rect 10410 4428 10416 4440
rect 10468 4428 10474 4480
rect 10686 4428 10692 4480
rect 10744 4428 10750 4480
rect 10778 4428 10784 4480
rect 10836 4468 10842 4480
rect 10965 4471 11023 4477
rect 10965 4468 10977 4471
rect 10836 4440 10977 4468
rect 10836 4428 10842 4440
rect 10965 4437 10977 4440
rect 11011 4437 11023 4471
rect 11146 4468 11152 4480
rect 11107 4440 11152 4468
rect 10965 4431 11023 4437
rect 11146 4428 11152 4440
rect 11204 4428 11210 4480
rect 12986 4428 12992 4480
rect 13044 4468 13050 4480
rect 13722 4468 13728 4480
rect 13044 4440 13728 4468
rect 13044 4428 13050 4440
rect 13722 4428 13728 4440
rect 13780 4428 13786 4480
rect 13814 4428 13820 4480
rect 13872 4468 13878 4480
rect 14093 4471 14151 4477
rect 14093 4468 14105 4471
rect 13872 4440 14105 4468
rect 13872 4428 13878 4440
rect 14093 4437 14105 4440
rect 14139 4437 14151 4471
rect 14093 4431 14151 4437
rect 14182 4428 14188 4480
rect 14240 4468 14246 4480
rect 16942 4468 16948 4480
rect 14240 4440 14285 4468
rect 16903 4440 16948 4468
rect 14240 4428 14246 4440
rect 16942 4428 16948 4440
rect 17000 4428 17006 4480
rect 18340 4468 18368 4564
rect 19337 4539 19395 4545
rect 19337 4505 19349 4539
rect 19383 4536 19395 4539
rect 19978 4536 19984 4548
rect 19383 4508 19984 4536
rect 19383 4505 19395 4508
rect 19337 4499 19395 4505
rect 19978 4496 19984 4508
rect 20036 4496 20042 4548
rect 19426 4468 19432 4480
rect 18340 4440 19432 4468
rect 19426 4428 19432 4440
rect 19484 4428 19490 4480
rect 1104 4378 21896 4400
rect 1104 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 4575 4378
rect 4627 4326 4639 4378
rect 4691 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 18308 4378
rect 18360 4326 18372 4378
rect 18424 4326 18436 4378
rect 18488 4326 18500 4378
rect 18552 4326 21896 4378
rect 1104 4304 21896 4326
rect 3694 4224 3700 4276
rect 3752 4264 3758 4276
rect 4157 4267 4215 4273
rect 4157 4264 4169 4267
rect 3752 4236 4169 4264
rect 3752 4224 3758 4236
rect 4157 4233 4169 4236
rect 4203 4233 4215 4267
rect 4157 4227 4215 4233
rect 4246 4224 4252 4276
rect 4304 4264 4310 4276
rect 4801 4267 4859 4273
rect 4801 4264 4813 4267
rect 4304 4236 4813 4264
rect 4304 4224 4310 4236
rect 4801 4233 4813 4236
rect 4847 4264 4859 4267
rect 4847 4236 5120 4264
rect 4847 4233 4859 4236
rect 4801 4227 4859 4233
rect 2774 4196 2780 4208
rect 2608 4168 2780 4196
rect 2406 4128 2412 4140
rect 2367 4100 2412 4128
rect 2406 4088 2412 4100
rect 2464 4088 2470 4140
rect 2608 4137 2636 4168
rect 2774 4156 2780 4168
rect 2832 4156 2838 4208
rect 4706 4156 4712 4208
rect 4764 4196 4770 4208
rect 4982 4196 4988 4208
rect 4764 4168 4988 4196
rect 4764 4156 4770 4168
rect 4982 4156 4988 4168
rect 5040 4156 5046 4208
rect 5092 4196 5120 4236
rect 5166 4224 5172 4276
rect 5224 4264 5230 4276
rect 6638 4264 6644 4276
rect 5224 4236 6644 4264
rect 5224 4224 5230 4236
rect 6638 4224 6644 4236
rect 6696 4224 6702 4276
rect 7098 4224 7104 4276
rect 7156 4264 7162 4276
rect 7156 4236 7880 4264
rect 7156 4224 7162 4236
rect 5442 4196 5448 4208
rect 5092 4168 5448 4196
rect 5442 4156 5448 4168
rect 5500 4156 5506 4208
rect 7852 4196 7880 4236
rect 8754 4224 8760 4276
rect 8812 4264 8818 4276
rect 12250 4264 12256 4276
rect 8812 4236 12256 4264
rect 8812 4224 8818 4236
rect 12250 4224 12256 4236
rect 12308 4224 12314 4276
rect 15102 4264 15108 4276
rect 12360 4236 13676 4264
rect 15063 4236 15108 4264
rect 12360 4208 12388 4236
rect 9490 4196 9496 4208
rect 5552 4168 6408 4196
rect 7852 4168 9496 4196
rect 2593 4131 2651 4137
rect 2593 4097 2605 4131
rect 2639 4097 2651 4131
rect 2593 4091 2651 4097
rect 4154 4088 4160 4140
rect 4212 4128 4218 4140
rect 4617 4131 4675 4137
rect 4617 4128 4629 4131
rect 4212 4100 4629 4128
rect 4212 4088 4218 4100
rect 4617 4097 4629 4100
rect 4663 4128 4675 4131
rect 5258 4128 5264 4140
rect 4663 4100 5264 4128
rect 4663 4097 4675 4100
rect 4617 4091 4675 4097
rect 5258 4088 5264 4100
rect 5316 4088 5322 4140
rect 5350 4088 5356 4140
rect 5408 4128 5414 4140
rect 5552 4137 5580 4168
rect 5537 4131 5595 4137
rect 5537 4128 5549 4131
rect 5408 4100 5549 4128
rect 5408 4088 5414 4100
rect 5537 4097 5549 4100
rect 5583 4097 5595 4131
rect 6270 4128 6276 4140
rect 6231 4100 6276 4128
rect 5537 4091 5595 4097
rect 6270 4088 6276 4100
rect 6328 4088 6334 4140
rect 6380 4137 6408 4168
rect 9490 4156 9496 4168
rect 9548 4196 9554 4208
rect 9677 4199 9735 4205
rect 9677 4196 9689 4199
rect 9548 4168 9689 4196
rect 9548 4156 9554 4168
rect 9677 4165 9689 4168
rect 9723 4165 9735 4199
rect 9677 4159 9735 4165
rect 9766 4156 9772 4208
rect 9824 4196 9830 4208
rect 10042 4196 10048 4208
rect 9824 4168 10048 4196
rect 9824 4156 9830 4168
rect 10042 4156 10048 4168
rect 10100 4156 10106 4208
rect 10502 4196 10508 4208
rect 10428 4168 10508 4196
rect 6365 4131 6423 4137
rect 6365 4097 6377 4131
rect 6411 4097 6423 4131
rect 6365 4091 6423 4097
rect 8294 4088 8300 4140
rect 8352 4128 8358 4140
rect 8481 4131 8539 4137
rect 8481 4128 8493 4131
rect 8352 4100 8493 4128
rect 8352 4088 8358 4100
rect 8481 4097 8493 4100
rect 8527 4128 8539 4131
rect 8938 4128 8944 4140
rect 8527 4100 8944 4128
rect 8527 4097 8539 4100
rect 8481 4091 8539 4097
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 9122 4128 9128 4140
rect 9083 4100 9128 4128
rect 9122 4088 9128 4100
rect 9180 4088 9186 4140
rect 10428 4137 10456 4168
rect 10502 4156 10508 4168
rect 10560 4156 10566 4208
rect 11698 4156 11704 4208
rect 11756 4196 11762 4208
rect 12342 4196 12348 4208
rect 11756 4168 11836 4196
rect 11756 4156 11762 4168
rect 11808 4137 11836 4168
rect 11900 4168 12348 4196
rect 11900 4137 11928 4168
rect 12342 4156 12348 4168
rect 12400 4156 12406 4208
rect 12526 4156 12532 4208
rect 12584 4196 12590 4208
rect 12710 4196 12716 4208
rect 12584 4168 12716 4196
rect 12584 4156 12590 4168
rect 12710 4156 12716 4168
rect 12768 4156 12774 4208
rect 12894 4196 12900 4208
rect 12855 4168 12900 4196
rect 12894 4156 12900 4168
rect 12952 4196 12958 4208
rect 13262 4196 13268 4208
rect 12952 4168 13268 4196
rect 12952 4156 12958 4168
rect 13262 4156 13268 4168
rect 13320 4156 13326 4208
rect 13648 4196 13676 4236
rect 15102 4224 15108 4236
rect 15160 4224 15166 4276
rect 17494 4264 17500 4276
rect 17407 4236 17500 4264
rect 17494 4224 17500 4236
rect 17552 4264 17558 4276
rect 18782 4264 18788 4276
rect 17552 4236 18788 4264
rect 17552 4224 17558 4236
rect 18782 4224 18788 4236
rect 18840 4224 18846 4276
rect 19426 4264 19432 4276
rect 19387 4236 19432 4264
rect 19426 4224 19432 4236
rect 19484 4224 19490 4276
rect 19521 4267 19579 4273
rect 19521 4233 19533 4267
rect 19567 4264 19579 4267
rect 19702 4264 19708 4276
rect 19567 4236 19708 4264
rect 19567 4233 19579 4236
rect 19521 4227 19579 4233
rect 19702 4224 19708 4236
rect 19760 4224 19766 4276
rect 13814 4196 13820 4208
rect 13648 4168 13820 4196
rect 9217 4131 9275 4137
rect 9217 4097 9229 4131
rect 9263 4097 9275 4131
rect 10413 4131 10471 4137
rect 9217 4091 9275 4097
rect 9508 4100 9812 4128
rect 2777 4063 2835 4069
rect 2777 4029 2789 4063
rect 2823 4060 2835 4063
rect 2866 4060 2872 4072
rect 2823 4032 2872 4060
rect 2823 4029 2835 4032
rect 2777 4023 2835 4029
rect 2866 4020 2872 4032
rect 2924 4020 2930 4072
rect 6917 4063 6975 4069
rect 6917 4029 6929 4063
rect 6963 4060 6975 4063
rect 7006 4060 7012 4072
rect 6963 4032 7012 4060
rect 6963 4029 6975 4032
rect 6917 4023 6975 4029
rect 7006 4020 7012 4032
rect 7064 4020 7070 4072
rect 7742 4020 7748 4072
rect 7800 4060 7806 4072
rect 9232 4060 9260 4091
rect 9508 4072 9536 4100
rect 7800 4032 9260 4060
rect 7800 4020 7806 4032
rect 9490 4020 9496 4072
rect 9548 4020 9554 4072
rect 9585 4063 9643 4069
rect 9585 4029 9597 4063
rect 9631 4060 9643 4063
rect 9674 4060 9680 4072
rect 9631 4032 9680 4060
rect 9631 4029 9643 4032
rect 9585 4023 9643 4029
rect 9674 4020 9680 4032
rect 9732 4020 9738 4072
rect 3044 3995 3102 4001
rect 3044 3961 3056 3995
rect 3090 3992 3102 3995
rect 4246 3992 4252 4004
rect 3090 3964 4252 3992
rect 3090 3961 3102 3964
rect 3044 3955 3102 3961
rect 4246 3952 4252 3964
rect 4304 3952 4310 4004
rect 5442 3992 5448 4004
rect 5403 3964 5448 3992
rect 5442 3952 5448 3964
rect 5500 3952 5506 4004
rect 5902 3952 5908 4004
rect 5960 3992 5966 4004
rect 5960 3964 6592 3992
rect 5960 3952 5966 3964
rect 1670 3884 1676 3936
rect 1728 3924 1734 3936
rect 1949 3927 2007 3933
rect 1949 3924 1961 3927
rect 1728 3896 1961 3924
rect 1728 3884 1734 3896
rect 1949 3893 1961 3896
rect 1995 3893 2007 3927
rect 2314 3924 2320 3936
rect 2275 3896 2320 3924
rect 1949 3887 2007 3893
rect 2314 3884 2320 3896
rect 2372 3884 2378 3936
rect 4982 3924 4988 3936
rect 4943 3896 4988 3924
rect 4982 3884 4988 3896
rect 5040 3884 5046 3936
rect 5258 3884 5264 3936
rect 5316 3924 5322 3936
rect 5353 3927 5411 3933
rect 5353 3924 5365 3927
rect 5316 3896 5365 3924
rect 5316 3884 5322 3896
rect 5353 3893 5365 3896
rect 5399 3893 5411 3927
rect 5810 3924 5816 3936
rect 5771 3896 5816 3924
rect 5353 3887 5411 3893
rect 5810 3884 5816 3896
rect 5868 3884 5874 3936
rect 6181 3927 6239 3933
rect 6181 3893 6193 3927
rect 6227 3924 6239 3927
rect 6454 3924 6460 3936
rect 6227 3896 6460 3924
rect 6227 3893 6239 3896
rect 6181 3887 6239 3893
rect 6454 3884 6460 3896
rect 6512 3884 6518 3936
rect 6564 3924 6592 3964
rect 6638 3952 6644 4004
rect 6696 3992 6702 4004
rect 7184 3995 7242 4001
rect 7184 3992 7196 3995
rect 6696 3964 7196 3992
rect 6696 3952 6702 3964
rect 7184 3961 7196 3964
rect 7230 3992 7242 3995
rect 8202 3992 8208 4004
rect 7230 3964 8208 3992
rect 7230 3961 7242 3964
rect 7184 3955 7242 3961
rect 8202 3952 8208 3964
rect 8260 3952 8266 4004
rect 9033 3995 9091 4001
rect 9033 3961 9045 3995
rect 9079 3992 9091 3995
rect 9784 3992 9812 4100
rect 10413 4097 10425 4131
rect 10459 4097 10471 4131
rect 10413 4091 10471 4097
rect 11793 4131 11851 4137
rect 11793 4097 11805 4131
rect 11839 4097 11851 4131
rect 11793 4091 11851 4097
rect 11885 4131 11943 4137
rect 11885 4097 11897 4131
rect 11931 4097 11943 4131
rect 11885 4091 11943 4097
rect 11974 4088 11980 4140
rect 12032 4128 12038 4140
rect 13648 4137 13676 4168
rect 13814 4156 13820 4168
rect 13872 4156 13878 4208
rect 14921 4199 14979 4205
rect 14921 4165 14933 4199
rect 14967 4165 14979 4199
rect 14921 4159 14979 4165
rect 12161 4131 12219 4137
rect 12161 4128 12173 4131
rect 12032 4100 12173 4128
rect 12032 4088 12038 4100
rect 12161 4097 12173 4100
rect 12207 4097 12219 4131
rect 12161 4091 12219 4097
rect 13633 4131 13691 4137
rect 13633 4097 13645 4131
rect 13679 4097 13691 4131
rect 14458 4128 14464 4140
rect 14419 4100 14464 4128
rect 13633 4091 13691 4097
rect 14458 4088 14464 4100
rect 14516 4088 14522 4140
rect 9858 4020 9864 4072
rect 9916 4060 9922 4072
rect 10229 4063 10287 4069
rect 10229 4060 10241 4063
rect 9916 4032 10241 4060
rect 9916 4020 9922 4032
rect 10229 4029 10241 4032
rect 10275 4029 10287 4063
rect 10229 4023 10287 4029
rect 10321 4063 10379 4069
rect 10321 4029 10333 4063
rect 10367 4060 10379 4063
rect 10594 4060 10600 4072
rect 10367 4032 10600 4060
rect 10367 4029 10379 4032
rect 10321 4023 10379 4029
rect 10594 4020 10600 4032
rect 10652 4020 10658 4072
rect 11146 4020 11152 4072
rect 11204 4060 11210 4072
rect 11701 4063 11759 4069
rect 11701 4060 11713 4063
rect 11204 4032 11713 4060
rect 11204 4020 11210 4032
rect 11701 4029 11713 4032
rect 11747 4029 11759 4063
rect 13354 4060 13360 4072
rect 13315 4032 13360 4060
rect 11701 4023 11759 4029
rect 13354 4020 13360 4032
rect 13412 4020 13418 4072
rect 13449 4063 13507 4069
rect 13449 4029 13461 4063
rect 13495 4060 13507 4063
rect 14182 4060 14188 4072
rect 13495 4032 14188 4060
rect 13495 4029 13507 4032
rect 13449 4023 13507 4029
rect 14182 4020 14188 4032
rect 14240 4020 14246 4072
rect 14550 4020 14556 4072
rect 14608 4060 14614 4072
rect 14737 4063 14795 4069
rect 14737 4060 14749 4063
rect 14608 4032 14749 4060
rect 14608 4020 14614 4032
rect 14737 4029 14749 4032
rect 14783 4029 14795 4063
rect 14936 4060 14964 4159
rect 15470 4156 15476 4208
rect 15528 4196 15534 4208
rect 15528 4168 16068 4196
rect 15528 4156 15534 4168
rect 16040 4140 16068 4168
rect 15562 4128 15568 4140
rect 15523 4100 15568 4128
rect 15562 4088 15568 4100
rect 15620 4088 15626 4140
rect 15749 4131 15807 4137
rect 15749 4097 15761 4131
rect 15795 4128 15807 4131
rect 15838 4128 15844 4140
rect 15795 4100 15844 4128
rect 15795 4097 15807 4100
rect 15749 4091 15807 4097
rect 15838 4088 15844 4100
rect 15896 4088 15902 4140
rect 16022 4088 16028 4140
rect 16080 4128 16086 4140
rect 16117 4131 16175 4137
rect 16117 4128 16129 4131
rect 16080 4100 16129 4128
rect 16080 4088 16086 4100
rect 16117 4097 16129 4100
rect 16163 4097 16175 4131
rect 16117 4091 16175 4097
rect 19518 4088 19524 4140
rect 19576 4128 19582 4140
rect 20073 4131 20131 4137
rect 20073 4128 20085 4131
rect 19576 4100 20085 4128
rect 19576 4088 19582 4100
rect 20073 4097 20085 4100
rect 20119 4097 20131 4131
rect 20073 4091 20131 4097
rect 21542 4088 21548 4140
rect 21600 4128 21606 4140
rect 22738 4128 22744 4140
rect 21600 4100 22744 4128
rect 21600 4088 21606 4100
rect 22738 4088 22744 4100
rect 22796 4088 22802 4140
rect 16390 4069 16396 4072
rect 16384 4060 16396 4069
rect 14936 4032 16252 4060
rect 16351 4032 16396 4060
rect 14737 4023 14795 4029
rect 12621 3995 12679 4001
rect 12621 3992 12633 3995
rect 9079 3964 9720 3992
rect 9784 3964 12633 3992
rect 9079 3961 9091 3964
rect 9033 3955 9091 3961
rect 7466 3924 7472 3936
rect 6564 3896 7472 3924
rect 7466 3884 7472 3896
rect 7524 3884 7530 3936
rect 7558 3884 7564 3936
rect 7616 3924 7622 3936
rect 8297 3927 8355 3933
rect 8297 3924 8309 3927
rect 7616 3896 8309 3924
rect 7616 3884 7622 3896
rect 8297 3893 8309 3896
rect 8343 3893 8355 3927
rect 8297 3887 8355 3893
rect 8665 3927 8723 3933
rect 8665 3893 8677 3927
rect 8711 3924 8723 3927
rect 8846 3924 8852 3936
rect 8711 3896 8852 3924
rect 8711 3893 8723 3896
rect 8665 3887 8723 3893
rect 8846 3884 8852 3896
rect 8904 3884 8910 3936
rect 8938 3884 8944 3936
rect 8996 3924 9002 3936
rect 9490 3924 9496 3936
rect 8996 3896 9496 3924
rect 8996 3884 9002 3896
rect 9490 3884 9496 3896
rect 9548 3884 9554 3936
rect 9692 3924 9720 3964
rect 12621 3961 12633 3964
rect 12667 3992 12679 3995
rect 12802 3992 12808 4004
rect 12667 3964 12808 3992
rect 12667 3961 12679 3964
rect 12621 3955 12679 3961
rect 12802 3952 12808 3964
rect 12860 3952 12866 4004
rect 14277 3995 14335 4001
rect 14277 3992 14289 3995
rect 13004 3964 14289 3992
rect 9766 3924 9772 3936
rect 9692 3896 9772 3924
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 9861 3927 9919 3933
rect 9861 3893 9873 3927
rect 9907 3924 9919 3927
rect 11238 3924 11244 3936
rect 9907 3896 11244 3924
rect 9907 3893 9919 3896
rect 9861 3887 9919 3893
rect 11238 3884 11244 3896
rect 11296 3884 11302 3936
rect 11333 3927 11391 3933
rect 11333 3893 11345 3927
rect 11379 3924 11391 3927
rect 12434 3924 12440 3936
rect 11379 3896 12440 3924
rect 11379 3893 11391 3896
rect 11333 3887 11391 3893
rect 12434 3884 12440 3896
rect 12492 3884 12498 3936
rect 12529 3927 12587 3933
rect 12529 3893 12541 3927
rect 12575 3924 12587 3927
rect 12894 3924 12900 3936
rect 12575 3896 12900 3924
rect 12575 3893 12587 3896
rect 12529 3887 12587 3893
rect 12894 3884 12900 3896
rect 12952 3884 12958 3936
rect 13004 3933 13032 3964
rect 14277 3961 14289 3964
rect 14323 3961 14335 3995
rect 15933 3995 15991 4001
rect 15933 3992 15945 3995
rect 14277 3955 14335 3961
rect 15488 3964 15945 3992
rect 15488 3936 15516 3964
rect 15933 3961 15945 3964
rect 15979 3961 15991 3995
rect 16224 3992 16252 4032
rect 16384 4023 16396 4032
rect 16390 4020 16396 4023
rect 16448 4020 16454 4072
rect 16666 4020 16672 4072
rect 16724 4060 16730 4072
rect 17954 4060 17960 4072
rect 16724 4032 17960 4060
rect 16724 4020 16730 4032
rect 17954 4020 17960 4032
rect 18012 4060 18018 4072
rect 18056 4063 18114 4069
rect 18056 4060 18068 4063
rect 18012 4032 18068 4060
rect 18012 4020 18018 4032
rect 18056 4029 18068 4032
rect 18102 4029 18114 4063
rect 18056 4023 18114 4029
rect 19426 4020 19432 4072
rect 19484 4060 19490 4072
rect 20714 4060 20720 4072
rect 19484 4032 20720 4060
rect 19484 4020 19490 4032
rect 20714 4020 20720 4032
rect 20772 4020 20778 4072
rect 17862 3992 17868 4004
rect 16224 3964 17724 3992
rect 17823 3964 17868 3992
rect 15933 3955 15991 3961
rect 12989 3927 13047 3933
rect 12989 3893 13001 3927
rect 13035 3893 13047 3927
rect 12989 3887 13047 3893
rect 13078 3884 13084 3936
rect 13136 3924 13142 3936
rect 13817 3927 13875 3933
rect 13817 3924 13829 3927
rect 13136 3896 13829 3924
rect 13136 3884 13142 3896
rect 13817 3893 13829 3896
rect 13863 3893 13875 3927
rect 14182 3924 14188 3936
rect 14143 3896 14188 3924
rect 13817 3887 13875 3893
rect 14182 3884 14188 3896
rect 14240 3884 14246 3936
rect 15470 3924 15476 3936
rect 15431 3896 15476 3924
rect 15470 3884 15476 3896
rect 15528 3884 15534 3936
rect 16114 3884 16120 3936
rect 16172 3924 16178 3936
rect 17589 3927 17647 3933
rect 17589 3924 17601 3927
rect 16172 3896 17601 3924
rect 16172 3884 16178 3896
rect 17589 3893 17601 3896
rect 17635 3893 17647 3927
rect 17696 3924 17724 3964
rect 17862 3952 17868 3964
rect 17920 3952 17926 4004
rect 18294 3995 18352 4001
rect 18294 3992 18306 3995
rect 18064 3964 18306 3992
rect 18064 3936 18092 3964
rect 18294 3961 18306 3964
rect 18340 3961 18352 3995
rect 18294 3955 18352 3961
rect 20622 3952 20628 4004
rect 20680 3992 20686 4004
rect 22278 3992 22284 4004
rect 20680 3964 22284 3992
rect 20680 3952 20686 3964
rect 22278 3952 22284 3964
rect 22336 3952 22342 4004
rect 17954 3924 17960 3936
rect 17696 3896 17960 3924
rect 17589 3887 17647 3893
rect 17954 3884 17960 3896
rect 18012 3884 18018 3936
rect 18046 3884 18052 3936
rect 18104 3884 18110 3936
rect 19334 3884 19340 3936
rect 19392 3924 19398 3936
rect 19702 3924 19708 3936
rect 19392 3896 19708 3924
rect 19392 3884 19398 3896
rect 19702 3884 19708 3896
rect 19760 3884 19766 3936
rect 19794 3884 19800 3936
rect 19852 3924 19858 3936
rect 19889 3927 19947 3933
rect 19889 3924 19901 3927
rect 19852 3896 19901 3924
rect 19852 3884 19858 3896
rect 19889 3893 19901 3896
rect 19935 3893 19947 3927
rect 19889 3887 19947 3893
rect 19978 3884 19984 3936
rect 20036 3924 20042 3936
rect 20349 3927 20407 3933
rect 20349 3924 20361 3927
rect 20036 3896 20361 3924
rect 20036 3884 20042 3896
rect 20349 3893 20361 3896
rect 20395 3893 20407 3927
rect 20349 3887 20407 3893
rect 1104 3834 21896 3856
rect 1104 3782 7912 3834
rect 7964 3782 7976 3834
rect 8028 3782 8040 3834
rect 8092 3782 8104 3834
rect 8156 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 15035 3834
rect 15087 3782 21896 3834
rect 1104 3760 21896 3782
rect 2314 3720 2320 3732
rect 2275 3692 2320 3720
rect 2314 3680 2320 3692
rect 2372 3680 2378 3732
rect 3145 3723 3203 3729
rect 3145 3689 3157 3723
rect 3191 3720 3203 3723
rect 3510 3720 3516 3732
rect 3191 3692 3516 3720
rect 3191 3689 3203 3692
rect 3145 3683 3203 3689
rect 3510 3680 3516 3692
rect 3568 3680 3574 3732
rect 3605 3723 3663 3729
rect 3605 3689 3617 3723
rect 3651 3720 3663 3723
rect 4798 3720 4804 3732
rect 3651 3692 4804 3720
rect 3651 3689 3663 3692
rect 3605 3683 3663 3689
rect 4798 3680 4804 3692
rect 4856 3680 4862 3732
rect 5445 3723 5503 3729
rect 5445 3689 5457 3723
rect 5491 3689 5503 3723
rect 5902 3720 5908 3732
rect 5863 3692 5908 3720
rect 5445 3683 5503 3689
rect 2777 3655 2835 3661
rect 2777 3621 2789 3655
rect 2823 3621 2835 3655
rect 2777 3615 2835 3621
rect 2498 3544 2504 3596
rect 2556 3584 2562 3596
rect 2685 3587 2743 3593
rect 2685 3584 2697 3587
rect 2556 3556 2697 3584
rect 2556 3544 2562 3556
rect 2685 3553 2697 3556
rect 2731 3553 2743 3587
rect 2792 3584 2820 3615
rect 3786 3612 3792 3664
rect 3844 3652 3850 3664
rect 3844 3624 4108 3652
rect 3844 3612 3850 3624
rect 3050 3584 3056 3596
rect 2792 3556 3056 3584
rect 2685 3547 2743 3553
rect 3050 3544 3056 3556
rect 3108 3544 3114 3596
rect 3513 3587 3571 3593
rect 3513 3553 3525 3587
rect 3559 3584 3571 3587
rect 3694 3584 3700 3596
rect 3559 3556 3700 3584
rect 3559 3553 3571 3556
rect 3513 3547 3571 3553
rect 3694 3544 3700 3556
rect 3752 3544 3758 3596
rect 4080 3593 4108 3624
rect 4154 3612 4160 3664
rect 4212 3652 4218 3664
rect 4310 3655 4368 3661
rect 4310 3652 4322 3655
rect 4212 3624 4322 3652
rect 4212 3612 4218 3624
rect 4310 3621 4322 3624
rect 4356 3621 4368 3655
rect 5460 3652 5488 3683
rect 5902 3680 5908 3692
rect 5960 3680 5966 3732
rect 6273 3723 6331 3729
rect 6273 3689 6285 3723
rect 6319 3720 6331 3723
rect 7374 3720 7380 3732
rect 6319 3692 7380 3720
rect 6319 3689 6331 3692
rect 6273 3683 6331 3689
rect 7374 3680 7380 3692
rect 7432 3680 7438 3732
rect 8113 3723 8171 3729
rect 8113 3689 8125 3723
rect 8159 3720 8171 3723
rect 8202 3720 8208 3732
rect 8159 3692 8208 3720
rect 8159 3689 8171 3692
rect 8113 3683 8171 3689
rect 8202 3680 8208 3692
rect 8260 3680 8266 3732
rect 8662 3680 8668 3732
rect 8720 3720 8726 3732
rect 8757 3723 8815 3729
rect 8757 3720 8769 3723
rect 8720 3692 8769 3720
rect 8720 3680 8726 3692
rect 8757 3689 8769 3692
rect 8803 3689 8815 3723
rect 9674 3720 9680 3732
rect 8757 3683 8815 3689
rect 9048 3692 9680 3720
rect 6730 3652 6736 3664
rect 5460 3624 6736 3652
rect 4310 3615 4368 3621
rect 6730 3612 6736 3624
rect 6788 3612 6794 3664
rect 6914 3612 6920 3664
rect 6972 3661 6978 3664
rect 6972 3655 7036 3661
rect 6972 3621 6990 3655
rect 7024 3621 7036 3655
rect 8570 3652 8576 3664
rect 8531 3624 8576 3652
rect 6972 3615 7036 3621
rect 6972 3612 6978 3615
rect 8570 3612 8576 3624
rect 8628 3652 8634 3664
rect 8938 3652 8944 3664
rect 8628 3624 8944 3652
rect 8628 3612 8634 3624
rect 8938 3612 8944 3624
rect 8996 3612 9002 3664
rect 4065 3587 4123 3593
rect 4065 3553 4077 3587
rect 4111 3553 4123 3587
rect 4065 3547 4123 3553
rect 7466 3544 7472 3596
rect 7524 3584 7530 3596
rect 8481 3587 8539 3593
rect 8481 3584 8493 3587
rect 7524 3556 8493 3584
rect 7524 3544 7530 3556
rect 8481 3553 8493 3556
rect 8527 3584 8539 3587
rect 9048 3584 9076 3692
rect 9674 3680 9680 3692
rect 9732 3680 9738 3732
rect 9858 3680 9864 3732
rect 9916 3720 9922 3732
rect 10226 3720 10232 3732
rect 9916 3692 10232 3720
rect 9916 3680 9922 3692
rect 10226 3680 10232 3692
rect 10284 3680 10290 3732
rect 10962 3680 10968 3732
rect 11020 3720 11026 3732
rect 11146 3720 11152 3732
rect 11020 3692 11152 3720
rect 11020 3680 11026 3692
rect 11146 3680 11152 3692
rect 11204 3680 11210 3732
rect 12897 3723 12955 3729
rect 12897 3689 12909 3723
rect 12943 3689 12955 3723
rect 12897 3683 12955 3689
rect 9214 3652 9220 3664
rect 9175 3624 9220 3652
rect 9214 3612 9220 3624
rect 9272 3612 9278 3664
rect 9398 3652 9404 3664
rect 9324 3624 9404 3652
rect 8527 3556 9076 3584
rect 9125 3587 9183 3593
rect 8527 3553 8539 3556
rect 8481 3547 8539 3553
rect 9125 3553 9137 3587
rect 9171 3584 9183 3587
rect 9324 3584 9352 3624
rect 9398 3612 9404 3624
rect 9456 3612 9462 3664
rect 12434 3652 12440 3664
rect 11532 3624 12440 3652
rect 9944 3587 10002 3593
rect 9944 3584 9956 3587
rect 9171 3556 9352 3584
rect 9416 3556 9956 3584
rect 9171 3553 9183 3556
rect 9125 3547 9183 3553
rect 2961 3519 3019 3525
rect 2961 3485 2973 3519
rect 3007 3485 3019 3519
rect 2961 3479 3019 3485
rect 3789 3519 3847 3525
rect 3789 3485 3801 3519
rect 3835 3485 3847 3519
rect 3789 3479 3847 3485
rect 2682 3408 2688 3460
rect 2740 3448 2746 3460
rect 2976 3448 3004 3479
rect 2740 3420 3004 3448
rect 2740 3408 2746 3420
rect 3510 3340 3516 3392
rect 3568 3380 3574 3392
rect 3804 3380 3832 3479
rect 5902 3476 5908 3528
rect 5960 3516 5966 3528
rect 6365 3519 6423 3525
rect 6365 3516 6377 3519
rect 5960 3488 6377 3516
rect 5960 3476 5966 3488
rect 6365 3485 6377 3488
rect 6411 3485 6423 3519
rect 6365 3479 6423 3485
rect 6549 3519 6607 3525
rect 6549 3485 6561 3519
rect 6595 3516 6607 3519
rect 6638 3516 6644 3528
rect 6595 3488 6644 3516
rect 6595 3485 6607 3488
rect 6549 3479 6607 3485
rect 6638 3476 6644 3488
rect 6696 3476 6702 3528
rect 9416 3525 9444 3556
rect 9944 3553 9956 3556
rect 9990 3584 10002 3587
rect 10962 3584 10968 3596
rect 9990 3556 10968 3584
rect 9990 3553 10002 3556
rect 9944 3547 10002 3553
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 11532 3593 11560 3624
rect 12434 3612 12440 3624
rect 12492 3652 12498 3664
rect 12618 3652 12624 3664
rect 12492 3624 12624 3652
rect 12492 3612 12498 3624
rect 12618 3612 12624 3624
rect 12676 3612 12682 3664
rect 12710 3612 12716 3664
rect 12768 3652 12774 3664
rect 12912 3652 12940 3683
rect 12986 3680 12992 3732
rect 13044 3720 13050 3732
rect 13449 3723 13507 3729
rect 13449 3720 13461 3723
rect 13044 3692 13461 3720
rect 13044 3680 13050 3692
rect 13449 3689 13461 3692
rect 13495 3689 13507 3723
rect 13449 3683 13507 3689
rect 14090 3680 14096 3732
rect 14148 3720 14154 3732
rect 14277 3723 14335 3729
rect 14277 3720 14289 3723
rect 14148 3692 14289 3720
rect 14148 3680 14154 3692
rect 14277 3689 14289 3692
rect 14323 3720 14335 3723
rect 15013 3723 15071 3729
rect 15013 3720 15025 3723
rect 14323 3692 15025 3720
rect 14323 3689 14335 3692
rect 14277 3683 14335 3689
rect 15013 3689 15025 3692
rect 15059 3720 15071 3723
rect 15194 3720 15200 3732
rect 15059 3692 15200 3720
rect 15059 3689 15071 3692
rect 15013 3683 15071 3689
rect 15194 3680 15200 3692
rect 15252 3680 15258 3732
rect 16301 3723 16359 3729
rect 16301 3689 16313 3723
rect 16347 3720 16359 3723
rect 16758 3720 16764 3732
rect 16347 3692 16764 3720
rect 16347 3689 16359 3692
rect 16301 3683 16359 3689
rect 16758 3680 16764 3692
rect 16816 3680 16822 3732
rect 18138 3680 18144 3732
rect 18196 3720 18202 3732
rect 18969 3723 19027 3729
rect 18969 3720 18981 3723
rect 18196 3692 18981 3720
rect 18196 3680 18202 3692
rect 18969 3689 18981 3692
rect 19015 3689 19027 3723
rect 19794 3720 19800 3732
rect 19755 3692 19800 3720
rect 18969 3683 19027 3689
rect 19794 3680 19800 3692
rect 19852 3680 19858 3732
rect 20165 3723 20223 3729
rect 20165 3689 20177 3723
rect 20211 3720 20223 3723
rect 20254 3720 20260 3732
rect 20211 3692 20260 3720
rect 20211 3689 20223 3692
rect 20165 3683 20223 3689
rect 20254 3680 20260 3692
rect 20312 3680 20318 3732
rect 14458 3652 14464 3664
rect 12768 3624 14464 3652
rect 12768 3612 12774 3624
rect 14458 3612 14464 3624
rect 14516 3612 14522 3664
rect 15286 3612 15292 3664
rect 15344 3652 15350 3664
rect 19429 3655 19487 3661
rect 19429 3652 19441 3655
rect 15344 3624 19441 3652
rect 15344 3612 15350 3624
rect 19429 3621 19441 3624
rect 19475 3621 19487 3655
rect 19429 3615 19487 3621
rect 11517 3587 11575 3593
rect 11517 3553 11529 3587
rect 11563 3553 11575 3587
rect 11517 3547 11575 3553
rect 11784 3587 11842 3593
rect 11784 3553 11796 3587
rect 11830 3584 11842 3587
rect 12342 3584 12348 3596
rect 11830 3556 12348 3584
rect 11830 3553 11842 3556
rect 11784 3547 11842 3553
rect 12342 3544 12348 3556
rect 12400 3544 12406 3596
rect 13354 3544 13360 3596
rect 13412 3584 13418 3596
rect 14182 3584 14188 3596
rect 13412 3556 13457 3584
rect 14143 3556 14188 3584
rect 13412 3544 13418 3556
rect 14182 3544 14188 3556
rect 14240 3544 14246 3596
rect 14642 3584 14648 3596
rect 14603 3556 14648 3584
rect 14642 3544 14648 3556
rect 14700 3584 14706 3596
rect 15102 3584 15108 3596
rect 14700 3556 15108 3584
rect 14700 3544 14706 3556
rect 15102 3544 15108 3556
rect 15160 3584 15166 3596
rect 15657 3587 15715 3593
rect 15657 3584 15669 3587
rect 15160 3556 15669 3584
rect 15160 3544 15166 3556
rect 15657 3553 15669 3556
rect 15703 3553 15715 3587
rect 16114 3584 16120 3596
rect 16075 3556 16120 3584
rect 15657 3547 15715 3553
rect 16114 3544 16120 3556
rect 16172 3544 16178 3596
rect 16936 3587 16994 3593
rect 16936 3584 16948 3587
rect 16500 3556 16948 3584
rect 6733 3519 6791 3525
rect 6733 3485 6745 3519
rect 6779 3485 6791 3519
rect 6733 3479 6791 3485
rect 9401 3519 9459 3525
rect 9401 3485 9413 3519
rect 9447 3485 9459 3519
rect 9401 3479 9459 3485
rect 4246 3380 4252 3392
rect 3568 3352 4252 3380
rect 3568 3340 3574 3352
rect 4246 3340 4252 3352
rect 4304 3340 4310 3392
rect 5813 3383 5871 3389
rect 5813 3349 5825 3383
rect 5859 3380 5871 3383
rect 6086 3380 6092 3392
rect 5859 3352 6092 3380
rect 5859 3349 5871 3352
rect 5813 3343 5871 3349
rect 6086 3340 6092 3352
rect 6144 3340 6150 3392
rect 6748 3380 6776 3479
rect 9490 3476 9496 3528
rect 9548 3516 9554 3528
rect 9677 3519 9735 3525
rect 9677 3516 9689 3519
rect 9548 3488 9689 3516
rect 9548 3476 9554 3488
rect 9677 3485 9689 3488
rect 9723 3485 9735 3519
rect 9677 3479 9735 3485
rect 10686 3476 10692 3528
rect 10744 3516 10750 3528
rect 11149 3519 11207 3525
rect 11149 3516 11161 3519
rect 10744 3488 11161 3516
rect 10744 3476 10750 3488
rect 11149 3485 11161 3488
rect 11195 3485 11207 3519
rect 11149 3479 11207 3485
rect 13633 3519 13691 3525
rect 13633 3485 13645 3519
rect 13679 3516 13691 3519
rect 13814 3516 13820 3528
rect 13679 3488 13820 3516
rect 13679 3485 13691 3488
rect 13633 3479 13691 3485
rect 13814 3476 13820 3488
rect 13872 3516 13878 3528
rect 14369 3519 14427 3525
rect 14369 3516 14381 3519
rect 13872 3488 14381 3516
rect 13872 3476 13878 3488
rect 14369 3485 14381 3488
rect 14415 3485 14427 3519
rect 15746 3516 15752 3528
rect 15707 3488 15752 3516
rect 14369 3479 14427 3485
rect 15746 3476 15752 3488
rect 15804 3476 15810 3528
rect 15838 3476 15844 3528
rect 15896 3516 15902 3528
rect 16500 3516 16528 3556
rect 16936 3553 16948 3556
rect 16982 3584 16994 3587
rect 17494 3584 17500 3596
rect 16982 3556 17500 3584
rect 16982 3553 16994 3556
rect 16936 3547 16994 3553
rect 17494 3544 17500 3556
rect 17552 3544 17558 3596
rect 17862 3544 17868 3596
rect 17920 3584 17926 3596
rect 18509 3587 18567 3593
rect 18509 3584 18521 3587
rect 17920 3556 18521 3584
rect 17920 3544 17926 3556
rect 18509 3553 18521 3556
rect 18555 3553 18567 3587
rect 19334 3584 19340 3596
rect 19295 3556 19340 3584
rect 18509 3547 18567 3553
rect 19334 3544 19340 3556
rect 19392 3544 19398 3596
rect 16666 3516 16672 3528
rect 15896 3488 16528 3516
rect 16627 3488 16672 3516
rect 15896 3476 15902 3488
rect 16666 3476 16672 3488
rect 16724 3476 16730 3528
rect 18598 3516 18604 3528
rect 18559 3488 18604 3516
rect 18598 3476 18604 3488
rect 18656 3476 18662 3528
rect 18782 3516 18788 3528
rect 18743 3488 18788 3516
rect 18782 3476 18788 3488
rect 18840 3476 18846 3528
rect 19518 3516 19524 3528
rect 19431 3488 19524 3516
rect 19518 3476 19524 3488
rect 19576 3476 19582 3528
rect 7834 3408 7840 3460
rect 7892 3448 7898 3460
rect 9508 3448 9536 3476
rect 15930 3448 15936 3460
rect 7892 3420 9536 3448
rect 12728 3420 15936 3448
rect 7892 3408 7898 3420
rect 7006 3380 7012 3392
rect 6748 3352 7012 3380
rect 7006 3340 7012 3352
rect 7064 3340 7070 3392
rect 8297 3383 8355 3389
rect 8297 3349 8309 3383
rect 8343 3380 8355 3383
rect 8662 3380 8668 3392
rect 8343 3352 8668 3380
rect 8343 3349 8355 3352
rect 8297 3343 8355 3349
rect 8662 3340 8668 3352
rect 8720 3380 8726 3392
rect 9306 3380 9312 3392
rect 8720 3352 9312 3380
rect 8720 3340 8726 3352
rect 9306 3340 9312 3352
rect 9364 3340 9370 3392
rect 9582 3340 9588 3392
rect 9640 3380 9646 3392
rect 10410 3380 10416 3392
rect 9640 3352 10416 3380
rect 9640 3340 9646 3352
rect 10410 3340 10416 3352
rect 10468 3380 10474 3392
rect 11057 3383 11115 3389
rect 11057 3380 11069 3383
rect 10468 3352 11069 3380
rect 10468 3340 10474 3352
rect 11057 3349 11069 3352
rect 11103 3349 11115 3383
rect 11057 3343 11115 3349
rect 11238 3340 11244 3392
rect 11296 3380 11302 3392
rect 12728 3380 12756 3420
rect 15930 3408 15936 3420
rect 15988 3408 15994 3460
rect 16022 3408 16028 3460
rect 16080 3448 16086 3460
rect 16684 3448 16712 3476
rect 19536 3448 19564 3476
rect 16080 3420 16712 3448
rect 18064 3420 19564 3448
rect 16080 3408 16086 3420
rect 18064 3392 18092 3420
rect 11296 3352 12756 3380
rect 11296 3340 11302 3352
rect 12986 3340 12992 3392
rect 13044 3380 13050 3392
rect 13817 3383 13875 3389
rect 13044 3352 13089 3380
rect 13044 3340 13050 3352
rect 13817 3349 13829 3383
rect 13863 3380 13875 3383
rect 13906 3380 13912 3392
rect 13863 3352 13912 3380
rect 13863 3349 13875 3352
rect 13817 3343 13875 3349
rect 13906 3340 13912 3352
rect 13964 3340 13970 3392
rect 14734 3340 14740 3392
rect 14792 3380 14798 3392
rect 14829 3383 14887 3389
rect 14829 3380 14841 3383
rect 14792 3352 14841 3380
rect 14792 3340 14798 3352
rect 14829 3349 14841 3352
rect 14875 3349 14887 3383
rect 15286 3380 15292 3392
rect 15247 3352 15292 3380
rect 14829 3343 14887 3349
rect 15286 3340 15292 3352
rect 15344 3340 15350 3392
rect 15746 3340 15752 3392
rect 15804 3380 15810 3392
rect 16485 3383 16543 3389
rect 16485 3380 16497 3383
rect 15804 3352 16497 3380
rect 15804 3340 15810 3352
rect 16485 3349 16497 3352
rect 16531 3349 16543 3383
rect 18046 3380 18052 3392
rect 18007 3352 18052 3380
rect 16485 3343 16543 3349
rect 18046 3340 18052 3352
rect 18104 3340 18110 3392
rect 18138 3340 18144 3392
rect 18196 3380 18202 3392
rect 18196 3352 18241 3380
rect 18196 3340 18202 3352
rect 18598 3340 18604 3392
rect 18656 3380 18662 3392
rect 20346 3380 20352 3392
rect 18656 3352 20352 3380
rect 18656 3340 18662 3352
rect 20346 3340 20352 3352
rect 20404 3340 20410 3392
rect 1104 3290 21896 3312
rect 1104 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 4575 3290
rect 4627 3238 4639 3290
rect 4691 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 18308 3290
rect 18360 3238 18372 3290
rect 18424 3238 18436 3290
rect 18488 3238 18500 3290
rect 18552 3238 21896 3290
rect 1104 3216 21896 3238
rect 2498 3176 2504 3188
rect 2459 3148 2504 3176
rect 2498 3136 2504 3148
rect 2556 3136 2562 3188
rect 2866 3136 2872 3188
rect 2924 3136 2930 3188
rect 3050 3136 3056 3188
rect 3108 3176 3114 3188
rect 3329 3179 3387 3185
rect 3329 3176 3341 3179
rect 3108 3148 3341 3176
rect 3108 3136 3114 3148
rect 3329 3145 3341 3148
rect 3375 3145 3387 3179
rect 3329 3139 3387 3145
rect 3694 3136 3700 3188
rect 3752 3176 3758 3188
rect 5534 3176 5540 3188
rect 3752 3148 5540 3176
rect 3752 3136 3758 3148
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 5902 3176 5908 3188
rect 5863 3148 5908 3176
rect 5902 3136 5908 3148
rect 5960 3136 5966 3188
rect 6546 3136 6552 3188
rect 6604 3176 6610 3188
rect 6822 3176 6828 3188
rect 6604 3148 6828 3176
rect 6604 3136 6610 3148
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 7742 3176 7748 3188
rect 6932 3148 7748 3176
rect 2884 3108 2912 3136
rect 6932 3120 6960 3148
rect 7742 3136 7748 3148
rect 7800 3176 7806 3188
rect 8389 3179 8447 3185
rect 8389 3176 8401 3179
rect 7800 3148 8401 3176
rect 7800 3136 7806 3148
rect 8389 3145 8401 3148
rect 8435 3145 8447 3179
rect 8389 3139 8447 3145
rect 9033 3179 9091 3185
rect 9033 3145 9045 3179
rect 9079 3176 9091 3179
rect 9122 3176 9128 3188
rect 9079 3148 9128 3176
rect 9079 3145 9091 3148
rect 9033 3139 9091 3145
rect 9122 3136 9128 3148
rect 9180 3136 9186 3188
rect 12342 3136 12348 3188
rect 12400 3176 12406 3188
rect 13817 3179 13875 3185
rect 13817 3176 13829 3179
rect 12400 3148 13829 3176
rect 12400 3136 12406 3148
rect 13817 3145 13829 3148
rect 13863 3145 13875 3179
rect 13817 3139 13875 3145
rect 15102 3136 15108 3188
rect 15160 3176 15166 3188
rect 16853 3179 16911 3185
rect 16853 3176 16865 3179
rect 15160 3148 16865 3176
rect 15160 3136 15166 3148
rect 16853 3145 16865 3148
rect 16899 3145 16911 3179
rect 17126 3176 17132 3188
rect 17087 3148 17132 3176
rect 16853 3139 16911 3145
rect 17126 3136 17132 3148
rect 17184 3136 17190 3188
rect 18141 3179 18199 3185
rect 18141 3145 18153 3179
rect 18187 3176 18199 3179
rect 19334 3176 19340 3188
rect 18187 3148 19340 3176
rect 18187 3145 18199 3148
rect 18141 3139 18199 3145
rect 19334 3136 19340 3148
rect 19392 3136 19398 3188
rect 19518 3136 19524 3188
rect 19576 3176 19582 3188
rect 19702 3176 19708 3188
rect 19576 3148 19708 3176
rect 19576 3136 19582 3148
rect 19702 3136 19708 3148
rect 19760 3136 19766 3188
rect 3786 3108 3792 3120
rect 2884 3080 3792 3108
rect 3786 3068 3792 3080
rect 3844 3108 3850 3120
rect 6914 3108 6920 3120
rect 3844 3080 4384 3108
rect 3844 3068 3850 3080
rect 3145 3043 3203 3049
rect 3145 3009 3157 3043
rect 3191 3040 3203 3043
rect 3510 3040 3516 3052
rect 3191 3012 3516 3040
rect 3191 3009 3203 3012
rect 3145 3003 3203 3009
rect 3510 3000 3516 3012
rect 3568 3040 3574 3052
rect 4356 3049 4384 3080
rect 6564 3080 6920 3108
rect 6564 3049 6592 3080
rect 6914 3068 6920 3080
rect 6972 3068 6978 3120
rect 10962 3068 10968 3120
rect 11020 3108 11026 3120
rect 11241 3111 11299 3117
rect 11241 3108 11253 3111
rect 11020 3080 11253 3108
rect 11020 3068 11026 3080
rect 11241 3077 11253 3080
rect 11287 3077 11299 3111
rect 11241 3071 11299 3077
rect 12434 3068 12440 3120
rect 12492 3068 12498 3120
rect 13446 3068 13452 3120
rect 13504 3108 13510 3120
rect 18966 3108 18972 3120
rect 13504 3080 18972 3108
rect 13504 3068 13510 3080
rect 18966 3068 18972 3080
rect 19024 3068 19030 3120
rect 19058 3068 19064 3120
rect 19116 3108 19122 3120
rect 20898 3108 20904 3120
rect 19116 3080 20904 3108
rect 19116 3068 19122 3080
rect 20898 3068 20904 3080
rect 20956 3068 20962 3120
rect 3881 3043 3939 3049
rect 3881 3040 3893 3043
rect 3568 3012 3893 3040
rect 3568 3000 3574 3012
rect 3881 3009 3893 3012
rect 3927 3009 3939 3043
rect 3881 3003 3939 3009
rect 4341 3043 4399 3049
rect 4341 3009 4353 3043
rect 4387 3009 4399 3043
rect 4341 3003 4399 3009
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3009 6607 3043
rect 9582 3040 9588 3052
rect 9543 3012 9588 3040
rect 6549 3003 6607 3009
rect 9582 3000 9588 3012
rect 9640 3000 9646 3052
rect 12069 3043 12127 3049
rect 12069 3009 12081 3043
rect 12115 3009 12127 3043
rect 12069 3003 12127 3009
rect 2409 2975 2467 2981
rect 2409 2941 2421 2975
rect 2455 2972 2467 2975
rect 2774 2972 2780 2984
rect 2455 2944 2780 2972
rect 2455 2941 2467 2944
rect 2409 2935 2467 2941
rect 2774 2932 2780 2944
rect 2832 2972 2838 2984
rect 2961 2975 3019 2981
rect 2961 2972 2973 2975
rect 2832 2944 2973 2972
rect 2832 2932 2838 2944
rect 2961 2941 2973 2944
rect 3007 2972 3019 2975
rect 3418 2972 3424 2984
rect 3007 2944 3424 2972
rect 3007 2941 3019 2944
rect 2961 2935 3019 2941
rect 3418 2932 3424 2944
rect 3476 2932 3482 2984
rect 3694 2972 3700 2984
rect 3655 2944 3700 2972
rect 3694 2932 3700 2944
rect 3752 2932 3758 2984
rect 3789 2975 3847 2981
rect 3789 2941 3801 2975
rect 3835 2972 3847 2975
rect 4154 2972 4160 2984
rect 3835 2944 4160 2972
rect 3835 2941 3847 2944
rect 3789 2935 3847 2941
rect 4154 2932 4160 2944
rect 4212 2932 4218 2984
rect 6362 2972 6368 2984
rect 6323 2944 6368 2972
rect 6362 2932 6368 2944
rect 6420 2932 6426 2984
rect 7006 2972 7012 2984
rect 6919 2944 7012 2972
rect 7006 2932 7012 2944
rect 7064 2972 7070 2984
rect 7834 2972 7840 2984
rect 7064 2944 7840 2972
rect 7064 2932 7070 2944
rect 7834 2932 7840 2944
rect 7892 2932 7898 2984
rect 8478 2972 8484 2984
rect 8439 2944 8484 2972
rect 8478 2932 8484 2944
rect 8536 2932 8542 2984
rect 8757 2975 8815 2981
rect 8757 2941 8769 2975
rect 8803 2972 8815 2975
rect 9122 2972 9128 2984
rect 8803 2944 9128 2972
rect 8803 2941 8815 2944
rect 8757 2935 8815 2941
rect 9122 2932 9128 2944
rect 9180 2932 9186 2984
rect 9493 2975 9551 2981
rect 9493 2972 9505 2975
rect 9407 2944 9505 2972
rect 3510 2864 3516 2916
rect 3568 2904 3574 2916
rect 4062 2904 4068 2916
rect 3568 2876 4068 2904
rect 3568 2864 3574 2876
rect 4062 2864 4068 2876
rect 4120 2904 4126 2916
rect 4249 2907 4307 2913
rect 4249 2904 4261 2907
rect 4120 2876 4261 2904
rect 4120 2864 4126 2876
rect 4249 2873 4261 2876
rect 4295 2873 4307 2907
rect 4249 2867 4307 2873
rect 4608 2907 4666 2913
rect 4608 2873 4620 2907
rect 4654 2904 4666 2907
rect 4706 2904 4712 2916
rect 4654 2876 4712 2904
rect 4654 2873 4666 2876
rect 4608 2867 4666 2873
rect 4706 2864 4712 2876
rect 4764 2864 4770 2916
rect 6273 2907 6331 2913
rect 6273 2873 6285 2907
rect 6319 2904 6331 2907
rect 6730 2904 6736 2916
rect 6319 2876 6736 2904
rect 6319 2873 6331 2876
rect 6273 2867 6331 2873
rect 6730 2864 6736 2876
rect 6788 2864 6794 2916
rect 6914 2904 6920 2916
rect 6875 2876 6920 2904
rect 6914 2864 6920 2876
rect 6972 2864 6978 2916
rect 7276 2907 7334 2913
rect 7276 2873 7288 2907
rect 7322 2904 7334 2907
rect 7558 2904 7564 2916
rect 7322 2876 7564 2904
rect 7322 2873 7334 2876
rect 7276 2867 7334 2873
rect 7558 2864 7564 2876
rect 7616 2864 7622 2916
rect 9030 2864 9036 2916
rect 9088 2904 9094 2916
rect 9407 2904 9435 2944
rect 9493 2941 9505 2944
rect 9539 2941 9551 2975
rect 9861 2975 9919 2981
rect 9861 2972 9873 2975
rect 9493 2935 9551 2941
rect 9646 2944 9873 2972
rect 9646 2916 9674 2944
rect 9861 2941 9873 2944
rect 9907 2941 9919 2975
rect 9861 2935 9919 2941
rect 10128 2975 10186 2981
rect 10128 2941 10140 2975
rect 10174 2972 10186 2975
rect 12084 2972 12112 3003
rect 12342 2972 12348 2984
rect 10174 2944 12348 2972
rect 10174 2941 10186 2944
rect 10128 2935 10186 2941
rect 12342 2932 12348 2944
rect 12400 2932 12406 2984
rect 12452 2981 12480 3068
rect 13538 3000 13544 3052
rect 13596 3040 13602 3052
rect 13596 3012 13952 3040
rect 13596 3000 13602 3012
rect 13924 2981 13952 3012
rect 14182 3000 14188 3052
rect 14240 3040 14246 3052
rect 15105 3043 15163 3049
rect 15105 3040 15117 3043
rect 14240 3012 15117 3040
rect 14240 3000 14246 3012
rect 15105 3009 15117 3012
rect 15151 3009 15163 3043
rect 15105 3003 15163 3009
rect 15657 3043 15715 3049
rect 15657 3009 15669 3043
rect 15703 3040 15715 3043
rect 16850 3040 16856 3052
rect 15703 3012 16856 3040
rect 15703 3009 15715 3012
rect 15657 3003 15715 3009
rect 16850 3000 16856 3012
rect 16908 3000 16914 3052
rect 17773 3043 17831 3049
rect 17773 3009 17785 3043
rect 17819 3040 17831 3043
rect 18046 3040 18052 3052
rect 17819 3012 18052 3040
rect 17819 3009 17831 3012
rect 17773 3003 17831 3009
rect 18046 3000 18052 3012
rect 18104 3000 18110 3052
rect 18782 3040 18788 3052
rect 18695 3012 18788 3040
rect 18782 3000 18788 3012
rect 18840 3040 18846 3052
rect 19521 3043 19579 3049
rect 19521 3040 19533 3043
rect 18840 3012 19533 3040
rect 18840 3000 18846 3012
rect 19521 3009 19533 3012
rect 19567 3009 19579 3043
rect 20254 3040 20260 3052
rect 19521 3003 19579 3009
rect 19720 3012 20260 3040
rect 12437 2975 12495 2981
rect 12437 2941 12449 2975
rect 12483 2941 12495 2975
rect 12437 2935 12495 2941
rect 13909 2975 13967 2981
rect 13909 2941 13921 2975
rect 13955 2941 13967 2975
rect 13909 2935 13967 2941
rect 14366 2932 14372 2984
rect 14424 2972 14430 2984
rect 14553 2975 14611 2981
rect 14553 2972 14565 2975
rect 14424 2944 14565 2972
rect 14424 2932 14430 2944
rect 14553 2941 14565 2944
rect 14599 2941 14611 2975
rect 15378 2972 15384 2984
rect 15339 2944 15384 2972
rect 14553 2935 14611 2941
rect 15378 2932 15384 2944
rect 15436 2932 15442 2984
rect 15930 2972 15936 2984
rect 15891 2944 15936 2972
rect 15930 2932 15936 2944
rect 15988 2932 15994 2984
rect 16485 2975 16543 2981
rect 16485 2941 16497 2975
rect 16531 2972 16543 2975
rect 16942 2972 16948 2984
rect 16531 2944 16948 2972
rect 16531 2941 16543 2944
rect 16485 2935 16543 2941
rect 16942 2932 16948 2944
rect 17000 2932 17006 2984
rect 17497 2975 17555 2981
rect 17497 2941 17509 2975
rect 17543 2972 17555 2975
rect 18138 2972 18144 2984
rect 17543 2944 18144 2972
rect 17543 2941 17555 2944
rect 17497 2935 17555 2941
rect 18138 2932 18144 2944
rect 18196 2932 18202 2984
rect 18509 2975 18567 2981
rect 18509 2941 18521 2975
rect 18555 2972 18567 2975
rect 19337 2975 19395 2981
rect 18555 2944 19288 2972
rect 18555 2941 18567 2944
rect 18509 2935 18567 2941
rect 9088 2876 9435 2904
rect 9088 2864 9094 2876
rect 9582 2864 9588 2916
rect 9640 2876 9674 2916
rect 11885 2907 11943 2913
rect 9640 2864 9646 2876
rect 11885 2873 11897 2907
rect 11931 2904 11943 2907
rect 12526 2904 12532 2916
rect 11931 2876 12532 2904
rect 11931 2873 11943 2876
rect 11885 2867 11943 2873
rect 12526 2864 12532 2876
rect 12584 2864 12590 2916
rect 12710 2913 12716 2916
rect 12704 2904 12716 2913
rect 12671 2876 12716 2904
rect 12704 2867 12716 2876
rect 12710 2864 12716 2867
rect 12768 2864 12774 2916
rect 12894 2864 12900 2916
rect 12952 2904 12958 2916
rect 14185 2907 14243 2913
rect 14185 2904 14197 2907
rect 12952 2876 14197 2904
rect 12952 2864 12958 2876
rect 14185 2873 14197 2876
rect 14231 2873 14243 2907
rect 14185 2867 14243 2873
rect 14829 2907 14887 2913
rect 14829 2873 14841 2907
rect 14875 2904 14887 2907
rect 15562 2904 15568 2916
rect 14875 2876 15568 2904
rect 14875 2873 14887 2876
rect 14829 2867 14887 2873
rect 15562 2864 15568 2876
rect 15620 2864 15626 2916
rect 16209 2907 16267 2913
rect 16209 2873 16221 2907
rect 16255 2904 16267 2907
rect 17218 2904 17224 2916
rect 16255 2876 17224 2904
rect 16255 2873 16267 2876
rect 16209 2867 16267 2873
rect 17218 2864 17224 2876
rect 17276 2864 17282 2916
rect 17589 2907 17647 2913
rect 17589 2873 17601 2907
rect 17635 2904 17647 2907
rect 17635 2876 19012 2904
rect 17635 2873 17647 2876
rect 17589 2867 17647 2873
rect 2866 2836 2872 2848
rect 2827 2808 2872 2836
rect 2866 2796 2872 2808
rect 2924 2796 2930 2848
rect 5442 2796 5448 2848
rect 5500 2836 5506 2848
rect 5721 2839 5779 2845
rect 5721 2836 5733 2839
rect 5500 2808 5733 2836
rect 5500 2796 5506 2808
rect 5721 2805 5733 2808
rect 5767 2805 5779 2839
rect 9398 2836 9404 2848
rect 9359 2808 9404 2836
rect 5721 2799 5779 2805
rect 9398 2796 9404 2808
rect 9456 2796 9462 2848
rect 11517 2839 11575 2845
rect 11517 2805 11529 2839
rect 11563 2836 11575 2839
rect 11790 2836 11796 2848
rect 11563 2808 11796 2836
rect 11563 2805 11575 2808
rect 11517 2799 11575 2805
rect 11790 2796 11796 2808
rect 11848 2796 11854 2848
rect 11977 2839 12035 2845
rect 11977 2805 11989 2839
rect 12023 2836 12035 2839
rect 13078 2836 13084 2848
rect 12023 2808 13084 2836
rect 12023 2805 12035 2808
rect 11977 2799 12035 2805
rect 13078 2796 13084 2808
rect 13136 2796 13142 2848
rect 13722 2796 13728 2848
rect 13780 2836 13786 2848
rect 15470 2836 15476 2848
rect 13780 2808 15476 2836
rect 13780 2796 13786 2808
rect 15470 2796 15476 2808
rect 15528 2796 15534 2848
rect 16482 2796 16488 2848
rect 16540 2836 16546 2848
rect 16669 2839 16727 2845
rect 16669 2836 16681 2839
rect 16540 2808 16681 2836
rect 16540 2796 16546 2808
rect 16669 2805 16681 2808
rect 16715 2805 16727 2839
rect 18598 2836 18604 2848
rect 18559 2808 18604 2836
rect 16669 2799 16727 2805
rect 18598 2796 18604 2808
rect 18656 2796 18662 2848
rect 18984 2845 19012 2876
rect 18969 2839 19027 2845
rect 18969 2805 18981 2839
rect 19015 2805 19027 2839
rect 19260 2836 19288 2944
rect 19337 2941 19349 2975
rect 19383 2972 19395 2975
rect 19720 2972 19748 3012
rect 20254 3000 20260 3012
rect 20312 3000 20318 3052
rect 19383 2944 19748 2972
rect 19383 2941 19395 2944
rect 19337 2935 19395 2941
rect 19794 2932 19800 2984
rect 19852 2972 19858 2984
rect 19852 2944 19897 2972
rect 19852 2932 19858 2944
rect 19978 2932 19984 2984
rect 20036 2932 20042 2984
rect 20070 2932 20076 2984
rect 20128 2972 20134 2984
rect 20165 2975 20223 2981
rect 20165 2972 20177 2975
rect 20128 2944 20177 2972
rect 20128 2932 20134 2944
rect 20165 2941 20177 2944
rect 20211 2941 20223 2975
rect 20165 2935 20223 2941
rect 20533 2975 20591 2981
rect 20533 2941 20545 2975
rect 20579 2972 20591 2975
rect 20901 2975 20959 2981
rect 20901 2972 20913 2975
rect 20579 2944 20913 2972
rect 20579 2941 20591 2944
rect 20533 2935 20591 2941
rect 20901 2941 20913 2944
rect 20947 2941 20959 2975
rect 20901 2935 20959 2941
rect 19429 2907 19487 2913
rect 19429 2873 19441 2907
rect 19475 2904 19487 2907
rect 19610 2904 19616 2916
rect 19475 2876 19616 2904
rect 19475 2873 19487 2876
rect 19429 2867 19487 2873
rect 19610 2864 19616 2876
rect 19668 2904 19674 2916
rect 19886 2904 19892 2916
rect 19668 2876 19892 2904
rect 19668 2864 19674 2876
rect 19886 2864 19892 2876
rect 19944 2864 19950 2916
rect 19996 2904 20024 2932
rect 20548 2904 20576 2935
rect 19996 2876 20576 2904
rect 19334 2836 19340 2848
rect 19260 2808 19340 2836
rect 18969 2799 19027 2805
rect 19334 2796 19340 2808
rect 19392 2796 19398 2848
rect 19794 2796 19800 2848
rect 19852 2836 19858 2848
rect 19981 2839 20039 2845
rect 19981 2836 19993 2839
rect 19852 2808 19993 2836
rect 19852 2796 19858 2808
rect 19981 2805 19993 2808
rect 20027 2805 20039 2839
rect 19981 2799 20039 2805
rect 20254 2796 20260 2848
rect 20312 2836 20318 2848
rect 20349 2839 20407 2845
rect 20349 2836 20361 2839
rect 20312 2808 20361 2836
rect 20312 2796 20318 2808
rect 20349 2805 20361 2808
rect 20395 2805 20407 2839
rect 20349 2799 20407 2805
rect 20622 2796 20628 2848
rect 20680 2836 20686 2848
rect 20717 2839 20775 2845
rect 20717 2836 20729 2839
rect 20680 2808 20729 2836
rect 20680 2796 20686 2808
rect 20717 2805 20729 2808
rect 20763 2805 20775 2839
rect 20717 2799 20775 2805
rect 1104 2746 21896 2768
rect 1104 2694 7912 2746
rect 7964 2694 7976 2746
rect 8028 2694 8040 2746
rect 8092 2694 8104 2746
rect 8156 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 15035 2746
rect 15087 2694 21896 2746
rect 1104 2672 21896 2694
rect 2866 2592 2872 2644
rect 2924 2632 2930 2644
rect 3329 2635 3387 2641
rect 3329 2632 3341 2635
rect 2924 2604 3341 2632
rect 2924 2592 2930 2604
rect 3329 2601 3341 2604
rect 3375 2601 3387 2635
rect 4154 2632 4160 2644
rect 4115 2604 4160 2632
rect 3329 2595 3387 2601
rect 4154 2592 4160 2604
rect 4212 2592 4218 2644
rect 4890 2592 4896 2644
rect 4948 2632 4954 2644
rect 4985 2635 5043 2641
rect 4985 2632 4997 2635
rect 4948 2604 4997 2632
rect 4948 2592 4954 2604
rect 4985 2601 4997 2604
rect 5031 2601 5043 2635
rect 4985 2595 5043 2601
rect 5353 2635 5411 2641
rect 5353 2601 5365 2635
rect 5399 2632 5411 2635
rect 5810 2632 5816 2644
rect 5399 2604 5816 2632
rect 5399 2601 5411 2604
rect 5353 2595 5411 2601
rect 5810 2592 5816 2604
rect 5868 2592 5874 2644
rect 5997 2635 6055 2641
rect 5997 2601 6009 2635
rect 6043 2601 6055 2635
rect 5997 2595 6055 2601
rect 5074 2564 5080 2576
rect 4540 2536 5080 2564
rect 3602 2456 3608 2508
rect 3660 2496 3666 2508
rect 4540 2505 4568 2536
rect 5074 2524 5080 2536
rect 5132 2524 5138 2576
rect 5534 2524 5540 2576
rect 5592 2564 5598 2576
rect 6012 2564 6040 2595
rect 6362 2592 6368 2644
rect 6420 2632 6426 2644
rect 7377 2635 7435 2641
rect 7377 2632 7389 2635
rect 6420 2604 7389 2632
rect 6420 2592 6426 2604
rect 7377 2601 7389 2604
rect 7423 2601 7435 2635
rect 7377 2595 7435 2601
rect 9309 2635 9367 2641
rect 9309 2601 9321 2635
rect 9355 2632 9367 2635
rect 9398 2632 9404 2644
rect 9355 2604 9404 2632
rect 9355 2601 9367 2604
rect 9309 2595 9367 2601
rect 9398 2592 9404 2604
rect 9456 2592 9462 2644
rect 9766 2632 9772 2644
rect 9727 2604 9772 2632
rect 9766 2592 9772 2604
rect 9824 2592 9830 2644
rect 10134 2592 10140 2644
rect 10192 2632 10198 2644
rect 10192 2604 10640 2632
rect 10192 2592 10198 2604
rect 5592 2536 6040 2564
rect 6457 2567 6515 2573
rect 5592 2524 5598 2536
rect 6457 2533 6469 2567
rect 6503 2564 6515 2567
rect 6914 2564 6920 2576
rect 6503 2536 6920 2564
rect 6503 2533 6515 2536
rect 6457 2527 6515 2533
rect 6914 2524 6920 2536
rect 6972 2524 6978 2576
rect 7558 2524 7564 2576
rect 7616 2564 7622 2576
rect 8573 2567 8631 2573
rect 7616 2536 8064 2564
rect 7616 2524 7622 2536
rect 4525 2499 4583 2505
rect 4525 2496 4537 2499
rect 3660 2468 4537 2496
rect 3660 2456 3666 2468
rect 4525 2465 4537 2468
rect 4571 2465 4583 2499
rect 4525 2459 4583 2465
rect 4982 2456 4988 2508
rect 5040 2496 5046 2508
rect 5445 2499 5503 2505
rect 5445 2496 5457 2499
rect 5040 2468 5457 2496
rect 5040 2456 5046 2468
rect 5445 2465 5457 2468
rect 5491 2465 5503 2499
rect 5445 2459 5503 2465
rect 5905 2499 5963 2505
rect 5905 2465 5917 2499
rect 5951 2496 5963 2499
rect 6362 2496 6368 2508
rect 5951 2468 6368 2496
rect 5951 2465 5963 2468
rect 5905 2459 5963 2465
rect 6362 2456 6368 2468
rect 6420 2456 6426 2508
rect 7009 2499 7067 2505
rect 7009 2465 7021 2499
rect 7055 2496 7067 2499
rect 7742 2496 7748 2508
rect 7055 2468 7748 2496
rect 7055 2465 7067 2468
rect 7009 2459 7067 2465
rect 7742 2456 7748 2468
rect 7800 2456 7806 2508
rect 8036 2496 8064 2536
rect 8573 2533 8585 2567
rect 8619 2564 8631 2567
rect 9674 2564 9680 2576
rect 8619 2536 9680 2564
rect 8619 2533 8631 2536
rect 8573 2527 8631 2533
rect 9674 2524 9680 2536
rect 9732 2524 9738 2576
rect 9950 2524 9956 2576
rect 10008 2564 10014 2576
rect 10229 2567 10287 2573
rect 10229 2564 10241 2567
rect 10008 2536 10241 2564
rect 10008 2524 10014 2536
rect 10229 2533 10241 2536
rect 10275 2533 10287 2567
rect 10229 2527 10287 2533
rect 9766 2496 9772 2508
rect 8036 2468 9772 2496
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 4617 2431 4675 2437
rect 4617 2428 4629 2431
rect 3292 2400 4629 2428
rect 3292 2388 3298 2400
rect 3694 2360 3700 2372
rect 3160 2332 3700 2360
rect 3160 2304 3188 2332
rect 3694 2320 3700 2332
rect 3752 2320 3758 2372
rect 3804 2304 3832 2400
rect 4617 2397 4629 2400
rect 4663 2397 4675 2431
rect 4617 2391 4675 2397
rect 4706 2388 4712 2440
rect 4764 2428 4770 2440
rect 4801 2431 4859 2437
rect 4801 2428 4813 2431
rect 4764 2400 4813 2428
rect 4764 2388 4770 2400
rect 4801 2397 4813 2400
rect 4847 2428 4859 2431
rect 4890 2428 4896 2440
rect 4847 2400 4896 2428
rect 4847 2397 4859 2400
rect 4801 2391 4859 2397
rect 4890 2388 4896 2400
rect 4948 2388 4954 2440
rect 5537 2431 5595 2437
rect 5537 2428 5549 2431
rect 5460 2400 5549 2428
rect 5460 2372 5488 2400
rect 5537 2397 5549 2400
rect 5583 2397 5595 2431
rect 5537 2391 5595 2397
rect 6549 2431 6607 2437
rect 6549 2397 6561 2431
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 4246 2320 4252 2372
rect 4304 2360 4310 2372
rect 5442 2360 5448 2372
rect 4304 2332 5448 2360
rect 4304 2320 4310 2332
rect 5442 2320 5448 2332
rect 5500 2320 5506 2372
rect 6564 2360 6592 2391
rect 7190 2388 7196 2440
rect 7248 2428 7254 2440
rect 8036 2437 8064 2468
rect 7837 2431 7895 2437
rect 7837 2428 7849 2431
rect 7248 2400 7849 2428
rect 7248 2388 7254 2400
rect 7837 2397 7849 2400
rect 7883 2397 7895 2431
rect 7837 2391 7895 2397
rect 8021 2431 8079 2437
rect 8021 2397 8033 2431
rect 8067 2397 8079 2431
rect 8662 2428 8668 2440
rect 8623 2400 8668 2428
rect 8021 2391 8079 2397
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 8864 2437 8892 2468
rect 9766 2456 9772 2468
rect 9824 2456 9830 2508
rect 10134 2496 10140 2508
rect 10095 2468 10140 2496
rect 10134 2456 10140 2468
rect 10192 2456 10198 2508
rect 10612 2505 10640 2604
rect 11146 2592 11152 2644
rect 11204 2632 11210 2644
rect 11425 2635 11483 2641
rect 11425 2632 11437 2635
rect 11204 2604 11437 2632
rect 11204 2592 11210 2604
rect 11425 2601 11437 2604
rect 11471 2601 11483 2635
rect 11425 2595 11483 2601
rect 12526 2592 12532 2644
rect 12584 2632 12590 2644
rect 12621 2635 12679 2641
rect 12621 2632 12633 2635
rect 12584 2604 12633 2632
rect 12584 2592 12590 2604
rect 12621 2601 12633 2604
rect 12667 2601 12679 2635
rect 12621 2595 12679 2601
rect 12986 2592 12992 2644
rect 13044 2632 13050 2644
rect 13081 2635 13139 2641
rect 13081 2632 13093 2635
rect 13044 2604 13093 2632
rect 13044 2592 13050 2604
rect 13081 2601 13093 2604
rect 13127 2601 13139 2635
rect 13081 2595 13139 2601
rect 16206 2592 16212 2644
rect 16264 2632 16270 2644
rect 16301 2635 16359 2641
rect 16301 2632 16313 2635
rect 16264 2604 16313 2632
rect 16264 2592 16270 2604
rect 16301 2601 16313 2604
rect 16347 2601 16359 2635
rect 16301 2595 16359 2601
rect 17037 2635 17095 2641
rect 17037 2601 17049 2635
rect 17083 2632 17095 2635
rect 17678 2632 17684 2644
rect 17083 2604 17684 2632
rect 17083 2601 17095 2604
rect 17037 2595 17095 2601
rect 12253 2567 12311 2573
rect 11624 2536 12112 2564
rect 11624 2505 11652 2536
rect 10597 2499 10655 2505
rect 10597 2465 10609 2499
rect 10643 2465 10655 2499
rect 10597 2459 10655 2465
rect 11609 2499 11667 2505
rect 11609 2465 11621 2499
rect 11655 2465 11667 2499
rect 11609 2459 11667 2465
rect 11790 2456 11796 2508
rect 11848 2496 11854 2508
rect 11977 2499 12035 2505
rect 11977 2496 11989 2499
rect 11848 2468 11989 2496
rect 11848 2456 11854 2468
rect 11977 2465 11989 2468
rect 12023 2465 12035 2499
rect 12084 2496 12112 2536
rect 12253 2533 12265 2567
rect 12299 2564 12311 2567
rect 12299 2536 13492 2564
rect 12299 2533 12311 2536
rect 12253 2527 12311 2533
rect 12894 2496 12900 2508
rect 12084 2468 12900 2496
rect 11977 2459 12035 2465
rect 12894 2456 12900 2468
rect 12952 2456 12958 2508
rect 13464 2505 13492 2536
rect 15028 2536 16252 2564
rect 12989 2499 13047 2505
rect 12989 2465 13001 2499
rect 13035 2496 13047 2499
rect 13449 2499 13507 2505
rect 13035 2468 13400 2496
rect 13035 2465 13047 2468
rect 12989 2459 13047 2465
rect 8849 2431 8907 2437
rect 8849 2397 8861 2431
rect 8895 2397 8907 2431
rect 10410 2428 10416 2440
rect 10371 2400 10416 2428
rect 8849 2391 8907 2397
rect 10410 2388 10416 2400
rect 10468 2388 10474 2440
rect 10873 2431 10931 2437
rect 10873 2397 10885 2431
rect 10919 2428 10931 2431
rect 12618 2428 12624 2440
rect 10919 2400 12624 2428
rect 10919 2397 10931 2400
rect 10873 2391 10931 2397
rect 12618 2388 12624 2400
rect 12676 2388 12682 2440
rect 12710 2388 12716 2440
rect 12768 2428 12774 2440
rect 13173 2431 13231 2437
rect 13173 2428 13185 2431
rect 12768 2400 13185 2428
rect 12768 2388 12774 2400
rect 13173 2397 13185 2400
rect 13219 2397 13231 2431
rect 13372 2428 13400 2468
rect 13449 2465 13461 2499
rect 13495 2465 13507 2499
rect 13814 2496 13820 2508
rect 13775 2468 13820 2496
rect 13449 2459 13507 2465
rect 13814 2456 13820 2468
rect 13872 2456 13878 2508
rect 14182 2496 14188 2508
rect 14143 2468 14188 2496
rect 14182 2456 14188 2468
rect 14240 2456 14246 2508
rect 14550 2496 14556 2508
rect 14511 2468 14556 2496
rect 14550 2456 14556 2468
rect 14608 2456 14614 2508
rect 14642 2456 14648 2508
rect 14700 2496 14706 2508
rect 15028 2505 15056 2536
rect 15013 2499 15071 2505
rect 15013 2496 15025 2499
rect 14700 2468 15025 2496
rect 14700 2456 14706 2468
rect 15013 2465 15025 2468
rect 15059 2465 15071 2499
rect 15013 2459 15071 2465
rect 15473 2499 15531 2505
rect 15473 2465 15485 2499
rect 15519 2465 15531 2499
rect 15473 2459 15531 2465
rect 13906 2428 13912 2440
rect 13372 2400 13912 2428
rect 13173 2391 13231 2397
rect 13906 2388 13912 2400
rect 13964 2388 13970 2440
rect 15488 2428 15516 2459
rect 15562 2456 15568 2508
rect 15620 2496 15626 2508
rect 16224 2505 16252 2536
rect 15841 2499 15899 2505
rect 15841 2496 15853 2499
rect 15620 2468 15853 2496
rect 15620 2456 15626 2468
rect 15841 2465 15853 2468
rect 15887 2465 15899 2499
rect 15841 2459 15899 2465
rect 16209 2499 16267 2505
rect 16209 2465 16221 2499
rect 16255 2465 16267 2499
rect 16316 2496 16344 2595
rect 17678 2592 17684 2604
rect 17736 2592 17742 2644
rect 19518 2592 19524 2644
rect 19576 2632 19582 2644
rect 19613 2635 19671 2641
rect 19613 2632 19625 2635
rect 19576 2604 19625 2632
rect 19576 2592 19582 2604
rect 19613 2601 19625 2604
rect 19659 2601 19671 2635
rect 20070 2632 20076 2644
rect 20031 2604 20076 2632
rect 19613 2595 19671 2601
rect 20070 2592 20076 2604
rect 20128 2592 20134 2644
rect 16390 2524 16396 2576
rect 16448 2564 16454 2576
rect 19245 2567 19303 2573
rect 19245 2564 19257 2567
rect 16448 2536 19257 2564
rect 16448 2524 16454 2536
rect 19245 2533 19257 2536
rect 19291 2533 19303 2567
rect 19245 2527 19303 2533
rect 16485 2499 16543 2505
rect 16485 2496 16497 2499
rect 16316 2468 16497 2496
rect 16209 2459 16267 2465
rect 16485 2465 16497 2468
rect 16531 2465 16543 2499
rect 16850 2496 16856 2508
rect 16811 2468 16856 2496
rect 16485 2459 16543 2465
rect 16850 2456 16856 2468
rect 16908 2456 16914 2508
rect 17218 2496 17224 2508
rect 17179 2468 17224 2496
rect 17218 2456 17224 2468
rect 17276 2456 17282 2508
rect 18325 2499 18383 2505
rect 18325 2496 18337 2499
rect 17972 2468 18337 2496
rect 15654 2428 15660 2440
rect 15488 2400 15660 2428
rect 15654 2388 15660 2400
rect 15712 2428 15718 2440
rect 16390 2428 16396 2440
rect 15712 2400 16396 2428
rect 15712 2388 15718 2400
rect 16390 2388 16396 2400
rect 16448 2388 16454 2440
rect 17972 2437 18000 2468
rect 18325 2465 18337 2468
rect 18371 2496 18383 2499
rect 18598 2496 18604 2508
rect 18371 2468 18604 2496
rect 18371 2465 18383 2468
rect 18325 2459 18383 2465
rect 18598 2456 18604 2468
rect 18656 2456 18662 2508
rect 18690 2456 18696 2508
rect 18748 2496 18754 2508
rect 19061 2499 19119 2505
rect 19061 2496 19073 2499
rect 18748 2468 19073 2496
rect 18748 2456 18754 2468
rect 19061 2465 19073 2468
rect 19107 2465 19119 2499
rect 19061 2459 19119 2465
rect 17773 2431 17831 2437
rect 17773 2428 17785 2431
rect 16592 2400 17785 2428
rect 5552 2332 6592 2360
rect 3142 2292 3148 2304
rect 3103 2264 3148 2292
rect 3142 2252 3148 2264
rect 3200 2252 3206 2304
rect 3602 2292 3608 2304
rect 3563 2264 3608 2292
rect 3602 2252 3608 2264
rect 3660 2252 3666 2304
rect 3786 2292 3792 2304
rect 3747 2264 3792 2292
rect 3786 2252 3792 2264
rect 3844 2252 3850 2304
rect 4890 2252 4896 2304
rect 4948 2292 4954 2304
rect 5350 2292 5356 2304
rect 4948 2264 5356 2292
rect 4948 2252 4954 2264
rect 5350 2252 5356 2264
rect 5408 2292 5414 2304
rect 5552 2292 5580 2332
rect 6730 2320 6736 2372
rect 6788 2360 6794 2372
rect 8205 2363 8263 2369
rect 8205 2360 8217 2363
rect 6788 2332 8217 2360
rect 6788 2320 6794 2332
rect 8205 2329 8217 2332
rect 8251 2329 8263 2363
rect 8205 2323 8263 2329
rect 9766 2320 9772 2372
rect 9824 2360 9830 2372
rect 10428 2360 10456 2388
rect 9824 2332 10456 2360
rect 9824 2320 9830 2332
rect 13538 2320 13544 2372
rect 13596 2360 13602 2372
rect 14001 2363 14059 2369
rect 14001 2360 14013 2363
rect 13596 2332 14013 2360
rect 13596 2320 13602 2332
rect 14001 2329 14013 2332
rect 14047 2329 14059 2363
rect 14001 2323 14059 2329
rect 15470 2320 15476 2372
rect 15528 2360 15534 2372
rect 16592 2360 16620 2400
rect 17773 2397 17785 2400
rect 17819 2428 17831 2431
rect 17957 2431 18015 2437
rect 17957 2428 17969 2431
rect 17819 2400 17969 2428
rect 17819 2397 17831 2400
rect 17773 2391 17831 2397
rect 17957 2397 17969 2400
rect 18003 2397 18015 2431
rect 17957 2391 18015 2397
rect 15528 2332 16620 2360
rect 16669 2363 16727 2369
rect 15528 2320 15534 2332
rect 16669 2329 16681 2363
rect 16715 2360 16727 2363
rect 17310 2360 17316 2372
rect 16715 2332 17316 2360
rect 16715 2329 16727 2332
rect 16669 2323 16727 2329
rect 17310 2320 17316 2332
rect 17368 2320 17374 2372
rect 17405 2363 17463 2369
rect 17405 2329 17417 2363
rect 17451 2360 17463 2363
rect 19334 2360 19340 2372
rect 17451 2332 19340 2360
rect 17451 2329 17463 2332
rect 17405 2323 17463 2329
rect 19334 2320 19340 2332
rect 19392 2320 19398 2372
rect 7190 2292 7196 2304
rect 5408 2264 5580 2292
rect 7151 2264 7196 2292
rect 5408 2252 5414 2264
rect 7190 2252 7196 2264
rect 7248 2252 7254 2304
rect 9030 2292 9036 2304
rect 8991 2264 9036 2292
rect 9030 2252 9036 2264
rect 9088 2252 9094 2304
rect 9585 2295 9643 2301
rect 9585 2261 9597 2295
rect 9631 2292 9643 2295
rect 9950 2292 9956 2304
rect 9631 2264 9956 2292
rect 9631 2261 9643 2264
rect 9585 2255 9643 2261
rect 9950 2252 9956 2264
rect 10008 2252 10014 2304
rect 10134 2252 10140 2304
rect 10192 2292 10198 2304
rect 10778 2292 10784 2304
rect 10192 2264 10784 2292
rect 10192 2252 10198 2264
rect 10778 2252 10784 2264
rect 10836 2292 10842 2304
rect 11149 2295 11207 2301
rect 11149 2292 11161 2295
rect 10836 2264 11161 2292
rect 10836 2252 10842 2264
rect 11149 2261 11161 2264
rect 11195 2261 11207 2295
rect 11149 2255 11207 2261
rect 11793 2295 11851 2301
rect 11793 2261 11805 2295
rect 11839 2292 11851 2295
rect 12710 2292 12716 2304
rect 11839 2264 12716 2292
rect 11839 2261 11851 2264
rect 11793 2255 11851 2261
rect 12710 2252 12716 2264
rect 12768 2252 12774 2304
rect 13078 2252 13084 2304
rect 13136 2292 13142 2304
rect 13633 2295 13691 2301
rect 13633 2292 13645 2295
rect 13136 2264 13645 2292
rect 13136 2252 13142 2264
rect 13633 2261 13645 2264
rect 13679 2261 13691 2295
rect 13633 2255 13691 2261
rect 14090 2252 14096 2304
rect 14148 2292 14154 2304
rect 14369 2295 14427 2301
rect 14369 2292 14381 2295
rect 14148 2264 14381 2292
rect 14148 2252 14154 2264
rect 14369 2261 14381 2264
rect 14415 2261 14427 2295
rect 14369 2255 14427 2261
rect 14458 2252 14464 2304
rect 14516 2292 14522 2304
rect 14737 2295 14795 2301
rect 14737 2292 14749 2295
rect 14516 2264 14749 2292
rect 14516 2252 14522 2264
rect 14737 2261 14749 2264
rect 14783 2261 14795 2295
rect 15194 2292 15200 2304
rect 15155 2264 15200 2292
rect 14737 2255 14795 2261
rect 15194 2252 15200 2264
rect 15252 2252 15258 2304
rect 15654 2292 15660 2304
rect 15615 2264 15660 2292
rect 15654 2252 15660 2264
rect 15712 2252 15718 2304
rect 16022 2292 16028 2304
rect 15983 2264 16028 2292
rect 16022 2252 16028 2264
rect 16080 2252 16086 2304
rect 16209 2295 16267 2301
rect 16209 2261 16221 2295
rect 16255 2292 16267 2295
rect 17586 2292 17592 2304
rect 16255 2264 17592 2292
rect 16255 2261 16267 2264
rect 16209 2255 16267 2261
rect 17586 2252 17592 2264
rect 17644 2252 17650 2304
rect 18509 2295 18567 2301
rect 18509 2261 18521 2295
rect 18555 2292 18567 2295
rect 18598 2292 18604 2304
rect 18555 2264 18604 2292
rect 18555 2261 18567 2264
rect 18509 2255 18567 2261
rect 18598 2252 18604 2264
rect 18656 2252 18662 2304
rect 18877 2295 18935 2301
rect 18877 2261 18889 2295
rect 18923 2292 18935 2295
rect 18966 2292 18972 2304
rect 18923 2264 18972 2292
rect 18923 2261 18935 2264
rect 18877 2255 18935 2261
rect 18966 2252 18972 2264
rect 19024 2252 19030 2304
rect 19518 2292 19524 2304
rect 19479 2264 19524 2292
rect 19518 2252 19524 2264
rect 19576 2252 19582 2304
rect 19886 2292 19892 2304
rect 19847 2264 19892 2292
rect 19886 2252 19892 2264
rect 19944 2252 19950 2304
rect 1104 2202 21896 2224
rect 1104 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 4575 2202
rect 4627 2150 4639 2202
rect 4691 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 18308 2202
rect 18360 2150 18372 2202
rect 18424 2150 18436 2202
rect 18488 2150 18500 2202
rect 18552 2150 21896 2202
rect 1104 2128 21896 2150
rect 1026 2048 1032 2100
rect 1084 2088 1090 2100
rect 6181 2091 6239 2097
rect 6181 2088 6193 2091
rect 1084 2060 6193 2088
rect 1084 2048 1090 2060
rect 6181 2057 6193 2060
rect 6227 2057 6239 2091
rect 6181 2051 6239 2057
rect 6914 2048 6920 2100
rect 6972 2088 6978 2100
rect 9214 2088 9220 2100
rect 6972 2060 9220 2088
rect 6972 2048 6978 2060
rect 9214 2048 9220 2060
rect 9272 2088 9278 2100
rect 9398 2088 9404 2100
rect 9272 2060 9404 2088
rect 9272 2048 9278 2060
rect 9398 2048 9404 2060
rect 9456 2048 9462 2100
rect 6362 1980 6368 2032
rect 6420 2020 6426 2032
rect 12250 2020 12256 2032
rect 6420 1992 12256 2020
rect 6420 1980 6426 1992
rect 12250 1980 12256 1992
rect 12308 1980 12314 2032
rect 12618 1980 12624 2032
rect 12676 2020 12682 2032
rect 14550 2020 14556 2032
rect 12676 1992 14556 2020
rect 12676 1980 12682 1992
rect 14550 1980 14556 1992
rect 14608 1980 14614 2032
rect 2682 1912 2688 1964
rect 2740 1952 2746 1964
rect 8662 1952 8668 1964
rect 2740 1924 8668 1952
rect 2740 1912 2746 1924
rect 8662 1912 8668 1924
rect 8720 1912 8726 1964
rect 1854 1844 1860 1896
rect 1912 1884 1918 1896
rect 7190 1884 7196 1896
rect 1912 1856 7196 1884
rect 1912 1844 1918 1856
rect 7190 1844 7196 1856
rect 7248 1844 7254 1896
rect 6181 1819 6239 1825
rect 6181 1785 6193 1819
rect 6227 1816 6239 1819
rect 9950 1816 9956 1828
rect 6227 1788 9956 1816
rect 6227 1785 6239 1788
rect 6181 1779 6239 1785
rect 9950 1776 9956 1788
rect 10008 1776 10014 1828
rect 566 1708 572 1760
rect 624 1748 630 1760
rect 9306 1748 9312 1760
rect 624 1720 9312 1748
rect 624 1708 630 1720
rect 9306 1708 9312 1720
rect 9364 1708 9370 1760
rect 198 1640 204 1692
rect 256 1680 262 1692
rect 9030 1680 9036 1692
rect 256 1652 9036 1680
rect 256 1640 262 1652
rect 9030 1640 9036 1652
rect 9088 1640 9094 1692
rect 3050 1572 3056 1624
rect 3108 1612 3114 1624
rect 7466 1612 7472 1624
rect 3108 1584 7472 1612
rect 3108 1572 3114 1584
rect 7466 1572 7472 1584
rect 7524 1572 7530 1624
rect 1394 1436 1400 1488
rect 1452 1476 1458 1488
rect 10134 1476 10140 1488
rect 1452 1448 10140 1476
rect 1452 1436 1458 1448
rect 10134 1436 10140 1448
rect 10192 1436 10198 1488
<< via1 >>
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 4575 20646 4627 20698
rect 4639 20646 4691 20698
rect 11378 20646 11430 20698
rect 11442 20646 11494 20698
rect 11506 20646 11558 20698
rect 11570 20646 11622 20698
rect 18308 20646 18360 20698
rect 18372 20646 18424 20698
rect 18436 20646 18488 20698
rect 18500 20646 18552 20698
rect 11704 20544 11756 20596
rect 18972 20587 19024 20596
rect 18972 20553 18981 20587
rect 18981 20553 19015 20587
rect 19015 20553 19024 20587
rect 18972 20544 19024 20553
rect 19340 20544 19392 20596
rect 20904 20544 20956 20596
rect 4344 20476 4396 20528
rect 5356 20476 5408 20528
rect 9864 20476 9916 20528
rect 20628 20476 20680 20528
rect 6644 20408 6696 20460
rect 22376 20408 22428 20460
rect 4344 20340 4396 20392
rect 5448 20272 5500 20324
rect 7840 20272 7892 20324
rect 13452 20272 13504 20324
rect 7288 20247 7340 20256
rect 7288 20213 7297 20247
rect 7297 20213 7331 20247
rect 7331 20213 7340 20247
rect 7288 20204 7340 20213
rect 19616 20204 19668 20256
rect 20720 20340 20772 20392
rect 20904 20340 20956 20392
rect 22744 20272 22796 20324
rect 21272 20204 21324 20256
rect 7912 20102 7964 20154
rect 7976 20102 8028 20154
rect 8040 20102 8092 20154
rect 8104 20102 8156 20154
rect 14843 20102 14895 20154
rect 14907 20102 14959 20154
rect 14971 20102 15023 20154
rect 15035 20102 15087 20154
rect 2872 20000 2924 20052
rect 3332 20000 3384 20052
rect 7380 20000 7432 20052
rect 7564 20000 7616 20052
rect 9036 20000 9088 20052
rect 10876 20000 10928 20052
rect 11244 20000 11296 20052
rect 12072 20000 12124 20052
rect 14004 20000 14056 20052
rect 15384 20000 15436 20052
rect 15844 20000 15896 20052
rect 18144 20000 18196 20052
rect 4068 19932 4120 19984
rect 19248 19932 19300 19984
rect 19432 19932 19484 19984
rect 19984 19975 20036 19984
rect 5540 19864 5592 19916
rect 6828 19864 6880 19916
rect 7380 19864 7432 19916
rect 4068 19839 4120 19848
rect 4068 19805 4077 19839
rect 4077 19805 4111 19839
rect 4111 19805 4120 19839
rect 4068 19796 4120 19805
rect 5264 19796 5316 19848
rect 8300 19839 8352 19848
rect 7564 19771 7616 19780
rect 7564 19737 7573 19771
rect 7573 19737 7607 19771
rect 7607 19737 7616 19771
rect 8300 19805 8309 19839
rect 8309 19805 8343 19839
rect 8343 19805 8352 19839
rect 8300 19796 8352 19805
rect 7564 19728 7616 19737
rect 8852 19728 8904 19780
rect 4988 19660 5040 19712
rect 7196 19703 7248 19712
rect 7196 19669 7205 19703
rect 7205 19669 7239 19703
rect 7239 19669 7248 19703
rect 7196 19660 7248 19669
rect 7656 19703 7708 19712
rect 7656 19669 7665 19703
rect 7665 19669 7699 19703
rect 7699 19669 7708 19703
rect 7656 19660 7708 19669
rect 8760 19703 8812 19712
rect 8760 19669 8769 19703
rect 8769 19669 8803 19703
rect 8803 19669 8812 19703
rect 8760 19660 8812 19669
rect 9680 19864 9732 19916
rect 9956 19864 10008 19916
rect 10876 19907 10928 19916
rect 10876 19873 10885 19907
rect 10885 19873 10919 19907
rect 10919 19873 10928 19907
rect 10876 19864 10928 19873
rect 12164 19907 12216 19916
rect 12164 19873 12173 19907
rect 12173 19873 12207 19907
rect 12207 19873 12216 19907
rect 12164 19864 12216 19873
rect 13084 19907 13136 19916
rect 13084 19873 13093 19907
rect 13093 19873 13127 19907
rect 13127 19873 13136 19907
rect 13084 19864 13136 19873
rect 14556 19907 14608 19916
rect 14556 19873 14565 19907
rect 14565 19873 14599 19907
rect 14599 19873 14608 19907
rect 14556 19864 14608 19873
rect 15200 19864 15252 19916
rect 16120 19864 16172 19916
rect 18972 19864 19024 19916
rect 19616 19864 19668 19916
rect 19984 19941 19993 19975
rect 19993 19941 20027 19975
rect 20027 19941 20036 19975
rect 19984 19932 20036 19941
rect 20536 19975 20588 19984
rect 20536 19941 20545 19975
rect 20545 19941 20579 19975
rect 20579 19941 20588 19975
rect 20536 19932 20588 19941
rect 20628 19932 20680 19984
rect 21640 19932 21692 19984
rect 19340 19796 19392 19848
rect 20628 19796 20680 19848
rect 12440 19728 12492 19780
rect 12256 19660 12308 19712
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 4575 19558 4627 19610
rect 4639 19558 4691 19610
rect 11378 19558 11430 19610
rect 11442 19558 11494 19610
rect 11506 19558 11558 19610
rect 11570 19558 11622 19610
rect 18308 19558 18360 19610
rect 18372 19558 18424 19610
rect 18436 19558 18488 19610
rect 18500 19558 18552 19610
rect 1952 19499 2004 19508
rect 1952 19465 1961 19499
rect 1961 19465 1995 19499
rect 1995 19465 2004 19499
rect 1952 19456 2004 19465
rect 4160 19456 4212 19508
rect 5264 19456 5316 19508
rect 5540 19456 5592 19508
rect 6644 19499 6696 19508
rect 6644 19465 6653 19499
rect 6653 19465 6687 19499
rect 6687 19465 6696 19499
rect 6644 19456 6696 19465
rect 204 19184 256 19236
rect 2136 19184 2188 19236
rect 3056 19116 3108 19168
rect 4344 19252 4396 19304
rect 5908 19252 5960 19304
rect 9128 19456 9180 19508
rect 15108 19499 15160 19508
rect 15108 19465 15117 19499
rect 15117 19465 15151 19499
rect 15151 19465 15160 19499
rect 15108 19456 15160 19465
rect 10140 19388 10192 19440
rect 10600 19388 10652 19440
rect 6920 19295 6972 19304
rect 6920 19261 6929 19295
rect 6929 19261 6963 19295
rect 6963 19261 6972 19295
rect 6920 19252 6972 19261
rect 8300 19252 8352 19304
rect 8760 19295 8812 19304
rect 8760 19261 8769 19295
rect 8769 19261 8803 19295
rect 8803 19261 8812 19295
rect 8760 19252 8812 19261
rect 4988 19184 5040 19236
rect 7012 19184 7064 19236
rect 7380 19184 7432 19236
rect 10876 19320 10928 19372
rect 10968 19363 11020 19372
rect 10968 19329 10977 19363
rect 10977 19329 11011 19363
rect 11011 19329 11020 19363
rect 10968 19320 11020 19329
rect 9680 19252 9732 19304
rect 9864 19252 9916 19304
rect 11980 19320 12032 19372
rect 13084 19320 13136 19372
rect 11704 19252 11756 19304
rect 12072 19252 12124 19304
rect 12992 19295 13044 19304
rect 11152 19184 11204 19236
rect 12992 19261 13001 19295
rect 13001 19261 13035 19295
rect 13035 19261 13044 19295
rect 12992 19252 13044 19261
rect 13360 19295 13412 19304
rect 13360 19261 13369 19295
rect 13369 19261 13403 19295
rect 13403 19261 13412 19295
rect 13360 19252 13412 19261
rect 13728 19295 13780 19304
rect 13728 19261 13737 19295
rect 13737 19261 13771 19295
rect 13771 19261 13780 19295
rect 13728 19252 13780 19261
rect 14188 19295 14240 19304
rect 14188 19261 14197 19295
rect 14197 19261 14231 19295
rect 14231 19261 14240 19295
rect 14188 19252 14240 19261
rect 14464 19252 14516 19304
rect 15568 19295 15620 19304
rect 4896 19116 4948 19168
rect 5080 19116 5132 19168
rect 5264 19116 5316 19168
rect 6736 19116 6788 19168
rect 6828 19116 6880 19168
rect 8392 19159 8444 19168
rect 8392 19125 8401 19159
rect 8401 19125 8435 19159
rect 8435 19125 8444 19159
rect 8852 19159 8904 19168
rect 8392 19116 8444 19125
rect 8852 19125 8861 19159
rect 8861 19125 8895 19159
rect 8895 19125 8904 19159
rect 8852 19116 8904 19125
rect 10140 19116 10192 19168
rect 10876 19159 10928 19168
rect 10876 19125 10885 19159
rect 10885 19125 10919 19159
rect 10919 19125 10928 19159
rect 15568 19261 15577 19295
rect 15577 19261 15611 19295
rect 15611 19261 15620 19295
rect 15568 19252 15620 19261
rect 16028 19252 16080 19304
rect 17132 19295 17184 19304
rect 15844 19227 15896 19236
rect 15844 19193 15853 19227
rect 15853 19193 15887 19227
rect 15887 19193 15896 19227
rect 15844 19184 15896 19193
rect 17132 19261 17141 19295
rect 17141 19261 17175 19295
rect 17175 19261 17184 19295
rect 17132 19252 17184 19261
rect 17592 19295 17644 19304
rect 17592 19261 17601 19295
rect 17601 19261 17635 19295
rect 17635 19261 17644 19295
rect 18972 19320 19024 19372
rect 21272 19363 21324 19372
rect 17592 19252 17644 19261
rect 18512 19295 18564 19304
rect 18512 19261 18521 19295
rect 18521 19261 18555 19295
rect 18555 19261 18564 19295
rect 18512 19252 18564 19261
rect 20168 19295 20220 19304
rect 10876 19116 10928 19125
rect 11336 19116 11388 19168
rect 12808 19116 12860 19168
rect 13268 19116 13320 19168
rect 13636 19116 13688 19168
rect 14372 19159 14424 19168
rect 14372 19125 14381 19159
rect 14381 19125 14415 19159
rect 14415 19125 14424 19159
rect 14372 19116 14424 19125
rect 14740 19159 14792 19168
rect 14740 19125 14749 19159
rect 14749 19125 14783 19159
rect 14783 19125 14792 19159
rect 14740 19116 14792 19125
rect 15292 19159 15344 19168
rect 15292 19125 15301 19159
rect 15301 19125 15335 19159
rect 15335 19125 15344 19159
rect 15292 19116 15344 19125
rect 16304 19159 16356 19168
rect 16304 19125 16313 19159
rect 16313 19125 16347 19159
rect 16347 19125 16356 19159
rect 16304 19116 16356 19125
rect 16672 19159 16724 19168
rect 16672 19125 16681 19159
rect 16681 19125 16715 19159
rect 16715 19125 16724 19159
rect 16672 19116 16724 19125
rect 16948 19159 17000 19168
rect 16948 19125 16957 19159
rect 16957 19125 16991 19159
rect 16991 19125 17000 19159
rect 16948 19116 17000 19125
rect 17408 19116 17460 19168
rect 17776 19159 17828 19168
rect 17776 19125 17785 19159
rect 17785 19125 17819 19159
rect 17819 19125 17828 19159
rect 17776 19116 17828 19125
rect 20168 19261 20177 19295
rect 20177 19261 20211 19295
rect 20211 19261 20220 19295
rect 20168 19252 20220 19261
rect 20444 19295 20496 19304
rect 20444 19261 20453 19295
rect 20453 19261 20487 19295
rect 20487 19261 20496 19295
rect 20444 19252 20496 19261
rect 20628 19252 20680 19304
rect 21272 19329 21281 19363
rect 21281 19329 21315 19363
rect 21315 19329 21324 19363
rect 21272 19320 21324 19329
rect 20996 19295 21048 19304
rect 20996 19261 21005 19295
rect 21005 19261 21039 19295
rect 21039 19261 21048 19295
rect 20996 19252 21048 19261
rect 18972 19184 19024 19236
rect 19524 19184 19576 19236
rect 19616 19184 19668 19236
rect 20076 19116 20128 19168
rect 7912 19014 7964 19066
rect 7976 19014 8028 19066
rect 8040 19014 8092 19066
rect 8104 19014 8156 19066
rect 14843 19014 14895 19066
rect 14907 19014 14959 19066
rect 14971 19014 15023 19066
rect 15035 19014 15087 19066
rect 1860 18912 1912 18964
rect 572 18844 624 18896
rect 5264 18912 5316 18964
rect 5448 18955 5500 18964
rect 5448 18921 5457 18955
rect 5457 18921 5491 18955
rect 5491 18921 5500 18955
rect 5448 18912 5500 18921
rect 5908 18955 5960 18964
rect 5908 18921 5917 18955
rect 5917 18921 5951 18955
rect 5951 18921 5960 18955
rect 5908 18912 5960 18921
rect 6368 18912 6420 18964
rect 7104 18912 7156 18964
rect 7656 18912 7708 18964
rect 10140 18955 10192 18964
rect 10140 18921 10149 18955
rect 10149 18921 10183 18955
rect 10183 18921 10192 18955
rect 10140 18912 10192 18921
rect 11612 18912 11664 18964
rect 13544 18912 13596 18964
rect 15568 18912 15620 18964
rect 19432 18912 19484 18964
rect 19800 18955 19852 18964
rect 19800 18921 19809 18955
rect 19809 18921 19843 18955
rect 19843 18921 19852 18955
rect 19800 18912 19852 18921
rect 20168 18912 20220 18964
rect 2228 18776 2280 18828
rect 2872 18776 2924 18828
rect 5816 18819 5868 18828
rect 5816 18785 5825 18819
rect 5825 18785 5859 18819
rect 5859 18785 5868 18819
rect 5816 18776 5868 18785
rect 6736 18844 6788 18896
rect 8852 18844 8904 18896
rect 17132 18844 17184 18896
rect 17868 18844 17920 18896
rect 6644 18819 6696 18828
rect 6644 18785 6653 18819
rect 6653 18785 6687 18819
rect 6687 18785 6696 18819
rect 6644 18776 6696 18785
rect 8392 18776 8444 18828
rect 2412 18708 2464 18760
rect 2688 18708 2740 18760
rect 4160 18751 4212 18760
rect 4160 18717 4169 18751
rect 4169 18717 4203 18751
rect 4203 18717 4212 18751
rect 4160 18708 4212 18717
rect 4988 18751 5040 18760
rect 1676 18640 1728 18692
rect 4068 18640 4120 18692
rect 4988 18717 4997 18751
rect 4997 18717 5031 18751
rect 5031 18717 5040 18751
rect 4988 18708 5040 18717
rect 5908 18640 5960 18692
rect 6184 18708 6236 18760
rect 6920 18751 6972 18760
rect 6920 18717 6929 18751
rect 6929 18717 6963 18751
rect 6963 18717 6972 18751
rect 6920 18708 6972 18717
rect 8116 18708 8168 18760
rect 8852 18751 8904 18760
rect 8852 18717 8861 18751
rect 8861 18717 8895 18751
rect 8895 18717 8904 18751
rect 8852 18708 8904 18717
rect 10232 18751 10284 18760
rect 10232 18717 10241 18751
rect 10241 18717 10275 18751
rect 10275 18717 10284 18751
rect 10232 18708 10284 18717
rect 11152 18776 11204 18828
rect 11244 18776 11296 18828
rect 12072 18776 12124 18828
rect 17592 18776 17644 18828
rect 18972 18844 19024 18896
rect 19248 18844 19300 18896
rect 7196 18640 7248 18692
rect 2504 18572 2556 18624
rect 3332 18572 3384 18624
rect 3792 18572 3844 18624
rect 4344 18615 4396 18624
rect 4344 18581 4353 18615
rect 4353 18581 4387 18615
rect 4387 18581 4396 18615
rect 4344 18572 4396 18581
rect 4988 18572 5040 18624
rect 8760 18640 8812 18692
rect 9864 18640 9916 18692
rect 10416 18572 10468 18624
rect 12992 18708 13044 18760
rect 18236 18751 18288 18760
rect 18236 18717 18245 18751
rect 18245 18717 18279 18751
rect 18279 18717 18288 18751
rect 18236 18708 18288 18717
rect 12072 18640 12124 18692
rect 13360 18640 13412 18692
rect 20720 18776 20772 18828
rect 22008 18844 22060 18896
rect 18788 18751 18840 18760
rect 18788 18717 18797 18751
rect 18797 18717 18831 18751
rect 18831 18717 18840 18751
rect 18788 18708 18840 18717
rect 19340 18751 19392 18760
rect 19340 18717 19349 18751
rect 19349 18717 19383 18751
rect 19383 18717 19392 18751
rect 19340 18708 19392 18717
rect 19800 18640 19852 18692
rect 11796 18572 11848 18624
rect 11980 18615 12032 18624
rect 11980 18581 11989 18615
rect 11989 18581 12023 18615
rect 12023 18581 12032 18615
rect 11980 18572 12032 18581
rect 13636 18615 13688 18624
rect 13636 18581 13645 18615
rect 13645 18581 13679 18615
rect 13679 18581 13688 18615
rect 13636 18572 13688 18581
rect 14188 18572 14240 18624
rect 14464 18615 14516 18624
rect 14464 18581 14473 18615
rect 14473 18581 14507 18615
rect 14507 18581 14516 18615
rect 14464 18572 14516 18581
rect 15568 18572 15620 18624
rect 16028 18572 16080 18624
rect 18604 18572 18656 18624
rect 20536 18572 20588 18624
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 4575 18470 4627 18522
rect 4639 18470 4691 18522
rect 11378 18470 11430 18522
rect 11442 18470 11494 18522
rect 11506 18470 11558 18522
rect 11570 18470 11622 18522
rect 18308 18470 18360 18522
rect 18372 18470 18424 18522
rect 18436 18470 18488 18522
rect 18500 18470 18552 18522
rect 2780 18368 2832 18420
rect 4160 18368 4212 18420
rect 4988 18368 5040 18420
rect 5816 18368 5868 18420
rect 7564 18368 7616 18420
rect 8116 18368 8168 18420
rect 8852 18368 8904 18420
rect 3056 18300 3108 18352
rect 940 18232 992 18284
rect 2136 18207 2188 18216
rect 2136 18173 2145 18207
rect 2145 18173 2179 18207
rect 2179 18173 2188 18207
rect 2136 18164 2188 18173
rect 2688 18164 2740 18216
rect 3148 18164 3200 18216
rect 2964 18096 3016 18148
rect 4620 18232 4672 18284
rect 5080 18232 5132 18284
rect 6092 18232 6144 18284
rect 4344 18207 4396 18216
rect 4344 18173 4353 18207
rect 4353 18173 4387 18207
rect 4387 18173 4396 18207
rect 4344 18164 4396 18173
rect 6276 18207 6328 18216
rect 6276 18173 6285 18207
rect 6285 18173 6319 18207
rect 6319 18173 6328 18207
rect 6276 18164 6328 18173
rect 7196 18300 7248 18352
rect 17040 18368 17092 18420
rect 18696 18411 18748 18420
rect 18696 18377 18705 18411
rect 18705 18377 18739 18411
rect 18739 18377 18748 18411
rect 18696 18368 18748 18377
rect 19708 18411 19760 18420
rect 19708 18377 19717 18411
rect 19717 18377 19751 18411
rect 19751 18377 19760 18411
rect 19708 18368 19760 18377
rect 20720 18368 20772 18420
rect 21456 18411 21508 18420
rect 21456 18377 21465 18411
rect 21465 18377 21499 18411
rect 21499 18377 21508 18411
rect 21456 18368 21508 18377
rect 6644 18232 6696 18284
rect 6920 18232 6972 18284
rect 11336 18300 11388 18352
rect 20168 18300 20220 18352
rect 8668 18207 8720 18216
rect 8668 18173 8677 18207
rect 8677 18173 8711 18207
rect 8711 18173 8720 18207
rect 8668 18164 8720 18173
rect 9864 18164 9916 18216
rect 10140 18207 10192 18216
rect 10140 18173 10149 18207
rect 10149 18173 10183 18207
rect 10183 18173 10192 18207
rect 10140 18164 10192 18173
rect 11796 18232 11848 18284
rect 12440 18275 12492 18284
rect 12440 18241 12449 18275
rect 12449 18241 12483 18275
rect 12483 18241 12492 18275
rect 12440 18232 12492 18241
rect 14556 18232 14608 18284
rect 10784 18164 10836 18216
rect 10968 18164 11020 18216
rect 11520 18164 11572 18216
rect 1952 18071 2004 18080
rect 1952 18037 1961 18071
rect 1961 18037 1995 18071
rect 1995 18037 2004 18071
rect 1952 18028 2004 18037
rect 2596 18028 2648 18080
rect 2872 18071 2924 18080
rect 2872 18037 2881 18071
rect 2881 18037 2915 18071
rect 2915 18037 2924 18071
rect 2872 18028 2924 18037
rect 3056 18071 3108 18080
rect 3056 18037 3065 18071
rect 3065 18037 3099 18071
rect 3099 18037 3108 18071
rect 3056 18028 3108 18037
rect 3884 18071 3936 18080
rect 3884 18037 3893 18071
rect 3893 18037 3927 18071
rect 3927 18037 3936 18071
rect 3884 18028 3936 18037
rect 4436 18096 4488 18148
rect 5632 18096 5684 18148
rect 8760 18096 8812 18148
rect 8852 18096 8904 18148
rect 10324 18096 10376 18148
rect 12164 18164 12216 18216
rect 13912 18207 13964 18216
rect 13912 18173 13921 18207
rect 13921 18173 13955 18207
rect 13955 18173 13964 18207
rect 13912 18164 13964 18173
rect 16488 18207 16540 18216
rect 16488 18173 16497 18207
rect 16497 18173 16531 18207
rect 16531 18173 16540 18207
rect 16488 18164 16540 18173
rect 18052 18164 18104 18216
rect 11980 18096 12032 18148
rect 20904 18096 20956 18148
rect 5264 18028 5316 18080
rect 7288 18028 7340 18080
rect 7748 18071 7800 18080
rect 7748 18037 7757 18071
rect 7757 18037 7791 18071
rect 7791 18037 7800 18071
rect 7748 18028 7800 18037
rect 8668 18028 8720 18080
rect 9312 18028 9364 18080
rect 10140 18028 10192 18080
rect 11152 18028 11204 18080
rect 12164 18028 12216 18080
rect 12808 18028 12860 18080
rect 19340 18071 19392 18080
rect 19340 18037 19349 18071
rect 19349 18037 19383 18071
rect 19383 18037 19392 18071
rect 19340 18028 19392 18037
rect 19984 18028 20036 18080
rect 7912 17926 7964 17978
rect 7976 17926 8028 17978
rect 8040 17926 8092 17978
rect 8104 17926 8156 17978
rect 14843 17926 14895 17978
rect 14907 17926 14959 17978
rect 14971 17926 15023 17978
rect 15035 17926 15087 17978
rect 1584 17867 1636 17876
rect 1584 17833 1593 17867
rect 1593 17833 1627 17867
rect 1627 17833 1636 17867
rect 1584 17824 1636 17833
rect 3056 17824 3108 17876
rect 3884 17824 3936 17876
rect 2136 17756 2188 17808
rect 4160 17824 4212 17876
rect 4436 17867 4488 17876
rect 4436 17833 4445 17867
rect 4445 17833 4479 17867
rect 4479 17833 4488 17867
rect 4436 17824 4488 17833
rect 4896 17867 4948 17876
rect 4896 17833 4905 17867
rect 4905 17833 4939 17867
rect 4939 17833 4948 17867
rect 4896 17824 4948 17833
rect 6092 17824 6144 17876
rect 6828 17824 6880 17876
rect 6920 17867 6972 17876
rect 6920 17833 6929 17867
rect 6929 17833 6963 17867
rect 6963 17833 6972 17867
rect 6920 17824 6972 17833
rect 8392 17824 8444 17876
rect 8852 17824 8904 17876
rect 9128 17824 9180 17876
rect 10232 17824 10284 17876
rect 10416 17867 10468 17876
rect 10416 17833 10425 17867
rect 10425 17833 10459 17867
rect 10459 17833 10468 17867
rect 10416 17824 10468 17833
rect 10876 17824 10928 17876
rect 11060 17824 11112 17876
rect 11520 17824 11572 17876
rect 11704 17824 11756 17876
rect 11980 17867 12032 17876
rect 11980 17833 11989 17867
rect 11989 17833 12023 17867
rect 12023 17833 12032 17867
rect 11980 17824 12032 17833
rect 13544 17867 13596 17876
rect 13544 17833 13553 17867
rect 13553 17833 13587 17867
rect 13587 17833 13596 17867
rect 13544 17824 13596 17833
rect 20076 17867 20128 17876
rect 20076 17833 20085 17867
rect 20085 17833 20119 17867
rect 20119 17833 20128 17867
rect 20076 17824 20128 17833
rect 21272 17824 21324 17876
rect 1400 17731 1452 17740
rect 1400 17697 1409 17731
rect 1409 17697 1443 17731
rect 1443 17697 1452 17731
rect 1400 17688 1452 17697
rect 4160 17688 4212 17740
rect 2136 17620 2188 17672
rect 2596 17620 2648 17672
rect 4896 17688 4948 17740
rect 6552 17688 6604 17740
rect 4620 17663 4672 17672
rect 2872 17552 2924 17604
rect 4620 17629 4629 17663
rect 4629 17629 4663 17663
rect 4663 17629 4672 17663
rect 4620 17620 4672 17629
rect 4988 17620 5040 17672
rect 5356 17663 5408 17672
rect 5356 17629 5365 17663
rect 5365 17629 5399 17663
rect 5399 17629 5408 17663
rect 5356 17620 5408 17629
rect 7656 17756 7708 17808
rect 7564 17688 7616 17740
rect 4068 17552 4120 17604
rect 10692 17756 10744 17808
rect 15292 17756 15344 17808
rect 15752 17756 15804 17808
rect 16488 17756 16540 17808
rect 11244 17731 11296 17740
rect 11244 17697 11253 17731
rect 11253 17697 11287 17731
rect 11287 17697 11296 17731
rect 11244 17688 11296 17697
rect 11796 17688 11848 17740
rect 13268 17688 13320 17740
rect 14188 17688 14240 17740
rect 15660 17731 15712 17740
rect 15660 17697 15669 17731
rect 15669 17697 15703 17731
rect 15703 17697 15712 17731
rect 15660 17688 15712 17697
rect 16212 17688 16264 17740
rect 8484 17663 8536 17672
rect 8484 17629 8493 17663
rect 8493 17629 8527 17663
rect 8527 17629 8536 17663
rect 8484 17620 8536 17629
rect 10784 17620 10836 17672
rect 11336 17663 11388 17672
rect 11336 17629 11345 17663
rect 11345 17629 11379 17663
rect 11379 17629 11388 17663
rect 11336 17620 11388 17629
rect 6828 17552 6880 17604
rect 8208 17552 8260 17604
rect 8392 17552 8444 17604
rect 9864 17552 9916 17604
rect 12164 17663 12216 17672
rect 12164 17629 12173 17663
rect 12173 17629 12207 17663
rect 12207 17629 12216 17663
rect 12164 17620 12216 17629
rect 15292 17620 15344 17672
rect 15384 17620 15436 17672
rect 15936 17663 15988 17672
rect 15936 17629 15945 17663
rect 15945 17629 15979 17663
rect 15979 17629 15988 17663
rect 15936 17620 15988 17629
rect 20720 17688 20772 17740
rect 20628 17620 20680 17672
rect 21548 17620 21600 17672
rect 17224 17552 17276 17604
rect 19708 17595 19760 17604
rect 19708 17561 19717 17595
rect 19717 17561 19751 17595
rect 19751 17561 19760 17595
rect 19708 17552 19760 17561
rect 22008 17595 22060 17604
rect 22008 17561 22017 17595
rect 22017 17561 22051 17595
rect 22051 17561 22060 17595
rect 22008 17552 22060 17561
rect 2228 17484 2280 17536
rect 2412 17484 2464 17536
rect 3240 17484 3292 17536
rect 3884 17484 3936 17536
rect 6736 17484 6788 17536
rect 7104 17484 7156 17536
rect 7656 17527 7708 17536
rect 7656 17493 7665 17527
rect 7665 17493 7699 17527
rect 7699 17493 7708 17527
rect 7656 17484 7708 17493
rect 7748 17484 7800 17536
rect 10140 17484 10192 17536
rect 10600 17484 10652 17536
rect 12256 17484 12308 17536
rect 13268 17484 13320 17536
rect 16580 17484 16632 17536
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 4575 17382 4627 17434
rect 4639 17382 4691 17434
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 18308 17382 18360 17434
rect 18372 17382 18424 17434
rect 18436 17382 18488 17434
rect 18500 17382 18552 17434
rect 5356 17280 5408 17332
rect 5908 17280 5960 17332
rect 6092 17280 6144 17332
rect 4068 17255 4120 17264
rect 4068 17221 4077 17255
rect 4077 17221 4111 17255
rect 4111 17221 4120 17255
rect 4068 17212 4120 17221
rect 4160 17255 4212 17264
rect 4160 17221 4169 17255
rect 4169 17221 4203 17255
rect 4203 17221 4212 17255
rect 4160 17212 4212 17221
rect 5540 17212 5592 17264
rect 6736 17280 6788 17332
rect 6920 17323 6972 17332
rect 6920 17289 6929 17323
rect 6929 17289 6963 17323
rect 6963 17289 6972 17323
rect 6920 17280 6972 17289
rect 7288 17280 7340 17332
rect 8668 17280 8720 17332
rect 9864 17323 9916 17332
rect 9864 17289 9873 17323
rect 9873 17289 9907 17323
rect 9907 17289 9916 17323
rect 9864 17280 9916 17289
rect 6368 17212 6420 17264
rect 2412 17144 2464 17196
rect 2228 17119 2280 17128
rect 2228 17085 2237 17119
rect 2237 17085 2271 17119
rect 2271 17085 2280 17119
rect 2228 17076 2280 17085
rect 3792 17144 3844 17196
rect 4712 17144 4764 17196
rect 4988 17144 5040 17196
rect 5632 17187 5684 17196
rect 5632 17153 5641 17187
rect 5641 17153 5675 17187
rect 5675 17153 5684 17187
rect 5632 17144 5684 17153
rect 6276 17144 6328 17196
rect 6552 17144 6604 17196
rect 7288 17144 7340 17196
rect 9220 17212 9272 17264
rect 9496 17212 9548 17264
rect 11980 17280 12032 17332
rect 15384 17323 15436 17332
rect 2688 17119 2740 17128
rect 2688 17085 2697 17119
rect 2697 17085 2731 17119
rect 2731 17085 2740 17119
rect 2688 17076 2740 17085
rect 3424 17076 3476 17128
rect 3976 17076 4028 17128
rect 5908 17076 5960 17128
rect 6184 17076 6236 17128
rect 6736 17076 6788 17128
rect 7840 17144 7892 17196
rect 8668 17187 8720 17196
rect 8668 17153 8677 17187
rect 8677 17153 8711 17187
rect 8711 17153 8720 17187
rect 8668 17144 8720 17153
rect 9588 17144 9640 17196
rect 9864 17144 9916 17196
rect 10784 17144 10836 17196
rect 11612 17187 11664 17196
rect 11612 17153 11621 17187
rect 11621 17153 11655 17187
rect 11655 17153 11664 17187
rect 11612 17144 11664 17153
rect 15384 17289 15393 17323
rect 15393 17289 15427 17323
rect 15427 17289 15436 17323
rect 15384 17280 15436 17289
rect 16212 17323 16264 17332
rect 16212 17289 16221 17323
rect 16221 17289 16255 17323
rect 16255 17289 16264 17323
rect 16212 17280 16264 17289
rect 20720 17280 20772 17332
rect 21640 17280 21692 17332
rect 15292 17255 15344 17264
rect 15292 17221 15301 17255
rect 15301 17221 15335 17255
rect 15335 17221 15344 17255
rect 15292 17212 15344 17221
rect 8484 17076 8536 17128
rect 9680 17119 9732 17128
rect 9680 17085 9689 17119
rect 9689 17085 9723 17119
rect 9723 17085 9732 17119
rect 9680 17076 9732 17085
rect 11060 17119 11112 17128
rect 11060 17085 11069 17119
rect 11069 17085 11103 17119
rect 11103 17085 11112 17119
rect 11060 17076 11112 17085
rect 11336 17076 11388 17128
rect 12440 17119 12492 17128
rect 12440 17085 12449 17119
rect 12449 17085 12483 17119
rect 12483 17085 12492 17119
rect 12440 17076 12492 17085
rect 13820 17076 13872 17128
rect 3240 17008 3292 17060
rect 3516 17008 3568 17060
rect 1400 16940 1452 16992
rect 4344 16940 4396 16992
rect 11704 17008 11756 17060
rect 13360 17008 13412 17060
rect 7104 16940 7156 16992
rect 8208 16983 8260 16992
rect 8208 16949 8217 16983
rect 8217 16949 8251 16983
rect 8251 16949 8260 16983
rect 8208 16940 8260 16949
rect 9496 16983 9548 16992
rect 9496 16949 9505 16983
rect 9505 16949 9539 16983
rect 9539 16949 9548 16983
rect 14280 17008 14332 17060
rect 16672 17144 16724 17196
rect 19524 17144 19576 17196
rect 15752 17076 15804 17128
rect 16580 17119 16632 17128
rect 16580 17085 16589 17119
rect 16589 17085 16623 17119
rect 16623 17085 16632 17119
rect 16580 17076 16632 17085
rect 19708 17076 19760 17128
rect 20444 17076 20496 17128
rect 19340 17008 19392 17060
rect 9496 16940 9548 16949
rect 14464 16940 14516 16992
rect 16764 16940 16816 16992
rect 21272 16940 21324 16992
rect 7912 16838 7964 16890
rect 7976 16838 8028 16890
rect 8040 16838 8092 16890
rect 8104 16838 8156 16890
rect 14843 16838 14895 16890
rect 14907 16838 14959 16890
rect 14971 16838 15023 16890
rect 15035 16838 15087 16890
rect 3700 16736 3752 16788
rect 6368 16736 6420 16788
rect 7380 16736 7432 16788
rect 8760 16779 8812 16788
rect 8760 16745 8769 16779
rect 8769 16745 8803 16779
rect 8803 16745 8812 16779
rect 8760 16736 8812 16745
rect 9956 16736 10008 16788
rect 10968 16736 11020 16788
rect 16764 16779 16816 16788
rect 2504 16668 2556 16720
rect 2688 16668 2740 16720
rect 4068 16668 4120 16720
rect 6092 16711 6144 16720
rect 6092 16677 6101 16711
rect 6101 16677 6135 16711
rect 6135 16677 6144 16711
rect 6092 16668 6144 16677
rect 1676 16600 1728 16652
rect 2596 16600 2648 16652
rect 5264 16600 5316 16652
rect 6644 16668 6696 16720
rect 8116 16668 8168 16720
rect 10508 16668 10560 16720
rect 16764 16745 16773 16779
rect 16773 16745 16807 16779
rect 16807 16745 16816 16779
rect 16764 16736 16816 16745
rect 17224 16779 17276 16788
rect 17224 16745 17233 16779
rect 17233 16745 17267 16779
rect 17267 16745 17276 16779
rect 17224 16736 17276 16745
rect 11612 16711 11664 16720
rect 6368 16600 6420 16652
rect 7564 16643 7616 16652
rect 4068 16532 4120 16584
rect 6276 16575 6328 16584
rect 6276 16541 6285 16575
rect 6285 16541 6319 16575
rect 6319 16541 6328 16575
rect 6276 16532 6328 16541
rect 7564 16609 7598 16643
rect 7598 16609 7616 16643
rect 7564 16600 7616 16609
rect 9128 16643 9180 16652
rect 9128 16609 9137 16643
rect 9137 16609 9171 16643
rect 9171 16609 9180 16643
rect 9128 16600 9180 16609
rect 7196 16532 7248 16584
rect 8484 16532 8536 16584
rect 3792 16507 3844 16516
rect 3792 16473 3801 16507
rect 3801 16473 3835 16507
rect 3835 16473 3844 16507
rect 3792 16464 3844 16473
rect 9680 16600 9732 16652
rect 11060 16600 11112 16652
rect 11612 16677 11621 16711
rect 11621 16677 11655 16711
rect 11655 16677 11664 16711
rect 11612 16668 11664 16677
rect 2504 16396 2556 16448
rect 3240 16439 3292 16448
rect 3240 16405 3249 16439
rect 3249 16405 3283 16439
rect 3283 16405 3292 16439
rect 3240 16396 3292 16405
rect 3332 16396 3384 16448
rect 5632 16439 5684 16448
rect 5632 16405 5641 16439
rect 5641 16405 5675 16439
rect 5675 16405 5684 16439
rect 5632 16396 5684 16405
rect 8760 16396 8812 16448
rect 9864 16464 9916 16516
rect 11336 16464 11388 16516
rect 12440 16643 12492 16652
rect 12440 16609 12449 16643
rect 12449 16609 12483 16643
rect 12483 16609 12492 16643
rect 13268 16643 13320 16652
rect 12440 16600 12492 16609
rect 13268 16609 13277 16643
rect 13277 16609 13311 16643
rect 13311 16609 13320 16643
rect 13268 16600 13320 16609
rect 12716 16575 12768 16584
rect 12716 16541 12725 16575
rect 12725 16541 12759 16575
rect 12759 16541 12768 16575
rect 12716 16532 12768 16541
rect 13360 16532 13412 16584
rect 12256 16464 12308 16516
rect 20444 16668 20496 16720
rect 13912 16600 13964 16652
rect 14464 16600 14516 16652
rect 15568 16643 15620 16652
rect 15568 16609 15602 16643
rect 15602 16609 15620 16643
rect 15568 16600 15620 16609
rect 15936 16600 15988 16652
rect 17132 16643 17184 16652
rect 14280 16575 14332 16584
rect 14280 16541 14289 16575
rect 14289 16541 14323 16575
rect 14323 16541 14332 16575
rect 14280 16532 14332 16541
rect 17132 16609 17141 16643
rect 17141 16609 17175 16643
rect 17175 16609 17184 16643
rect 17132 16600 17184 16609
rect 20812 16600 20864 16652
rect 12808 16396 12860 16448
rect 16672 16507 16724 16516
rect 16672 16473 16681 16507
rect 16681 16473 16715 16507
rect 16715 16473 16724 16507
rect 16672 16464 16724 16473
rect 15936 16396 15988 16448
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 4575 16294 4627 16346
rect 4639 16294 4691 16346
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 18308 16294 18360 16346
rect 18372 16294 18424 16346
rect 18436 16294 18488 16346
rect 18500 16294 18552 16346
rect 1584 16235 1636 16244
rect 1584 16201 1593 16235
rect 1593 16201 1627 16235
rect 1627 16201 1636 16235
rect 1584 16192 1636 16201
rect 2320 16235 2372 16244
rect 2320 16201 2329 16235
rect 2329 16201 2363 16235
rect 2363 16201 2372 16235
rect 2320 16192 2372 16201
rect 2780 16192 2832 16244
rect 2872 16235 2924 16244
rect 2872 16201 2881 16235
rect 2881 16201 2915 16235
rect 2915 16201 2924 16235
rect 2872 16192 2924 16201
rect 3056 16192 3108 16244
rect 4252 16192 4304 16244
rect 4804 16235 4856 16244
rect 4804 16201 4813 16235
rect 4813 16201 4847 16235
rect 4847 16201 4856 16235
rect 4804 16192 4856 16201
rect 5264 16192 5316 16244
rect 2596 16124 2648 16176
rect 3240 16056 3292 16108
rect 4068 16124 4120 16176
rect 7196 16192 7248 16244
rect 7564 16192 7616 16244
rect 8760 16192 8812 16244
rect 8116 16124 8168 16176
rect 10692 16192 10744 16244
rect 15476 16192 15528 16244
rect 15568 16192 15620 16244
rect 19064 16192 19116 16244
rect 20996 16235 21048 16244
rect 20996 16201 21005 16235
rect 21005 16201 21039 16235
rect 21039 16201 21048 16235
rect 20996 16192 21048 16201
rect 21364 16235 21416 16244
rect 21364 16201 21373 16235
rect 21373 16201 21407 16235
rect 21407 16201 21416 16235
rect 21364 16192 21416 16201
rect 17500 16124 17552 16176
rect 20168 16124 20220 16176
rect 1400 16031 1452 16040
rect 1400 15997 1409 16031
rect 1409 15997 1443 16031
rect 1443 15997 1452 16031
rect 1400 15988 1452 15997
rect 1768 16031 1820 16040
rect 1768 15997 1777 16031
rect 1777 15997 1811 16031
rect 1811 15997 1820 16031
rect 1768 15988 1820 15997
rect 3332 15988 3384 16040
rect 4804 15988 4856 16040
rect 9128 16056 9180 16108
rect 9312 16056 9364 16108
rect 11152 16056 11204 16108
rect 12348 16056 12400 16108
rect 3056 15920 3108 15972
rect 3976 15920 4028 15972
rect 4252 15920 4304 15972
rect 5356 15920 5408 15972
rect 5908 15920 5960 15972
rect 1952 15895 2004 15904
rect 1952 15861 1961 15895
rect 1961 15861 1995 15895
rect 1995 15861 2004 15895
rect 1952 15852 2004 15861
rect 3240 15895 3292 15904
rect 3240 15861 3249 15895
rect 3249 15861 3283 15895
rect 3283 15861 3292 15895
rect 3240 15852 3292 15861
rect 4436 15852 4488 15904
rect 5264 15852 5316 15904
rect 6736 15920 6788 15972
rect 8208 15920 8260 15972
rect 12072 15988 12124 16040
rect 17040 16056 17092 16108
rect 12532 15988 12584 16040
rect 12716 16031 12768 16040
rect 12716 15997 12750 16031
rect 12750 15997 12768 16031
rect 12716 15988 12768 15997
rect 13912 15988 13964 16040
rect 9864 15963 9916 15972
rect 9864 15929 9898 15963
rect 9898 15929 9916 15963
rect 9864 15920 9916 15929
rect 7104 15852 7156 15904
rect 8760 15895 8812 15904
rect 8760 15861 8769 15895
rect 8769 15861 8803 15895
rect 8803 15861 8812 15895
rect 8760 15852 8812 15861
rect 8944 15852 8996 15904
rect 10048 15852 10100 15904
rect 11152 15852 11204 15904
rect 12348 15920 12400 15972
rect 12808 15920 12860 15972
rect 15292 15988 15344 16040
rect 15936 16031 15988 16040
rect 15936 15997 15945 16031
rect 15945 15997 15979 16031
rect 15979 15997 15988 16031
rect 15936 15988 15988 15997
rect 16672 15988 16724 16040
rect 16304 15920 16356 15972
rect 13360 15852 13412 15904
rect 13820 15895 13872 15904
rect 13820 15861 13829 15895
rect 13829 15861 13863 15895
rect 13863 15861 13872 15895
rect 13820 15852 13872 15861
rect 14004 15895 14056 15904
rect 14004 15861 14013 15895
rect 14013 15861 14047 15895
rect 14047 15861 14056 15895
rect 14004 15852 14056 15861
rect 17040 15852 17092 15904
rect 17408 15895 17460 15904
rect 17408 15861 17417 15895
rect 17417 15861 17451 15895
rect 17451 15861 17460 15895
rect 17408 15852 17460 15861
rect 7912 15750 7964 15802
rect 7976 15750 8028 15802
rect 8040 15750 8092 15802
rect 8104 15750 8156 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 15035 15750 15087 15802
rect 1676 15648 1728 15700
rect 1400 15580 1452 15632
rect 2596 15648 2648 15700
rect 4436 15691 4488 15700
rect 4436 15657 4445 15691
rect 4445 15657 4479 15691
rect 4479 15657 4488 15691
rect 4436 15648 4488 15657
rect 3516 15580 3568 15632
rect 5632 15648 5684 15700
rect 6368 15648 6420 15700
rect 7380 15648 7432 15700
rect 9220 15691 9272 15700
rect 8760 15580 8812 15632
rect 1584 15351 1636 15360
rect 1584 15317 1593 15351
rect 1593 15317 1627 15351
rect 1627 15317 1636 15351
rect 1584 15308 1636 15317
rect 2504 15512 2556 15564
rect 4160 15512 4212 15564
rect 5264 15512 5316 15564
rect 5540 15512 5592 15564
rect 7104 15512 7156 15564
rect 8116 15555 8168 15564
rect 8116 15521 8125 15555
rect 8125 15521 8159 15555
rect 8159 15521 8168 15555
rect 8116 15512 8168 15521
rect 9220 15657 9229 15691
rect 9229 15657 9263 15691
rect 9263 15657 9272 15691
rect 9220 15648 9272 15657
rect 9864 15648 9916 15700
rect 12164 15648 12216 15700
rect 12440 15648 12492 15700
rect 13268 15648 13320 15700
rect 13544 15691 13596 15700
rect 13544 15657 13553 15691
rect 13553 15657 13587 15691
rect 13587 15657 13596 15691
rect 13544 15648 13596 15657
rect 13728 15648 13780 15700
rect 14096 15648 14148 15700
rect 9312 15580 9364 15632
rect 9956 15555 10008 15564
rect 9956 15521 9990 15555
rect 9990 15521 10008 15555
rect 11980 15580 12032 15632
rect 12072 15580 12124 15632
rect 15660 15648 15712 15700
rect 17408 15648 17460 15700
rect 19340 15648 19392 15700
rect 21088 15691 21140 15700
rect 12624 15555 12676 15564
rect 9956 15512 10008 15521
rect 4988 15487 5040 15496
rect 4988 15453 4997 15487
rect 4997 15453 5031 15487
rect 5031 15453 5040 15487
rect 5908 15487 5960 15496
rect 4988 15444 5040 15453
rect 5908 15453 5917 15487
rect 5917 15453 5951 15487
rect 5951 15453 5960 15487
rect 5908 15444 5960 15453
rect 6736 15487 6788 15496
rect 6736 15453 6745 15487
rect 6745 15453 6779 15487
rect 6779 15453 6788 15487
rect 6736 15444 6788 15453
rect 6828 15444 6880 15496
rect 7380 15487 7432 15496
rect 7380 15453 7389 15487
rect 7389 15453 7423 15487
rect 7423 15453 7432 15487
rect 7380 15444 7432 15453
rect 7472 15487 7524 15496
rect 7472 15453 7481 15487
rect 7481 15453 7515 15487
rect 7515 15453 7524 15487
rect 7472 15444 7524 15453
rect 8760 15444 8812 15496
rect 8944 15444 8996 15496
rect 6368 15376 6420 15428
rect 4988 15308 5040 15360
rect 5356 15308 5408 15360
rect 9128 15376 9180 15428
rect 6736 15308 6788 15360
rect 8208 15308 8260 15360
rect 11152 15376 11204 15428
rect 11244 15351 11296 15360
rect 11244 15317 11253 15351
rect 11253 15317 11287 15351
rect 11287 15317 11296 15351
rect 11244 15308 11296 15317
rect 12624 15521 12633 15555
rect 12633 15521 12667 15555
rect 12667 15521 12676 15555
rect 12624 15512 12676 15521
rect 14004 15512 14056 15564
rect 14280 15555 14332 15564
rect 14280 15521 14289 15555
rect 14289 15521 14323 15555
rect 14323 15521 14332 15555
rect 14280 15512 14332 15521
rect 11888 15487 11940 15496
rect 11888 15453 11897 15487
rect 11897 15453 11931 15487
rect 11931 15453 11940 15487
rect 11888 15444 11940 15453
rect 12716 15487 12768 15496
rect 12716 15453 12725 15487
rect 12725 15453 12759 15487
rect 12759 15453 12768 15487
rect 12716 15444 12768 15453
rect 12900 15487 12952 15496
rect 12900 15453 12909 15487
rect 12909 15453 12943 15487
rect 12943 15453 12952 15487
rect 13728 15487 13780 15496
rect 12900 15444 12952 15453
rect 13728 15453 13737 15487
rect 13737 15453 13771 15487
rect 13771 15453 13780 15487
rect 13728 15444 13780 15453
rect 17132 15580 17184 15632
rect 17224 15623 17276 15632
rect 17224 15589 17233 15623
rect 17233 15589 17267 15623
rect 17267 15589 17276 15623
rect 17224 15580 17276 15589
rect 15476 15512 15528 15564
rect 16856 15512 16908 15564
rect 20812 15580 20864 15632
rect 21088 15657 21097 15691
rect 21097 15657 21131 15691
rect 21131 15657 21140 15691
rect 21088 15648 21140 15657
rect 21456 15691 21508 15700
rect 21456 15657 21465 15691
rect 21465 15657 21499 15691
rect 21499 15657 21508 15691
rect 21456 15648 21508 15657
rect 18144 15555 18196 15564
rect 15844 15444 15896 15496
rect 13820 15376 13872 15428
rect 14004 15376 14056 15428
rect 15292 15376 15344 15428
rect 16304 15444 16356 15496
rect 18144 15521 18153 15555
rect 18153 15521 18187 15555
rect 18187 15521 18196 15555
rect 18144 15512 18196 15521
rect 17040 15444 17092 15496
rect 16856 15376 16908 15428
rect 17960 15376 18012 15428
rect 18696 15376 18748 15428
rect 19156 15308 19208 15360
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 4575 15206 4627 15258
rect 4639 15206 4691 15258
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 18308 15206 18360 15258
rect 18372 15206 18424 15258
rect 18436 15206 18488 15258
rect 18500 15206 18552 15258
rect 3240 15104 3292 15156
rect 3976 15147 4028 15156
rect 3976 15113 3985 15147
rect 3985 15113 4019 15147
rect 4019 15113 4028 15147
rect 3976 15104 4028 15113
rect 1768 15079 1820 15088
rect 1768 15045 1777 15079
rect 1777 15045 1811 15079
rect 1811 15045 1820 15079
rect 1768 15036 1820 15045
rect 2596 15011 2648 15020
rect 2596 14977 2605 15011
rect 2605 14977 2639 15011
rect 2639 14977 2648 15011
rect 2596 14968 2648 14977
rect 4160 14968 4212 15020
rect 5080 15104 5132 15156
rect 6368 15147 6420 15156
rect 6368 15113 6377 15147
rect 6377 15113 6411 15147
rect 6411 15113 6420 15147
rect 6368 15104 6420 15113
rect 6736 15104 6788 15156
rect 7748 15104 7800 15156
rect 5908 15036 5960 15088
rect 7472 15036 7524 15088
rect 4804 15011 4856 15020
rect 4804 14977 4813 15011
rect 4813 14977 4847 15011
rect 4847 14977 4856 15011
rect 4804 14968 4856 14977
rect 8024 15036 8076 15088
rect 8208 15036 8260 15088
rect 7932 15011 7984 15020
rect 7932 14977 7941 15011
rect 7941 14977 7975 15011
rect 7975 14977 7984 15011
rect 7932 14968 7984 14977
rect 8392 14968 8444 15020
rect 1584 14943 1636 14952
rect 1584 14909 1593 14943
rect 1593 14909 1627 14943
rect 1627 14909 1636 14943
rect 4344 14943 4396 14952
rect 1584 14900 1636 14909
rect 4344 14909 4353 14943
rect 4353 14909 4387 14943
rect 4387 14909 4396 14943
rect 4344 14900 4396 14909
rect 5356 14900 5408 14952
rect 7564 14900 7616 14952
rect 9956 15104 10008 15156
rect 10600 15104 10652 15156
rect 11888 15104 11940 15156
rect 15936 15104 15988 15156
rect 16580 15104 16632 15156
rect 17960 15104 18012 15156
rect 20996 15147 21048 15156
rect 20996 15113 21005 15147
rect 21005 15113 21039 15147
rect 21039 15113 21048 15147
rect 20996 15104 21048 15113
rect 11244 15036 11296 15088
rect 12072 15036 12124 15088
rect 13728 15036 13780 15088
rect 16304 15036 16356 15088
rect 10876 14968 10928 15020
rect 12164 15011 12216 15020
rect 12164 14977 12173 15011
rect 12173 14977 12207 15011
rect 12207 14977 12216 15011
rect 12164 14968 12216 14977
rect 14280 14968 14332 15020
rect 15384 15011 15436 15020
rect 15384 14977 15393 15011
rect 15393 14977 15427 15011
rect 15427 14977 15436 15011
rect 15384 14968 15436 14977
rect 9128 14900 9180 14952
rect 9864 14900 9916 14952
rect 2596 14764 2648 14816
rect 3056 14764 3108 14816
rect 6092 14832 6144 14884
rect 8944 14832 8996 14884
rect 12072 14900 12124 14952
rect 12532 14900 12584 14952
rect 13176 14900 13228 14952
rect 15844 14943 15896 14952
rect 15844 14909 15853 14943
rect 15853 14909 15887 14943
rect 15887 14909 15896 14943
rect 15844 14900 15896 14909
rect 11336 14832 11388 14884
rect 12808 14832 12860 14884
rect 16120 14832 16172 14884
rect 17316 14968 17368 15020
rect 20168 15011 20220 15020
rect 20168 14977 20177 15011
rect 20177 14977 20211 15011
rect 20211 14977 20220 15011
rect 20168 14968 20220 14977
rect 16396 14900 16448 14952
rect 17960 14900 18012 14952
rect 20812 14943 20864 14952
rect 20812 14909 20821 14943
rect 20821 14909 20855 14943
rect 20855 14909 20864 14943
rect 20812 14900 20864 14909
rect 18880 14832 18932 14884
rect 3424 14764 3476 14816
rect 3608 14807 3660 14816
rect 3608 14773 3617 14807
rect 3617 14773 3651 14807
rect 3651 14773 3660 14807
rect 3608 14764 3660 14773
rect 5172 14764 5224 14816
rect 6736 14764 6788 14816
rect 7288 14807 7340 14816
rect 7288 14773 7297 14807
rect 7297 14773 7331 14807
rect 7331 14773 7340 14807
rect 7288 14764 7340 14773
rect 8668 14764 8720 14816
rect 10140 14764 10192 14816
rect 10416 14764 10468 14816
rect 11980 14807 12032 14816
rect 11980 14773 11989 14807
rect 11989 14773 12023 14807
rect 12023 14773 12032 14807
rect 11980 14764 12032 14773
rect 14096 14764 14148 14816
rect 15292 14807 15344 14816
rect 15292 14773 15301 14807
rect 15301 14773 15335 14807
rect 15335 14773 15344 14807
rect 15292 14764 15344 14773
rect 16028 14764 16080 14816
rect 19524 14807 19576 14816
rect 19524 14773 19533 14807
rect 19533 14773 19567 14807
rect 19567 14773 19576 14807
rect 21180 14807 21232 14816
rect 19524 14764 19576 14773
rect 21180 14773 21189 14807
rect 21189 14773 21223 14807
rect 21223 14773 21232 14807
rect 21180 14764 21232 14773
rect 7912 14662 7964 14714
rect 7976 14662 8028 14714
rect 8040 14662 8092 14714
rect 8104 14662 8156 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 15035 14662 15087 14714
rect 1860 14603 1912 14612
rect 1860 14569 1869 14603
rect 1869 14569 1903 14603
rect 1903 14569 1912 14603
rect 1860 14560 1912 14569
rect 3056 14560 3108 14612
rect 3608 14560 3660 14612
rect 3792 14603 3844 14612
rect 3792 14569 3801 14603
rect 3801 14569 3835 14603
rect 3835 14569 3844 14603
rect 3792 14560 3844 14569
rect 3976 14560 4028 14612
rect 4344 14560 4396 14612
rect 5724 14560 5776 14612
rect 5816 14560 5868 14612
rect 6552 14603 6604 14612
rect 6552 14569 6561 14603
rect 6561 14569 6595 14603
rect 6595 14569 6604 14603
rect 6552 14560 6604 14569
rect 7012 14560 7064 14612
rect 7288 14560 7340 14612
rect 9864 14603 9916 14612
rect 1676 14467 1728 14476
rect 1676 14433 1685 14467
rect 1685 14433 1719 14467
rect 1719 14433 1728 14467
rect 1676 14424 1728 14433
rect 2044 14467 2096 14476
rect 2044 14433 2053 14467
rect 2053 14433 2087 14467
rect 2087 14433 2096 14467
rect 2044 14424 2096 14433
rect 2688 14424 2740 14476
rect 6828 14492 6880 14544
rect 9864 14569 9873 14603
rect 9873 14569 9907 14603
rect 9907 14569 9916 14603
rect 9864 14560 9916 14569
rect 10232 14603 10284 14612
rect 10232 14569 10241 14603
rect 10241 14569 10275 14603
rect 10275 14569 10284 14603
rect 10232 14560 10284 14569
rect 3792 14424 3844 14476
rect 4804 14424 4856 14476
rect 8208 14492 8260 14544
rect 10784 14560 10836 14612
rect 11060 14603 11112 14612
rect 11060 14569 11069 14603
rect 11069 14569 11103 14603
rect 11103 14569 11112 14603
rect 11060 14560 11112 14569
rect 11152 14560 11204 14612
rect 11796 14560 11848 14612
rect 12440 14560 12492 14612
rect 13544 14560 13596 14612
rect 7840 14467 7892 14476
rect 7840 14433 7874 14467
rect 7874 14433 7892 14467
rect 7840 14424 7892 14433
rect 8116 14424 8168 14476
rect 14280 14560 14332 14612
rect 15844 14560 15896 14612
rect 19524 14560 19576 14612
rect 9036 14424 9088 14476
rect 2320 14399 2372 14408
rect 2320 14365 2329 14399
rect 2329 14365 2363 14399
rect 2363 14365 2372 14399
rect 2320 14356 2372 14365
rect 2596 14288 2648 14340
rect 1400 14220 1452 14272
rect 4160 14356 4212 14408
rect 5816 14356 5868 14408
rect 6000 14399 6052 14408
rect 6000 14365 6009 14399
rect 6009 14365 6043 14399
rect 6043 14365 6052 14399
rect 6000 14356 6052 14365
rect 6184 14399 6236 14408
rect 6184 14365 6193 14399
rect 6193 14365 6227 14399
rect 6227 14365 6236 14399
rect 6184 14356 6236 14365
rect 7196 14399 7248 14408
rect 7196 14365 7205 14399
rect 7205 14365 7239 14399
rect 7239 14365 7248 14399
rect 7196 14356 7248 14365
rect 7472 14356 7524 14408
rect 9956 14399 10008 14408
rect 9956 14365 9965 14399
rect 9965 14365 9999 14399
rect 9999 14365 10008 14399
rect 9956 14356 10008 14365
rect 10876 14399 10928 14408
rect 10876 14365 10885 14399
rect 10885 14365 10919 14399
rect 10919 14365 10928 14399
rect 10876 14356 10928 14365
rect 10968 14356 11020 14408
rect 5908 14288 5960 14340
rect 8944 14331 8996 14340
rect 8944 14297 8953 14331
rect 8953 14297 8987 14331
rect 8987 14297 8996 14331
rect 8944 14288 8996 14297
rect 9404 14288 9456 14340
rect 10600 14288 10652 14340
rect 15384 14492 15436 14544
rect 16028 14492 16080 14544
rect 19432 14535 19484 14544
rect 19432 14501 19441 14535
rect 19441 14501 19475 14535
rect 19475 14501 19484 14535
rect 21088 14603 21140 14612
rect 21088 14569 21097 14603
rect 21097 14569 21131 14603
rect 21131 14569 21140 14603
rect 21088 14560 21140 14569
rect 21456 14603 21508 14612
rect 21456 14569 21465 14603
rect 21465 14569 21499 14603
rect 21499 14569 21508 14603
rect 21456 14560 21508 14569
rect 19432 14492 19484 14501
rect 20812 14492 20864 14544
rect 21180 14492 21232 14544
rect 12532 14424 12584 14476
rect 13728 14424 13780 14476
rect 16672 14424 16724 14476
rect 17592 14424 17644 14476
rect 18604 14424 18656 14476
rect 19156 14424 19208 14476
rect 21088 14424 21140 14476
rect 12992 14399 13044 14408
rect 12992 14365 13001 14399
rect 13001 14365 13035 14399
rect 13035 14365 13044 14399
rect 12992 14356 13044 14365
rect 13084 14399 13136 14408
rect 13084 14365 13093 14399
rect 13093 14365 13127 14399
rect 13127 14365 13136 14399
rect 13084 14356 13136 14365
rect 16580 14356 16632 14408
rect 17316 14356 17368 14408
rect 12624 14288 12676 14340
rect 18880 14331 18932 14340
rect 18880 14297 18889 14331
rect 18889 14297 18923 14331
rect 18923 14297 18932 14331
rect 18880 14288 18932 14297
rect 20352 14356 20404 14408
rect 3056 14220 3108 14272
rect 3608 14220 3660 14272
rect 5172 14263 5224 14272
rect 5172 14229 5181 14263
rect 5181 14229 5215 14263
rect 5215 14229 5224 14263
rect 5172 14220 5224 14229
rect 5540 14263 5592 14272
rect 5540 14229 5549 14263
rect 5549 14229 5583 14263
rect 5583 14229 5592 14263
rect 5540 14220 5592 14229
rect 9220 14220 9272 14272
rect 10784 14220 10836 14272
rect 13820 14220 13872 14272
rect 14372 14220 14424 14272
rect 16396 14220 16448 14272
rect 16948 14220 17000 14272
rect 17776 14220 17828 14272
rect 18972 14263 19024 14272
rect 18972 14229 18981 14263
rect 18981 14229 19015 14263
rect 19015 14229 19024 14263
rect 18972 14220 19024 14229
rect 21088 14220 21140 14272
rect 21456 14220 21508 14272
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 4575 14118 4627 14170
rect 4639 14118 4691 14170
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 18308 14118 18360 14170
rect 18372 14118 18424 14170
rect 18436 14118 18488 14170
rect 18500 14118 18552 14170
rect 1768 14059 1820 14068
rect 1768 14025 1777 14059
rect 1777 14025 1811 14059
rect 1811 14025 1820 14059
rect 1768 14016 1820 14025
rect 1584 13855 1636 13864
rect 1584 13821 1593 13855
rect 1593 13821 1627 13855
rect 1627 13821 1636 13855
rect 1584 13812 1636 13821
rect 5632 14016 5684 14068
rect 5816 14059 5868 14068
rect 5816 14025 5825 14059
rect 5825 14025 5859 14059
rect 5859 14025 5868 14059
rect 5816 14016 5868 14025
rect 7012 14016 7064 14068
rect 7104 14016 7156 14068
rect 2596 13948 2648 14000
rect 5908 13948 5960 14000
rect 8944 14016 8996 14068
rect 10968 14016 11020 14068
rect 13176 14016 13228 14068
rect 10508 13991 10560 14000
rect 6184 13880 6236 13932
rect 7380 13923 7432 13932
rect 7380 13889 7389 13923
rect 7389 13889 7423 13923
rect 7423 13889 7432 13923
rect 7380 13880 7432 13889
rect 7472 13880 7524 13932
rect 2596 13855 2648 13864
rect 2596 13821 2605 13855
rect 2605 13821 2639 13855
rect 2639 13821 2648 13855
rect 2596 13812 2648 13821
rect 3976 13812 4028 13864
rect 4528 13812 4580 13864
rect 6552 13812 6604 13864
rect 7104 13812 7156 13864
rect 8116 13855 8168 13864
rect 8116 13821 8125 13855
rect 8125 13821 8159 13855
rect 8159 13821 8168 13855
rect 8116 13812 8168 13821
rect 3240 13744 3292 13796
rect 4160 13744 4212 13796
rect 5816 13676 5868 13728
rect 5908 13719 5960 13728
rect 5908 13685 5917 13719
rect 5917 13685 5951 13719
rect 5951 13685 5960 13719
rect 5908 13676 5960 13685
rect 6092 13676 6144 13728
rect 9036 13880 9088 13932
rect 9404 13880 9456 13932
rect 8852 13812 8904 13864
rect 9220 13812 9272 13864
rect 9864 13880 9916 13932
rect 10140 13923 10192 13932
rect 10140 13889 10149 13923
rect 10149 13889 10183 13923
rect 10183 13889 10192 13923
rect 10140 13880 10192 13889
rect 10508 13957 10517 13991
rect 10517 13957 10551 13991
rect 10551 13957 10560 13991
rect 10508 13948 10560 13957
rect 10048 13812 10100 13864
rect 12256 13948 12308 14000
rect 13820 14016 13872 14068
rect 15292 14016 15344 14068
rect 14740 13948 14792 14000
rect 15384 13948 15436 14000
rect 15752 13948 15804 14000
rect 17592 14059 17644 14068
rect 17592 14025 17601 14059
rect 17601 14025 17635 14059
rect 17635 14025 17644 14059
rect 17592 14016 17644 14025
rect 17960 14016 18012 14068
rect 18144 14016 18196 14068
rect 19064 14016 19116 14068
rect 20996 14059 21048 14068
rect 15292 13880 15344 13932
rect 16396 13923 16448 13932
rect 16396 13889 16405 13923
rect 16405 13889 16439 13923
rect 16439 13889 16448 13923
rect 16396 13880 16448 13889
rect 11796 13812 11848 13864
rect 8944 13744 8996 13796
rect 10324 13744 10376 13796
rect 11060 13744 11112 13796
rect 11612 13787 11664 13796
rect 11612 13753 11621 13787
rect 11621 13753 11655 13787
rect 11655 13753 11664 13787
rect 11612 13744 11664 13753
rect 11888 13744 11940 13796
rect 12256 13744 12308 13796
rect 14096 13812 14148 13864
rect 15476 13812 15528 13864
rect 15844 13812 15896 13864
rect 15936 13812 15988 13864
rect 19340 13948 19392 14000
rect 20996 14025 21005 14059
rect 21005 14025 21039 14059
rect 21039 14025 21048 14059
rect 20996 14016 21048 14025
rect 18604 13923 18656 13932
rect 18604 13889 18613 13923
rect 18613 13889 18647 13923
rect 18647 13889 18656 13923
rect 18604 13880 18656 13889
rect 18880 13880 18932 13932
rect 13912 13744 13964 13796
rect 18696 13812 18748 13864
rect 18972 13812 19024 13864
rect 20536 13855 20588 13864
rect 7380 13676 7432 13728
rect 8760 13676 8812 13728
rect 8852 13676 8904 13728
rect 12440 13719 12492 13728
rect 12440 13685 12449 13719
rect 12449 13685 12483 13719
rect 12483 13685 12492 13719
rect 12440 13676 12492 13685
rect 13176 13719 13228 13728
rect 13176 13685 13185 13719
rect 13185 13685 13219 13719
rect 13219 13685 13228 13719
rect 13176 13676 13228 13685
rect 13728 13676 13780 13728
rect 17960 13744 18012 13796
rect 20536 13821 20545 13855
rect 20545 13821 20579 13855
rect 20579 13821 20588 13855
rect 20536 13812 20588 13821
rect 21272 13855 21324 13864
rect 21272 13821 21281 13855
rect 21281 13821 21315 13855
rect 21315 13821 21324 13855
rect 21272 13812 21324 13821
rect 14096 13676 14148 13728
rect 15384 13719 15436 13728
rect 15384 13685 15393 13719
rect 15393 13685 15427 13719
rect 15427 13685 15436 13719
rect 15384 13676 15436 13685
rect 15476 13719 15528 13728
rect 15476 13685 15485 13719
rect 15485 13685 15519 13719
rect 15519 13685 15528 13719
rect 15476 13676 15528 13685
rect 15752 13676 15804 13728
rect 16488 13676 16540 13728
rect 17592 13676 17644 13728
rect 7912 13574 7964 13626
rect 7976 13574 8028 13626
rect 8040 13574 8092 13626
rect 8104 13574 8156 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 15035 13574 15087 13626
rect 2412 13515 2464 13524
rect 2412 13481 2421 13515
rect 2421 13481 2455 13515
rect 2455 13481 2464 13515
rect 2412 13472 2464 13481
rect 2780 13515 2832 13524
rect 2780 13481 2789 13515
rect 2789 13481 2823 13515
rect 2823 13481 2832 13515
rect 2780 13472 2832 13481
rect 3792 13472 3844 13524
rect 4160 13472 4212 13524
rect 5356 13472 5408 13524
rect 6092 13515 6144 13524
rect 6092 13481 6101 13515
rect 6101 13481 6135 13515
rect 6135 13481 6144 13515
rect 6092 13472 6144 13481
rect 6184 13472 6236 13524
rect 6552 13472 6604 13524
rect 7012 13472 7064 13524
rect 4528 13404 4580 13456
rect 5816 13404 5868 13456
rect 8300 13472 8352 13524
rect 9496 13515 9548 13524
rect 9496 13481 9505 13515
rect 9505 13481 9539 13515
rect 9539 13481 9548 13515
rect 9496 13472 9548 13481
rect 9680 13515 9732 13524
rect 9680 13481 9689 13515
rect 9689 13481 9723 13515
rect 9723 13481 9732 13515
rect 9680 13472 9732 13481
rect 10508 13472 10560 13524
rect 13176 13472 13228 13524
rect 14556 13472 14608 13524
rect 15476 13472 15528 13524
rect 16120 13515 16172 13524
rect 16120 13481 16129 13515
rect 16129 13481 16163 13515
rect 16163 13481 16172 13515
rect 16120 13472 16172 13481
rect 16488 13515 16540 13524
rect 16488 13481 16497 13515
rect 16497 13481 16531 13515
rect 16531 13481 16540 13515
rect 16488 13472 16540 13481
rect 17040 13515 17092 13524
rect 17040 13481 17049 13515
rect 17049 13481 17083 13515
rect 17083 13481 17092 13515
rect 17040 13472 17092 13481
rect 21088 13515 21140 13524
rect 21088 13481 21097 13515
rect 21097 13481 21131 13515
rect 21131 13481 21140 13515
rect 21088 13472 21140 13481
rect 1768 13336 1820 13388
rect 1492 13268 1544 13320
rect 2320 13336 2372 13388
rect 3792 13336 3844 13388
rect 4160 13336 4212 13388
rect 4344 13379 4396 13388
rect 4344 13345 4378 13379
rect 4378 13345 4396 13379
rect 4344 13336 4396 13345
rect 3056 13243 3108 13252
rect 3056 13209 3065 13243
rect 3065 13209 3099 13243
rect 3099 13209 3108 13243
rect 3056 13200 3108 13209
rect 3976 13268 4028 13320
rect 6184 13336 6236 13388
rect 4344 13132 4396 13184
rect 6184 13132 6236 13184
rect 6552 13311 6604 13320
rect 6552 13277 6561 13311
rect 6561 13277 6595 13311
rect 6595 13277 6604 13311
rect 7748 13404 7800 13456
rect 8484 13404 8536 13456
rect 8208 13336 8260 13388
rect 6552 13268 6604 13277
rect 7564 13132 7616 13184
rect 8300 13175 8352 13184
rect 8300 13141 8309 13175
rect 8309 13141 8343 13175
rect 8343 13141 8352 13175
rect 9864 13404 9916 13456
rect 10324 13404 10376 13456
rect 13728 13404 13780 13456
rect 14004 13447 14056 13456
rect 14004 13413 14013 13447
rect 14013 13413 14047 13447
rect 14047 13413 14056 13447
rect 14004 13404 14056 13413
rect 14096 13404 14148 13456
rect 14280 13404 14332 13456
rect 11612 13336 11664 13388
rect 11796 13379 11848 13388
rect 11796 13345 11830 13379
rect 11830 13345 11848 13379
rect 11796 13336 11848 13345
rect 9036 13268 9088 13320
rect 10140 13268 10192 13320
rect 10600 13268 10652 13320
rect 14832 13404 14884 13456
rect 14648 13336 14700 13388
rect 15936 13404 15988 13456
rect 15108 13336 15160 13388
rect 18052 13336 18104 13388
rect 18788 13336 18840 13388
rect 14832 13311 14884 13320
rect 9864 13200 9916 13252
rect 10416 13200 10468 13252
rect 10876 13200 10928 13252
rect 14832 13277 14841 13311
rect 14841 13277 14875 13311
rect 14875 13277 14884 13311
rect 14832 13268 14884 13277
rect 14924 13311 14976 13320
rect 14924 13277 14933 13311
rect 14933 13277 14967 13311
rect 14967 13277 14976 13311
rect 14924 13268 14976 13277
rect 15292 13268 15344 13320
rect 12716 13200 12768 13252
rect 16028 13268 16080 13320
rect 16396 13268 16448 13320
rect 8300 13132 8352 13141
rect 9036 13132 9088 13184
rect 9312 13175 9364 13184
rect 9312 13141 9321 13175
rect 9321 13141 9355 13175
rect 9355 13141 9364 13175
rect 9312 13132 9364 13141
rect 12808 13132 12860 13184
rect 16212 13200 16264 13252
rect 17684 13268 17736 13320
rect 18604 13268 18656 13320
rect 19432 13268 19484 13320
rect 18880 13200 18932 13252
rect 13636 13132 13688 13184
rect 13728 13132 13780 13184
rect 14188 13132 14240 13184
rect 19892 13132 19944 13184
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 4575 13030 4627 13082
rect 4639 13030 4691 13082
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 18308 13030 18360 13082
rect 18372 13030 18424 13082
rect 18436 13030 18488 13082
rect 18500 13030 18552 13082
rect 3240 12971 3292 12980
rect 3240 12937 3249 12971
rect 3249 12937 3283 12971
rect 3283 12937 3292 12971
rect 3240 12928 3292 12937
rect 3792 12971 3844 12980
rect 3792 12937 3801 12971
rect 3801 12937 3835 12971
rect 3835 12937 3844 12971
rect 3792 12928 3844 12937
rect 4804 12971 4856 12980
rect 4804 12937 4813 12971
rect 4813 12937 4847 12971
rect 4847 12937 4856 12971
rect 4804 12928 4856 12937
rect 5632 12928 5684 12980
rect 6000 12928 6052 12980
rect 7104 12928 7156 12980
rect 8576 12928 8628 12980
rect 9128 12928 9180 12980
rect 11796 12971 11848 12980
rect 4620 12860 4672 12912
rect 5080 12860 5132 12912
rect 3516 12792 3568 12844
rect 4252 12792 4304 12844
rect 5356 12835 5408 12844
rect 1860 12767 1912 12776
rect 1860 12733 1869 12767
rect 1869 12733 1903 12767
rect 1903 12733 1912 12767
rect 1860 12724 1912 12733
rect 2596 12724 2648 12776
rect 5356 12801 5365 12835
rect 5365 12801 5399 12835
rect 5399 12801 5408 12835
rect 5356 12792 5408 12801
rect 5632 12792 5684 12844
rect 6368 12792 6420 12844
rect 6552 12835 6604 12844
rect 6552 12801 6561 12835
rect 6561 12801 6595 12835
rect 6595 12801 6604 12835
rect 6552 12792 6604 12801
rect 7380 12835 7432 12844
rect 7380 12801 7389 12835
rect 7389 12801 7423 12835
rect 7423 12801 7432 12835
rect 7380 12792 7432 12801
rect 8668 12792 8720 12844
rect 10140 12860 10192 12912
rect 9128 12835 9180 12844
rect 9128 12801 9137 12835
rect 9137 12801 9171 12835
rect 9171 12801 9180 12835
rect 9128 12792 9180 12801
rect 9496 12792 9548 12844
rect 11796 12937 11805 12971
rect 11805 12937 11839 12971
rect 11839 12937 11848 12971
rect 11796 12928 11848 12937
rect 12440 12928 12492 12980
rect 14648 12971 14700 12980
rect 13912 12860 13964 12912
rect 14648 12937 14657 12971
rect 14657 12937 14691 12971
rect 14691 12937 14700 12971
rect 14648 12928 14700 12937
rect 14832 12928 14884 12980
rect 15384 12928 15436 12980
rect 17684 12928 17736 12980
rect 18052 12928 18104 12980
rect 20996 12971 21048 12980
rect 20996 12937 21005 12971
rect 21005 12937 21039 12971
rect 21039 12937 21048 12971
rect 20996 12928 21048 12937
rect 13636 12792 13688 12844
rect 14004 12792 14056 12844
rect 14556 12860 14608 12912
rect 19432 12903 19484 12912
rect 19432 12869 19441 12903
rect 19441 12869 19475 12903
rect 19475 12869 19484 12903
rect 19432 12860 19484 12869
rect 16028 12792 16080 12844
rect 2504 12656 2556 12708
rect 3516 12656 3568 12708
rect 4160 12631 4212 12640
rect 4160 12597 4169 12631
rect 4169 12597 4203 12631
rect 4203 12597 4212 12631
rect 4160 12588 4212 12597
rect 4804 12724 4856 12776
rect 4988 12724 5040 12776
rect 5080 12724 5132 12776
rect 5908 12724 5960 12776
rect 4988 12588 5040 12640
rect 5540 12588 5592 12640
rect 5724 12631 5776 12640
rect 5724 12597 5733 12631
rect 5733 12597 5767 12631
rect 5767 12597 5776 12631
rect 8484 12724 8536 12776
rect 9312 12724 9364 12776
rect 10048 12724 10100 12776
rect 10508 12724 10560 12776
rect 7380 12656 7432 12708
rect 14096 12724 14148 12776
rect 14556 12724 14608 12776
rect 17316 12724 17368 12776
rect 6276 12631 6328 12640
rect 5724 12588 5776 12597
rect 6276 12597 6285 12631
rect 6285 12597 6319 12631
rect 6319 12597 6328 12631
rect 6276 12588 6328 12597
rect 6552 12588 6604 12640
rect 6828 12588 6880 12640
rect 6920 12588 6972 12640
rect 7288 12631 7340 12640
rect 7288 12597 7297 12631
rect 7297 12597 7331 12631
rect 7331 12597 7340 12631
rect 7288 12588 7340 12597
rect 7564 12588 7616 12640
rect 8760 12588 8812 12640
rect 9128 12588 9180 12640
rect 10876 12656 10928 12708
rect 11428 12656 11480 12708
rect 11244 12588 11296 12640
rect 11888 12631 11940 12640
rect 11888 12597 11897 12631
rect 11897 12597 11931 12631
rect 11931 12597 11940 12631
rect 13912 12656 13964 12708
rect 15476 12656 15528 12708
rect 16672 12656 16724 12708
rect 16948 12656 17000 12708
rect 19892 12767 19944 12776
rect 19892 12733 19901 12767
rect 19901 12733 19935 12767
rect 19935 12733 19944 12767
rect 19892 12724 19944 12733
rect 20260 12724 20312 12776
rect 18696 12656 18748 12708
rect 19340 12656 19392 12708
rect 11888 12588 11940 12597
rect 12532 12588 12584 12640
rect 12900 12631 12952 12640
rect 12900 12597 12909 12631
rect 12909 12597 12943 12631
rect 12943 12597 12952 12631
rect 12900 12588 12952 12597
rect 13820 12588 13872 12640
rect 14004 12588 14056 12640
rect 15936 12588 15988 12640
rect 16764 12588 16816 12640
rect 7912 12486 7964 12538
rect 7976 12486 8028 12538
rect 8040 12486 8092 12538
rect 8104 12486 8156 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 15035 12486 15087 12538
rect 1676 12427 1728 12436
rect 1676 12393 1685 12427
rect 1685 12393 1719 12427
rect 1719 12393 1728 12427
rect 1676 12384 1728 12393
rect 1768 12384 1820 12436
rect 4160 12384 4212 12436
rect 4344 12384 4396 12436
rect 3976 12316 4028 12368
rect 1492 12291 1544 12300
rect 1492 12257 1501 12291
rect 1501 12257 1535 12291
rect 1535 12257 1544 12291
rect 1492 12248 1544 12257
rect 2228 12291 2280 12300
rect 2228 12257 2237 12291
rect 2237 12257 2271 12291
rect 2271 12257 2280 12291
rect 2228 12248 2280 12257
rect 4252 12248 4304 12300
rect 2504 12223 2556 12232
rect 2504 12189 2513 12223
rect 2513 12189 2547 12223
rect 2547 12189 2556 12223
rect 2504 12180 2556 12189
rect 3240 12223 3292 12232
rect 3240 12189 3249 12223
rect 3249 12189 3283 12223
rect 3283 12189 3292 12223
rect 3240 12180 3292 12189
rect 2688 12112 2740 12164
rect 3976 12044 4028 12096
rect 6184 12316 6236 12368
rect 7472 12384 7524 12436
rect 8484 12384 8536 12436
rect 8668 12384 8720 12436
rect 10048 12384 10100 12436
rect 11428 12427 11480 12436
rect 11428 12393 11437 12427
rect 11437 12393 11471 12427
rect 11471 12393 11480 12427
rect 11428 12384 11480 12393
rect 8300 12359 8352 12368
rect 8300 12325 8334 12359
rect 8334 12325 8352 12359
rect 8300 12316 8352 12325
rect 8944 12316 8996 12368
rect 9772 12316 9824 12368
rect 11888 12384 11940 12436
rect 12440 12384 12492 12436
rect 16764 12427 16816 12436
rect 16764 12393 16773 12427
rect 16773 12393 16807 12427
rect 16807 12393 16816 12427
rect 16764 12384 16816 12393
rect 16948 12427 17000 12436
rect 16948 12393 16957 12427
rect 16957 12393 16991 12427
rect 16991 12393 17000 12427
rect 16948 12384 17000 12393
rect 17132 12384 17184 12436
rect 17684 12384 17736 12436
rect 18788 12427 18840 12436
rect 18788 12393 18797 12427
rect 18797 12393 18831 12427
rect 18831 12393 18840 12427
rect 18788 12384 18840 12393
rect 19432 12384 19484 12436
rect 6092 12291 6144 12300
rect 6092 12257 6126 12291
rect 6126 12257 6144 12291
rect 6092 12248 6144 12257
rect 7472 12291 7524 12300
rect 7472 12257 7481 12291
rect 7481 12257 7515 12291
rect 7515 12257 7524 12291
rect 7472 12248 7524 12257
rect 9128 12248 9180 12300
rect 12532 12316 12584 12368
rect 12808 12316 12860 12368
rect 14188 12316 14240 12368
rect 15660 12316 15712 12368
rect 20260 12359 20312 12368
rect 11428 12248 11480 12300
rect 11704 12248 11756 12300
rect 13912 12248 13964 12300
rect 14280 12248 14332 12300
rect 17316 12291 17368 12300
rect 17316 12257 17325 12291
rect 17325 12257 17359 12291
rect 17359 12257 17368 12291
rect 17316 12248 17368 12257
rect 17592 12291 17644 12300
rect 17592 12257 17626 12291
rect 17626 12257 17644 12291
rect 17592 12248 17644 12257
rect 20260 12325 20269 12359
rect 20269 12325 20303 12359
rect 20303 12325 20312 12359
rect 20260 12316 20312 12325
rect 5080 12223 5132 12232
rect 5080 12189 5089 12223
rect 5089 12189 5123 12223
rect 5123 12189 5132 12223
rect 5816 12223 5868 12232
rect 5080 12180 5132 12189
rect 5816 12189 5825 12223
rect 5825 12189 5859 12223
rect 5859 12189 5868 12223
rect 5816 12180 5868 12189
rect 8024 12223 8076 12232
rect 8024 12189 8033 12223
rect 8033 12189 8067 12223
rect 8067 12189 8076 12223
rect 8024 12180 8076 12189
rect 9404 12180 9456 12232
rect 9864 12180 9916 12232
rect 10232 12180 10284 12232
rect 10600 12223 10652 12232
rect 10600 12189 10609 12223
rect 10609 12189 10643 12223
rect 10643 12189 10652 12223
rect 10600 12180 10652 12189
rect 10876 12180 10928 12232
rect 11152 12180 11204 12232
rect 11888 12180 11940 12232
rect 12532 12180 12584 12232
rect 14740 12180 14792 12232
rect 15292 12223 15344 12232
rect 15292 12189 15301 12223
rect 15301 12189 15335 12223
rect 15335 12189 15344 12223
rect 15292 12180 15344 12189
rect 16672 12180 16724 12232
rect 17132 12180 17184 12232
rect 4896 12044 4948 12096
rect 5356 12044 5408 12096
rect 5540 12044 5592 12096
rect 7196 12087 7248 12096
rect 7196 12053 7205 12087
rect 7205 12053 7239 12087
rect 7239 12053 7248 12087
rect 7196 12044 7248 12053
rect 7288 12044 7340 12096
rect 7840 12044 7892 12096
rect 8944 12044 8996 12096
rect 12440 12044 12492 12096
rect 14648 12112 14700 12164
rect 18696 12155 18748 12164
rect 18696 12121 18705 12155
rect 18705 12121 18739 12155
rect 18739 12121 18748 12155
rect 18696 12112 18748 12121
rect 13912 12044 13964 12096
rect 14832 12087 14884 12096
rect 14832 12053 14841 12087
rect 14841 12053 14875 12087
rect 14875 12053 14884 12087
rect 14832 12044 14884 12053
rect 16028 12044 16080 12096
rect 16212 12044 16264 12096
rect 16580 12044 16632 12096
rect 16764 12044 16816 12096
rect 17040 12044 17092 12096
rect 20076 12044 20128 12096
rect 22008 12019 22060 12028
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 4575 11942 4627 11994
rect 4639 11942 4691 11994
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 18308 11942 18360 11994
rect 18372 11942 18424 11994
rect 18436 11942 18488 11994
rect 18500 11942 18552 11994
rect 22008 11985 22017 12019
rect 22017 11985 22051 12019
rect 22051 11985 22060 12019
rect 22008 11976 22060 11985
rect 1860 11840 1912 11892
rect 2504 11840 2556 11892
rect 3148 11883 3200 11892
rect 3148 11849 3157 11883
rect 3157 11849 3191 11883
rect 3191 11849 3200 11883
rect 3148 11840 3200 11849
rect 3240 11840 3292 11892
rect 4252 11883 4304 11892
rect 4252 11849 4261 11883
rect 4261 11849 4295 11883
rect 4295 11849 4304 11883
rect 4252 11840 4304 11849
rect 3884 11772 3936 11824
rect 6368 11840 6420 11892
rect 6920 11883 6972 11892
rect 6920 11849 6929 11883
rect 6929 11849 6963 11883
rect 6963 11849 6972 11883
rect 6920 11840 6972 11849
rect 7380 11840 7432 11892
rect 8760 11883 8812 11892
rect 8760 11849 8769 11883
rect 8769 11849 8803 11883
rect 8803 11849 8812 11883
rect 8760 11840 8812 11849
rect 10140 11883 10192 11892
rect 10140 11849 10149 11883
rect 10149 11849 10183 11883
rect 10183 11849 10192 11883
rect 10140 11840 10192 11849
rect 6460 11772 6512 11824
rect 7196 11772 7248 11824
rect 3700 11704 3752 11756
rect 6920 11704 6972 11756
rect 2780 11636 2832 11688
rect 4344 11636 4396 11688
rect 4988 11636 5040 11688
rect 2136 11568 2188 11620
rect 2688 11568 2740 11620
rect 6368 11636 6420 11688
rect 7564 11747 7616 11756
rect 7564 11713 7573 11747
rect 7573 11713 7607 11747
rect 7607 11713 7616 11747
rect 7564 11704 7616 11713
rect 7288 11636 7340 11688
rect 8300 11704 8352 11756
rect 5816 11568 5868 11620
rect 7840 11568 7892 11620
rect 8760 11568 8812 11620
rect 3792 11543 3844 11552
rect 3792 11509 3801 11543
rect 3801 11509 3835 11543
rect 3835 11509 3844 11543
rect 3792 11500 3844 11509
rect 4160 11500 4212 11552
rect 4620 11543 4672 11552
rect 4620 11509 4629 11543
rect 4629 11509 4663 11543
rect 4663 11509 4672 11543
rect 4620 11500 4672 11509
rect 4804 11500 4856 11552
rect 5080 11543 5132 11552
rect 5080 11509 5089 11543
rect 5089 11509 5123 11543
rect 5123 11509 5132 11543
rect 5080 11500 5132 11509
rect 6184 11500 6236 11552
rect 6644 11543 6696 11552
rect 6644 11509 6653 11543
rect 6653 11509 6687 11543
rect 6687 11509 6696 11543
rect 6644 11500 6696 11509
rect 7472 11543 7524 11552
rect 7472 11509 7481 11543
rect 7481 11509 7515 11543
rect 7515 11509 7524 11543
rect 7472 11500 7524 11509
rect 8208 11500 8260 11552
rect 8300 11543 8352 11552
rect 8300 11509 8309 11543
rect 8309 11509 8343 11543
rect 8343 11509 8352 11543
rect 10048 11772 10100 11824
rect 9496 11704 9548 11756
rect 9772 11704 9824 11756
rect 10508 11840 10560 11892
rect 10692 11840 10744 11892
rect 11060 11840 11112 11892
rect 11244 11840 11296 11892
rect 13636 11840 13688 11892
rect 15200 11840 15252 11892
rect 15660 11840 15712 11892
rect 17592 11883 17644 11892
rect 11428 11772 11480 11824
rect 12532 11772 12584 11824
rect 12440 11704 12492 11756
rect 14832 11704 14884 11756
rect 15476 11704 15528 11756
rect 15660 11704 15712 11756
rect 17592 11849 17601 11883
rect 17601 11849 17635 11883
rect 17635 11849 17644 11883
rect 17592 11840 17644 11849
rect 19340 11840 19392 11892
rect 20996 11883 21048 11892
rect 20996 11849 21005 11883
rect 21005 11849 21039 11883
rect 21039 11849 21048 11883
rect 20996 11840 21048 11849
rect 21364 11883 21416 11892
rect 21364 11849 21373 11883
rect 21373 11849 21407 11883
rect 21407 11849 21416 11883
rect 21364 11840 21416 11849
rect 18972 11815 19024 11824
rect 18972 11781 18981 11815
rect 18981 11781 19015 11815
rect 19015 11781 19024 11815
rect 18972 11772 19024 11781
rect 19432 11772 19484 11824
rect 18696 11747 18748 11756
rect 18696 11713 18705 11747
rect 18705 11713 18739 11747
rect 18739 11713 18748 11747
rect 18696 11704 18748 11713
rect 11152 11568 11204 11620
rect 11796 11611 11848 11620
rect 11796 11577 11805 11611
rect 11805 11577 11839 11611
rect 11839 11577 11848 11611
rect 11796 11568 11848 11577
rect 9680 11543 9732 11552
rect 8300 11500 8352 11509
rect 9680 11509 9689 11543
rect 9689 11509 9723 11543
rect 9723 11509 9732 11543
rect 9680 11500 9732 11509
rect 10048 11500 10100 11552
rect 10324 11500 10376 11552
rect 10876 11500 10928 11552
rect 11428 11500 11480 11552
rect 11980 11636 12032 11688
rect 13360 11636 13412 11688
rect 15292 11636 15344 11688
rect 20536 11636 20588 11688
rect 21180 11679 21232 11688
rect 21180 11645 21189 11679
rect 21189 11645 21223 11679
rect 21223 11645 21232 11679
rect 21180 11636 21232 11645
rect 12440 11568 12492 11620
rect 13544 11568 13596 11620
rect 13912 11568 13964 11620
rect 17500 11568 17552 11620
rect 20260 11568 20312 11620
rect 12808 11543 12860 11552
rect 12808 11509 12817 11543
rect 12817 11509 12851 11543
rect 12851 11509 12860 11543
rect 12808 11500 12860 11509
rect 14188 11500 14240 11552
rect 15200 11500 15252 11552
rect 15752 11543 15804 11552
rect 15752 11509 15761 11543
rect 15761 11509 15795 11543
rect 15795 11509 15804 11543
rect 15752 11500 15804 11509
rect 16948 11500 17000 11552
rect 17776 11543 17828 11552
rect 17776 11509 17785 11543
rect 17785 11509 17819 11543
rect 17819 11509 17828 11543
rect 17776 11500 17828 11509
rect 7912 11398 7964 11450
rect 7976 11398 8028 11450
rect 8040 11398 8092 11450
rect 8104 11398 8156 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 15035 11398 15087 11450
rect 1584 11339 1636 11348
rect 1584 11305 1593 11339
rect 1593 11305 1627 11339
rect 1627 11305 1636 11339
rect 1584 11296 1636 11305
rect 2688 11296 2740 11348
rect 4620 11296 4672 11348
rect 4988 11339 5040 11348
rect 4988 11305 4997 11339
rect 4997 11305 5031 11339
rect 5031 11305 5040 11339
rect 4988 11296 5040 11305
rect 6460 11296 6512 11348
rect 6644 11296 6696 11348
rect 3424 11228 3476 11280
rect 1676 11160 1728 11212
rect 1860 11160 1912 11212
rect 2872 11160 2924 11212
rect 3700 11160 3752 11212
rect 3240 11092 3292 11144
rect 3976 11092 4028 11144
rect 4712 11160 4764 11212
rect 5540 11160 5592 11212
rect 4988 11092 5040 11144
rect 3148 11024 3200 11076
rect 6092 11092 6144 11144
rect 6000 11024 6052 11076
rect 6092 10999 6144 11008
rect 6092 10965 6101 10999
rect 6101 10965 6135 10999
rect 6135 10965 6144 10999
rect 6092 10956 6144 10965
rect 7472 11296 7524 11348
rect 8208 11296 8260 11348
rect 8944 11296 8996 11348
rect 9956 11296 10008 11348
rect 10600 11296 10652 11348
rect 12532 11296 12584 11348
rect 12808 11296 12860 11348
rect 14096 11296 14148 11348
rect 7472 11160 7524 11212
rect 10140 11228 10192 11280
rect 10508 11228 10560 11280
rect 9772 11203 9824 11212
rect 7564 11135 7616 11144
rect 7564 11101 7573 11135
rect 7573 11101 7607 11135
rect 7607 11101 7616 11135
rect 7564 11092 7616 11101
rect 8668 11092 8720 11144
rect 7380 11024 7432 11076
rect 9772 11169 9781 11203
rect 9781 11169 9815 11203
rect 9815 11169 9824 11203
rect 9772 11160 9824 11169
rect 9496 11135 9548 11144
rect 9496 11101 9505 11135
rect 9505 11101 9539 11135
rect 9539 11101 9548 11135
rect 9496 11092 9548 11101
rect 9680 11092 9732 11144
rect 12256 11160 12308 11212
rect 12440 11160 12492 11212
rect 13544 11228 13596 11280
rect 14004 11228 14056 11280
rect 14648 11228 14700 11280
rect 15752 11228 15804 11280
rect 18144 11228 18196 11280
rect 11152 11092 11204 11144
rect 13820 11160 13872 11212
rect 14740 11203 14792 11212
rect 14740 11169 14749 11203
rect 14749 11169 14783 11203
rect 14783 11169 14792 11203
rect 14740 11160 14792 11169
rect 15108 11160 15160 11212
rect 13360 11092 13412 11144
rect 14188 11135 14240 11144
rect 14188 11101 14197 11135
rect 14197 11101 14231 11135
rect 14231 11101 14240 11135
rect 17132 11160 17184 11212
rect 17316 11203 17368 11212
rect 17316 11169 17325 11203
rect 17325 11169 17359 11203
rect 17359 11169 17368 11203
rect 17316 11160 17368 11169
rect 18236 11203 18288 11212
rect 18236 11169 18245 11203
rect 18245 11169 18279 11203
rect 18279 11169 18288 11203
rect 18236 11160 18288 11169
rect 14188 11092 14240 11101
rect 15936 11135 15988 11144
rect 15936 11101 15945 11135
rect 15945 11101 15979 11135
rect 15979 11101 15988 11135
rect 15936 11092 15988 11101
rect 16120 11092 16172 11144
rect 15108 11024 15160 11076
rect 15292 11067 15344 11076
rect 15292 11033 15301 11067
rect 15301 11033 15335 11067
rect 15335 11033 15344 11067
rect 15292 11024 15344 11033
rect 16212 11024 16264 11076
rect 16948 11067 17000 11076
rect 16948 11033 16957 11067
rect 16957 11033 16991 11067
rect 16991 11033 17000 11067
rect 16948 11024 17000 11033
rect 7656 10956 7708 11008
rect 7932 10956 7984 11008
rect 8300 10956 8352 11008
rect 8668 10956 8720 11008
rect 9220 10999 9272 11008
rect 9220 10965 9229 10999
rect 9229 10965 9263 10999
rect 9263 10965 9272 10999
rect 9220 10956 9272 10965
rect 16764 10956 16816 11008
rect 18604 11092 18656 11144
rect 19156 11135 19208 11144
rect 19156 11101 19165 11135
rect 19165 11101 19199 11135
rect 19199 11101 19208 11135
rect 19156 11092 19208 11101
rect 20444 11160 20496 11212
rect 17500 11024 17552 11076
rect 18604 10956 18656 11008
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 4575 10854 4627 10906
rect 4639 10854 4691 10906
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 18308 10854 18360 10906
rect 18372 10854 18424 10906
rect 18436 10854 18488 10906
rect 18500 10854 18552 10906
rect 2228 10752 2280 10804
rect 3700 10795 3752 10804
rect 3700 10761 3709 10795
rect 3709 10761 3743 10795
rect 3743 10761 3752 10795
rect 3700 10752 3752 10761
rect 3792 10752 3844 10804
rect 4804 10752 4856 10804
rect 5080 10752 5132 10804
rect 5632 10752 5684 10804
rect 6276 10752 6328 10804
rect 7012 10752 7064 10804
rect 8668 10752 8720 10804
rect 9680 10752 9732 10804
rect 10968 10752 11020 10804
rect 11152 10752 11204 10804
rect 2136 10659 2188 10668
rect 2136 10625 2145 10659
rect 2145 10625 2179 10659
rect 2179 10625 2188 10659
rect 2136 10616 2188 10625
rect 4344 10659 4396 10668
rect 4344 10625 4353 10659
rect 4353 10625 4387 10659
rect 4387 10625 4396 10659
rect 4344 10616 4396 10625
rect 4988 10616 5040 10668
rect 5448 10616 5500 10668
rect 3884 10548 3936 10600
rect 5724 10616 5776 10668
rect 6092 10616 6144 10668
rect 6368 10659 6420 10668
rect 6368 10625 6377 10659
rect 6377 10625 6411 10659
rect 6411 10625 6420 10659
rect 6368 10616 6420 10625
rect 9312 10684 9364 10736
rect 8944 10616 8996 10668
rect 9496 10616 9548 10668
rect 9588 10616 9640 10668
rect 12532 10752 12584 10804
rect 13176 10752 13228 10804
rect 11796 10684 11848 10736
rect 12440 10684 12492 10736
rect 14648 10684 14700 10736
rect 17316 10752 17368 10804
rect 18144 10752 18196 10804
rect 15936 10684 15988 10736
rect 19156 10684 19208 10736
rect 5816 10548 5868 10600
rect 7472 10548 7524 10600
rect 7932 10548 7984 10600
rect 8208 10548 8260 10600
rect 9772 10548 9824 10600
rect 9864 10548 9916 10600
rect 11060 10548 11112 10600
rect 11336 10548 11388 10600
rect 12440 10548 12492 10600
rect 13544 10616 13596 10668
rect 14188 10616 14240 10668
rect 15200 10548 15252 10600
rect 2688 10480 2740 10532
rect 4988 10480 5040 10532
rect 1860 10455 1912 10464
rect 1860 10421 1869 10455
rect 1869 10421 1903 10455
rect 1903 10421 1912 10455
rect 1860 10412 1912 10421
rect 2044 10412 2096 10464
rect 5080 10455 5132 10464
rect 5080 10421 5089 10455
rect 5089 10421 5123 10455
rect 5123 10421 5132 10455
rect 5080 10412 5132 10421
rect 6000 10480 6052 10532
rect 6184 10480 6236 10532
rect 8944 10480 8996 10532
rect 10048 10480 10100 10532
rect 10324 10480 10376 10532
rect 6828 10412 6880 10464
rect 7196 10412 7248 10464
rect 9680 10412 9732 10464
rect 11060 10412 11112 10464
rect 11888 10412 11940 10464
rect 11980 10412 12032 10464
rect 12532 10412 12584 10464
rect 13452 10480 13504 10532
rect 15292 10480 15344 10532
rect 15936 10591 15988 10600
rect 15936 10557 15945 10591
rect 15945 10557 15979 10591
rect 15979 10557 15988 10591
rect 15936 10548 15988 10557
rect 17868 10616 17920 10668
rect 18696 10659 18748 10668
rect 16212 10591 16264 10600
rect 16212 10557 16246 10591
rect 16246 10557 16264 10591
rect 16212 10548 16264 10557
rect 16764 10548 16816 10600
rect 18696 10625 18705 10659
rect 18705 10625 18739 10659
rect 18739 10625 18748 10659
rect 18696 10616 18748 10625
rect 18788 10616 18840 10668
rect 19892 10659 19944 10668
rect 19892 10625 19901 10659
rect 19901 10625 19935 10659
rect 19935 10625 19944 10659
rect 19892 10616 19944 10625
rect 20444 10659 20496 10668
rect 20444 10625 20453 10659
rect 20453 10625 20487 10659
rect 20487 10625 20496 10659
rect 20444 10616 20496 10625
rect 18144 10480 18196 10532
rect 19432 10548 19484 10600
rect 21180 10616 21232 10668
rect 20352 10480 20404 10532
rect 13636 10412 13688 10464
rect 14004 10455 14056 10464
rect 14004 10421 14013 10455
rect 14013 10421 14047 10455
rect 14047 10421 14056 10455
rect 14004 10412 14056 10421
rect 14188 10412 14240 10464
rect 14740 10412 14792 10464
rect 15752 10412 15804 10464
rect 16856 10412 16908 10464
rect 17500 10412 17552 10464
rect 19708 10455 19760 10464
rect 19708 10421 19717 10455
rect 19717 10421 19751 10455
rect 19751 10421 19760 10455
rect 19708 10412 19760 10421
rect 20444 10412 20496 10464
rect 7912 10310 7964 10362
rect 7976 10310 8028 10362
rect 8040 10310 8092 10362
rect 8104 10310 8156 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 15035 10310 15087 10362
rect 2044 10251 2096 10260
rect 2044 10217 2053 10251
rect 2053 10217 2087 10251
rect 2087 10217 2096 10251
rect 2044 10208 2096 10217
rect 3148 10251 3200 10260
rect 3148 10217 3157 10251
rect 3157 10217 3191 10251
rect 3191 10217 3200 10251
rect 3148 10208 3200 10217
rect 4160 10208 4212 10260
rect 4896 10208 4948 10260
rect 5632 10208 5684 10260
rect 6092 10251 6144 10260
rect 6092 10217 6101 10251
rect 6101 10217 6135 10251
rect 6135 10217 6144 10251
rect 6092 10208 6144 10217
rect 8300 10208 8352 10260
rect 8484 10208 8536 10260
rect 11336 10251 11388 10260
rect 6460 10140 6512 10192
rect 7012 10140 7064 10192
rect 7196 10140 7248 10192
rect 2412 10115 2464 10124
rect 2412 10081 2421 10115
rect 2421 10081 2455 10115
rect 2455 10081 2464 10115
rect 2412 10072 2464 10081
rect 3332 10072 3384 10124
rect 3792 10072 3844 10124
rect 5540 10072 5592 10124
rect 6736 10072 6788 10124
rect 6920 10072 6972 10124
rect 7472 10115 7524 10124
rect 7472 10081 7481 10115
rect 7481 10081 7515 10115
rect 7515 10081 7524 10115
rect 7472 10072 7524 10081
rect 7656 10072 7708 10124
rect 8852 10140 8904 10192
rect 8760 10072 8812 10124
rect 10140 10140 10192 10192
rect 11336 10217 11345 10251
rect 11345 10217 11379 10251
rect 11379 10217 11388 10251
rect 11336 10208 11388 10217
rect 11520 10208 11572 10260
rect 11980 10208 12032 10260
rect 12072 10208 12124 10260
rect 12348 10208 12400 10260
rect 11704 10140 11756 10192
rect 13820 10208 13872 10260
rect 14188 10208 14240 10260
rect 14648 10251 14700 10260
rect 14648 10217 14657 10251
rect 14657 10217 14691 10251
rect 14691 10217 14700 10251
rect 14648 10208 14700 10217
rect 15292 10251 15344 10260
rect 15292 10217 15301 10251
rect 15301 10217 15335 10251
rect 15335 10217 15344 10251
rect 15292 10208 15344 10217
rect 16120 10251 16172 10260
rect 2504 10047 2556 10056
rect 2504 10013 2513 10047
rect 2513 10013 2547 10047
rect 2547 10013 2556 10047
rect 2504 10004 2556 10013
rect 2872 10004 2924 10056
rect 4804 10047 4856 10056
rect 4804 10013 4813 10047
rect 4813 10013 4847 10047
rect 4847 10013 4856 10047
rect 4804 10004 4856 10013
rect 5448 10004 5500 10056
rect 5908 10047 5960 10056
rect 5908 10013 5917 10047
rect 5917 10013 5951 10047
rect 5951 10013 5960 10047
rect 5908 10004 5960 10013
rect 6828 10047 6880 10056
rect 6828 10013 6837 10047
rect 6837 10013 6871 10047
rect 6871 10013 6880 10047
rect 6828 10004 6880 10013
rect 3332 9936 3384 9988
rect 3516 9936 3568 9988
rect 7748 10047 7800 10056
rect 7748 10013 7757 10047
rect 7757 10013 7791 10047
rect 7791 10013 7800 10047
rect 7748 10004 7800 10013
rect 8208 10004 8260 10056
rect 9496 10072 9548 10124
rect 11888 10072 11940 10124
rect 8300 9936 8352 9988
rect 9220 10047 9272 10056
rect 9220 10013 9229 10047
rect 9229 10013 9263 10047
rect 9263 10013 9272 10047
rect 9220 10004 9272 10013
rect 9588 10004 9640 10056
rect 9312 9936 9364 9988
rect 11980 10004 12032 10056
rect 15752 10183 15804 10192
rect 15752 10149 15761 10183
rect 15761 10149 15795 10183
rect 15795 10149 15804 10183
rect 15752 10140 15804 10149
rect 16120 10217 16129 10251
rect 16129 10217 16163 10251
rect 16163 10217 16172 10251
rect 16120 10208 16172 10217
rect 16488 10251 16540 10260
rect 16488 10217 16497 10251
rect 16497 10217 16531 10251
rect 16531 10217 16540 10251
rect 16488 10208 16540 10217
rect 18420 10208 18472 10260
rect 18696 10208 18748 10260
rect 16028 10140 16080 10192
rect 12348 10072 12400 10124
rect 13268 10072 13320 10124
rect 14188 10072 14240 10124
rect 15476 10072 15528 10124
rect 17684 10183 17736 10192
rect 17684 10149 17696 10183
rect 17696 10149 17736 10183
rect 16396 10072 16448 10124
rect 17684 10140 17736 10149
rect 18788 10072 18840 10124
rect 19892 10072 19944 10124
rect 20352 10072 20404 10124
rect 13544 10004 13596 10056
rect 13636 9936 13688 9988
rect 14832 9936 14884 9988
rect 15016 9936 15068 9988
rect 15476 9936 15528 9988
rect 16856 10004 16908 10056
rect 3700 9868 3752 9920
rect 7196 9868 7248 9920
rect 8208 9868 8260 9920
rect 9864 9868 9916 9920
rect 11888 9868 11940 9920
rect 12072 9868 12124 9920
rect 15752 9868 15804 9920
rect 15936 9868 15988 9920
rect 16212 9868 16264 9920
rect 16764 9868 16816 9920
rect 16948 9911 17000 9920
rect 16948 9877 16957 9911
rect 16957 9877 16991 9911
rect 16991 9877 17000 9911
rect 16948 9868 17000 9877
rect 18420 10004 18472 10056
rect 18972 10004 19024 10056
rect 18604 9868 18656 9920
rect 19156 9911 19208 9920
rect 19156 9877 19165 9911
rect 19165 9877 19199 9911
rect 19199 9877 19208 9911
rect 19156 9868 19208 9877
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 4575 9766 4627 9818
rect 4639 9766 4691 9818
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 18308 9766 18360 9818
rect 18372 9766 18424 9818
rect 18436 9766 18488 9818
rect 18500 9766 18552 9818
rect 1860 9664 1912 9716
rect 2412 9707 2464 9716
rect 2412 9673 2421 9707
rect 2421 9673 2455 9707
rect 2455 9673 2464 9707
rect 2412 9664 2464 9673
rect 2964 9664 3016 9716
rect 3516 9664 3568 9716
rect 4804 9664 4856 9716
rect 8576 9664 8628 9716
rect 8760 9664 8812 9716
rect 9496 9664 9548 9716
rect 10140 9707 10192 9716
rect 4712 9596 4764 9648
rect 5540 9596 5592 9648
rect 10140 9673 10149 9707
rect 10149 9673 10183 9707
rect 10183 9673 10192 9707
rect 10140 9664 10192 9673
rect 12164 9664 12216 9716
rect 12532 9707 12584 9716
rect 12532 9673 12541 9707
rect 12541 9673 12575 9707
rect 12575 9673 12584 9707
rect 12532 9664 12584 9673
rect 13360 9664 13412 9716
rect 12348 9596 12400 9648
rect 2872 9528 2924 9580
rect 3056 9571 3108 9580
rect 3056 9537 3065 9571
rect 3065 9537 3099 9571
rect 3099 9537 3108 9571
rect 3056 9528 3108 9537
rect 2688 9460 2740 9512
rect 3148 9460 3200 9512
rect 4252 9528 4304 9580
rect 4804 9571 4856 9580
rect 4804 9537 4813 9571
rect 4813 9537 4847 9571
rect 4847 9537 4856 9571
rect 4804 9528 4856 9537
rect 8760 9571 8812 9580
rect 5448 9460 5500 9512
rect 5540 9460 5592 9512
rect 6460 9460 6512 9512
rect 8760 9537 8769 9571
rect 8769 9537 8803 9571
rect 8803 9537 8812 9571
rect 8760 9528 8812 9537
rect 10048 9528 10100 9580
rect 12624 9528 12676 9580
rect 13728 9596 13780 9648
rect 14740 9596 14792 9648
rect 13176 9571 13228 9580
rect 13176 9537 13185 9571
rect 13185 9537 13219 9571
rect 13219 9537 13228 9571
rect 13176 9528 13228 9537
rect 13544 9528 13596 9580
rect 7748 9460 7800 9512
rect 9588 9460 9640 9512
rect 1308 9324 1360 9376
rect 6644 9392 6696 9444
rect 7932 9392 7984 9444
rect 1584 9324 1636 9376
rect 2136 9324 2188 9376
rect 3332 9324 3384 9376
rect 3700 9324 3752 9376
rect 4620 9367 4672 9376
rect 4620 9333 4629 9367
rect 4629 9333 4663 9367
rect 4663 9333 4672 9367
rect 4620 9324 4672 9333
rect 4712 9367 4764 9376
rect 4712 9333 4721 9367
rect 4721 9333 4755 9367
rect 4755 9333 4764 9367
rect 4712 9324 4764 9333
rect 5080 9324 5132 9376
rect 5172 9324 5224 9376
rect 5816 9324 5868 9376
rect 6092 9324 6144 9376
rect 6276 9367 6328 9376
rect 6276 9333 6285 9367
rect 6285 9333 6319 9367
rect 6319 9333 6328 9367
rect 6276 9324 6328 9333
rect 8392 9367 8444 9376
rect 8392 9333 8401 9367
rect 8401 9333 8435 9367
rect 8435 9333 8444 9367
rect 8576 9367 8628 9376
rect 8392 9324 8444 9333
rect 8576 9333 8585 9367
rect 8585 9333 8619 9367
rect 8619 9333 8628 9367
rect 8576 9324 8628 9333
rect 8760 9324 8812 9376
rect 8944 9324 8996 9376
rect 10048 9392 10100 9444
rect 10508 9392 10560 9444
rect 11980 9460 12032 9512
rect 11336 9392 11388 9444
rect 11704 9392 11756 9444
rect 12164 9460 12216 9512
rect 13636 9460 13688 9512
rect 13912 9528 13964 9580
rect 15016 9528 15068 9580
rect 14096 9460 14148 9512
rect 16396 9664 16448 9716
rect 16672 9596 16724 9648
rect 19616 9664 19668 9716
rect 20444 9707 20496 9716
rect 20444 9673 20453 9707
rect 20453 9673 20487 9707
rect 20487 9673 20496 9707
rect 20444 9664 20496 9673
rect 20812 9664 20864 9716
rect 21456 9664 21508 9716
rect 20352 9639 20404 9648
rect 15200 9528 15252 9580
rect 15476 9571 15528 9580
rect 15476 9537 15485 9571
rect 15485 9537 15519 9571
rect 15519 9537 15528 9571
rect 15476 9528 15528 9537
rect 15752 9528 15804 9580
rect 16212 9528 16264 9580
rect 16580 9528 16632 9580
rect 16764 9528 16816 9580
rect 16856 9528 16908 9580
rect 20352 9605 20361 9639
rect 20361 9605 20395 9639
rect 20395 9605 20404 9639
rect 20352 9596 20404 9605
rect 21640 9596 21692 9648
rect 21824 9596 21876 9648
rect 12716 9324 12768 9376
rect 12900 9367 12952 9376
rect 12900 9333 12909 9367
rect 12909 9333 12943 9367
rect 12943 9333 12952 9367
rect 12900 9324 12952 9333
rect 13636 9324 13688 9376
rect 15844 9324 15896 9376
rect 16212 9324 16264 9376
rect 18604 9460 18656 9512
rect 18972 9503 19024 9512
rect 18972 9469 18981 9503
rect 18981 9469 19015 9503
rect 19015 9469 19024 9503
rect 18972 9460 19024 9469
rect 20168 9528 20220 9580
rect 20904 9460 20956 9512
rect 21916 9460 21968 9512
rect 16396 9392 16448 9444
rect 16580 9324 16632 9376
rect 16948 9367 17000 9376
rect 16948 9333 16957 9367
rect 16957 9333 16991 9367
rect 16991 9333 17000 9367
rect 17408 9367 17460 9376
rect 16948 9324 17000 9333
rect 17408 9333 17417 9367
rect 17417 9333 17451 9367
rect 17451 9333 17460 9367
rect 17408 9324 17460 9333
rect 19708 9392 19760 9444
rect 18512 9367 18564 9376
rect 18512 9333 18521 9367
rect 18521 9333 18555 9367
rect 18555 9333 18564 9367
rect 18512 9324 18564 9333
rect 18880 9324 18932 9376
rect 18972 9324 19024 9376
rect 20904 9367 20956 9376
rect 20904 9333 20913 9367
rect 20913 9333 20947 9367
rect 20947 9333 20956 9367
rect 20904 9324 20956 9333
rect 7912 9222 7964 9274
rect 7976 9222 8028 9274
rect 8040 9222 8092 9274
rect 8104 9222 8156 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 15035 9222 15087 9274
rect 1584 9163 1636 9172
rect 1584 9129 1593 9163
rect 1593 9129 1627 9163
rect 1627 9129 1636 9163
rect 1584 9120 1636 9129
rect 2504 9120 2556 9172
rect 2872 9163 2924 9172
rect 2872 9129 2881 9163
rect 2881 9129 2915 9163
rect 2915 9129 2924 9163
rect 2872 9120 2924 9129
rect 3424 9120 3476 9172
rect 4620 9120 4672 9172
rect 5448 9163 5500 9172
rect 4804 9052 4856 9104
rect 5448 9129 5457 9163
rect 5457 9129 5491 9163
rect 5491 9129 5500 9163
rect 5448 9120 5500 9129
rect 6276 9120 6328 9172
rect 8208 9120 8260 9172
rect 5632 9052 5684 9104
rect 1492 8916 1544 8968
rect 2412 8916 2464 8968
rect 2872 8916 2924 8968
rect 3056 8959 3108 8968
rect 3056 8925 3065 8959
rect 3065 8925 3099 8959
rect 3099 8925 3108 8959
rect 3056 8916 3108 8925
rect 2504 8780 2556 8832
rect 3148 8780 3200 8832
rect 3884 8984 3936 9036
rect 6460 9052 6512 9104
rect 7288 9052 7340 9104
rect 8024 9052 8076 9104
rect 8484 9052 8536 9104
rect 9036 9052 9088 9104
rect 10140 9120 10192 9172
rect 10600 9120 10652 9172
rect 6828 8984 6880 9036
rect 7380 9027 7432 9036
rect 7380 8993 7389 9027
rect 7389 8993 7423 9027
rect 7423 8993 7432 9027
rect 7380 8984 7432 8993
rect 7472 8984 7524 9036
rect 8208 8984 8260 9036
rect 8300 8984 8352 9036
rect 5080 8916 5132 8968
rect 5540 8916 5592 8968
rect 5080 8780 5132 8832
rect 5632 8823 5684 8832
rect 5632 8789 5641 8823
rect 5641 8789 5675 8823
rect 5675 8789 5684 8823
rect 5632 8780 5684 8789
rect 5724 8780 5776 8832
rect 7012 8848 7064 8900
rect 8208 8848 8260 8900
rect 7288 8780 7340 8832
rect 7932 8823 7984 8832
rect 7932 8789 7941 8823
rect 7941 8789 7975 8823
rect 7975 8789 7984 8823
rect 7932 8780 7984 8789
rect 9864 9052 9916 9104
rect 10324 9052 10376 9104
rect 10508 9052 10560 9104
rect 10968 9120 11020 9172
rect 11336 9120 11388 9172
rect 12900 9120 12952 9172
rect 13084 9095 13136 9104
rect 13084 9061 13093 9095
rect 13093 9061 13127 9095
rect 13127 9061 13136 9095
rect 14740 9120 14792 9172
rect 15200 9120 15252 9172
rect 15752 9120 15804 9172
rect 17132 9163 17184 9172
rect 17132 9129 17141 9163
rect 17141 9129 17175 9163
rect 17175 9129 17184 9163
rect 17132 9120 17184 9129
rect 17408 9120 17460 9172
rect 18512 9120 18564 9172
rect 20168 9163 20220 9172
rect 20168 9129 20177 9163
rect 20177 9129 20211 9163
rect 20211 9129 20220 9163
rect 20168 9120 20220 9129
rect 13084 9052 13136 9061
rect 9864 8916 9916 8968
rect 10140 8959 10192 8968
rect 10140 8925 10149 8959
rect 10149 8925 10183 8959
rect 10183 8925 10192 8959
rect 10140 8916 10192 8925
rect 9496 8780 9548 8832
rect 9588 8780 9640 8832
rect 10416 8984 10468 9036
rect 11428 8984 11480 9036
rect 11888 8984 11940 9036
rect 13728 9052 13780 9104
rect 14188 9052 14240 9104
rect 14556 9052 14608 9104
rect 15844 9052 15896 9104
rect 13636 9027 13688 9036
rect 13636 8993 13645 9027
rect 13645 8993 13679 9027
rect 13679 8993 13688 9027
rect 13636 8984 13688 8993
rect 15752 8984 15804 9036
rect 16488 8984 16540 9036
rect 19248 9052 19300 9104
rect 10876 8916 10928 8968
rect 12256 8916 12308 8968
rect 12532 8916 12584 8968
rect 12808 8916 12860 8968
rect 13452 8916 13504 8968
rect 14188 8916 14240 8968
rect 17500 8916 17552 8968
rect 17684 8959 17736 8968
rect 17684 8925 17693 8959
rect 17693 8925 17727 8959
rect 17727 8925 17736 8959
rect 17684 8916 17736 8925
rect 18052 8916 18104 8968
rect 19340 8984 19392 9036
rect 10416 8848 10468 8900
rect 10692 8848 10744 8900
rect 12808 8780 12860 8832
rect 13452 8780 13504 8832
rect 14648 8780 14700 8832
rect 14832 8891 14884 8900
rect 14832 8857 14841 8891
rect 14841 8857 14875 8891
rect 14875 8857 14884 8891
rect 14832 8848 14884 8857
rect 15936 8780 15988 8832
rect 16856 8780 16908 8832
rect 17960 8780 18012 8832
rect 18604 8780 18656 8832
rect 19524 8780 19576 8832
rect 20444 8780 20496 8832
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 4575 8678 4627 8730
rect 4639 8678 4691 8730
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 18308 8678 18360 8730
rect 18372 8678 18424 8730
rect 18436 8678 18488 8730
rect 18500 8678 18552 8730
rect 3148 8576 3200 8628
rect 4804 8576 4856 8628
rect 5908 8576 5960 8628
rect 6920 8576 6972 8628
rect 7472 8576 7524 8628
rect 2872 8508 2924 8560
rect 6828 8508 6880 8560
rect 1952 8372 2004 8424
rect 2688 8440 2740 8492
rect 6184 8440 6236 8492
rect 8760 8576 8812 8628
rect 10140 8576 10192 8628
rect 12716 8576 12768 8628
rect 13268 8619 13320 8628
rect 13268 8585 13277 8619
rect 13277 8585 13311 8619
rect 13311 8585 13320 8619
rect 13268 8576 13320 8585
rect 9588 8508 9640 8560
rect 11888 8508 11940 8560
rect 16396 8576 16448 8628
rect 16488 8576 16540 8628
rect 17500 8576 17552 8628
rect 18972 8576 19024 8628
rect 19156 8576 19208 8628
rect 19340 8576 19392 8628
rect 20904 8576 20956 8628
rect 8392 8440 8444 8492
rect 8484 8483 8536 8492
rect 8484 8449 8493 8483
rect 8493 8449 8527 8483
rect 8527 8449 8536 8483
rect 8484 8440 8536 8449
rect 10048 8440 10100 8492
rect 10508 8483 10560 8492
rect 2780 8372 2832 8424
rect 3884 8372 3936 8424
rect 6460 8372 6512 8424
rect 7012 8415 7064 8424
rect 7012 8381 7021 8415
rect 7021 8381 7055 8415
rect 7055 8381 7064 8415
rect 7012 8372 7064 8381
rect 7380 8372 7432 8424
rect 9772 8372 9824 8424
rect 10508 8449 10517 8483
rect 10517 8449 10551 8483
rect 10551 8449 10560 8483
rect 10508 8440 10560 8449
rect 12440 8440 12492 8492
rect 13084 8483 13136 8492
rect 2044 8304 2096 8356
rect 3056 8304 3108 8356
rect 5448 8304 5500 8356
rect 7288 8304 7340 8356
rect 7472 8304 7524 8356
rect 7656 8304 7708 8356
rect 8024 8304 8076 8356
rect 9496 8304 9548 8356
rect 10692 8304 10744 8356
rect 10968 8304 11020 8356
rect 3976 8236 4028 8288
rect 6092 8236 6144 8288
rect 6276 8279 6328 8288
rect 6276 8245 6285 8279
rect 6285 8245 6319 8279
rect 6319 8245 6328 8279
rect 6276 8236 6328 8245
rect 6460 8236 6512 8288
rect 7380 8279 7432 8288
rect 7380 8245 7389 8279
rect 7389 8245 7423 8279
rect 7423 8245 7432 8279
rect 7380 8236 7432 8245
rect 8852 8236 8904 8288
rect 9036 8236 9088 8288
rect 12348 8372 12400 8424
rect 12808 8415 12860 8424
rect 12808 8381 12817 8415
rect 12817 8381 12851 8415
rect 12851 8381 12860 8415
rect 12808 8372 12860 8381
rect 13084 8449 13093 8483
rect 13093 8449 13127 8483
rect 13127 8449 13136 8483
rect 13084 8440 13136 8449
rect 13268 8440 13320 8492
rect 15200 8483 15252 8492
rect 15200 8449 15209 8483
rect 15209 8449 15243 8483
rect 15243 8449 15252 8483
rect 15200 8440 15252 8449
rect 16764 8440 16816 8492
rect 16856 8372 16908 8424
rect 11888 8304 11940 8356
rect 14648 8304 14700 8356
rect 15936 8304 15988 8356
rect 17684 8440 17736 8492
rect 17132 8415 17184 8424
rect 17132 8381 17141 8415
rect 17141 8381 17175 8415
rect 17175 8381 17184 8415
rect 17132 8372 17184 8381
rect 19524 8508 19576 8560
rect 19616 8508 19668 8560
rect 18604 8483 18656 8492
rect 18604 8449 18613 8483
rect 18613 8449 18647 8483
rect 18647 8449 18656 8483
rect 18604 8440 18656 8449
rect 19156 8440 19208 8492
rect 21088 8483 21140 8492
rect 21088 8449 21097 8483
rect 21097 8449 21131 8483
rect 21131 8449 21140 8483
rect 21088 8440 21140 8449
rect 18512 8415 18564 8424
rect 18512 8381 18521 8415
rect 18521 8381 18555 8415
rect 18555 8381 18564 8415
rect 18512 8372 18564 8381
rect 18696 8372 18748 8424
rect 19984 8304 20036 8356
rect 12256 8279 12308 8288
rect 12256 8245 12265 8279
rect 12265 8245 12299 8279
rect 12299 8245 12308 8279
rect 12256 8236 12308 8245
rect 12808 8236 12860 8288
rect 13912 8236 13964 8288
rect 14740 8236 14792 8288
rect 16764 8236 16816 8288
rect 16856 8236 16908 8288
rect 17408 8236 17460 8288
rect 18144 8236 18196 8288
rect 19616 8236 19668 8288
rect 20076 8279 20128 8288
rect 20076 8245 20085 8279
rect 20085 8245 20119 8279
rect 20119 8245 20128 8279
rect 20076 8236 20128 8245
rect 20720 8236 20772 8288
rect 21456 8279 21508 8288
rect 21456 8245 21465 8279
rect 21465 8245 21499 8279
rect 21499 8245 21508 8279
rect 21456 8236 21508 8245
rect 7912 8134 7964 8186
rect 7976 8134 8028 8186
rect 8040 8134 8092 8186
rect 8104 8134 8156 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 15035 8134 15087 8186
rect 1492 8075 1544 8084
rect 1492 8041 1501 8075
rect 1501 8041 1535 8075
rect 1535 8041 1544 8075
rect 1492 8032 1544 8041
rect 2872 8032 2924 8084
rect 5172 8032 5224 8084
rect 6276 8032 6328 8084
rect 6736 8075 6788 8084
rect 6736 8041 6745 8075
rect 6745 8041 6779 8075
rect 6779 8041 6788 8075
rect 6736 8032 6788 8041
rect 7380 8032 7432 8084
rect 8300 8032 8352 8084
rect 3608 7964 3660 8016
rect 6644 7964 6696 8016
rect 7196 8007 7248 8016
rect 7196 7973 7205 8007
rect 7205 7973 7239 8007
rect 7239 7973 7248 8007
rect 7196 7964 7248 7973
rect 8668 7964 8720 8016
rect 8944 8032 8996 8084
rect 10324 8032 10376 8084
rect 9128 8007 9180 8016
rect 9128 7973 9137 8007
rect 9137 7973 9171 8007
rect 9171 7973 9180 8007
rect 11244 8032 11296 8084
rect 11336 8032 11388 8084
rect 11980 8032 12032 8084
rect 12440 8075 12492 8084
rect 12440 8041 12449 8075
rect 12449 8041 12483 8075
rect 12483 8041 12492 8075
rect 12440 8032 12492 8041
rect 12808 8032 12860 8084
rect 9128 7964 9180 7973
rect 2688 7896 2740 7948
rect 5080 7896 5132 7948
rect 6920 7896 6972 7948
rect 1676 7871 1728 7880
rect 1676 7837 1685 7871
rect 1685 7837 1719 7871
rect 1719 7837 1728 7871
rect 1676 7828 1728 7837
rect 3608 7871 3660 7880
rect 3608 7837 3617 7871
rect 3617 7837 3651 7871
rect 3651 7837 3660 7871
rect 3608 7828 3660 7837
rect 3056 7803 3108 7812
rect 3056 7769 3065 7803
rect 3065 7769 3099 7803
rect 3099 7769 3108 7803
rect 3056 7760 3108 7769
rect 3148 7735 3200 7744
rect 3148 7701 3157 7735
rect 3157 7701 3191 7735
rect 3191 7701 3200 7735
rect 3148 7692 3200 7701
rect 3700 7692 3752 7744
rect 5816 7760 5868 7812
rect 6828 7828 6880 7880
rect 7748 7896 7800 7948
rect 8300 7939 8352 7948
rect 7288 7871 7340 7880
rect 6736 7760 6788 7812
rect 7288 7837 7297 7871
rect 7297 7837 7331 7871
rect 7331 7837 7340 7871
rect 7288 7828 7340 7837
rect 8300 7905 8309 7939
rect 8309 7905 8343 7939
rect 8343 7905 8352 7939
rect 8300 7896 8352 7905
rect 9588 7896 9640 7948
rect 9956 7896 10008 7948
rect 7012 7760 7064 7812
rect 9496 7828 9548 7880
rect 10692 7896 10744 7948
rect 11060 7896 11112 7948
rect 12624 7939 12676 7948
rect 12624 7905 12633 7939
rect 12633 7905 12667 7939
rect 12667 7905 12676 7939
rect 12624 7896 12676 7905
rect 14648 8032 14700 8084
rect 18236 8032 18288 8084
rect 18972 8032 19024 8084
rect 19340 8032 19392 8084
rect 19984 8075 20036 8084
rect 19984 8041 19993 8075
rect 19993 8041 20027 8075
rect 20027 8041 20036 8075
rect 19984 8032 20036 8041
rect 20260 8032 20312 8084
rect 14556 7964 14608 8016
rect 15200 7964 15252 8016
rect 16672 8007 16724 8016
rect 16672 7973 16681 8007
rect 16681 7973 16715 8007
rect 16715 7973 16724 8007
rect 16672 7964 16724 7973
rect 13544 7896 13596 7948
rect 13912 7939 13964 7948
rect 13912 7905 13921 7939
rect 13921 7905 13955 7939
rect 13955 7905 13964 7939
rect 13912 7896 13964 7905
rect 14188 7896 14240 7948
rect 16488 7896 16540 7948
rect 17960 7939 18012 7948
rect 7748 7760 7800 7812
rect 8484 7760 8536 7812
rect 8944 7760 8996 7812
rect 9312 7760 9364 7812
rect 9864 7760 9916 7812
rect 10968 7871 11020 7880
rect 10968 7837 10977 7871
rect 10977 7837 11011 7871
rect 11011 7837 11020 7871
rect 10968 7828 11020 7837
rect 12348 7828 12400 7880
rect 13636 7828 13688 7880
rect 14004 7871 14056 7880
rect 14004 7837 14013 7871
rect 14013 7837 14047 7871
rect 14047 7837 14056 7871
rect 14004 7828 14056 7837
rect 14096 7871 14148 7880
rect 14096 7837 14105 7871
rect 14105 7837 14139 7871
rect 14139 7837 14148 7871
rect 14096 7828 14148 7837
rect 14740 7828 14792 7880
rect 15476 7828 15528 7880
rect 15936 7871 15988 7880
rect 15936 7837 15945 7871
rect 15945 7837 15979 7871
rect 15979 7837 15988 7871
rect 15936 7828 15988 7837
rect 5080 7692 5132 7744
rect 6460 7692 6512 7744
rect 8760 7692 8812 7744
rect 9772 7735 9824 7744
rect 9772 7701 9781 7735
rect 9781 7701 9815 7735
rect 9815 7701 9824 7735
rect 10692 7760 10744 7812
rect 16304 7828 16356 7880
rect 17960 7905 17969 7939
rect 17969 7905 18003 7939
rect 18003 7905 18012 7939
rect 17960 7896 18012 7905
rect 18604 7896 18656 7948
rect 19340 7896 19392 7948
rect 9772 7692 9824 7701
rect 10324 7692 10376 7744
rect 16948 7760 17000 7812
rect 12348 7735 12400 7744
rect 12348 7701 12357 7735
rect 12357 7701 12391 7735
rect 12391 7701 12400 7735
rect 12348 7692 12400 7701
rect 12992 7692 13044 7744
rect 13912 7692 13964 7744
rect 14556 7692 14608 7744
rect 15568 7692 15620 7744
rect 17684 7871 17736 7880
rect 17684 7837 17693 7871
rect 17693 7837 17727 7871
rect 17727 7837 17736 7871
rect 17684 7828 17736 7837
rect 19064 7828 19116 7880
rect 20904 7828 20956 7880
rect 21088 7828 21140 7880
rect 19616 7803 19668 7812
rect 19616 7769 19625 7803
rect 19625 7769 19659 7803
rect 19659 7769 19668 7803
rect 19616 7760 19668 7769
rect 20720 7760 20772 7812
rect 19156 7692 19208 7744
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 4575 7590 4627 7642
rect 4639 7590 4691 7642
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 18308 7590 18360 7642
rect 18372 7590 18424 7642
rect 18436 7590 18488 7642
rect 18500 7590 18552 7642
rect 3608 7488 3660 7540
rect 1676 7284 1728 7336
rect 3884 7352 3936 7404
rect 5448 7420 5500 7472
rect 6184 7420 6236 7472
rect 5172 7352 5224 7404
rect 2596 7216 2648 7268
rect 2688 7148 2740 7200
rect 4804 7284 4856 7336
rect 5356 7327 5408 7336
rect 5356 7293 5365 7327
rect 5365 7293 5399 7327
rect 5399 7293 5408 7327
rect 5356 7284 5408 7293
rect 5448 7284 5500 7336
rect 7380 7395 7432 7404
rect 7380 7361 7389 7395
rect 7389 7361 7423 7395
rect 7423 7361 7432 7395
rect 7380 7352 7432 7361
rect 7012 7284 7064 7336
rect 7104 7284 7156 7336
rect 8024 7488 8076 7540
rect 8300 7488 8352 7540
rect 10048 7488 10100 7540
rect 10508 7488 10560 7540
rect 10692 7531 10744 7540
rect 10692 7497 10701 7531
rect 10701 7497 10735 7531
rect 10735 7497 10744 7531
rect 10692 7488 10744 7497
rect 10876 7531 10928 7540
rect 10876 7497 10885 7531
rect 10885 7497 10919 7531
rect 10919 7497 10928 7531
rect 10876 7488 10928 7497
rect 12072 7488 12124 7540
rect 9312 7420 9364 7472
rect 13084 7488 13136 7540
rect 13728 7488 13780 7540
rect 14648 7488 14700 7540
rect 9496 7352 9548 7404
rect 9772 7352 9824 7404
rect 10048 7352 10100 7404
rect 10232 7395 10284 7404
rect 10232 7361 10241 7395
rect 10241 7361 10275 7395
rect 10275 7361 10284 7395
rect 10232 7352 10284 7361
rect 10692 7352 10744 7404
rect 11060 7352 11112 7404
rect 12992 7420 13044 7472
rect 4344 7216 4396 7268
rect 4988 7191 5040 7200
rect 4988 7157 4997 7191
rect 4997 7157 5031 7191
rect 5031 7157 5040 7191
rect 4988 7148 5040 7157
rect 5632 7216 5684 7268
rect 6092 7216 6144 7268
rect 7748 7284 7800 7336
rect 11244 7284 11296 7336
rect 12624 7352 12676 7404
rect 13636 7352 13688 7404
rect 13728 7395 13780 7404
rect 13728 7361 13737 7395
rect 13737 7361 13771 7395
rect 13771 7361 13780 7395
rect 13728 7352 13780 7361
rect 14096 7352 14148 7404
rect 16580 7488 16632 7540
rect 16672 7488 16724 7540
rect 16856 7488 16908 7540
rect 17132 7531 17184 7540
rect 17132 7497 17141 7531
rect 17141 7497 17175 7531
rect 17175 7497 17184 7531
rect 17132 7488 17184 7497
rect 17500 7488 17552 7540
rect 17776 7488 17828 7540
rect 18052 7531 18104 7540
rect 18052 7497 18061 7531
rect 18061 7497 18095 7531
rect 18095 7497 18104 7531
rect 18052 7488 18104 7497
rect 18604 7488 18656 7540
rect 19800 7488 19852 7540
rect 20076 7488 20128 7540
rect 19432 7420 19484 7472
rect 15568 7352 15620 7404
rect 16488 7352 16540 7404
rect 16856 7395 16908 7404
rect 16396 7284 16448 7336
rect 16856 7361 16865 7395
rect 16865 7361 16899 7395
rect 16899 7361 16908 7395
rect 16856 7352 16908 7361
rect 17040 7352 17092 7404
rect 18604 7395 18656 7404
rect 18604 7361 18613 7395
rect 18613 7361 18647 7395
rect 18647 7361 18656 7395
rect 18604 7352 18656 7361
rect 20812 7420 20864 7472
rect 17776 7284 17828 7336
rect 7564 7216 7616 7268
rect 8024 7216 8076 7268
rect 9036 7216 9088 7268
rect 10416 7259 10468 7268
rect 10416 7225 10425 7259
rect 10425 7225 10459 7259
rect 10459 7225 10468 7259
rect 10416 7216 10468 7225
rect 10784 7216 10836 7268
rect 11520 7216 11572 7268
rect 8300 7148 8352 7200
rect 9956 7191 10008 7200
rect 9956 7157 9965 7191
rect 9965 7157 9999 7191
rect 9999 7157 10008 7191
rect 9956 7148 10008 7157
rect 10048 7148 10100 7200
rect 11428 7148 11480 7200
rect 12072 7191 12124 7200
rect 12072 7157 12081 7191
rect 12081 7157 12115 7191
rect 12115 7157 12124 7191
rect 12624 7216 12676 7268
rect 16764 7216 16816 7268
rect 17408 7216 17460 7268
rect 19800 7352 19852 7404
rect 20904 7395 20956 7404
rect 20904 7361 20913 7395
rect 20913 7361 20947 7395
rect 20947 7361 20956 7395
rect 20904 7352 20956 7361
rect 19340 7284 19392 7336
rect 20352 7284 20404 7336
rect 20444 7284 20496 7336
rect 20812 7284 20864 7336
rect 20076 7216 20128 7268
rect 20168 7216 20220 7268
rect 12808 7191 12860 7200
rect 12072 7148 12124 7157
rect 12808 7157 12817 7191
rect 12817 7157 12851 7191
rect 12851 7157 12860 7191
rect 12808 7148 12860 7157
rect 13728 7148 13780 7200
rect 14096 7191 14148 7200
rect 14096 7157 14105 7191
rect 14105 7157 14139 7191
rect 14139 7157 14148 7191
rect 14096 7148 14148 7157
rect 14464 7191 14516 7200
rect 14464 7157 14473 7191
rect 14473 7157 14507 7191
rect 14507 7157 14516 7191
rect 14464 7148 14516 7157
rect 14648 7148 14700 7200
rect 16028 7148 16080 7200
rect 16304 7148 16356 7200
rect 16580 7148 16632 7200
rect 16672 7148 16724 7200
rect 19340 7148 19392 7200
rect 19524 7191 19576 7200
rect 19524 7157 19533 7191
rect 19533 7157 19567 7191
rect 19567 7157 19576 7191
rect 19524 7148 19576 7157
rect 19984 7191 20036 7200
rect 19984 7157 19993 7191
rect 19993 7157 20027 7191
rect 20027 7157 20036 7191
rect 19984 7148 20036 7157
rect 20720 7191 20772 7200
rect 20720 7157 20729 7191
rect 20729 7157 20763 7191
rect 20763 7157 20772 7191
rect 20720 7148 20772 7157
rect 20812 7191 20864 7200
rect 20812 7157 20821 7191
rect 20821 7157 20855 7191
rect 20855 7157 20864 7191
rect 20812 7148 20864 7157
rect 7912 7046 7964 7098
rect 7976 7046 8028 7098
rect 8040 7046 8092 7098
rect 8104 7046 8156 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 15035 7046 15087 7098
rect 2412 6944 2464 6996
rect 3056 6944 3108 6996
rect 7012 6987 7064 6996
rect 7012 6953 7021 6987
rect 7021 6953 7055 6987
rect 7055 6953 7064 6987
rect 7012 6944 7064 6953
rect 7196 6944 7248 6996
rect 9956 6944 10008 6996
rect 10324 6987 10376 6996
rect 10324 6953 10333 6987
rect 10333 6953 10367 6987
rect 10367 6953 10376 6987
rect 10324 6944 10376 6953
rect 11520 6987 11572 6996
rect 11520 6953 11529 6987
rect 11529 6953 11563 6987
rect 11563 6953 11572 6987
rect 11520 6944 11572 6953
rect 1768 6808 1820 6860
rect 2504 6876 2556 6928
rect 3424 6876 3476 6928
rect 3700 6876 3752 6928
rect 4068 6876 4120 6928
rect 11704 6944 11756 6996
rect 12900 6944 12952 6996
rect 14556 6987 14608 6996
rect 1676 6783 1728 6792
rect 1676 6749 1685 6783
rect 1685 6749 1719 6783
rect 1719 6749 1728 6783
rect 1676 6740 1728 6749
rect 2596 6783 2648 6792
rect 1952 6715 2004 6724
rect 1952 6681 1961 6715
rect 1961 6681 1995 6715
rect 1995 6681 2004 6715
rect 1952 6672 2004 6681
rect 2596 6749 2605 6783
rect 2605 6749 2639 6783
rect 2639 6749 2648 6783
rect 2596 6740 2648 6749
rect 1308 6604 1360 6656
rect 5172 6808 5224 6860
rect 5816 6851 5868 6860
rect 5816 6817 5850 6851
rect 5850 6817 5868 6851
rect 5816 6808 5868 6817
rect 6184 6808 6236 6860
rect 3056 6740 3108 6792
rect 3424 6783 3476 6792
rect 3424 6749 3433 6783
rect 3433 6749 3467 6783
rect 3467 6749 3476 6783
rect 3424 6740 3476 6749
rect 3884 6740 3936 6792
rect 7656 6808 7708 6860
rect 5448 6647 5500 6656
rect 5448 6613 5457 6647
rect 5457 6613 5491 6647
rect 5491 6613 5500 6647
rect 5448 6604 5500 6613
rect 6920 6647 6972 6656
rect 6920 6613 6929 6647
rect 6929 6613 6963 6647
rect 6963 6613 6972 6647
rect 6920 6604 6972 6613
rect 7840 6783 7892 6792
rect 7380 6672 7432 6724
rect 7840 6749 7849 6783
rect 7849 6749 7883 6783
rect 7883 6749 7892 6783
rect 7840 6740 7892 6749
rect 8024 6783 8076 6792
rect 8024 6749 8033 6783
rect 8033 6749 8067 6783
rect 8067 6749 8076 6783
rect 8024 6740 8076 6749
rect 8208 6740 8260 6792
rect 8668 6808 8720 6860
rect 9404 6740 9456 6792
rect 10324 6740 10376 6792
rect 14556 6953 14565 6987
rect 14565 6953 14599 6987
rect 14599 6953 14608 6987
rect 14556 6944 14608 6953
rect 15200 6944 15252 6996
rect 16028 6944 16080 6996
rect 16488 6944 16540 6996
rect 17132 6944 17184 6996
rect 18144 6944 18196 6996
rect 19524 6944 19576 6996
rect 19800 6944 19852 6996
rect 20076 6987 20128 6996
rect 20076 6953 20085 6987
rect 20085 6953 20119 6987
rect 20119 6953 20128 6987
rect 20076 6944 20128 6953
rect 12348 6808 12400 6860
rect 16304 6876 16356 6928
rect 17592 6876 17644 6928
rect 18512 6876 18564 6928
rect 19432 6876 19484 6928
rect 8116 6672 8168 6724
rect 8300 6672 8352 6724
rect 10600 6672 10652 6724
rect 10968 6672 11020 6724
rect 8484 6604 8536 6656
rect 9036 6604 9088 6656
rect 10324 6604 10376 6656
rect 13360 6740 13412 6792
rect 13636 6783 13688 6792
rect 13636 6749 13645 6783
rect 13645 6749 13679 6783
rect 13679 6749 13688 6783
rect 14004 6808 14056 6860
rect 14832 6783 14884 6792
rect 13636 6740 13688 6749
rect 14464 6672 14516 6724
rect 14832 6749 14841 6783
rect 14841 6749 14875 6783
rect 14875 6749 14884 6783
rect 14832 6740 14884 6749
rect 15752 6740 15804 6792
rect 16120 6740 16172 6792
rect 17224 6808 17276 6860
rect 17408 6851 17460 6860
rect 17408 6817 17417 6851
rect 17417 6817 17451 6851
rect 17451 6817 17460 6851
rect 17408 6808 17460 6817
rect 17040 6740 17092 6792
rect 17224 6672 17276 6724
rect 18144 6740 18196 6792
rect 18604 6740 18656 6792
rect 19156 6740 19208 6792
rect 20904 6740 20956 6792
rect 18880 6715 18932 6724
rect 18880 6681 18889 6715
rect 18889 6681 18923 6715
rect 18923 6681 18932 6715
rect 18880 6672 18932 6681
rect 19248 6672 19300 6724
rect 21088 6715 21140 6724
rect 21088 6681 21097 6715
rect 21097 6681 21131 6715
rect 21131 6681 21140 6715
rect 21088 6672 21140 6681
rect 12992 6647 13044 6656
rect 12992 6613 13001 6647
rect 13001 6613 13035 6647
rect 13035 6613 13044 6647
rect 12992 6604 13044 6613
rect 13636 6604 13688 6656
rect 14004 6604 14056 6656
rect 14188 6647 14240 6656
rect 14188 6613 14197 6647
rect 14197 6613 14231 6647
rect 14231 6613 14240 6647
rect 14188 6604 14240 6613
rect 15476 6604 15528 6656
rect 16120 6604 16172 6656
rect 17776 6604 17828 6656
rect 18604 6604 18656 6656
rect 18696 6604 18748 6656
rect 19984 6604 20036 6656
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 4575 6502 4627 6554
rect 4639 6502 4691 6554
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 18308 6502 18360 6554
rect 18372 6502 18424 6554
rect 18436 6502 18488 6554
rect 18500 6502 18552 6554
rect 2044 6443 2096 6452
rect 2044 6409 2053 6443
rect 2053 6409 2087 6443
rect 2087 6409 2096 6443
rect 2044 6400 2096 6409
rect 4344 6400 4396 6452
rect 5264 6400 5316 6452
rect 2596 6332 2648 6384
rect 3792 6307 3844 6316
rect 3792 6273 3801 6307
rect 3801 6273 3835 6307
rect 3835 6273 3844 6307
rect 3792 6264 3844 6273
rect 4988 6264 5040 6316
rect 5448 6332 5500 6384
rect 6000 6332 6052 6384
rect 6920 6264 6972 6316
rect 1676 6196 1728 6248
rect 3516 6196 3568 6248
rect 6368 6239 6420 6248
rect 6368 6205 6377 6239
rect 6377 6205 6411 6239
rect 6411 6205 6420 6239
rect 6368 6196 6420 6205
rect 7380 6307 7432 6316
rect 7380 6273 7389 6307
rect 7389 6273 7423 6307
rect 7423 6273 7432 6307
rect 7380 6264 7432 6273
rect 9588 6400 9640 6452
rect 10692 6443 10744 6452
rect 10692 6409 10701 6443
rect 10701 6409 10735 6443
rect 10735 6409 10744 6443
rect 10692 6400 10744 6409
rect 8208 6332 8260 6384
rect 11428 6332 11480 6384
rect 8392 6264 8444 6316
rect 10784 6264 10836 6316
rect 12532 6400 12584 6452
rect 13360 6443 13412 6452
rect 13360 6409 13369 6443
rect 13369 6409 13403 6443
rect 13403 6409 13412 6443
rect 13360 6400 13412 6409
rect 14096 6400 14148 6452
rect 14188 6400 14240 6452
rect 13544 6332 13596 6384
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 12716 6264 12768 6316
rect 12992 6307 13044 6316
rect 12992 6273 13001 6307
rect 13001 6273 13035 6307
rect 13035 6273 13044 6307
rect 15292 6400 15344 6452
rect 18144 6443 18196 6452
rect 16764 6332 16816 6384
rect 12992 6264 13044 6273
rect 1492 6128 1544 6180
rect 1768 6103 1820 6112
rect 1768 6069 1777 6103
rect 1777 6069 1811 6103
rect 1811 6069 1820 6103
rect 1768 6060 1820 6069
rect 3056 6128 3108 6180
rect 3700 6128 3752 6180
rect 4160 6128 4212 6180
rect 2688 6060 2740 6112
rect 3148 6103 3200 6112
rect 3148 6069 3157 6103
rect 3157 6069 3191 6103
rect 3191 6069 3200 6103
rect 3148 6060 3200 6069
rect 3516 6103 3568 6112
rect 3516 6069 3525 6103
rect 3525 6069 3559 6103
rect 3559 6069 3568 6103
rect 3516 6060 3568 6069
rect 4344 6060 4396 6112
rect 5908 6103 5960 6112
rect 5908 6069 5917 6103
rect 5917 6069 5951 6103
rect 5951 6069 5960 6103
rect 5908 6060 5960 6069
rect 6276 6103 6328 6112
rect 6276 6069 6285 6103
rect 6285 6069 6319 6103
rect 6319 6069 6328 6103
rect 6276 6060 6328 6069
rect 7840 6128 7892 6180
rect 8116 6171 8168 6180
rect 8116 6137 8125 6171
rect 8125 6137 8159 6171
rect 8159 6137 8168 6171
rect 8116 6128 8168 6137
rect 10324 6128 10376 6180
rect 11152 6196 11204 6248
rect 12624 6128 12676 6180
rect 18144 6409 18153 6443
rect 18153 6409 18187 6443
rect 18187 6409 18196 6443
rect 18144 6400 18196 6409
rect 20904 6400 20956 6452
rect 17960 6332 18012 6384
rect 18696 6332 18748 6384
rect 17224 6307 17276 6316
rect 17224 6273 17233 6307
rect 17233 6273 17267 6307
rect 17267 6273 17276 6307
rect 17224 6264 17276 6273
rect 17408 6307 17460 6316
rect 17408 6273 17417 6307
rect 17417 6273 17451 6307
rect 17451 6273 17460 6307
rect 17408 6264 17460 6273
rect 20352 6332 20404 6384
rect 21088 6332 21140 6384
rect 7656 6103 7708 6112
rect 7656 6069 7665 6103
rect 7665 6069 7699 6103
rect 7699 6069 7708 6103
rect 7656 6060 7708 6069
rect 7748 6060 7800 6112
rect 8760 6060 8812 6112
rect 9220 6060 9272 6112
rect 9864 6060 9916 6112
rect 10048 6103 10100 6112
rect 10048 6069 10057 6103
rect 10057 6069 10091 6103
rect 10091 6069 10100 6103
rect 10048 6060 10100 6069
rect 10968 6060 11020 6112
rect 12440 6060 12492 6112
rect 14832 6196 14884 6248
rect 16120 6239 16172 6248
rect 16120 6205 16129 6239
rect 16129 6205 16163 6239
rect 16163 6205 16172 6239
rect 16120 6196 16172 6205
rect 14004 6128 14056 6180
rect 15844 6128 15896 6180
rect 17684 6128 17736 6180
rect 20076 6128 20128 6180
rect 13636 6103 13688 6112
rect 13636 6069 13645 6103
rect 13645 6069 13679 6103
rect 13679 6069 13688 6103
rect 13636 6060 13688 6069
rect 13912 6060 13964 6112
rect 15200 6060 15252 6112
rect 16856 6060 16908 6112
rect 17040 6103 17092 6112
rect 17040 6069 17049 6103
rect 17049 6069 17083 6103
rect 17083 6069 17092 6103
rect 17040 6060 17092 6069
rect 18144 6060 18196 6112
rect 7912 5958 7964 6010
rect 7976 5958 8028 6010
rect 8040 5958 8092 6010
rect 8104 5958 8156 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 15035 5958 15087 6010
rect 2320 5899 2372 5908
rect 2320 5865 2329 5899
rect 2329 5865 2363 5899
rect 2363 5865 2372 5899
rect 2320 5856 2372 5865
rect 3148 5856 3200 5908
rect 4068 5856 4120 5908
rect 1860 5788 1912 5840
rect 5540 5788 5592 5840
rect 6276 5856 6328 5908
rect 7012 5856 7064 5908
rect 7748 5856 7800 5908
rect 8576 5899 8628 5908
rect 8576 5865 8585 5899
rect 8585 5865 8619 5899
rect 8619 5865 8628 5899
rect 8576 5856 8628 5865
rect 9680 5856 9732 5908
rect 10692 5856 10744 5908
rect 11980 5856 12032 5908
rect 1676 5763 1728 5772
rect 1676 5729 1685 5763
rect 1685 5729 1719 5763
rect 1719 5729 1728 5763
rect 1676 5720 1728 5729
rect 3976 5720 4028 5772
rect 2964 5652 3016 5704
rect 7012 5720 7064 5772
rect 7840 5720 7892 5772
rect 14648 5856 14700 5908
rect 15844 5856 15896 5908
rect 15936 5856 15988 5908
rect 16672 5856 16724 5908
rect 17040 5856 17092 5908
rect 17316 5856 17368 5908
rect 17592 5899 17644 5908
rect 17592 5865 17601 5899
rect 17601 5865 17635 5899
rect 17635 5865 17644 5899
rect 17592 5856 17644 5865
rect 17776 5856 17828 5908
rect 18144 5856 18196 5908
rect 20076 5899 20128 5908
rect 20076 5865 20085 5899
rect 20085 5865 20119 5899
rect 20119 5865 20128 5899
rect 20076 5856 20128 5865
rect 12992 5788 13044 5840
rect 9496 5720 9548 5772
rect 10324 5720 10376 5772
rect 12440 5720 12492 5772
rect 12624 5720 12676 5772
rect 13728 5720 13780 5772
rect 3056 5584 3108 5636
rect 3516 5584 3568 5636
rect 3700 5584 3752 5636
rect 3884 5584 3936 5636
rect 5356 5652 5408 5704
rect 6828 5695 6880 5704
rect 6828 5661 6837 5695
rect 6837 5661 6871 5695
rect 6871 5661 6880 5695
rect 6828 5652 6880 5661
rect 7288 5695 7340 5704
rect 7288 5661 7297 5695
rect 7297 5661 7331 5695
rect 7331 5661 7340 5695
rect 7288 5652 7340 5661
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 8576 5652 8628 5704
rect 9036 5695 9088 5704
rect 9036 5661 9045 5695
rect 9045 5661 9079 5695
rect 9079 5661 9088 5695
rect 9036 5652 9088 5661
rect 6184 5584 6236 5636
rect 6736 5584 6788 5636
rect 9404 5652 9456 5704
rect 11704 5695 11756 5704
rect 11704 5661 11713 5695
rect 11713 5661 11747 5695
rect 11747 5661 11756 5695
rect 11704 5652 11756 5661
rect 10968 5584 11020 5636
rect 15476 5720 15528 5772
rect 17132 5763 17184 5772
rect 17132 5729 17141 5763
rect 17141 5729 17175 5763
rect 17175 5729 17184 5763
rect 17132 5720 17184 5729
rect 17408 5720 17460 5772
rect 5724 5559 5776 5568
rect 5724 5525 5733 5559
rect 5733 5525 5767 5559
rect 5767 5525 5776 5559
rect 5724 5516 5776 5525
rect 6276 5559 6328 5568
rect 6276 5525 6285 5559
rect 6285 5525 6319 5559
rect 6319 5525 6328 5559
rect 6276 5516 6328 5525
rect 7748 5559 7800 5568
rect 7748 5525 7757 5559
rect 7757 5525 7791 5559
rect 7791 5525 7800 5559
rect 7748 5516 7800 5525
rect 8024 5516 8076 5568
rect 8760 5516 8812 5568
rect 9496 5559 9548 5568
rect 9496 5525 9505 5559
rect 9505 5525 9539 5559
rect 9539 5525 9548 5559
rect 9496 5516 9548 5525
rect 9588 5516 9640 5568
rect 10692 5516 10744 5568
rect 10784 5516 10836 5568
rect 11244 5516 11296 5568
rect 14556 5584 14608 5636
rect 15292 5652 15344 5704
rect 17224 5652 17276 5704
rect 13912 5559 13964 5568
rect 13912 5525 13921 5559
rect 13921 5525 13955 5559
rect 13955 5525 13964 5559
rect 13912 5516 13964 5525
rect 15108 5516 15160 5568
rect 15476 5516 15528 5568
rect 16672 5516 16724 5568
rect 19984 5788 20036 5840
rect 20536 5788 20588 5840
rect 18696 5763 18748 5772
rect 18696 5729 18705 5763
rect 18705 5729 18739 5763
rect 18739 5729 18748 5763
rect 18696 5720 18748 5729
rect 19524 5720 19576 5772
rect 20168 5763 20220 5772
rect 20168 5729 20177 5763
rect 20177 5729 20211 5763
rect 20211 5729 20220 5763
rect 20168 5720 20220 5729
rect 22008 5559 22060 5568
rect 22008 5525 22017 5559
rect 22017 5525 22051 5559
rect 22051 5525 22060 5559
rect 22008 5516 22060 5525
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 4575 5414 4627 5466
rect 4639 5414 4691 5466
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 18308 5414 18360 5466
rect 18372 5414 18424 5466
rect 18436 5414 18488 5466
rect 18500 5414 18552 5466
rect 3056 5312 3108 5364
rect 3884 5312 3936 5364
rect 4344 5312 4396 5364
rect 5540 5355 5592 5364
rect 5540 5321 5549 5355
rect 5549 5321 5583 5355
rect 5583 5321 5592 5355
rect 5540 5312 5592 5321
rect 7012 5355 7064 5364
rect 7012 5321 7021 5355
rect 7021 5321 7055 5355
rect 7055 5321 7064 5355
rect 7012 5312 7064 5321
rect 7104 5312 7156 5364
rect 7840 5312 7892 5364
rect 8392 5312 8444 5364
rect 8668 5244 8720 5296
rect 9404 5312 9456 5364
rect 5356 5219 5408 5228
rect 5356 5185 5365 5219
rect 5365 5185 5399 5219
rect 5399 5185 5408 5219
rect 5356 5176 5408 5185
rect 5908 5176 5960 5228
rect 6184 5219 6236 5228
rect 6184 5185 6193 5219
rect 6193 5185 6227 5219
rect 6227 5185 6236 5219
rect 6184 5176 6236 5185
rect 7104 5176 7156 5228
rect 7380 5176 7432 5228
rect 7748 5176 7800 5228
rect 7932 5219 7984 5228
rect 7932 5185 7941 5219
rect 7941 5185 7975 5219
rect 7975 5185 7984 5219
rect 7932 5176 7984 5185
rect 1400 5108 1452 5160
rect 2780 5040 2832 5092
rect 2872 5040 2924 5092
rect 3792 5108 3844 5160
rect 10784 5312 10836 5364
rect 11704 5312 11756 5364
rect 11980 5312 12032 5364
rect 12716 5312 12768 5364
rect 14556 5312 14608 5364
rect 16580 5355 16632 5364
rect 11336 5244 11388 5296
rect 12256 5244 12308 5296
rect 12900 5244 12952 5296
rect 10784 5176 10836 5228
rect 10968 5176 11020 5228
rect 11980 5219 12032 5228
rect 11980 5185 11989 5219
rect 11989 5185 12023 5219
rect 12023 5185 12032 5219
rect 11980 5176 12032 5185
rect 13084 5219 13136 5228
rect 13084 5185 13093 5219
rect 13093 5185 13127 5219
rect 13127 5185 13136 5219
rect 13084 5176 13136 5185
rect 13912 5176 13964 5228
rect 14740 5176 14792 5228
rect 14832 5219 14884 5228
rect 14832 5185 14841 5219
rect 14841 5185 14875 5219
rect 14875 5185 14884 5219
rect 16580 5321 16589 5355
rect 16589 5321 16623 5355
rect 16623 5321 16632 5355
rect 16580 5312 16632 5321
rect 17132 5312 17184 5364
rect 19064 5312 19116 5364
rect 19524 5355 19576 5364
rect 19524 5321 19533 5355
rect 19533 5321 19567 5355
rect 19567 5321 19576 5355
rect 19524 5312 19576 5321
rect 20168 5312 20220 5364
rect 16672 5244 16724 5296
rect 14832 5176 14884 5185
rect 16580 5176 16632 5228
rect 16764 5176 16816 5228
rect 17592 5244 17644 5296
rect 18144 5244 18196 5296
rect 17408 5176 17460 5228
rect 19708 5244 19760 5296
rect 20076 5244 20128 5296
rect 11796 5151 11848 5160
rect 11796 5117 11805 5151
rect 11805 5117 11839 5151
rect 11839 5117 11848 5151
rect 11796 5108 11848 5117
rect 12440 5108 12492 5160
rect 13176 5108 13228 5160
rect 13728 5108 13780 5160
rect 15200 5108 15252 5160
rect 16856 5108 16908 5160
rect 17316 5108 17368 5160
rect 17868 5108 17920 5160
rect 18052 5108 18104 5160
rect 18696 5108 18748 5160
rect 3700 5040 3752 5092
rect 4252 5040 4304 5092
rect 6276 5040 6328 5092
rect 6644 5083 6696 5092
rect 6644 5049 6653 5083
rect 6653 5049 6687 5083
rect 6687 5049 6696 5083
rect 6644 5040 6696 5049
rect 3424 4972 3476 5024
rect 5724 4972 5776 5024
rect 7380 5015 7432 5024
rect 7380 4981 7389 5015
rect 7389 4981 7423 5015
rect 7423 4981 7432 5015
rect 7380 4972 7432 4981
rect 7656 5040 7708 5092
rect 8024 5040 8076 5092
rect 8760 5083 8812 5092
rect 8760 5049 8769 5083
rect 8769 5049 8803 5083
rect 8803 5049 8812 5083
rect 8760 5040 8812 5049
rect 9220 5040 9272 5092
rect 9680 4972 9732 5024
rect 10508 5015 10560 5024
rect 10508 4981 10517 5015
rect 10517 4981 10551 5015
rect 10551 4981 10560 5015
rect 10508 4972 10560 4981
rect 10600 5015 10652 5024
rect 10600 4981 10609 5015
rect 10609 4981 10643 5015
rect 10643 4981 10652 5015
rect 10876 5040 10928 5092
rect 12256 5040 12308 5092
rect 10600 4972 10652 4981
rect 11244 4972 11296 5024
rect 11704 4972 11756 5024
rect 12532 4972 12584 5024
rect 12716 5040 12768 5092
rect 13912 5040 13964 5092
rect 13360 5015 13412 5024
rect 13360 4981 13369 5015
rect 13369 4981 13403 5015
rect 13403 4981 13412 5015
rect 13360 4972 13412 4981
rect 13728 5015 13780 5024
rect 13728 4981 13737 5015
rect 13737 4981 13771 5015
rect 13771 4981 13780 5015
rect 13728 4972 13780 4981
rect 14004 4972 14056 5024
rect 15016 5040 15068 5092
rect 15292 5040 15344 5092
rect 18328 5040 18380 5092
rect 16120 4972 16172 5024
rect 17868 4972 17920 5024
rect 19984 5015 20036 5024
rect 19984 4981 19993 5015
rect 19993 4981 20027 5015
rect 20027 4981 20036 5015
rect 19984 4972 20036 4981
rect 7912 4870 7964 4922
rect 7976 4870 8028 4922
rect 8040 4870 8092 4922
rect 8104 4870 8156 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 15035 4870 15087 4922
rect 2780 4811 2832 4820
rect 2780 4777 2789 4811
rect 2789 4777 2823 4811
rect 2823 4777 2832 4811
rect 4068 4811 4120 4820
rect 2780 4768 2832 4777
rect 4068 4777 4077 4811
rect 4077 4777 4111 4811
rect 4111 4777 4120 4811
rect 4068 4768 4120 4777
rect 7104 4768 7156 4820
rect 8392 4811 8444 4820
rect 8392 4777 8401 4811
rect 8401 4777 8435 4811
rect 8435 4777 8444 4811
rect 8392 4768 8444 4777
rect 8760 4811 8812 4820
rect 8760 4777 8769 4811
rect 8769 4777 8803 4811
rect 8803 4777 8812 4811
rect 8760 4768 8812 4777
rect 9128 4811 9180 4820
rect 9128 4777 9137 4811
rect 9137 4777 9171 4811
rect 9171 4777 9180 4811
rect 9128 4768 9180 4777
rect 10048 4768 10100 4820
rect 10416 4768 10468 4820
rect 11336 4768 11388 4820
rect 11796 4768 11848 4820
rect 12256 4811 12308 4820
rect 12256 4777 12265 4811
rect 12265 4777 12299 4811
rect 12299 4777 12308 4811
rect 12256 4768 12308 4777
rect 12440 4811 12492 4820
rect 12440 4777 12449 4811
rect 12449 4777 12483 4811
rect 12483 4777 12492 4811
rect 12440 4768 12492 4777
rect 1308 4700 1360 4752
rect 1400 4675 1452 4684
rect 1400 4641 1409 4675
rect 1409 4641 1443 4675
rect 1443 4641 1452 4675
rect 1400 4632 1452 4641
rect 2688 4700 2740 4752
rect 3516 4675 3568 4684
rect 3516 4641 3525 4675
rect 3525 4641 3559 4675
rect 3559 4641 3568 4675
rect 3516 4632 3568 4641
rect 3700 4700 3752 4752
rect 5172 4675 5224 4684
rect 5172 4641 5181 4675
rect 5181 4641 5215 4675
rect 5215 4641 5224 4675
rect 5172 4632 5224 4641
rect 10508 4700 10560 4752
rect 7472 4675 7524 4684
rect 2412 4496 2464 4548
rect 2964 4471 3016 4480
rect 2964 4437 2973 4471
rect 2973 4437 3007 4471
rect 3007 4437 3016 4471
rect 2964 4428 3016 4437
rect 3700 4607 3752 4616
rect 3700 4573 3709 4607
rect 3709 4573 3743 4607
rect 3743 4573 3752 4607
rect 3700 4564 3752 4573
rect 5356 4607 5408 4616
rect 5356 4573 5365 4607
rect 5365 4573 5399 4607
rect 5399 4573 5408 4607
rect 7472 4641 7481 4675
rect 7481 4641 7515 4675
rect 7515 4641 7524 4675
rect 7472 4632 7524 4641
rect 5356 4564 5408 4573
rect 7564 4564 7616 4616
rect 8208 4564 8260 4616
rect 8668 4632 8720 4684
rect 8852 4564 8904 4616
rect 9128 4632 9180 4684
rect 4896 4496 4948 4548
rect 8576 4496 8628 4548
rect 9128 4496 9180 4548
rect 4252 4428 4304 4480
rect 4804 4471 4856 4480
rect 4804 4437 4813 4471
rect 4813 4437 4847 4471
rect 4847 4437 4856 4471
rect 4804 4428 4856 4437
rect 5356 4428 5408 4480
rect 8484 4428 8536 4480
rect 9496 4632 9548 4684
rect 12348 4700 12400 4752
rect 15568 4768 15620 4820
rect 16396 4768 16448 4820
rect 17868 4768 17920 4820
rect 13084 4700 13136 4752
rect 14096 4700 14148 4752
rect 14648 4743 14700 4752
rect 14648 4709 14657 4743
rect 14657 4709 14691 4743
rect 14691 4709 14700 4743
rect 14648 4700 14700 4709
rect 9680 4564 9732 4616
rect 10692 4632 10744 4684
rect 10876 4675 10928 4684
rect 10876 4641 10885 4675
rect 10885 4641 10919 4675
rect 10919 4641 10928 4675
rect 10876 4632 10928 4641
rect 10324 4607 10376 4616
rect 10324 4573 10333 4607
rect 10333 4573 10367 4607
rect 10367 4573 10376 4607
rect 10324 4564 10376 4573
rect 10784 4564 10836 4616
rect 11152 4564 11204 4616
rect 11980 4564 12032 4616
rect 9588 4496 9640 4548
rect 14004 4632 14056 4684
rect 12624 4564 12676 4616
rect 14740 4607 14792 4616
rect 14740 4573 14749 4607
rect 14749 4573 14783 4607
rect 14783 4573 14792 4607
rect 14740 4564 14792 4573
rect 13912 4496 13964 4548
rect 15476 4700 15528 4752
rect 16672 4700 16724 4752
rect 15108 4632 15160 4684
rect 17132 4632 17184 4684
rect 18236 4632 18288 4684
rect 19156 4700 19208 4752
rect 15200 4564 15252 4616
rect 15476 4607 15528 4616
rect 15476 4573 15485 4607
rect 15485 4573 15519 4607
rect 15519 4573 15528 4607
rect 15476 4564 15528 4573
rect 18144 4607 18196 4616
rect 18144 4573 18153 4607
rect 18153 4573 18187 4607
rect 18187 4573 18196 4607
rect 18144 4564 18196 4573
rect 18328 4607 18380 4616
rect 18328 4573 18337 4607
rect 18337 4573 18371 4607
rect 18371 4573 18380 4607
rect 18328 4564 18380 4573
rect 19524 4632 19576 4684
rect 19708 4675 19760 4684
rect 19708 4641 19717 4675
rect 19717 4641 19751 4675
rect 19751 4641 19760 4675
rect 19708 4632 19760 4641
rect 19432 4564 19484 4616
rect 16580 4496 16632 4548
rect 18236 4496 18288 4548
rect 10416 4428 10468 4480
rect 10692 4428 10744 4480
rect 10784 4428 10836 4480
rect 11152 4471 11204 4480
rect 11152 4437 11161 4471
rect 11161 4437 11195 4471
rect 11195 4437 11204 4471
rect 11152 4428 11204 4437
rect 12992 4428 13044 4480
rect 13728 4428 13780 4480
rect 13820 4428 13872 4480
rect 14188 4471 14240 4480
rect 14188 4437 14197 4471
rect 14197 4437 14231 4471
rect 14231 4437 14240 4471
rect 16948 4471 17000 4480
rect 14188 4428 14240 4437
rect 16948 4437 16957 4471
rect 16957 4437 16991 4471
rect 16991 4437 17000 4471
rect 16948 4428 17000 4437
rect 19984 4496 20036 4548
rect 19432 4428 19484 4480
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 4575 4326 4627 4378
rect 4639 4326 4691 4378
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 18308 4326 18360 4378
rect 18372 4326 18424 4378
rect 18436 4326 18488 4378
rect 18500 4326 18552 4378
rect 3700 4224 3752 4276
rect 4252 4224 4304 4276
rect 2412 4131 2464 4140
rect 2412 4097 2421 4131
rect 2421 4097 2455 4131
rect 2455 4097 2464 4131
rect 2412 4088 2464 4097
rect 2780 4156 2832 4208
rect 4712 4156 4764 4208
rect 4988 4156 5040 4208
rect 5172 4224 5224 4276
rect 6644 4224 6696 4276
rect 7104 4224 7156 4276
rect 5448 4156 5500 4208
rect 8760 4224 8812 4276
rect 12256 4224 12308 4276
rect 15108 4267 15160 4276
rect 4160 4088 4212 4140
rect 5264 4088 5316 4140
rect 5356 4088 5408 4140
rect 6276 4131 6328 4140
rect 6276 4097 6285 4131
rect 6285 4097 6319 4131
rect 6319 4097 6328 4131
rect 6276 4088 6328 4097
rect 9496 4156 9548 4208
rect 9772 4156 9824 4208
rect 10048 4156 10100 4208
rect 8300 4088 8352 4140
rect 8944 4088 8996 4140
rect 9128 4131 9180 4140
rect 9128 4097 9137 4131
rect 9137 4097 9171 4131
rect 9171 4097 9180 4131
rect 9128 4088 9180 4097
rect 10508 4156 10560 4208
rect 11704 4156 11756 4208
rect 12348 4156 12400 4208
rect 12532 4156 12584 4208
rect 12716 4156 12768 4208
rect 12900 4199 12952 4208
rect 12900 4165 12909 4199
rect 12909 4165 12943 4199
rect 12943 4165 12952 4199
rect 12900 4156 12952 4165
rect 13268 4156 13320 4208
rect 15108 4233 15117 4267
rect 15117 4233 15151 4267
rect 15151 4233 15160 4267
rect 15108 4224 15160 4233
rect 17500 4267 17552 4276
rect 17500 4233 17509 4267
rect 17509 4233 17543 4267
rect 17543 4233 17552 4267
rect 17500 4224 17552 4233
rect 18788 4224 18840 4276
rect 19432 4267 19484 4276
rect 19432 4233 19441 4267
rect 19441 4233 19475 4267
rect 19475 4233 19484 4267
rect 19432 4224 19484 4233
rect 19708 4224 19760 4276
rect 2872 4020 2924 4072
rect 7012 4020 7064 4072
rect 7748 4020 7800 4072
rect 9496 4020 9548 4072
rect 9680 4020 9732 4072
rect 4252 3952 4304 4004
rect 5448 3995 5500 4004
rect 5448 3961 5457 3995
rect 5457 3961 5491 3995
rect 5491 3961 5500 3995
rect 5448 3952 5500 3961
rect 5908 3952 5960 4004
rect 1676 3884 1728 3936
rect 2320 3927 2372 3936
rect 2320 3893 2329 3927
rect 2329 3893 2363 3927
rect 2363 3893 2372 3927
rect 2320 3884 2372 3893
rect 4988 3927 5040 3936
rect 4988 3893 4997 3927
rect 4997 3893 5031 3927
rect 5031 3893 5040 3927
rect 4988 3884 5040 3893
rect 5264 3884 5316 3936
rect 5816 3927 5868 3936
rect 5816 3893 5825 3927
rect 5825 3893 5859 3927
rect 5859 3893 5868 3927
rect 5816 3884 5868 3893
rect 6460 3884 6512 3936
rect 6644 3952 6696 4004
rect 8208 3952 8260 4004
rect 11980 4088 12032 4140
rect 13820 4156 13872 4208
rect 14464 4131 14516 4140
rect 14464 4097 14473 4131
rect 14473 4097 14507 4131
rect 14507 4097 14516 4131
rect 14464 4088 14516 4097
rect 9864 4020 9916 4072
rect 10600 4020 10652 4072
rect 11152 4020 11204 4072
rect 13360 4063 13412 4072
rect 13360 4029 13369 4063
rect 13369 4029 13403 4063
rect 13403 4029 13412 4063
rect 13360 4020 13412 4029
rect 14188 4020 14240 4072
rect 14556 4020 14608 4072
rect 15476 4156 15528 4208
rect 15568 4131 15620 4140
rect 15568 4097 15577 4131
rect 15577 4097 15611 4131
rect 15611 4097 15620 4131
rect 15568 4088 15620 4097
rect 15844 4088 15896 4140
rect 16028 4088 16080 4140
rect 19524 4088 19576 4140
rect 21548 4088 21600 4140
rect 22744 4088 22796 4140
rect 16396 4063 16448 4072
rect 7472 3884 7524 3936
rect 7564 3884 7616 3936
rect 8852 3884 8904 3936
rect 8944 3884 8996 3936
rect 9496 3884 9548 3936
rect 12808 3952 12860 4004
rect 9772 3884 9824 3936
rect 11244 3884 11296 3936
rect 12440 3884 12492 3936
rect 12900 3884 12952 3936
rect 16396 4029 16430 4063
rect 16430 4029 16448 4063
rect 16396 4020 16448 4029
rect 16672 4020 16724 4072
rect 17960 4020 18012 4072
rect 19432 4020 19484 4072
rect 20720 4020 20772 4072
rect 17868 3995 17920 4004
rect 13084 3884 13136 3936
rect 14188 3927 14240 3936
rect 14188 3893 14197 3927
rect 14197 3893 14231 3927
rect 14231 3893 14240 3927
rect 14188 3884 14240 3893
rect 15476 3927 15528 3936
rect 15476 3893 15485 3927
rect 15485 3893 15519 3927
rect 15519 3893 15528 3927
rect 15476 3884 15528 3893
rect 16120 3884 16172 3936
rect 17868 3961 17877 3995
rect 17877 3961 17911 3995
rect 17911 3961 17920 3995
rect 17868 3952 17920 3961
rect 20628 3952 20680 4004
rect 22284 3952 22336 4004
rect 17960 3884 18012 3936
rect 18052 3884 18104 3936
rect 19340 3884 19392 3936
rect 19708 3884 19760 3936
rect 19800 3884 19852 3936
rect 19984 3927 20036 3936
rect 19984 3893 19993 3927
rect 19993 3893 20027 3927
rect 20027 3893 20036 3927
rect 19984 3884 20036 3893
rect 7912 3782 7964 3834
rect 7976 3782 8028 3834
rect 8040 3782 8092 3834
rect 8104 3782 8156 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 15035 3782 15087 3834
rect 2320 3723 2372 3732
rect 2320 3689 2329 3723
rect 2329 3689 2363 3723
rect 2363 3689 2372 3723
rect 2320 3680 2372 3689
rect 3516 3680 3568 3732
rect 4804 3680 4856 3732
rect 5908 3723 5960 3732
rect 2504 3544 2556 3596
rect 3792 3612 3844 3664
rect 3056 3544 3108 3596
rect 3700 3544 3752 3596
rect 4160 3612 4212 3664
rect 5908 3689 5917 3723
rect 5917 3689 5951 3723
rect 5951 3689 5960 3723
rect 5908 3680 5960 3689
rect 7380 3680 7432 3732
rect 8208 3680 8260 3732
rect 8668 3680 8720 3732
rect 6736 3612 6788 3664
rect 6920 3612 6972 3664
rect 8576 3655 8628 3664
rect 8576 3621 8585 3655
rect 8585 3621 8619 3655
rect 8619 3621 8628 3655
rect 8576 3612 8628 3621
rect 8944 3612 8996 3664
rect 7472 3544 7524 3596
rect 9680 3680 9732 3732
rect 9864 3680 9916 3732
rect 10232 3680 10284 3732
rect 10968 3680 11020 3732
rect 11152 3680 11204 3732
rect 9220 3655 9272 3664
rect 9220 3621 9229 3655
rect 9229 3621 9263 3655
rect 9263 3621 9272 3655
rect 9220 3612 9272 3621
rect 9404 3612 9456 3664
rect 2688 3408 2740 3460
rect 3516 3340 3568 3392
rect 5908 3476 5960 3528
rect 6644 3476 6696 3528
rect 10968 3544 11020 3596
rect 12440 3612 12492 3664
rect 12624 3612 12676 3664
rect 12716 3612 12768 3664
rect 12992 3680 13044 3732
rect 14096 3680 14148 3732
rect 15200 3680 15252 3732
rect 16764 3680 16816 3732
rect 18144 3680 18196 3732
rect 19800 3723 19852 3732
rect 19800 3689 19809 3723
rect 19809 3689 19843 3723
rect 19843 3689 19852 3723
rect 19800 3680 19852 3689
rect 20260 3680 20312 3732
rect 14464 3612 14516 3664
rect 15292 3612 15344 3664
rect 12348 3544 12400 3596
rect 13360 3587 13412 3596
rect 13360 3553 13369 3587
rect 13369 3553 13403 3587
rect 13403 3553 13412 3587
rect 14188 3587 14240 3596
rect 13360 3544 13412 3553
rect 14188 3553 14197 3587
rect 14197 3553 14231 3587
rect 14231 3553 14240 3587
rect 14188 3544 14240 3553
rect 14648 3587 14700 3596
rect 14648 3553 14657 3587
rect 14657 3553 14691 3587
rect 14691 3553 14700 3587
rect 14648 3544 14700 3553
rect 15108 3544 15160 3596
rect 16120 3587 16172 3596
rect 16120 3553 16129 3587
rect 16129 3553 16163 3587
rect 16163 3553 16172 3587
rect 16120 3544 16172 3553
rect 4252 3340 4304 3392
rect 6092 3340 6144 3392
rect 9496 3476 9548 3528
rect 10692 3476 10744 3528
rect 13820 3476 13872 3528
rect 15752 3519 15804 3528
rect 15752 3485 15761 3519
rect 15761 3485 15795 3519
rect 15795 3485 15804 3519
rect 15752 3476 15804 3485
rect 15844 3519 15896 3528
rect 15844 3485 15853 3519
rect 15853 3485 15887 3519
rect 15887 3485 15896 3519
rect 17500 3544 17552 3596
rect 17868 3544 17920 3596
rect 19340 3587 19392 3596
rect 19340 3553 19349 3587
rect 19349 3553 19383 3587
rect 19383 3553 19392 3587
rect 19340 3544 19392 3553
rect 16672 3519 16724 3528
rect 15844 3476 15896 3485
rect 16672 3485 16681 3519
rect 16681 3485 16715 3519
rect 16715 3485 16724 3519
rect 16672 3476 16724 3485
rect 18604 3519 18656 3528
rect 18604 3485 18613 3519
rect 18613 3485 18647 3519
rect 18647 3485 18656 3519
rect 18604 3476 18656 3485
rect 18788 3519 18840 3528
rect 18788 3485 18797 3519
rect 18797 3485 18831 3519
rect 18831 3485 18840 3519
rect 18788 3476 18840 3485
rect 19524 3519 19576 3528
rect 19524 3485 19533 3519
rect 19533 3485 19567 3519
rect 19567 3485 19576 3519
rect 19524 3476 19576 3485
rect 7840 3408 7892 3460
rect 7012 3340 7064 3392
rect 8668 3340 8720 3392
rect 9312 3340 9364 3392
rect 9588 3340 9640 3392
rect 10416 3340 10468 3392
rect 11244 3340 11296 3392
rect 15936 3408 15988 3460
rect 16028 3408 16080 3460
rect 12992 3383 13044 3392
rect 12992 3349 13001 3383
rect 13001 3349 13035 3383
rect 13035 3349 13044 3383
rect 12992 3340 13044 3349
rect 13912 3340 13964 3392
rect 14740 3340 14792 3392
rect 15292 3383 15344 3392
rect 15292 3349 15301 3383
rect 15301 3349 15335 3383
rect 15335 3349 15344 3383
rect 15292 3340 15344 3349
rect 15752 3340 15804 3392
rect 18052 3383 18104 3392
rect 18052 3349 18061 3383
rect 18061 3349 18095 3383
rect 18095 3349 18104 3383
rect 18052 3340 18104 3349
rect 18144 3383 18196 3392
rect 18144 3349 18153 3383
rect 18153 3349 18187 3383
rect 18187 3349 18196 3383
rect 18144 3340 18196 3349
rect 18604 3340 18656 3392
rect 20352 3383 20404 3392
rect 20352 3349 20361 3383
rect 20361 3349 20395 3383
rect 20395 3349 20404 3383
rect 20352 3340 20404 3349
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 4575 3238 4627 3290
rect 4639 3238 4691 3290
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 18308 3238 18360 3290
rect 18372 3238 18424 3290
rect 18436 3238 18488 3290
rect 18500 3238 18552 3290
rect 2504 3179 2556 3188
rect 2504 3145 2513 3179
rect 2513 3145 2547 3179
rect 2547 3145 2556 3179
rect 2504 3136 2556 3145
rect 2872 3136 2924 3188
rect 3056 3136 3108 3188
rect 3700 3136 3752 3188
rect 5540 3136 5592 3188
rect 5908 3179 5960 3188
rect 5908 3145 5917 3179
rect 5917 3145 5951 3179
rect 5951 3145 5960 3179
rect 5908 3136 5960 3145
rect 6552 3136 6604 3188
rect 6828 3136 6880 3188
rect 7748 3136 7800 3188
rect 9128 3136 9180 3188
rect 12348 3136 12400 3188
rect 15108 3136 15160 3188
rect 17132 3179 17184 3188
rect 17132 3145 17141 3179
rect 17141 3145 17175 3179
rect 17175 3145 17184 3179
rect 17132 3136 17184 3145
rect 19340 3136 19392 3188
rect 19524 3136 19576 3188
rect 19708 3136 19760 3188
rect 3792 3068 3844 3120
rect 3516 3000 3568 3052
rect 6920 3068 6972 3120
rect 10968 3068 11020 3120
rect 12440 3068 12492 3120
rect 13452 3068 13504 3120
rect 18972 3068 19024 3120
rect 19064 3068 19116 3120
rect 20904 3068 20956 3120
rect 9588 3043 9640 3052
rect 9588 3009 9597 3043
rect 9597 3009 9631 3043
rect 9631 3009 9640 3043
rect 9588 3000 9640 3009
rect 2780 2932 2832 2984
rect 3424 2932 3476 2984
rect 3700 2975 3752 2984
rect 3700 2941 3709 2975
rect 3709 2941 3743 2975
rect 3743 2941 3752 2975
rect 3700 2932 3752 2941
rect 4160 2932 4212 2984
rect 6368 2975 6420 2984
rect 6368 2941 6377 2975
rect 6377 2941 6411 2975
rect 6411 2941 6420 2975
rect 6368 2932 6420 2941
rect 7012 2975 7064 2984
rect 7012 2941 7021 2975
rect 7021 2941 7055 2975
rect 7055 2941 7064 2975
rect 7012 2932 7064 2941
rect 7840 2932 7892 2984
rect 8484 2975 8536 2984
rect 8484 2941 8493 2975
rect 8493 2941 8527 2975
rect 8527 2941 8536 2975
rect 8484 2932 8536 2941
rect 9128 2932 9180 2984
rect 3516 2864 3568 2916
rect 4068 2864 4120 2916
rect 4712 2864 4764 2916
rect 6736 2864 6788 2916
rect 6920 2907 6972 2916
rect 6920 2873 6929 2907
rect 6929 2873 6963 2907
rect 6963 2873 6972 2907
rect 6920 2864 6972 2873
rect 7564 2864 7616 2916
rect 9036 2864 9088 2916
rect 12348 2932 12400 2984
rect 13544 3000 13596 3052
rect 14188 3000 14240 3052
rect 16856 3000 16908 3052
rect 18052 3000 18104 3052
rect 18788 3043 18840 3052
rect 18788 3009 18797 3043
rect 18797 3009 18831 3043
rect 18831 3009 18840 3043
rect 18788 3000 18840 3009
rect 14372 2932 14424 2984
rect 15384 2975 15436 2984
rect 15384 2941 15393 2975
rect 15393 2941 15427 2975
rect 15427 2941 15436 2975
rect 15384 2932 15436 2941
rect 15936 2975 15988 2984
rect 15936 2941 15945 2975
rect 15945 2941 15979 2975
rect 15979 2941 15988 2975
rect 15936 2932 15988 2941
rect 16948 2932 17000 2984
rect 18144 2932 18196 2984
rect 9588 2864 9640 2916
rect 12532 2864 12584 2916
rect 12716 2907 12768 2916
rect 12716 2873 12750 2907
rect 12750 2873 12768 2907
rect 12716 2864 12768 2873
rect 12900 2864 12952 2916
rect 15568 2864 15620 2916
rect 17224 2864 17276 2916
rect 2872 2839 2924 2848
rect 2872 2805 2881 2839
rect 2881 2805 2915 2839
rect 2915 2805 2924 2839
rect 2872 2796 2924 2805
rect 5448 2796 5500 2848
rect 9404 2839 9456 2848
rect 9404 2805 9413 2839
rect 9413 2805 9447 2839
rect 9447 2805 9456 2839
rect 9404 2796 9456 2805
rect 11796 2796 11848 2848
rect 13084 2796 13136 2848
rect 13728 2796 13780 2848
rect 15476 2796 15528 2848
rect 16488 2796 16540 2848
rect 18604 2839 18656 2848
rect 18604 2805 18613 2839
rect 18613 2805 18647 2839
rect 18647 2805 18656 2839
rect 18604 2796 18656 2805
rect 20260 3000 20312 3052
rect 19800 2975 19852 2984
rect 19800 2941 19809 2975
rect 19809 2941 19843 2975
rect 19843 2941 19852 2975
rect 19800 2932 19852 2941
rect 19984 2932 20036 2984
rect 20076 2932 20128 2984
rect 19616 2864 19668 2916
rect 19892 2864 19944 2916
rect 19340 2796 19392 2848
rect 19800 2796 19852 2848
rect 20260 2796 20312 2848
rect 20628 2796 20680 2848
rect 7912 2694 7964 2746
rect 7976 2694 8028 2746
rect 8040 2694 8092 2746
rect 8104 2694 8156 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 15035 2694 15087 2746
rect 2872 2592 2924 2644
rect 4160 2635 4212 2644
rect 4160 2601 4169 2635
rect 4169 2601 4203 2635
rect 4203 2601 4212 2635
rect 4160 2592 4212 2601
rect 4896 2592 4948 2644
rect 5816 2592 5868 2644
rect 3608 2456 3660 2508
rect 5080 2524 5132 2576
rect 5540 2524 5592 2576
rect 6368 2592 6420 2644
rect 9404 2592 9456 2644
rect 9772 2635 9824 2644
rect 9772 2601 9781 2635
rect 9781 2601 9815 2635
rect 9815 2601 9824 2635
rect 9772 2592 9824 2601
rect 10140 2592 10192 2644
rect 6920 2524 6972 2576
rect 7564 2524 7616 2576
rect 4988 2456 5040 2508
rect 6368 2499 6420 2508
rect 6368 2465 6377 2499
rect 6377 2465 6411 2499
rect 6411 2465 6420 2499
rect 6368 2456 6420 2465
rect 7748 2499 7800 2508
rect 7748 2465 7757 2499
rect 7757 2465 7791 2499
rect 7791 2465 7800 2499
rect 7748 2456 7800 2465
rect 9680 2524 9732 2576
rect 9956 2524 10008 2576
rect 3240 2388 3292 2440
rect 3700 2320 3752 2372
rect 4712 2388 4764 2440
rect 4896 2388 4948 2440
rect 4252 2320 4304 2372
rect 5448 2320 5500 2372
rect 7196 2388 7248 2440
rect 8668 2431 8720 2440
rect 8668 2397 8677 2431
rect 8677 2397 8711 2431
rect 8711 2397 8720 2431
rect 8668 2388 8720 2397
rect 9772 2456 9824 2508
rect 10140 2499 10192 2508
rect 10140 2465 10149 2499
rect 10149 2465 10183 2499
rect 10183 2465 10192 2499
rect 10140 2456 10192 2465
rect 11152 2592 11204 2644
rect 12532 2592 12584 2644
rect 12992 2592 13044 2644
rect 16212 2592 16264 2644
rect 11796 2456 11848 2508
rect 12900 2456 12952 2508
rect 10416 2431 10468 2440
rect 10416 2397 10425 2431
rect 10425 2397 10459 2431
rect 10459 2397 10468 2431
rect 10416 2388 10468 2397
rect 12624 2388 12676 2440
rect 12716 2388 12768 2440
rect 13820 2499 13872 2508
rect 13820 2465 13829 2499
rect 13829 2465 13863 2499
rect 13863 2465 13872 2499
rect 13820 2456 13872 2465
rect 14188 2499 14240 2508
rect 14188 2465 14197 2499
rect 14197 2465 14231 2499
rect 14231 2465 14240 2499
rect 14188 2456 14240 2465
rect 14556 2499 14608 2508
rect 14556 2465 14565 2499
rect 14565 2465 14599 2499
rect 14599 2465 14608 2499
rect 14556 2456 14608 2465
rect 14648 2456 14700 2508
rect 13912 2388 13964 2440
rect 15568 2456 15620 2508
rect 17684 2592 17736 2644
rect 19524 2592 19576 2644
rect 20076 2635 20128 2644
rect 20076 2601 20085 2635
rect 20085 2601 20119 2635
rect 20119 2601 20128 2635
rect 20076 2592 20128 2601
rect 16396 2524 16448 2576
rect 16856 2499 16908 2508
rect 16856 2465 16865 2499
rect 16865 2465 16899 2499
rect 16899 2465 16908 2499
rect 16856 2456 16908 2465
rect 17224 2499 17276 2508
rect 17224 2465 17233 2499
rect 17233 2465 17267 2499
rect 17267 2465 17276 2499
rect 17224 2456 17276 2465
rect 15660 2388 15712 2440
rect 16396 2388 16448 2440
rect 18604 2456 18656 2508
rect 18696 2499 18748 2508
rect 18696 2465 18705 2499
rect 18705 2465 18739 2499
rect 18739 2465 18748 2499
rect 18696 2456 18748 2465
rect 3148 2295 3200 2304
rect 3148 2261 3157 2295
rect 3157 2261 3191 2295
rect 3191 2261 3200 2295
rect 3148 2252 3200 2261
rect 3608 2295 3660 2304
rect 3608 2261 3617 2295
rect 3617 2261 3651 2295
rect 3651 2261 3660 2295
rect 3608 2252 3660 2261
rect 3792 2295 3844 2304
rect 3792 2261 3801 2295
rect 3801 2261 3835 2295
rect 3835 2261 3844 2295
rect 3792 2252 3844 2261
rect 4896 2252 4948 2304
rect 5356 2252 5408 2304
rect 6736 2320 6788 2372
rect 9772 2320 9824 2372
rect 13544 2320 13596 2372
rect 15476 2320 15528 2372
rect 17316 2320 17368 2372
rect 19340 2320 19392 2372
rect 7196 2295 7248 2304
rect 7196 2261 7205 2295
rect 7205 2261 7239 2295
rect 7239 2261 7248 2295
rect 7196 2252 7248 2261
rect 9036 2295 9088 2304
rect 9036 2261 9045 2295
rect 9045 2261 9079 2295
rect 9079 2261 9088 2295
rect 9036 2252 9088 2261
rect 9956 2252 10008 2304
rect 10140 2252 10192 2304
rect 10784 2252 10836 2304
rect 12716 2252 12768 2304
rect 13084 2252 13136 2304
rect 14096 2252 14148 2304
rect 14464 2252 14516 2304
rect 15200 2295 15252 2304
rect 15200 2261 15209 2295
rect 15209 2261 15243 2295
rect 15243 2261 15252 2295
rect 15200 2252 15252 2261
rect 15660 2295 15712 2304
rect 15660 2261 15669 2295
rect 15669 2261 15703 2295
rect 15703 2261 15712 2295
rect 15660 2252 15712 2261
rect 16028 2295 16080 2304
rect 16028 2261 16037 2295
rect 16037 2261 16071 2295
rect 16071 2261 16080 2295
rect 16028 2252 16080 2261
rect 17592 2295 17644 2304
rect 17592 2261 17601 2295
rect 17601 2261 17635 2295
rect 17635 2261 17644 2295
rect 17592 2252 17644 2261
rect 18604 2252 18656 2304
rect 18972 2252 19024 2304
rect 19524 2295 19576 2304
rect 19524 2261 19533 2295
rect 19533 2261 19567 2295
rect 19567 2261 19576 2295
rect 19524 2252 19576 2261
rect 19892 2295 19944 2304
rect 19892 2261 19901 2295
rect 19901 2261 19935 2295
rect 19935 2261 19944 2295
rect 19892 2252 19944 2261
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 4575 2150 4627 2202
rect 4639 2150 4691 2202
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 18308 2150 18360 2202
rect 18372 2150 18424 2202
rect 18436 2150 18488 2202
rect 18500 2150 18552 2202
rect 1032 2048 1084 2100
rect 6920 2048 6972 2100
rect 9220 2048 9272 2100
rect 9404 2048 9456 2100
rect 6368 1980 6420 2032
rect 12256 1980 12308 2032
rect 12624 1980 12676 2032
rect 14556 1980 14608 2032
rect 2688 1912 2740 1964
rect 8668 1912 8720 1964
rect 1860 1844 1912 1896
rect 7196 1844 7248 1896
rect 9956 1776 10008 1828
rect 572 1708 624 1760
rect 9312 1708 9364 1760
rect 204 1640 256 1692
rect 9036 1640 9088 1692
rect 3056 1572 3108 1624
rect 7472 1572 7524 1624
rect 1400 1436 1452 1488
rect 10140 1436 10192 1488
<< metal2 >>
rect 202 22200 258 23000
rect 570 22200 626 23000
rect 938 22200 994 23000
rect 1306 22200 1362 23000
rect 1674 22200 1730 23000
rect 2042 22200 2098 23000
rect 2502 22200 2558 23000
rect 2870 22200 2926 23000
rect 3238 22200 3294 23000
rect 3514 22672 3570 22681
rect 3514 22607 3570 22616
rect 216 19242 244 22200
rect 204 19236 256 19242
rect 204 19178 256 19184
rect 584 18902 612 22200
rect 572 18896 624 18902
rect 572 18838 624 18844
rect 952 18290 980 22200
rect 1320 18601 1348 22200
rect 1688 18698 1716 22200
rect 1950 20224 2006 20233
rect 1950 20159 2006 20168
rect 1858 19680 1914 19689
rect 1858 19615 1914 19624
rect 1872 18970 1900 19615
rect 1964 19514 1992 20159
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 1860 18964 1912 18970
rect 1860 18906 1912 18912
rect 2056 18816 2084 22200
rect 2136 19236 2188 19242
rect 2136 19178 2188 19184
rect 2148 19009 2176 19178
rect 2134 19000 2190 19009
rect 2134 18935 2190 18944
rect 2228 18828 2280 18834
rect 2056 18788 2228 18816
rect 2228 18770 2280 18776
rect 2412 18760 2464 18766
rect 2412 18702 2464 18708
rect 1676 18692 1728 18698
rect 1676 18634 1728 18640
rect 1306 18592 1362 18601
rect 1306 18527 1362 18536
rect 1582 18456 1638 18465
rect 1582 18391 1638 18400
rect 940 18284 992 18290
rect 940 18226 992 18232
rect 1596 17882 1624 18391
rect 2136 18216 2188 18222
rect 2136 18158 2188 18164
rect 1952 18080 2004 18086
rect 1950 18048 1952 18057
rect 2004 18048 2006 18057
rect 1950 17983 2006 17992
rect 1584 17876 1636 17882
rect 1584 17818 1636 17824
rect 2148 17814 2176 18158
rect 2136 17808 2188 17814
rect 2424 17785 2452 18702
rect 2516 18630 2544 22200
rect 2884 20058 2912 22200
rect 2872 20052 2924 20058
rect 2872 19994 2924 20000
rect 2594 19272 2650 19281
rect 2594 19207 2650 19216
rect 2504 18624 2556 18630
rect 2502 18592 2504 18601
rect 2556 18592 2558 18601
rect 2502 18527 2558 18536
rect 2608 18086 2636 19207
rect 3056 19168 3108 19174
rect 2962 19136 3018 19145
rect 3056 19110 3108 19116
rect 2962 19071 3018 19080
rect 2778 18864 2834 18873
rect 2778 18799 2834 18808
rect 2872 18828 2924 18834
rect 2688 18760 2740 18766
rect 2688 18702 2740 18708
rect 2700 18222 2728 18702
rect 2792 18426 2820 18799
rect 2976 18816 3004 19071
rect 2924 18788 3004 18816
rect 2872 18770 2924 18776
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 2688 18216 2740 18222
rect 2688 18158 2740 18164
rect 2596 18080 2648 18086
rect 2596 18022 2648 18028
rect 2136 17750 2188 17756
rect 2410 17776 2466 17785
rect 1400 17740 1452 17746
rect 2410 17711 2466 17720
rect 1400 17682 1452 17688
rect 1412 16998 1440 17682
rect 2136 17672 2188 17678
rect 1674 17640 1730 17649
rect 2136 17614 2188 17620
rect 2596 17672 2648 17678
rect 2596 17614 2648 17620
rect 1674 17575 1730 17584
rect 1582 17232 1638 17241
rect 1582 17167 1638 17176
rect 1400 16992 1452 16998
rect 1400 16934 1452 16940
rect 1596 16250 1624 17167
rect 1688 16658 1716 17575
rect 1676 16652 1728 16658
rect 1676 16594 1728 16600
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1766 16144 1822 16153
rect 1766 16079 1822 16088
rect 1780 16046 1808 16079
rect 1400 16040 1452 16046
rect 1400 15982 1452 15988
rect 1768 16040 1820 16046
rect 1768 15982 1820 15988
rect 1412 15638 1440 15982
rect 1952 15904 2004 15910
rect 1950 15872 1952 15881
rect 2004 15872 2006 15881
rect 1950 15807 2006 15816
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 1400 15632 1452 15638
rect 1400 15574 1452 15580
rect 1584 15360 1636 15366
rect 1584 15302 1636 15308
rect 1596 14958 1624 15302
rect 1584 14952 1636 14958
rect 1584 14894 1636 14900
rect 1688 14482 1716 15642
rect 1768 15088 1820 15094
rect 1766 15056 1768 15065
rect 1820 15056 1822 15065
rect 1766 14991 1822 15000
rect 1858 14648 1914 14657
rect 1858 14583 1860 14592
rect 1912 14583 1914 14592
rect 2042 14648 2098 14657
rect 2042 14583 2098 14592
rect 1860 14554 1912 14560
rect 2056 14482 2084 14583
rect 1676 14476 1728 14482
rect 1676 14418 1728 14424
rect 2044 14476 2096 14482
rect 2044 14418 2096 14424
rect 1582 14376 1638 14385
rect 1582 14311 1638 14320
rect 1400 14272 1452 14278
rect 1400 14214 1452 14220
rect 1412 9897 1440 14214
rect 1596 13870 1624 14311
rect 1766 14240 1822 14249
rect 1766 14175 1822 14184
rect 1780 14074 1808 14175
rect 1768 14068 1820 14074
rect 1768 14010 1820 14016
rect 1584 13864 1636 13870
rect 1584 13806 1636 13812
rect 1768 13388 1820 13394
rect 1768 13330 1820 13336
rect 1492 13320 1544 13326
rect 1492 13262 1544 13268
rect 1504 12306 1532 13262
rect 1674 12880 1730 12889
rect 1674 12815 1730 12824
rect 1688 12442 1716 12815
rect 1780 12442 1808 13330
rect 2148 13274 2176 17614
rect 2228 17536 2280 17542
rect 2228 17478 2280 17484
rect 2412 17536 2464 17542
rect 2412 17478 2464 17484
rect 2240 17134 2268 17478
rect 2424 17202 2452 17478
rect 2412 17196 2464 17202
rect 2412 17138 2464 17144
rect 2228 17128 2280 17134
rect 2228 17070 2280 17076
rect 2504 16720 2556 16726
rect 2504 16662 2556 16668
rect 2516 16454 2544 16662
rect 2608 16658 2636 17614
rect 2700 17218 2728 18158
rect 2976 18154 3004 18788
rect 3068 18358 3096 19110
rect 3146 18592 3202 18601
rect 3146 18527 3202 18536
rect 3056 18352 3108 18358
rect 3056 18294 3108 18300
rect 3160 18222 3188 18527
rect 3148 18216 3200 18222
rect 3148 18158 3200 18164
rect 2964 18148 3016 18154
rect 2964 18090 3016 18096
rect 2872 18080 2924 18086
rect 2870 18048 2872 18057
rect 3056 18080 3108 18086
rect 2924 18048 2926 18057
rect 3056 18022 3108 18028
rect 2870 17983 2926 17992
rect 3068 17882 3096 18022
rect 3056 17876 3108 17882
rect 3056 17818 3108 17824
rect 2872 17604 2924 17610
rect 2872 17546 2924 17552
rect 2700 17190 2820 17218
rect 2688 17128 2740 17134
rect 2688 17070 2740 17076
rect 2700 16726 2728 17070
rect 2792 16969 2820 17190
rect 2778 16960 2834 16969
rect 2778 16895 2834 16904
rect 2778 16824 2834 16833
rect 2778 16759 2834 16768
rect 2688 16720 2740 16726
rect 2688 16662 2740 16668
rect 2596 16652 2648 16658
rect 2596 16594 2648 16600
rect 2504 16448 2556 16454
rect 2504 16390 2556 16396
rect 2318 16280 2374 16289
rect 2318 16215 2320 16224
rect 2372 16215 2374 16224
rect 2320 16186 2372 16192
rect 2516 15570 2544 16390
rect 2608 16182 2636 16594
rect 2792 16250 2820 16759
rect 2884 16250 2912 17546
rect 3160 17513 3188 18158
rect 3252 17542 3280 22200
rect 3422 21856 3478 21865
rect 3422 21791 3478 21800
rect 3332 20052 3384 20058
rect 3332 19994 3384 20000
rect 3344 18630 3372 19994
rect 3332 18624 3384 18630
rect 3332 18566 3384 18572
rect 3436 18193 3464 21791
rect 3528 18737 3556 22607
rect 3606 22200 3662 23000
rect 3790 22264 3846 22273
rect 3514 18728 3570 18737
rect 3514 18663 3570 18672
rect 3422 18184 3478 18193
rect 3422 18119 3478 18128
rect 3240 17536 3292 17542
rect 3146 17504 3202 17513
rect 3240 17478 3292 17484
rect 3146 17439 3202 17448
rect 3620 17354 3648 22200
rect 3790 22199 3846 22208
rect 3974 22200 4030 23000
rect 4342 22200 4398 23000
rect 4802 22200 4858 23000
rect 5170 22200 5226 23000
rect 5538 22200 5594 23000
rect 5906 22200 5962 23000
rect 6274 22200 6330 23000
rect 6642 22200 6698 23000
rect 7102 22200 7158 23000
rect 7470 22200 7526 23000
rect 7838 22200 7894 23000
rect 8206 22200 8262 23000
rect 8574 22200 8630 23000
rect 8942 22200 8998 23000
rect 9402 22200 9458 23000
rect 9770 22200 9826 23000
rect 10138 22200 10194 23000
rect 10506 22200 10562 23000
rect 10874 22200 10930 23000
rect 11242 22200 11298 23000
rect 11702 22200 11758 23000
rect 12070 22200 12126 23000
rect 12438 22200 12494 23000
rect 12806 22200 12862 23000
rect 13174 22200 13230 23000
rect 13542 22200 13598 23000
rect 14002 22200 14058 23000
rect 14370 22200 14426 23000
rect 14738 22200 14794 23000
rect 15106 22200 15162 23000
rect 15474 22200 15530 23000
rect 15842 22200 15898 23000
rect 16302 22200 16358 23000
rect 16670 22200 16726 23000
rect 17038 22200 17094 23000
rect 17406 22200 17462 23000
rect 17774 22200 17830 23000
rect 18142 22200 18198 23000
rect 18602 22200 18658 23000
rect 18970 22200 19026 23000
rect 19154 22264 19210 22273
rect 3698 21448 3754 21457
rect 3698 21383 3754 21392
rect 3712 18329 3740 21383
rect 3804 18873 3832 22199
rect 3882 20632 3938 20641
rect 3882 20567 3938 20576
rect 3896 19281 3924 20567
rect 3882 19272 3938 19281
rect 3882 19207 3938 19216
rect 3790 18864 3846 18873
rect 3790 18799 3846 18808
rect 3792 18624 3844 18630
rect 3792 18566 3844 18572
rect 3698 18320 3754 18329
rect 3698 18255 3754 18264
rect 2976 17326 3648 17354
rect 2780 16244 2832 16250
rect 2780 16186 2832 16192
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 2596 16176 2648 16182
rect 2596 16118 2648 16124
rect 2608 15706 2636 16118
rect 2596 15700 2648 15706
rect 2596 15642 2648 15648
rect 2504 15564 2556 15570
rect 2504 15506 2556 15512
rect 2320 14408 2372 14414
rect 2320 14350 2372 14356
rect 2332 13394 2360 14350
rect 2516 13852 2544 15506
rect 2608 15026 2636 15642
rect 2596 15020 2648 15026
rect 2596 14962 2648 14968
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 2608 14346 2636 14758
rect 2688 14476 2740 14482
rect 2688 14418 2740 14424
rect 2596 14340 2648 14346
rect 2596 14282 2648 14288
rect 2700 14090 2728 14418
rect 2608 14062 2728 14090
rect 2608 14006 2636 14062
rect 2596 14000 2648 14006
rect 2596 13942 2648 13948
rect 2596 13864 2648 13870
rect 2516 13824 2596 13852
rect 2596 13806 2648 13812
rect 2778 13832 2834 13841
rect 2412 13524 2464 13530
rect 2412 13466 2464 13472
rect 2424 13433 2452 13466
rect 2410 13424 2466 13433
rect 2320 13388 2372 13394
rect 2410 13359 2466 13368
rect 2320 13330 2372 13336
rect 2148 13246 2360 13274
rect 1860 12776 1912 12782
rect 1860 12718 1912 12724
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 1768 12436 1820 12442
rect 1768 12378 1820 12384
rect 1492 12300 1544 12306
rect 1492 12242 1544 12248
rect 1582 12064 1638 12073
rect 1582 11999 1638 12008
rect 1596 11354 1624 11999
rect 1872 11898 1900 12718
rect 2228 12300 2280 12306
rect 2228 12242 2280 12248
rect 1860 11892 1912 11898
rect 1860 11834 1912 11840
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 1872 11218 1900 11834
rect 2136 11620 2188 11626
rect 2136 11562 2188 11568
rect 1676 11212 1728 11218
rect 1676 11154 1728 11160
rect 1860 11212 1912 11218
rect 1860 11154 1912 11160
rect 1398 9888 1454 9897
rect 1398 9823 1454 9832
rect 1308 9376 1360 9382
rect 1308 9318 1360 9324
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1320 6662 1348 9318
rect 1596 9178 1624 9318
rect 1584 9172 1636 9178
rect 1584 9114 1636 9120
rect 1688 9092 1716 11154
rect 2148 10674 2176 11562
rect 2240 10810 2268 12242
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 1860 10464 1912 10470
rect 1860 10406 1912 10412
rect 2044 10464 2096 10470
rect 2044 10406 2096 10412
rect 1872 9722 1900 10406
rect 2056 10266 2084 10406
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 1860 9716 1912 9722
rect 1860 9658 1912 9664
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 1688 9064 1900 9092
rect 1492 8968 1544 8974
rect 1492 8910 1544 8916
rect 1504 8090 1532 8910
rect 1492 8084 1544 8090
rect 1492 8026 1544 8032
rect 1308 6656 1360 6662
rect 1308 6598 1360 6604
rect 1320 4758 1348 6598
rect 1504 6186 1532 8026
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 1688 7342 1716 7822
rect 1676 7336 1728 7342
rect 1676 7278 1728 7284
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1688 6254 1716 6734
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1492 6180 1544 6186
rect 1492 6122 1544 6128
rect 1780 6118 1808 6802
rect 1768 6112 1820 6118
rect 1768 6054 1820 6060
rect 1676 5772 1728 5778
rect 1676 5714 1728 5720
rect 1400 5160 1452 5166
rect 1400 5102 1452 5108
rect 1308 4752 1360 4758
rect 1308 4694 1360 4700
rect 1032 2100 1084 2106
rect 1032 2042 1084 2048
rect 572 1760 624 1766
rect 572 1702 624 1708
rect 204 1692 256 1698
rect 204 1634 256 1640
rect 216 800 244 1634
rect 584 800 612 1702
rect 1044 800 1072 2042
rect 1320 1465 1348 4694
rect 1412 4690 1440 5102
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 1688 3942 1716 5714
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 1780 2281 1808 6054
rect 1872 5846 1900 9064
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 1964 6730 1992 8366
rect 2044 8356 2096 8362
rect 2044 8298 2096 8304
rect 1952 6724 2004 6730
rect 1952 6666 2004 6672
rect 2056 6458 2084 8298
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 1860 5840 1912 5846
rect 1860 5782 1912 5788
rect 1766 2272 1822 2281
rect 1766 2207 1822 2216
rect 1860 1896 1912 1902
rect 2148 1873 2176 9318
rect 2332 5914 2360 13246
rect 2608 12782 2636 13806
rect 2778 13767 2834 13776
rect 2792 13530 2820 13767
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2596 12776 2648 12782
rect 2596 12718 2648 12724
rect 2504 12708 2556 12714
rect 2504 12650 2556 12656
rect 2516 12238 2544 12650
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 2516 11898 2544 12174
rect 2688 12164 2740 12170
rect 2688 12106 2740 12112
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 2700 11626 2728 12106
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2688 11620 2740 11626
rect 2688 11562 2740 11568
rect 2700 11354 2728 11562
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2688 10532 2740 10538
rect 2688 10474 2740 10480
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 2424 9722 2452 10066
rect 2504 10056 2556 10062
rect 2504 9998 2556 10004
rect 2412 9716 2464 9722
rect 2412 9658 2464 9664
rect 2516 9178 2544 9998
rect 2700 9518 2728 10474
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2412 8968 2464 8974
rect 2412 8910 2464 8916
rect 2424 7002 2452 8910
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 2412 6996 2464 7002
rect 2412 6938 2464 6944
rect 2516 6934 2544 8774
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2700 7954 2728 8434
rect 2792 8430 2820 11630
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 2884 10062 2912 11154
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 2884 9586 2912 9998
rect 2976 9722 3004 17326
rect 3804 17202 3832 18566
rect 3884 18080 3936 18086
rect 3884 18022 3936 18028
rect 3896 17882 3924 18022
rect 3884 17876 3936 17882
rect 3884 17818 3936 17824
rect 3884 17536 3936 17542
rect 3884 17478 3936 17484
rect 3792 17196 3844 17202
rect 3792 17138 3844 17144
rect 3424 17128 3476 17134
rect 3424 17070 3476 17076
rect 3240 17060 3292 17066
rect 3240 17002 3292 17008
rect 3252 16454 3280 17002
rect 3240 16448 3292 16454
rect 3240 16390 3292 16396
rect 3332 16448 3384 16454
rect 3332 16390 3384 16396
rect 3056 16244 3108 16250
rect 3056 16186 3108 16192
rect 3068 15978 3096 16186
rect 3252 16114 3280 16390
rect 3240 16108 3292 16114
rect 3240 16050 3292 16056
rect 3344 16046 3372 16390
rect 3332 16040 3384 16046
rect 3332 15982 3384 15988
rect 3056 15972 3108 15978
rect 3056 15914 3108 15920
rect 3240 15904 3292 15910
rect 3436 15858 3464 17070
rect 3516 17060 3568 17066
rect 3516 17002 3568 17008
rect 3240 15846 3292 15852
rect 3252 15162 3280 15846
rect 3344 15830 3464 15858
rect 3240 15156 3292 15162
rect 3240 15098 3292 15104
rect 3056 14816 3108 14822
rect 3056 14758 3108 14764
rect 3068 14618 3096 14758
rect 3056 14612 3108 14618
rect 3056 14554 3108 14560
rect 3068 14278 3096 14554
rect 3056 14272 3108 14278
rect 3056 14214 3108 14220
rect 3240 13796 3292 13802
rect 3240 13738 3292 13744
rect 3054 13288 3110 13297
rect 3054 13223 3056 13232
rect 3108 13223 3110 13232
rect 3056 13194 3108 13200
rect 3252 12986 3280 13738
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 3146 12472 3202 12481
rect 3146 12407 3202 12416
rect 3160 11898 3188 12407
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3252 11898 3280 12174
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 3344 11529 3372 15830
rect 3528 15638 3556 17002
rect 3700 16788 3752 16794
rect 3700 16730 3752 16736
rect 3516 15632 3568 15638
rect 3712 15609 3740 16730
rect 3792 16516 3844 16522
rect 3792 16458 3844 16464
rect 3804 16153 3832 16458
rect 3790 16144 3846 16153
rect 3790 16079 3846 16088
rect 3516 15574 3568 15580
rect 3698 15600 3754 15609
rect 3424 14816 3476 14822
rect 3424 14758 3476 14764
rect 3330 11520 3386 11529
rect 3330 11455 3386 11464
rect 3436 11370 3464 14758
rect 3528 12850 3556 15574
rect 3698 15535 3754 15544
rect 3790 15464 3846 15473
rect 3790 15399 3846 15408
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 3620 14618 3648 14758
rect 3804 14618 3832 15399
rect 3608 14612 3660 14618
rect 3608 14554 3660 14560
rect 3792 14612 3844 14618
rect 3792 14554 3844 14560
rect 3792 14476 3844 14482
rect 3792 14418 3844 14424
rect 3608 14272 3660 14278
rect 3608 14214 3660 14220
rect 3516 12844 3568 12850
rect 3516 12786 3568 12792
rect 3516 12708 3568 12714
rect 3516 12650 3568 12656
rect 3344 11342 3464 11370
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 3148 11076 3200 11082
rect 3148 11018 3200 11024
rect 3160 10266 3188 11018
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2884 8974 2912 9114
rect 3068 8974 3096 9522
rect 3160 9518 3188 10202
rect 3148 9512 3200 9518
rect 3148 9454 3200 9460
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 3160 8838 3188 9454
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 2872 8560 2924 8566
rect 2872 8502 2924 8508
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2884 8090 2912 8502
rect 3056 8356 3108 8362
rect 3056 8298 3108 8304
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 2596 7268 2648 7274
rect 2596 7210 2648 7216
rect 2504 6928 2556 6934
rect 2504 6870 2556 6876
rect 2608 6798 2636 7210
rect 2700 7206 2728 7890
rect 3068 7818 3096 8298
rect 3056 7812 3108 7818
rect 3056 7754 3108 7760
rect 3160 7750 3188 8570
rect 3148 7744 3200 7750
rect 2870 7712 2926 7721
rect 3148 7686 3200 7692
rect 2870 7647 2926 7656
rect 2688 7200 2740 7206
rect 2688 7142 2740 7148
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2608 6390 2636 6734
rect 2596 6384 2648 6390
rect 2596 6326 2648 6332
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2700 5760 2728 6054
rect 2700 5732 2820 5760
rect 2792 5556 2820 5732
rect 2884 5681 2912 7647
rect 3056 6996 3108 7002
rect 3056 6938 3108 6944
rect 3068 6798 3096 6938
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 3068 6186 3096 6734
rect 3056 6180 3108 6186
rect 3056 6122 3108 6128
rect 3068 5794 3096 6122
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 3160 5914 3188 6054
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 3068 5766 3188 5794
rect 2964 5704 3016 5710
rect 2870 5672 2926 5681
rect 2964 5646 3016 5652
rect 2870 5607 2926 5616
rect 2976 5556 3004 5646
rect 3056 5636 3108 5642
rect 3056 5578 3108 5584
rect 2792 5528 3004 5556
rect 2780 5092 2832 5098
rect 2780 5034 2832 5040
rect 2872 5092 2924 5098
rect 2872 5034 2924 5040
rect 2792 4826 2820 5034
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2688 4752 2740 4758
rect 2688 4694 2740 4700
rect 2412 4548 2464 4554
rect 2412 4490 2464 4496
rect 2424 4146 2452 4490
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 2332 3738 2360 3878
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 2504 3596 2556 3602
rect 2504 3538 2556 3544
rect 2516 3194 2544 3538
rect 2700 3466 2728 4694
rect 2792 4214 2820 4762
rect 2780 4208 2832 4214
rect 2780 4150 2832 4156
rect 2884 4078 2912 5034
rect 2976 4486 3004 5528
rect 3068 5370 3096 5578
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 2964 4480 3016 4486
rect 2964 4422 3016 4428
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 2688 3460 2740 3466
rect 2688 3402 2740 3408
rect 2884 3194 2912 4014
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 2976 3097 3004 4422
rect 3056 3596 3108 3602
rect 3056 3538 3108 3544
rect 3068 3194 3096 3538
rect 3056 3188 3108 3194
rect 3056 3130 3108 3136
rect 2962 3088 3018 3097
rect 2962 3023 3018 3032
rect 2780 2984 2832 2990
rect 3160 2938 3188 5766
rect 2780 2926 2832 2932
rect 2226 2816 2282 2825
rect 2226 2751 2282 2760
rect 1860 1838 1912 1844
rect 2134 1864 2190 1873
rect 1400 1488 1452 1494
rect 1306 1456 1362 1465
rect 1400 1430 1452 1436
rect 1306 1391 1362 1400
rect 1412 800 1440 1430
rect 1872 800 1900 1838
rect 2134 1799 2190 1808
rect 2240 800 2268 2751
rect 2792 2689 2820 2926
rect 2976 2910 3188 2938
rect 2872 2848 2924 2854
rect 2872 2790 2924 2796
rect 2778 2680 2834 2689
rect 2884 2650 2912 2790
rect 2778 2615 2834 2624
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 2688 1964 2740 1970
rect 2688 1906 2740 1912
rect 2700 800 2728 1906
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1398 0 1454 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2686 0 2742 800
rect 2976 649 3004 2910
rect 3252 2446 3280 11086
rect 3344 10130 3372 11342
rect 3424 11280 3476 11286
rect 3424 11222 3476 11228
rect 3332 10124 3384 10130
rect 3332 10066 3384 10072
rect 3332 9988 3384 9994
rect 3332 9930 3384 9936
rect 3344 9382 3372 9930
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 3436 9178 3464 11222
rect 3528 9994 3556 12650
rect 3516 9988 3568 9994
rect 3516 9930 3568 9936
rect 3516 9716 3568 9722
rect 3516 9658 3568 9664
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3422 8936 3478 8945
rect 3422 8871 3478 8880
rect 3436 6934 3464 8871
rect 3424 6928 3476 6934
rect 3424 6870 3476 6876
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 3436 5030 3464 6734
rect 3528 6254 3556 9658
rect 3620 9489 3648 14214
rect 3804 13530 3832 14418
rect 3792 13524 3844 13530
rect 3792 13466 3844 13472
rect 3792 13388 3844 13394
rect 3792 13330 3844 13336
rect 3804 12986 3832 13330
rect 3792 12980 3844 12986
rect 3792 12922 3844 12928
rect 3896 11937 3924 17478
rect 3988 17134 4016 22200
rect 4066 21040 4122 21049
rect 4066 20975 4122 20984
rect 4080 19990 4108 20975
rect 4356 20534 4384 22200
rect 4421 20700 4717 20720
rect 4477 20698 4501 20700
rect 4557 20698 4581 20700
rect 4637 20698 4661 20700
rect 4499 20646 4501 20698
rect 4563 20646 4575 20698
rect 4637 20646 4639 20698
rect 4477 20644 4501 20646
rect 4557 20644 4581 20646
rect 4637 20644 4661 20646
rect 4421 20624 4717 20644
rect 4344 20528 4396 20534
rect 4344 20470 4396 20476
rect 4344 20392 4396 20398
rect 4344 20334 4396 20340
rect 4068 19984 4120 19990
rect 4068 19926 4120 19932
rect 4068 19848 4120 19854
rect 4120 19796 4200 19802
rect 4068 19790 4200 19796
rect 4080 19774 4200 19790
rect 4172 19514 4200 19774
rect 4160 19508 4212 19514
rect 4160 19450 4212 19456
rect 4172 19394 4200 19450
rect 4172 19366 4292 19394
rect 4158 19000 4214 19009
rect 4158 18935 4214 18944
rect 4172 18766 4200 18935
rect 4160 18760 4212 18766
rect 4160 18702 4212 18708
rect 4068 18692 4120 18698
rect 4068 18634 4120 18640
rect 4080 17864 4108 18634
rect 4158 18456 4214 18465
rect 4158 18391 4160 18400
rect 4212 18391 4214 18400
rect 4160 18362 4212 18368
rect 4160 17876 4212 17882
rect 4080 17836 4160 17864
rect 4160 17818 4212 17824
rect 4160 17740 4212 17746
rect 4160 17682 4212 17688
rect 4068 17604 4120 17610
rect 4068 17546 4120 17552
rect 4080 17270 4108 17546
rect 4172 17270 4200 17682
rect 4068 17264 4120 17270
rect 4068 17206 4120 17212
rect 4160 17264 4212 17270
rect 4160 17206 4212 17212
rect 3976 17128 4028 17134
rect 3976 17070 4028 17076
rect 4080 16726 4108 17206
rect 4068 16720 4120 16726
rect 4068 16662 4120 16668
rect 4068 16584 4120 16590
rect 4264 16572 4292 19366
rect 4356 19310 4384 20334
rect 4421 19612 4717 19632
rect 4477 19610 4501 19612
rect 4557 19610 4581 19612
rect 4637 19610 4661 19612
rect 4499 19558 4501 19610
rect 4563 19558 4575 19610
rect 4637 19558 4639 19610
rect 4477 19556 4501 19558
rect 4557 19556 4581 19558
rect 4637 19556 4661 19558
rect 4421 19536 4717 19556
rect 4344 19304 4396 19310
rect 4344 19246 4396 19252
rect 4344 18624 4396 18630
rect 4344 18566 4396 18572
rect 4356 18222 4384 18566
rect 4421 18524 4717 18544
rect 4477 18522 4501 18524
rect 4557 18522 4581 18524
rect 4637 18522 4661 18524
rect 4499 18470 4501 18522
rect 4563 18470 4575 18522
rect 4637 18470 4639 18522
rect 4477 18468 4501 18470
rect 4557 18468 4581 18470
rect 4637 18468 4661 18470
rect 4421 18448 4717 18468
rect 4620 18284 4672 18290
rect 4620 18226 4672 18232
rect 4344 18216 4396 18222
rect 4344 18158 4396 18164
rect 4436 18148 4488 18154
rect 4436 18090 4488 18096
rect 4448 17882 4476 18090
rect 4436 17876 4488 17882
rect 4436 17818 4488 17824
rect 4632 17678 4660 18226
rect 4620 17672 4672 17678
rect 4620 17614 4672 17620
rect 4421 17436 4717 17456
rect 4477 17434 4501 17436
rect 4557 17434 4581 17436
rect 4637 17434 4661 17436
rect 4499 17382 4501 17434
rect 4563 17382 4575 17434
rect 4637 17382 4639 17434
rect 4477 17380 4501 17382
rect 4557 17380 4581 17382
rect 4637 17380 4661 17382
rect 4421 17360 4717 17380
rect 4816 17354 4844 22200
rect 4988 19712 5040 19718
rect 4988 19654 5040 19660
rect 5000 19242 5028 19654
rect 4988 19236 5040 19242
rect 4988 19178 5040 19184
rect 4896 19168 4948 19174
rect 4896 19110 4948 19116
rect 4908 17882 4936 19110
rect 5000 18766 5028 19178
rect 5080 19168 5132 19174
rect 5080 19110 5132 19116
rect 4988 18760 5040 18766
rect 4988 18702 5040 18708
rect 4988 18624 5040 18630
rect 4988 18566 5040 18572
rect 5000 18426 5028 18566
rect 4988 18420 5040 18426
rect 4988 18362 5040 18368
rect 4896 17876 4948 17882
rect 4896 17818 4948 17824
rect 5000 17762 5028 18362
rect 5092 18290 5120 19110
rect 5080 18284 5132 18290
rect 5080 18226 5132 18232
rect 4908 17746 5028 17762
rect 4896 17740 5028 17746
rect 4948 17734 5028 17740
rect 4896 17682 4948 17688
rect 4988 17672 5040 17678
rect 4988 17614 5040 17620
rect 4816 17326 4936 17354
rect 4712 17196 4764 17202
rect 4764 17156 4844 17184
rect 4712 17138 4764 17144
rect 4344 16992 4396 16998
rect 4344 16934 4396 16940
rect 4120 16544 4292 16572
rect 4068 16526 4120 16532
rect 4080 16182 4108 16526
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 4068 16176 4120 16182
rect 4068 16118 4120 16124
rect 3976 15972 4028 15978
rect 3976 15914 4028 15920
rect 3988 15162 4016 15914
rect 3976 15156 4028 15162
rect 3976 15098 4028 15104
rect 3974 14648 4030 14657
rect 3974 14583 3976 14592
rect 4028 14583 4030 14592
rect 3976 14554 4028 14560
rect 3976 13864 4028 13870
rect 4080 13852 4108 16118
rect 4264 15978 4292 16186
rect 4252 15972 4304 15978
rect 4252 15914 4304 15920
rect 4160 15564 4212 15570
rect 4160 15506 4212 15512
rect 4172 15026 4200 15506
rect 4160 15020 4212 15026
rect 4160 14962 4212 14968
rect 4172 14414 4200 14962
rect 4356 14958 4384 16934
rect 4421 16348 4717 16368
rect 4477 16346 4501 16348
rect 4557 16346 4581 16348
rect 4637 16346 4661 16348
rect 4499 16294 4501 16346
rect 4563 16294 4575 16346
rect 4637 16294 4639 16346
rect 4477 16292 4501 16294
rect 4557 16292 4581 16294
rect 4637 16292 4661 16294
rect 4421 16272 4717 16292
rect 4816 16250 4844 17156
rect 4804 16244 4856 16250
rect 4804 16186 4856 16192
rect 4804 16040 4856 16046
rect 4804 15982 4856 15988
rect 4436 15904 4488 15910
rect 4436 15846 4488 15852
rect 4448 15706 4476 15846
rect 4436 15700 4488 15706
rect 4436 15642 4488 15648
rect 4421 15260 4717 15280
rect 4477 15258 4501 15260
rect 4557 15258 4581 15260
rect 4637 15258 4661 15260
rect 4499 15206 4501 15258
rect 4563 15206 4575 15258
rect 4637 15206 4639 15258
rect 4477 15204 4501 15206
rect 4557 15204 4581 15206
rect 4637 15204 4661 15206
rect 4421 15184 4717 15204
rect 4816 15026 4844 15982
rect 4804 15020 4856 15026
rect 4804 14962 4856 14968
rect 4344 14952 4396 14958
rect 4344 14894 4396 14900
rect 4356 14618 4384 14894
rect 4344 14612 4396 14618
rect 4344 14554 4396 14560
rect 4804 14476 4856 14482
rect 4804 14418 4856 14424
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 4421 14172 4717 14192
rect 4477 14170 4501 14172
rect 4557 14170 4581 14172
rect 4637 14170 4661 14172
rect 4499 14118 4501 14170
rect 4563 14118 4575 14170
rect 4637 14118 4639 14170
rect 4477 14116 4501 14118
rect 4557 14116 4581 14118
rect 4637 14116 4661 14118
rect 4421 14096 4717 14116
rect 4028 13824 4108 13852
rect 4528 13864 4580 13870
rect 3976 13806 4028 13812
rect 4528 13806 4580 13812
rect 3988 13326 4016 13806
rect 4160 13796 4212 13802
rect 4160 13738 4212 13744
rect 4172 13530 4200 13738
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 4172 13394 4200 13466
rect 4540 13462 4568 13806
rect 4528 13456 4580 13462
rect 4528 13398 4580 13404
rect 4160 13388 4212 13394
rect 4344 13388 4396 13394
rect 4160 13330 4212 13336
rect 4264 13348 4344 13376
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 3988 12374 4016 13262
rect 4264 12850 4292 13348
rect 4344 13330 4396 13336
rect 4344 13184 4396 13190
rect 4344 13126 4396 13132
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4172 12442 4200 12582
rect 4356 12442 4384 13126
rect 4421 13084 4717 13104
rect 4477 13082 4501 13084
rect 4557 13082 4581 13084
rect 4637 13082 4661 13084
rect 4499 13030 4501 13082
rect 4563 13030 4575 13082
rect 4637 13030 4639 13082
rect 4477 13028 4501 13030
rect 4557 13028 4581 13030
rect 4637 13028 4661 13030
rect 4421 13008 4717 13028
rect 4816 12986 4844 14418
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4620 12912 4672 12918
rect 4620 12854 4672 12860
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 3976 12368 4028 12374
rect 3976 12310 4028 12316
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 3882 11928 3938 11937
rect 3882 11863 3938 11872
rect 3884 11824 3936 11830
rect 3884 11766 3936 11772
rect 3700 11756 3752 11762
rect 3700 11698 3752 11704
rect 3712 11218 3740 11698
rect 3896 11665 3924 11766
rect 3882 11656 3938 11665
rect 3882 11591 3938 11600
rect 3792 11552 3844 11558
rect 3792 11494 3844 11500
rect 3700 11212 3752 11218
rect 3700 11154 3752 11160
rect 3712 10810 3740 11154
rect 3804 10810 3832 11494
rect 3988 11150 4016 12038
rect 4264 11898 4292 12242
rect 4632 12152 4660 12854
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4356 12124 4660 12152
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4356 11778 4384 12124
rect 4421 11996 4717 12016
rect 4477 11994 4501 11996
rect 4557 11994 4581 11996
rect 4637 11994 4661 11996
rect 4499 11942 4501 11994
rect 4563 11942 4575 11994
rect 4637 11942 4639 11994
rect 4477 11940 4501 11942
rect 4557 11940 4581 11942
rect 4637 11940 4661 11942
rect 4421 11920 4717 11940
rect 4264 11750 4384 11778
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 3700 10804 3752 10810
rect 3700 10746 3752 10752
rect 3792 10804 3844 10810
rect 3792 10746 3844 10752
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3792 10124 3844 10130
rect 3792 10066 3844 10072
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 3606 9480 3662 9489
rect 3606 9415 3662 9424
rect 3620 8022 3648 9415
rect 3712 9382 3740 9862
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 3608 8016 3660 8022
rect 3608 7958 3660 7964
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 3620 7546 3648 7822
rect 3712 7750 3740 9318
rect 3700 7744 3752 7750
rect 3804 7721 3832 10066
rect 3896 9042 3924 10542
rect 4172 10266 4200 11494
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 4158 10024 4214 10033
rect 4158 9959 4214 9968
rect 3884 9036 3936 9042
rect 3884 8978 3936 8984
rect 3884 8424 3936 8430
rect 3884 8366 3936 8372
rect 3700 7686 3752 7692
rect 3790 7712 3846 7721
rect 3608 7540 3660 7546
rect 3608 7482 3660 7488
rect 3712 7426 3740 7686
rect 3790 7647 3846 7656
rect 3620 7398 3740 7426
rect 3896 7410 3924 8366
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3988 7449 4016 8230
rect 4066 7848 4122 7857
rect 4066 7783 4122 7792
rect 3974 7440 4030 7449
rect 3884 7404 3936 7410
rect 3516 6248 3568 6254
rect 3516 6190 3568 6196
rect 3516 6112 3568 6118
rect 3516 6054 3568 6060
rect 3528 5642 3556 6054
rect 3516 5636 3568 5642
rect 3516 5578 3568 5584
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 3516 4684 3568 4690
rect 3516 4626 3568 4632
rect 3528 3738 3556 4626
rect 3516 3732 3568 3738
rect 3516 3674 3568 3680
rect 3620 3618 3648 7398
rect 3974 7375 4030 7384
rect 3884 7346 3936 7352
rect 3700 6928 3752 6934
rect 3700 6870 3752 6876
rect 3712 6186 3740 6870
rect 3896 6798 3924 7346
rect 4080 6934 4108 7783
rect 4068 6928 4120 6934
rect 4068 6870 4120 6876
rect 3884 6792 3936 6798
rect 4172 6780 4200 9959
rect 4264 9586 4292 11750
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 4816 11642 4844 12718
rect 4908 12102 4936 17326
rect 5000 17202 5028 17614
rect 4988 17196 5040 17202
rect 4988 17138 5040 17144
rect 5000 15502 5028 17138
rect 4988 15496 5040 15502
rect 5040 15456 5120 15484
rect 4988 15438 5040 15444
rect 4988 15360 5040 15366
rect 4988 15302 5040 15308
rect 5000 12782 5028 15302
rect 5092 15162 5120 15456
rect 5080 15156 5132 15162
rect 5080 15098 5132 15104
rect 5184 14906 5212 22200
rect 5356 20528 5408 20534
rect 5356 20470 5408 20476
rect 5264 19848 5316 19854
rect 5264 19790 5316 19796
rect 5276 19514 5304 19790
rect 5264 19508 5316 19514
rect 5264 19450 5316 19456
rect 5264 19168 5316 19174
rect 5264 19110 5316 19116
rect 5276 18970 5304 19110
rect 5264 18964 5316 18970
rect 5264 18906 5316 18912
rect 5264 18080 5316 18086
rect 5264 18022 5316 18028
rect 5276 16658 5304 18022
rect 5368 17762 5396 20470
rect 5448 20324 5500 20330
rect 5448 20266 5500 20272
rect 5460 18970 5488 20266
rect 5552 20074 5580 22200
rect 5552 20046 5764 20074
rect 5540 19916 5592 19922
rect 5540 19858 5592 19864
rect 5552 19514 5580 19858
rect 5540 19508 5592 19514
rect 5540 19450 5592 19456
rect 5448 18964 5500 18970
rect 5448 18906 5500 18912
rect 5632 18148 5684 18154
rect 5632 18090 5684 18096
rect 5368 17734 5488 17762
rect 5356 17672 5408 17678
rect 5356 17614 5408 17620
rect 5368 17338 5396 17614
rect 5356 17332 5408 17338
rect 5356 17274 5408 17280
rect 5264 16652 5316 16658
rect 5264 16594 5316 16600
rect 5276 16250 5304 16594
rect 5264 16244 5316 16250
rect 5264 16186 5316 16192
rect 5356 15972 5408 15978
rect 5356 15914 5408 15920
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 5276 15570 5304 15846
rect 5264 15564 5316 15570
rect 5264 15506 5316 15512
rect 5092 14878 5212 14906
rect 5092 12918 5120 14878
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5184 14278 5212 14758
rect 5172 14272 5224 14278
rect 5172 14214 5224 14220
rect 5080 12912 5132 12918
rect 5080 12854 5132 12860
rect 4988 12776 5040 12782
rect 4988 12718 5040 12724
rect 5080 12776 5132 12782
rect 5080 12718 5132 12724
rect 4988 12640 5040 12646
rect 4988 12582 5040 12588
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 5000 11694 5028 12582
rect 5092 12238 5120 12718
rect 5080 12232 5132 12238
rect 5080 12174 5132 12180
rect 5078 12064 5134 12073
rect 5078 11999 5134 12008
rect 4988 11688 5040 11694
rect 4356 10674 4384 11630
rect 4816 11614 4936 11642
rect 4988 11630 5040 11636
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 4632 11354 4660 11494
rect 4710 11384 4766 11393
rect 4620 11348 4672 11354
rect 4710 11319 4766 11328
rect 4620 11290 4672 11296
rect 4724 11218 4752 11319
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4421 10908 4717 10928
rect 4477 10906 4501 10908
rect 4557 10906 4581 10908
rect 4637 10906 4661 10908
rect 4499 10854 4501 10906
rect 4563 10854 4575 10906
rect 4637 10854 4639 10906
rect 4477 10852 4501 10854
rect 4557 10852 4581 10854
rect 4637 10852 4661 10854
rect 4421 10832 4717 10852
rect 4816 10810 4844 11494
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 4252 9580 4304 9586
rect 4252 9522 4304 9528
rect 4356 7392 4384 10610
rect 4908 10266 4936 11614
rect 5000 11354 5028 11630
rect 5092 11558 5120 11999
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 5092 11393 5120 11494
rect 5078 11384 5134 11393
rect 4988 11348 5040 11354
rect 5078 11319 5134 11328
rect 4988 11290 5040 11296
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 5000 10674 5028 11086
rect 5080 10804 5132 10810
rect 5080 10746 5132 10752
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 4988 10532 5040 10538
rect 4988 10474 5040 10480
rect 4896 10260 4948 10266
rect 4896 10202 4948 10208
rect 5000 10146 5028 10474
rect 5092 10470 5120 10746
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 4908 10118 5028 10146
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 4421 9820 4717 9840
rect 4477 9818 4501 9820
rect 4557 9818 4581 9820
rect 4637 9818 4661 9820
rect 4499 9766 4501 9818
rect 4563 9766 4575 9818
rect 4637 9766 4639 9818
rect 4477 9764 4501 9766
rect 4557 9764 4581 9766
rect 4637 9764 4661 9766
rect 4421 9744 4717 9764
rect 4816 9722 4844 9998
rect 4804 9716 4856 9722
rect 4804 9658 4856 9664
rect 4712 9648 4764 9654
rect 4712 9590 4764 9596
rect 4724 9382 4752 9590
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4632 9178 4660 9318
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4816 9110 4844 9522
rect 4804 9104 4856 9110
rect 4804 9046 4856 9052
rect 4421 8732 4717 8752
rect 4477 8730 4501 8732
rect 4557 8730 4581 8732
rect 4637 8730 4661 8732
rect 4499 8678 4501 8730
rect 4563 8678 4575 8730
rect 4637 8678 4639 8730
rect 4477 8676 4501 8678
rect 4557 8676 4581 8678
rect 4637 8676 4661 8678
rect 4421 8656 4717 8676
rect 4816 8634 4844 9046
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 4421 7644 4717 7664
rect 4477 7642 4501 7644
rect 4557 7642 4581 7644
rect 4637 7642 4661 7644
rect 4499 7590 4501 7642
rect 4563 7590 4575 7642
rect 4637 7590 4639 7642
rect 4477 7588 4501 7590
rect 4557 7588 4581 7590
rect 4637 7588 4661 7590
rect 4421 7568 4717 7588
rect 4080 6752 4200 6780
rect 4264 7364 4384 7392
rect 4080 6746 4108 6752
rect 3884 6734 3936 6740
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 3700 6180 3752 6186
rect 3700 6122 3752 6128
rect 3700 5636 3752 5642
rect 3700 5578 3752 5584
rect 3712 5098 3740 5578
rect 3804 5166 3832 6258
rect 3896 5642 3924 6734
rect 3988 6718 4108 6746
rect 3988 6089 4016 6718
rect 4066 6488 4122 6497
rect 4066 6423 4122 6432
rect 3974 6080 4030 6089
rect 3974 6015 4030 6024
rect 4080 5914 4108 6423
rect 4160 6180 4212 6186
rect 4160 6122 4212 6128
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 3976 5772 4028 5778
rect 4028 5732 4108 5760
rect 3976 5714 4028 5720
rect 3884 5636 3936 5642
rect 3884 5578 3936 5584
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3700 5092 3752 5098
rect 3700 5034 3752 5040
rect 3712 4758 3740 5034
rect 3700 4752 3752 4758
rect 3700 4694 3752 4700
rect 3700 4616 3752 4622
rect 3700 4558 3752 4564
rect 3712 4282 3740 4558
rect 3700 4276 3752 4282
rect 3700 4218 3752 4224
rect 3436 3590 3648 3618
rect 3792 3664 3844 3670
rect 3792 3606 3844 3612
rect 3700 3596 3752 3602
rect 3436 2990 3464 3590
rect 3700 3538 3752 3544
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3528 3058 3556 3334
rect 3712 3194 3740 3538
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 3804 3126 3832 3606
rect 3792 3120 3844 3126
rect 3792 3062 3844 3068
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 3700 2984 3752 2990
rect 3700 2926 3752 2932
rect 3516 2916 3568 2922
rect 3516 2858 3568 2864
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3148 2304 3200 2310
rect 3148 2246 3200 2252
rect 3160 1873 3188 2246
rect 3146 1864 3202 1873
rect 3146 1799 3202 1808
rect 3056 1624 3108 1630
rect 3056 1566 3108 1572
rect 3068 800 3096 1566
rect 3528 800 3556 2858
rect 3608 2508 3660 2514
rect 3608 2450 3660 2456
rect 3620 2310 3648 2450
rect 3712 2378 3740 2926
rect 3700 2372 3752 2378
rect 3700 2314 3752 2320
rect 3608 2304 3660 2310
rect 3608 2246 3660 2252
rect 3792 2304 3844 2310
rect 3792 2246 3844 2252
rect 3620 1057 3648 2246
rect 3606 1048 3662 1057
rect 3606 983 3662 992
rect 2962 640 3018 649
rect 2962 575 3018 584
rect 3054 0 3110 800
rect 3514 0 3570 800
rect 3804 241 3832 2246
rect 3896 800 3924 5306
rect 4080 4826 4108 5732
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4172 4146 4200 6122
rect 4264 5817 4292 7364
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4344 7268 4396 7274
rect 4344 7210 4396 7216
rect 4356 6458 4384 7210
rect 4421 6556 4717 6576
rect 4477 6554 4501 6556
rect 4557 6554 4581 6556
rect 4637 6554 4661 6556
rect 4499 6502 4501 6554
rect 4563 6502 4575 6554
rect 4637 6502 4639 6554
rect 4477 6500 4501 6502
rect 4557 6500 4581 6502
rect 4637 6500 4661 6502
rect 4421 6480 4717 6500
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4250 5808 4306 5817
rect 4250 5743 4306 5752
rect 4356 5370 4384 6054
rect 4421 5468 4717 5488
rect 4477 5466 4501 5468
rect 4557 5466 4581 5468
rect 4637 5466 4661 5468
rect 4499 5414 4501 5466
rect 4563 5414 4575 5466
rect 4637 5414 4639 5466
rect 4477 5412 4501 5414
rect 4557 5412 4581 5414
rect 4637 5412 4661 5414
rect 4421 5392 4717 5412
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4816 5250 4844 7278
rect 4356 5222 4844 5250
rect 4252 5092 4304 5098
rect 4252 5034 4304 5040
rect 4264 4486 4292 5034
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4250 4312 4306 4321
rect 4250 4247 4252 4256
rect 4304 4247 4306 4256
rect 4252 4218 4304 4224
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4252 4004 4304 4010
rect 4252 3946 4304 3952
rect 4160 3664 4212 3670
rect 4080 3624 4160 3652
rect 4080 2922 4108 3624
rect 4160 3606 4212 3612
rect 4264 3398 4292 3946
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 4068 2916 4120 2922
rect 4068 2858 4120 2864
rect 4172 2650 4200 2926
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 4264 2378 4292 3334
rect 4252 2372 4304 2378
rect 4252 2314 4304 2320
rect 4356 800 4384 5222
rect 4908 4842 4936 10118
rect 5184 9874 5212 14214
rect 5276 12345 5304 15506
rect 5368 15366 5396 15914
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 5356 14952 5408 14958
rect 5354 14920 5356 14929
rect 5408 14920 5410 14929
rect 5354 14855 5410 14864
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 5368 12850 5396 13466
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 5262 12336 5318 12345
rect 5262 12271 5318 12280
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 5092 9846 5212 9874
rect 5092 9602 5120 9846
rect 5092 9574 5304 9602
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 5092 8974 5120 9318
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 5092 7954 5120 8774
rect 5184 8090 5212 9318
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 5080 7948 5132 7954
rect 5080 7890 5132 7896
rect 5092 7750 5120 7890
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 5000 6322 5028 7142
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 4908 4814 5028 4842
rect 4896 4548 4948 4554
rect 4896 4490 4948 4496
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4421 4380 4717 4400
rect 4477 4378 4501 4380
rect 4557 4378 4581 4380
rect 4637 4378 4661 4380
rect 4499 4326 4501 4378
rect 4563 4326 4575 4378
rect 4637 4326 4639 4378
rect 4477 4324 4501 4326
rect 4557 4324 4581 4326
rect 4637 4324 4661 4326
rect 4421 4304 4717 4324
rect 4712 4208 4764 4214
rect 4712 4150 4764 4156
rect 4724 3618 4752 4150
rect 4816 3738 4844 4422
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4724 3590 4844 3618
rect 4421 3292 4717 3312
rect 4477 3290 4501 3292
rect 4557 3290 4581 3292
rect 4637 3290 4661 3292
rect 4499 3238 4501 3290
rect 4563 3238 4575 3290
rect 4637 3238 4639 3290
rect 4477 3236 4501 3238
rect 4557 3236 4581 3238
rect 4637 3236 4661 3238
rect 4421 3216 4717 3236
rect 4712 2916 4764 2922
rect 4712 2858 4764 2864
rect 4724 2446 4752 2858
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 4421 2204 4717 2224
rect 4477 2202 4501 2204
rect 4557 2202 4581 2204
rect 4637 2202 4661 2204
rect 4499 2150 4501 2202
rect 4563 2150 4575 2202
rect 4637 2150 4639 2202
rect 4477 2148 4501 2150
rect 4557 2148 4581 2150
rect 4637 2148 4661 2150
rect 4421 2128 4717 2148
rect 4816 800 4844 3590
rect 4908 2650 4936 4490
rect 5000 4214 5028 4814
rect 4988 4208 5040 4214
rect 4988 4150 5040 4156
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 4896 2644 4948 2650
rect 4896 2586 4948 2592
rect 5000 2514 5028 3878
rect 5092 2582 5120 7686
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5184 6866 5212 7346
rect 5172 6860 5224 6866
rect 5172 6802 5224 6808
rect 5184 6497 5212 6802
rect 5170 6488 5226 6497
rect 5276 6458 5304 9574
rect 5368 8072 5396 12038
rect 5460 11393 5488 17734
rect 5540 17264 5592 17270
rect 5540 17206 5592 17212
rect 5552 15570 5580 17206
rect 5644 17202 5672 18090
rect 5632 17196 5684 17202
rect 5632 17138 5684 17144
rect 5632 16448 5684 16454
rect 5632 16390 5684 16396
rect 5644 15706 5672 16390
rect 5632 15700 5684 15706
rect 5632 15642 5684 15648
rect 5540 15564 5592 15570
rect 5540 15506 5592 15512
rect 5736 14770 5764 20046
rect 5920 19310 5948 22200
rect 5908 19304 5960 19310
rect 5908 19246 5960 19252
rect 5906 19000 5962 19009
rect 5906 18935 5908 18944
rect 5960 18935 5962 18944
rect 5908 18906 5960 18912
rect 5816 18828 5868 18834
rect 5816 18770 5868 18776
rect 5828 18426 5856 18770
rect 6184 18760 6236 18766
rect 6184 18702 6236 18708
rect 5908 18692 5960 18698
rect 5908 18634 5960 18640
rect 5816 18420 5868 18426
rect 5816 18362 5868 18368
rect 5920 17338 5948 18634
rect 6092 18284 6144 18290
rect 6092 18226 6144 18232
rect 6104 17882 6132 18226
rect 6092 17876 6144 17882
rect 6092 17818 6144 17824
rect 5908 17332 5960 17338
rect 5908 17274 5960 17280
rect 6092 17332 6144 17338
rect 6092 17274 6144 17280
rect 5906 17232 5962 17241
rect 5906 17167 5962 17176
rect 5920 17134 5948 17167
rect 5908 17128 5960 17134
rect 6104 17105 6132 17274
rect 6196 17134 6224 18702
rect 6288 18465 6316 22200
rect 6656 20618 6684 22200
rect 6472 20590 6684 20618
rect 6368 18964 6420 18970
rect 6368 18906 6420 18912
rect 6274 18456 6330 18465
rect 6274 18391 6330 18400
rect 6276 18216 6328 18222
rect 6380 18204 6408 18906
rect 6328 18176 6408 18204
rect 6276 18158 6328 18164
rect 6368 17264 6420 17270
rect 6368 17206 6420 17212
rect 6276 17196 6328 17202
rect 6276 17138 6328 17144
rect 6184 17128 6236 17134
rect 5908 17070 5960 17076
rect 6090 17096 6146 17105
rect 6184 17070 6236 17076
rect 6090 17031 6146 17040
rect 6104 16726 6132 17031
rect 6092 16720 6144 16726
rect 6092 16662 6144 16668
rect 6288 16590 6316 17138
rect 6380 16794 6408 17206
rect 6368 16788 6420 16794
rect 6368 16730 6420 16736
rect 6368 16652 6420 16658
rect 6368 16594 6420 16600
rect 6276 16584 6328 16590
rect 6276 16526 6328 16532
rect 5908 15972 5960 15978
rect 5908 15914 5960 15920
rect 5920 15502 5948 15914
rect 5908 15496 5960 15502
rect 5908 15438 5960 15444
rect 5920 15094 5948 15438
rect 5908 15088 5960 15094
rect 5908 15030 5960 15036
rect 6288 14929 6316 16526
rect 6380 15706 6408 16594
rect 6368 15700 6420 15706
rect 6368 15642 6420 15648
rect 6368 15428 6420 15434
rect 6368 15370 6420 15376
rect 6380 15162 6408 15370
rect 6368 15156 6420 15162
rect 6368 15098 6420 15104
rect 6274 14920 6330 14929
rect 6092 14884 6144 14890
rect 6274 14855 6330 14864
rect 6092 14826 6144 14832
rect 5736 14742 5856 14770
rect 5828 14618 5856 14742
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5552 12646 5580 14214
rect 5632 14068 5684 14074
rect 5632 14010 5684 14016
rect 5644 12986 5672 14010
rect 5632 12980 5684 12986
rect 5736 12968 5764 14554
rect 5816 14408 5868 14414
rect 5816 14350 5868 14356
rect 6000 14408 6052 14414
rect 6000 14350 6052 14356
rect 5828 14074 5856 14350
rect 5908 14340 5960 14346
rect 5908 14282 5960 14288
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 5920 14006 5948 14282
rect 5908 14000 5960 14006
rect 5908 13942 5960 13948
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 5908 13728 5960 13734
rect 5908 13670 5960 13676
rect 5828 13462 5856 13670
rect 5816 13456 5868 13462
rect 5816 13398 5868 13404
rect 5736 12940 5856 12968
rect 5632 12922 5684 12928
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5446 11384 5502 11393
rect 5446 11319 5502 11328
rect 5552 11218 5580 12038
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5644 10810 5672 12786
rect 5724 12640 5776 12646
rect 5722 12608 5724 12617
rect 5776 12608 5778 12617
rect 5722 12543 5778 12552
rect 5828 12322 5856 12940
rect 5920 12782 5948 13670
rect 6012 12986 6040 14350
rect 6104 13818 6132 14826
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 6196 13938 6224 14350
rect 6184 13932 6236 13938
rect 6184 13874 6236 13880
rect 6104 13790 6224 13818
rect 6092 13728 6144 13734
rect 6092 13670 6144 13676
rect 6104 13530 6132 13670
rect 6196 13530 6224 13790
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6196 13394 6224 13466
rect 6184 13388 6236 13394
rect 6184 13330 6236 13336
rect 6184 13184 6236 13190
rect 6184 13126 6236 13132
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 5908 12776 5960 12782
rect 5908 12718 5960 12724
rect 6196 12374 6224 13126
rect 6380 12850 6408 15098
rect 6368 12844 6420 12850
rect 6368 12786 6420 12792
rect 6276 12640 6328 12646
rect 6276 12582 6328 12588
rect 5736 12294 5856 12322
rect 6184 12368 6236 12374
rect 6184 12310 6236 12316
rect 6092 12300 6144 12306
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5460 10062 5488 10610
rect 5644 10266 5672 10746
rect 5736 10674 5764 12294
rect 6092 12242 6144 12248
rect 5816 12232 5868 12238
rect 5816 12174 5868 12180
rect 5828 11626 5856 12174
rect 6104 11665 6132 12242
rect 6090 11656 6146 11665
rect 5816 11620 5868 11626
rect 6090 11591 6146 11600
rect 5816 11562 5868 11568
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 5632 10260 5684 10266
rect 5632 10202 5684 10208
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 5460 9518 5488 9998
rect 5552 9654 5580 10066
rect 5736 9897 5764 10610
rect 5828 10606 5856 11562
rect 6104 11150 6132 11591
rect 6184 11552 6236 11558
rect 6184 11494 6236 11500
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6000 11076 6052 11082
rect 6000 11018 6052 11024
rect 5906 10840 5962 10849
rect 5906 10775 5962 10784
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5920 10441 5948 10775
rect 6012 10538 6040 11018
rect 6092 11008 6144 11014
rect 6092 10950 6144 10956
rect 6104 10674 6132 10950
rect 6092 10668 6144 10674
rect 6092 10610 6144 10616
rect 6196 10538 6224 11494
rect 6288 10810 6316 12582
rect 6366 12336 6422 12345
rect 6366 12271 6422 12280
rect 6380 11898 6408 12271
rect 6368 11892 6420 11898
rect 6368 11834 6420 11840
rect 6472 11830 6500 20590
rect 6644 20460 6696 20466
rect 6644 20402 6696 20408
rect 6656 19514 6684 20402
rect 7116 20346 7144 22200
rect 7484 20482 7512 22200
rect 7484 20454 7604 20482
rect 7116 20318 7512 20346
rect 7288 20256 7340 20262
rect 7288 20198 7340 20204
rect 6828 19916 6880 19922
rect 6828 19858 6880 19864
rect 6644 19508 6696 19514
rect 6644 19450 6696 19456
rect 6840 19174 6868 19858
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 6920 19304 6972 19310
rect 7208 19258 7236 19654
rect 6920 19246 6972 19252
rect 6736 19168 6788 19174
rect 6736 19110 6788 19116
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6748 18902 6776 19110
rect 6736 18896 6788 18902
rect 6736 18838 6788 18844
rect 6644 18828 6696 18834
rect 6644 18770 6696 18776
rect 6656 18290 6684 18770
rect 6840 18714 6868 19110
rect 6932 18850 6960 19246
rect 7024 19242 7236 19258
rect 7012 19236 7236 19242
rect 7064 19230 7236 19236
rect 7012 19178 7064 19184
rect 7102 19000 7158 19009
rect 7102 18935 7104 18944
rect 7156 18935 7158 18944
rect 7104 18906 7156 18912
rect 6932 18822 7144 18850
rect 6920 18760 6972 18766
rect 6840 18708 6920 18714
rect 6840 18702 6972 18708
rect 6840 18686 6960 18702
rect 6840 18306 6868 18686
rect 7116 18465 7144 18822
rect 7208 18698 7236 19230
rect 7196 18692 7248 18698
rect 7196 18634 7248 18640
rect 7102 18456 7158 18465
rect 7102 18391 7158 18400
rect 6840 18290 6960 18306
rect 6644 18284 6696 18290
rect 6644 18226 6696 18232
rect 6840 18284 6972 18290
rect 6840 18278 6920 18284
rect 6840 17882 6868 18278
rect 6920 18226 6972 18232
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6552 17740 6604 17746
rect 6552 17682 6604 17688
rect 6564 17649 6592 17682
rect 6550 17640 6606 17649
rect 6550 17575 6606 17584
rect 6828 17604 6880 17610
rect 6828 17546 6880 17552
rect 6736 17536 6788 17542
rect 6736 17478 6788 17484
rect 6748 17338 6776 17478
rect 6736 17332 6788 17338
rect 6736 17274 6788 17280
rect 6550 17232 6606 17241
rect 6840 17218 6868 17546
rect 6932 17338 6960 17818
rect 7116 17626 7144 18391
rect 7208 18358 7236 18634
rect 7196 18352 7248 18358
rect 7196 18294 7248 18300
rect 7300 18086 7328 20198
rect 7380 20052 7432 20058
rect 7380 19994 7432 20000
rect 7392 19922 7420 19994
rect 7380 19916 7432 19922
rect 7380 19858 7432 19864
rect 7380 19236 7432 19242
rect 7380 19178 7432 19184
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7116 17598 7236 17626
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 6550 17167 6552 17176
rect 6604 17167 6606 17176
rect 6656 17190 6868 17218
rect 6552 17138 6604 17144
rect 6656 16726 6684 17190
rect 6736 17128 6788 17134
rect 6736 17070 6788 17076
rect 6644 16720 6696 16726
rect 6644 16662 6696 16668
rect 6748 16572 6776 17070
rect 7116 16998 7144 17478
rect 7104 16992 7156 16998
rect 6918 16960 6974 16969
rect 7104 16934 7156 16940
rect 6918 16895 6974 16904
rect 6656 16544 6776 16572
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 6564 13870 6592 14554
rect 6552 13864 6604 13870
rect 6552 13806 6604 13812
rect 6550 13696 6606 13705
rect 6550 13631 6606 13640
rect 6564 13530 6592 13631
rect 6552 13524 6604 13530
rect 6552 13466 6604 13472
rect 6552 13320 6604 13326
rect 6550 13288 6552 13297
rect 6604 13288 6606 13297
rect 6550 13223 6606 13232
rect 6656 12889 6684 16544
rect 6736 15972 6788 15978
rect 6736 15914 6788 15920
rect 6748 15502 6776 15914
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 6828 15496 6880 15502
rect 6828 15438 6880 15444
rect 6736 15360 6788 15366
rect 6736 15302 6788 15308
rect 6748 15162 6776 15302
rect 6736 15156 6788 15162
rect 6736 15098 6788 15104
rect 6736 14816 6788 14822
rect 6840 14804 6868 15438
rect 6788 14776 6868 14804
rect 6736 14758 6788 14764
rect 6642 12880 6698 12889
rect 6552 12844 6604 12850
rect 6642 12815 6698 12824
rect 6552 12786 6604 12792
rect 6564 12730 6592 12786
rect 6564 12702 6684 12730
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6460 11824 6512 11830
rect 6460 11766 6512 11772
rect 6368 11688 6420 11694
rect 6368 11630 6420 11636
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 6380 10674 6408 11630
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6472 11121 6500 11290
rect 6458 11112 6514 11121
rect 6458 11047 6514 11056
rect 6458 10976 6514 10985
rect 6458 10911 6514 10920
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 6000 10532 6052 10538
rect 6000 10474 6052 10480
rect 6184 10532 6236 10538
rect 6184 10474 6236 10480
rect 5906 10432 5962 10441
rect 5906 10367 5962 10376
rect 5998 10296 6054 10305
rect 5998 10231 6054 10240
rect 6092 10260 6144 10266
rect 5908 10056 5960 10062
rect 5908 9998 5960 10004
rect 5722 9888 5778 9897
rect 5722 9823 5778 9832
rect 5722 9752 5778 9761
rect 5722 9687 5778 9696
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 5460 9178 5488 9454
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5552 9058 5580 9454
rect 5460 9030 5580 9058
rect 5632 9104 5684 9110
rect 5632 9046 5684 9052
rect 5460 8362 5488 9030
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5368 8044 5488 8072
rect 5354 7984 5410 7993
rect 5354 7919 5410 7928
rect 5368 7342 5396 7919
rect 5460 7478 5488 8044
rect 5552 7732 5580 8910
rect 5644 8838 5672 9046
rect 5736 8838 5764 9687
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5632 8832 5684 8838
rect 5632 8774 5684 8780
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5644 7857 5672 8774
rect 5630 7848 5686 7857
rect 5630 7783 5686 7792
rect 5552 7704 5672 7732
rect 5448 7472 5500 7478
rect 5448 7414 5500 7420
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5460 6662 5488 7278
rect 5644 7274 5672 7704
rect 5632 7268 5684 7274
rect 5632 7210 5684 7216
rect 5736 6712 5764 8774
rect 5828 7818 5856 9318
rect 5920 8634 5948 9998
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 5816 7812 5868 7818
rect 5816 7754 5868 7760
rect 5816 6860 5868 6866
rect 5920 6848 5948 8570
rect 5868 6820 5948 6848
rect 5816 6802 5868 6808
rect 5644 6684 5764 6712
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5170 6423 5226 6432
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 5460 6390 5488 6598
rect 5448 6384 5500 6390
rect 5448 6326 5500 6332
rect 5540 5840 5592 5846
rect 5540 5782 5592 5788
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 5368 5234 5396 5646
rect 5552 5370 5580 5782
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5184 4282 5212 4626
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5368 4486 5396 4558
rect 5356 4480 5408 4486
rect 5356 4422 5408 4428
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 5080 2576 5132 2582
rect 5080 2518 5132 2524
rect 4988 2508 5040 2514
rect 4988 2450 5040 2456
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 4908 2310 4936 2382
rect 4896 2304 4948 2310
rect 4896 2246 4948 2252
rect 5184 800 5212 4218
rect 5262 4176 5318 4185
rect 5368 4146 5396 4422
rect 5446 4312 5502 4321
rect 5446 4247 5502 4256
rect 5460 4214 5488 4247
rect 5448 4208 5500 4214
rect 5448 4150 5500 4156
rect 5262 4111 5264 4120
rect 5316 4111 5318 4120
rect 5356 4140 5408 4146
rect 5264 4082 5316 4088
rect 5356 4082 5408 4088
rect 5276 3942 5304 4082
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 5368 2310 5396 4082
rect 5460 4010 5488 4150
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5448 2848 5500 2854
rect 5448 2790 5500 2796
rect 5460 2378 5488 2790
rect 5552 2582 5580 3130
rect 5540 2576 5592 2582
rect 5540 2518 5592 2524
rect 5448 2372 5500 2378
rect 5448 2314 5500 2320
rect 5356 2304 5408 2310
rect 5356 2246 5408 2252
rect 5644 800 5672 6684
rect 6012 6390 6040 10231
rect 6092 10202 6144 10208
rect 6104 9761 6132 10202
rect 6472 10198 6500 10911
rect 6460 10192 6512 10198
rect 6460 10134 6512 10140
rect 6090 9752 6146 9761
rect 6090 9687 6146 9696
rect 6366 9752 6422 9761
rect 6366 9687 6422 9696
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6104 8786 6132 9318
rect 6288 9178 6316 9318
rect 6276 9172 6328 9178
rect 6276 9114 6328 9120
rect 6104 8758 6224 8786
rect 6090 8664 6146 8673
rect 6090 8599 6146 8608
rect 6104 8294 6132 8599
rect 6196 8498 6224 8758
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 6276 8288 6328 8294
rect 6276 8230 6328 8236
rect 6288 8090 6316 8230
rect 6276 8084 6328 8090
rect 6276 8026 6328 8032
rect 6184 7472 6236 7478
rect 6184 7414 6236 7420
rect 6274 7440 6330 7449
rect 6092 7268 6144 7274
rect 6092 7210 6144 7216
rect 6000 6384 6052 6390
rect 6000 6326 6052 6332
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5736 5030 5764 5510
rect 5920 5234 5948 6054
rect 5908 5228 5960 5234
rect 5908 5170 5960 5176
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5736 4593 5764 4966
rect 5722 4584 5778 4593
rect 5722 4519 5778 4528
rect 5908 4004 5960 4010
rect 5908 3946 5960 3952
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 5828 2650 5856 3878
rect 5920 3738 5948 3946
rect 5908 3732 5960 3738
rect 5908 3674 5960 3680
rect 5908 3528 5960 3534
rect 5908 3470 5960 3476
rect 5920 3194 5948 3470
rect 6012 3369 6040 6326
rect 6104 3398 6132 7210
rect 6196 6866 6224 7414
rect 6274 7375 6330 7384
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6288 6118 6316 7375
rect 6380 6474 6408 9687
rect 6460 9512 6512 9518
rect 6460 9454 6512 9460
rect 6472 9110 6500 9454
rect 6460 9104 6512 9110
rect 6460 9046 6512 9052
rect 6472 8430 6500 9046
rect 6460 8424 6512 8430
rect 6460 8366 6512 8372
rect 6472 8294 6500 8366
rect 6460 8288 6512 8294
rect 6460 8230 6512 8236
rect 6460 7744 6512 7750
rect 6460 7686 6512 7692
rect 6472 7041 6500 7686
rect 6458 7032 6514 7041
rect 6458 6967 6514 6976
rect 6380 6446 6500 6474
rect 6366 6352 6422 6361
rect 6366 6287 6422 6296
rect 6380 6254 6408 6287
rect 6368 6248 6420 6254
rect 6368 6190 6420 6196
rect 6276 6112 6328 6118
rect 6472 6100 6500 6446
rect 6276 6054 6328 6060
rect 6380 6072 6500 6100
rect 6288 5914 6316 6054
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6184 5636 6236 5642
rect 6184 5578 6236 5584
rect 6196 5234 6224 5578
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6288 5098 6316 5510
rect 6276 5092 6328 5098
rect 6276 5034 6328 5040
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 6288 3641 6316 4082
rect 6274 3632 6330 3641
rect 6274 3567 6330 3576
rect 6092 3392 6144 3398
rect 5998 3360 6054 3369
rect 6380 3380 6408 6072
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 6472 3505 6500 3878
rect 6458 3496 6514 3505
rect 6458 3431 6514 3440
rect 6380 3352 6500 3380
rect 6092 3334 6144 3340
rect 5998 3295 6054 3304
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 6012 800 6040 3295
rect 6104 3233 6132 3334
rect 6090 3224 6146 3233
rect 6090 3159 6146 3168
rect 6368 2984 6420 2990
rect 6368 2926 6420 2932
rect 6380 2650 6408 2926
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 6368 2508 6420 2514
rect 6368 2450 6420 2456
rect 6380 2038 6408 2450
rect 6368 2032 6420 2038
rect 6368 1974 6420 1980
rect 6472 800 6500 3352
rect 6564 3194 6592 12582
rect 6656 11558 6684 12702
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6642 11384 6698 11393
rect 6642 11319 6644 11328
rect 6696 11319 6698 11328
rect 6644 11290 6696 11296
rect 6748 11234 6776 14758
rect 6828 14544 6880 14550
rect 6828 14486 6880 14492
rect 6840 12646 6868 14486
rect 6932 12646 6960 16895
rect 7208 16590 7236 17598
rect 7288 17332 7340 17338
rect 7288 17274 7340 17280
rect 7300 17202 7328 17274
rect 7288 17196 7340 17202
rect 7288 17138 7340 17144
rect 7392 16794 7420 19178
rect 7380 16788 7432 16794
rect 7380 16730 7432 16736
rect 7196 16584 7248 16590
rect 7196 16526 7248 16532
rect 7208 16250 7236 16526
rect 7196 16244 7248 16250
rect 7196 16186 7248 16192
rect 7104 15904 7156 15910
rect 7104 15846 7156 15852
rect 7116 15688 7144 15846
rect 7024 15660 7144 15688
rect 7380 15700 7432 15706
rect 7024 14618 7052 15660
rect 7380 15642 7432 15648
rect 7104 15564 7156 15570
rect 7104 15506 7156 15512
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 7116 14074 7144 15506
rect 7392 15502 7420 15642
rect 7484 15586 7512 20318
rect 7576 20058 7604 20454
rect 7852 20330 7880 22200
rect 7840 20324 7892 20330
rect 7840 20266 7892 20272
rect 7886 20156 8182 20176
rect 7942 20154 7966 20156
rect 8022 20154 8046 20156
rect 8102 20154 8126 20156
rect 7964 20102 7966 20154
rect 8028 20102 8040 20154
rect 8102 20102 8104 20154
rect 7942 20100 7966 20102
rect 8022 20100 8046 20102
rect 8102 20100 8126 20102
rect 7886 20080 8182 20100
rect 7564 20052 7616 20058
rect 7564 19994 7616 20000
rect 7564 19780 7616 19786
rect 7564 19722 7616 19728
rect 7576 19145 7604 19722
rect 7656 19712 7708 19718
rect 7656 19654 7708 19660
rect 7562 19136 7618 19145
rect 7562 19071 7618 19080
rect 7576 18426 7604 19071
rect 7668 18970 7696 19654
rect 8220 19417 8248 22200
rect 8300 19848 8352 19854
rect 8300 19790 8352 19796
rect 8206 19408 8262 19417
rect 8206 19343 8262 19352
rect 8312 19310 8340 19790
rect 8588 19417 8616 22200
rect 8852 19780 8904 19786
rect 8852 19722 8904 19728
rect 8760 19712 8812 19718
rect 8760 19654 8812 19660
rect 8574 19408 8630 19417
rect 8574 19343 8630 19352
rect 8772 19310 8800 19654
rect 8300 19304 8352 19310
rect 8300 19246 8352 19252
rect 8760 19304 8812 19310
rect 8760 19246 8812 19252
rect 7886 19068 8182 19088
rect 7942 19066 7966 19068
rect 8022 19066 8046 19068
rect 8102 19066 8126 19068
rect 7964 19014 7966 19066
rect 8028 19014 8040 19066
rect 8102 19014 8104 19066
rect 7942 19012 7966 19014
rect 8022 19012 8046 19014
rect 8102 19012 8126 19014
rect 7886 18992 8182 19012
rect 7656 18964 7708 18970
rect 7656 18906 7708 18912
rect 8116 18760 8168 18766
rect 8116 18702 8168 18708
rect 8312 18714 8340 19246
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 8404 18834 8432 19110
rect 8392 18828 8444 18834
rect 8392 18770 8444 18776
rect 7654 18592 7710 18601
rect 7654 18527 7710 18536
rect 7564 18420 7616 18426
rect 7564 18362 7616 18368
rect 7562 18048 7618 18057
rect 7562 17983 7618 17992
rect 7576 17746 7604 17983
rect 7668 17814 7696 18527
rect 8128 18426 8156 18702
rect 8312 18686 8432 18714
rect 8772 18698 8800 19246
rect 8864 19174 8892 19722
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 8864 18902 8892 19110
rect 8852 18896 8904 18902
rect 8852 18838 8904 18844
rect 8852 18760 8904 18766
rect 8852 18702 8904 18708
rect 8116 18420 8168 18426
rect 8116 18362 8168 18368
rect 7748 18080 7800 18086
rect 7748 18022 7800 18028
rect 7656 17808 7708 17814
rect 7656 17750 7708 17756
rect 7564 17740 7616 17746
rect 7564 17682 7616 17688
rect 7668 17542 7696 17750
rect 7760 17542 7788 18022
rect 7886 17980 8182 18000
rect 7942 17978 7966 17980
rect 8022 17978 8046 17980
rect 8102 17978 8126 17980
rect 7964 17926 7966 17978
rect 8028 17926 8040 17978
rect 8102 17926 8104 17978
rect 7942 17924 7966 17926
rect 8022 17924 8046 17926
rect 8102 17924 8126 17926
rect 7886 17904 8182 17924
rect 8404 17882 8432 18686
rect 8760 18692 8812 18698
rect 8760 18634 8812 18640
rect 8666 18456 8722 18465
rect 8864 18426 8892 18702
rect 8666 18391 8722 18400
rect 8852 18420 8904 18426
rect 8680 18222 8708 18391
rect 8852 18362 8904 18368
rect 8668 18216 8720 18222
rect 8668 18158 8720 18164
rect 8680 18086 8708 18158
rect 8864 18154 8892 18362
rect 8760 18148 8812 18154
rect 8760 18090 8812 18096
rect 8852 18148 8904 18154
rect 8852 18090 8904 18096
rect 8668 18080 8720 18086
rect 8668 18022 8720 18028
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8484 17672 8536 17678
rect 8484 17614 8536 17620
rect 8208 17604 8260 17610
rect 8208 17546 8260 17552
rect 8392 17604 8444 17610
rect 8392 17546 8444 17552
rect 7656 17536 7708 17542
rect 7654 17504 7656 17513
rect 7748 17536 7800 17542
rect 7708 17504 7710 17513
rect 7748 17478 7800 17484
rect 7654 17439 7710 17448
rect 8220 17377 8248 17546
rect 8206 17368 8262 17377
rect 8206 17303 8262 17312
rect 7840 17196 7892 17202
rect 7760 17156 7840 17184
rect 7564 16652 7616 16658
rect 7564 16594 7616 16600
rect 7576 16250 7604 16594
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 7484 15558 7696 15586
rect 7380 15496 7432 15502
rect 7380 15438 7432 15444
rect 7472 15496 7524 15502
rect 7472 15438 7524 15444
rect 7484 15094 7512 15438
rect 7472 15088 7524 15094
rect 7472 15030 7524 15036
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7300 14618 7328 14758
rect 7288 14612 7340 14618
rect 7288 14554 7340 14560
rect 7484 14414 7512 15030
rect 7564 14952 7616 14958
rect 7564 14894 7616 14900
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 7472 14408 7524 14414
rect 7472 14350 7524 14356
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 7104 14068 7156 14074
rect 7104 14010 7156 14016
rect 7024 13530 7052 14010
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7012 13524 7064 13530
rect 7012 13466 7064 13472
rect 7116 12986 7144 13806
rect 7208 13569 7236 14350
rect 7484 13938 7512 14350
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7392 13734 7420 13874
rect 7380 13728 7432 13734
rect 7380 13670 7432 13676
rect 7194 13560 7250 13569
rect 7194 13495 7250 13504
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7392 12850 7420 13670
rect 7576 13546 7604 14894
rect 7484 13518 7604 13546
rect 7484 13138 7512 13518
rect 7564 13184 7616 13190
rect 7484 13132 7564 13138
rect 7484 13126 7616 13132
rect 7484 13110 7604 13126
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 7380 12708 7432 12714
rect 7380 12650 7432 12656
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7300 12102 7328 12582
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 6918 11928 6974 11937
rect 6918 11863 6920 11872
rect 6972 11863 6974 11872
rect 6920 11834 6972 11840
rect 7208 11830 7236 12038
rect 7392 11898 7420 12650
rect 7484 12442 7512 13110
rect 7564 12640 7616 12646
rect 7564 12582 7616 12588
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7196 11824 7248 11830
rect 7102 11792 7158 11801
rect 6920 11756 6972 11762
rect 7196 11766 7248 11772
rect 7102 11727 7158 11736
rect 6920 11698 6972 11704
rect 6656 11206 6776 11234
rect 6656 9450 6684 11206
rect 6826 10568 6882 10577
rect 6826 10503 6882 10512
rect 6840 10470 6868 10503
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6932 10130 6960 11698
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 7024 10198 7052 10746
rect 7012 10192 7064 10198
rect 7012 10134 7064 10140
rect 6736 10124 6788 10130
rect 6736 10066 6788 10072
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6644 9444 6696 9450
rect 6644 9386 6696 9392
rect 6656 8945 6684 9386
rect 6642 8936 6698 8945
rect 6642 8871 6698 8880
rect 6748 8090 6776 10066
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6840 9042 6868 9998
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6840 8566 6868 8978
rect 7012 8900 7064 8906
rect 7012 8842 7064 8848
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6644 8016 6696 8022
rect 6644 7958 6696 7964
rect 6656 6769 6684 7958
rect 6840 7886 6868 8502
rect 6932 7954 6960 8570
rect 7024 8430 7052 8842
rect 7012 8424 7064 8430
rect 7012 8366 7064 8372
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 7024 7818 7052 8366
rect 6736 7812 6788 7818
rect 6736 7754 6788 7760
rect 7012 7812 7064 7818
rect 7012 7754 7064 7760
rect 6642 6760 6698 6769
rect 6642 6695 6698 6704
rect 6748 5642 6776 7754
rect 7116 7342 7144 11727
rect 7288 11688 7340 11694
rect 7484 11642 7512 12242
rect 7576 11762 7604 12582
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 7288 11630 7340 11636
rect 7300 11529 7328 11630
rect 7392 11614 7512 11642
rect 7286 11520 7342 11529
rect 7286 11455 7342 11464
rect 7286 11384 7342 11393
rect 7286 11319 7342 11328
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 7208 10198 7236 10406
rect 7196 10192 7248 10198
rect 7196 10134 7248 10140
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7208 8022 7236 9862
rect 7300 9110 7328 11319
rect 7392 11082 7420 11614
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7484 11354 7512 11494
rect 7668 11393 7696 15558
rect 7760 15162 7788 17156
rect 7840 17138 7892 17144
rect 8206 17096 8262 17105
rect 8206 17031 8262 17040
rect 8220 16998 8248 17031
rect 8208 16992 8260 16998
rect 8208 16934 8260 16940
rect 7886 16892 8182 16912
rect 7942 16890 7966 16892
rect 8022 16890 8046 16892
rect 8102 16890 8126 16892
rect 7964 16838 7966 16890
rect 8028 16838 8040 16890
rect 8102 16838 8104 16890
rect 7942 16836 7966 16838
rect 8022 16836 8046 16838
rect 8102 16836 8126 16838
rect 7886 16816 8182 16836
rect 8116 16720 8168 16726
rect 8116 16662 8168 16668
rect 8128 16182 8156 16662
rect 8404 16436 8432 17546
rect 8496 17134 8524 17614
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 8680 17202 8708 17274
rect 8668 17196 8720 17202
rect 8668 17138 8720 17144
rect 8484 17128 8536 17134
rect 8484 17070 8536 17076
rect 8496 16590 8524 17070
rect 8772 16794 8800 18090
rect 8852 17876 8904 17882
rect 8852 17818 8904 17824
rect 8760 16788 8812 16794
rect 8760 16730 8812 16736
rect 8484 16584 8536 16590
rect 8484 16526 8536 16532
rect 8760 16448 8812 16454
rect 8404 16408 8524 16436
rect 8116 16176 8168 16182
rect 8116 16118 8168 16124
rect 8208 15972 8260 15978
rect 8208 15914 8260 15920
rect 7886 15804 8182 15824
rect 7942 15802 7966 15804
rect 8022 15802 8046 15804
rect 8102 15802 8126 15804
rect 7964 15750 7966 15802
rect 8028 15750 8040 15802
rect 8102 15750 8104 15802
rect 7942 15748 7966 15750
rect 8022 15748 8046 15750
rect 8102 15748 8126 15750
rect 7886 15728 8182 15748
rect 8114 15600 8170 15609
rect 8036 15544 8114 15552
rect 8036 15524 8116 15544
rect 7748 15156 7800 15162
rect 7748 15098 7800 15104
rect 7760 14464 7788 15098
rect 8036 15094 8064 15524
rect 8168 15535 8170 15544
rect 8116 15506 8168 15512
rect 8220 15366 8248 15914
rect 8208 15360 8260 15366
rect 8208 15302 8260 15308
rect 8024 15088 8076 15094
rect 8024 15030 8076 15036
rect 8208 15088 8260 15094
rect 8208 15030 8260 15036
rect 7932 15020 7984 15026
rect 7932 14962 7984 14968
rect 7944 14929 7972 14962
rect 7930 14920 7986 14929
rect 7930 14855 7986 14864
rect 7886 14716 8182 14736
rect 7942 14714 7966 14716
rect 8022 14714 8046 14716
rect 8102 14714 8126 14716
rect 7964 14662 7966 14714
rect 8028 14662 8040 14714
rect 8102 14662 8104 14714
rect 7942 14660 7966 14662
rect 8022 14660 8046 14662
rect 8102 14660 8126 14662
rect 7886 14640 8182 14660
rect 8220 14550 8248 15030
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8208 14544 8260 14550
rect 8208 14486 8260 14492
rect 7840 14476 7892 14482
rect 7760 14436 7840 14464
rect 7840 14418 7892 14424
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 8128 14113 8156 14418
rect 8114 14104 8170 14113
rect 8114 14039 8170 14048
rect 8116 13864 8168 13870
rect 8114 13832 8116 13841
rect 8168 13832 8170 13841
rect 8114 13767 8170 13776
rect 7886 13628 8182 13648
rect 7942 13626 7966 13628
rect 8022 13626 8046 13628
rect 8102 13626 8126 13628
rect 7964 13574 7966 13626
rect 8028 13574 8040 13626
rect 8102 13574 8104 13626
rect 7942 13572 7966 13574
rect 8022 13572 8046 13574
rect 8102 13572 8126 13574
rect 7886 13552 8182 13572
rect 7748 13456 7800 13462
rect 7748 13398 7800 13404
rect 7654 11384 7710 11393
rect 7472 11348 7524 11354
rect 7654 11319 7710 11328
rect 7472 11290 7524 11296
rect 7472 11212 7524 11218
rect 7472 11154 7524 11160
rect 7484 11121 7512 11154
rect 7564 11144 7616 11150
rect 7470 11112 7526 11121
rect 7380 11076 7432 11082
rect 7564 11086 7616 11092
rect 7470 11047 7526 11056
rect 7380 11018 7432 11024
rect 7288 9104 7340 9110
rect 7288 9046 7340 9052
rect 7392 9042 7420 11018
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 7484 10441 7512 10542
rect 7470 10432 7526 10441
rect 7470 10367 7526 10376
rect 7472 10124 7524 10130
rect 7472 10066 7524 10072
rect 7484 9042 7512 10066
rect 7380 9036 7432 9042
rect 7380 8978 7432 8984
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7470 8936 7526 8945
rect 7470 8871 7526 8880
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7300 8362 7328 8774
rect 7484 8634 7512 8871
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7576 8514 7604 11086
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 7668 10130 7696 10950
rect 7760 10146 7788 13398
rect 8220 13394 8248 14486
rect 8404 13954 8432 14962
rect 8496 14532 8524 16408
rect 8760 16390 8812 16396
rect 8772 16250 8800 16390
rect 8760 16244 8812 16250
rect 8760 16186 8812 16192
rect 8760 15904 8812 15910
rect 8760 15846 8812 15852
rect 8772 15638 8800 15846
rect 8760 15632 8812 15638
rect 8760 15574 8812 15580
rect 8772 15502 8800 15533
rect 8760 15496 8812 15502
rect 8758 15464 8760 15473
rect 8812 15464 8814 15473
rect 8758 15399 8814 15408
rect 8668 14816 8720 14822
rect 8668 14758 8720 14764
rect 8496 14504 8616 14532
rect 8404 13926 8524 13954
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8312 13433 8340 13466
rect 8496 13462 8524 13926
rect 8484 13456 8536 13462
rect 8298 13424 8354 13433
rect 8208 13388 8260 13394
rect 8484 13398 8536 13404
rect 8298 13359 8354 13368
rect 8208 13330 8260 13336
rect 7886 12540 8182 12560
rect 7942 12538 7966 12540
rect 8022 12538 8046 12540
rect 8102 12538 8126 12540
rect 7964 12486 7966 12538
rect 8028 12486 8040 12538
rect 8102 12486 8104 12538
rect 7942 12484 7966 12486
rect 8022 12484 8046 12486
rect 8102 12484 8126 12486
rect 7886 12464 8182 12484
rect 8024 12232 8076 12238
rect 8220 12220 8248 13330
rect 8300 13184 8352 13190
rect 8588 13138 8616 14504
rect 8680 14113 8708 14758
rect 8666 14104 8722 14113
rect 8666 14039 8722 14048
rect 8772 13818 8800 15399
rect 8864 14929 8892 17818
rect 8956 16425 8984 22200
rect 9036 20052 9088 20058
rect 9036 19994 9088 20000
rect 8942 16416 8998 16425
rect 8942 16351 8998 16360
rect 8942 16144 8998 16153
rect 8942 16079 8998 16088
rect 8956 15910 8984 16079
rect 8944 15904 8996 15910
rect 8944 15846 8996 15852
rect 8944 15496 8996 15502
rect 8944 15438 8996 15444
rect 8850 14920 8906 14929
rect 8956 14890 8984 15438
rect 8850 14855 8906 14864
rect 8944 14884 8996 14890
rect 8944 14826 8996 14832
rect 8956 14346 8984 14826
rect 9048 14482 9076 19994
rect 9128 19508 9180 19514
rect 9128 19450 9180 19456
rect 9140 17882 9168 19450
rect 9312 18080 9364 18086
rect 9312 18022 9364 18028
rect 9128 17876 9180 17882
rect 9128 17818 9180 17824
rect 9220 17264 9272 17270
rect 9220 17206 9272 17212
rect 9128 16652 9180 16658
rect 9128 16594 9180 16600
rect 9140 16289 9168 16594
rect 9126 16280 9182 16289
rect 9126 16215 9182 16224
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 9140 15434 9168 16050
rect 9232 15706 9260 17206
rect 9324 16114 9352 18022
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 9220 15700 9272 15706
rect 9220 15642 9272 15648
rect 9312 15632 9364 15638
rect 9310 15600 9312 15609
rect 9364 15600 9366 15609
rect 9310 15535 9366 15544
rect 9128 15428 9180 15434
rect 9128 15370 9180 15376
rect 9140 14958 9168 15370
rect 9128 14952 9180 14958
rect 9128 14894 9180 14900
rect 9218 14920 9274 14929
rect 9218 14855 9274 14864
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 8944 14340 8996 14346
rect 8944 14282 8996 14288
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 8680 13790 8800 13818
rect 8852 13864 8904 13870
rect 8852 13806 8904 13812
rect 8680 13376 8708 13790
rect 8864 13734 8892 13806
rect 8956 13802 8984 14010
rect 9048 13938 9076 14418
rect 9232 14362 9260 14855
rect 9416 14464 9444 22200
rect 9680 19916 9732 19922
rect 9680 19858 9732 19864
rect 9692 19310 9720 19858
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9496 17264 9548 17270
rect 9494 17232 9496 17241
rect 9548 17232 9550 17241
rect 9494 17167 9550 17176
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9140 14334 9260 14362
rect 9324 14436 9444 14464
rect 9036 13932 9088 13938
rect 9036 13874 9088 13880
rect 8944 13796 8996 13802
rect 8944 13738 8996 13744
rect 8760 13728 8812 13734
rect 8758 13696 8760 13705
rect 8852 13728 8904 13734
rect 8812 13696 8814 13705
rect 8852 13670 8904 13676
rect 8758 13631 8814 13640
rect 8864 13569 8892 13670
rect 8850 13560 8906 13569
rect 8850 13495 8906 13504
rect 8680 13348 8800 13376
rect 8300 13126 8352 13132
rect 8312 12889 8340 13126
rect 8404 13110 8616 13138
rect 8298 12880 8354 12889
rect 8298 12815 8354 12824
rect 8312 12374 8340 12815
rect 8300 12368 8352 12374
rect 8300 12310 8352 12316
rect 8076 12192 8248 12220
rect 8024 12174 8076 12180
rect 7840 12096 7892 12102
rect 7840 12038 7892 12044
rect 7852 11626 7880 12038
rect 8312 11762 8340 12310
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 7840 11620 7892 11626
rect 7840 11562 7892 11568
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 7886 11452 8182 11472
rect 7942 11450 7966 11452
rect 8022 11450 8046 11452
rect 8102 11450 8126 11452
rect 7964 11398 7966 11450
rect 8028 11398 8040 11450
rect 8102 11398 8104 11450
rect 7942 11396 7966 11398
rect 8022 11396 8046 11398
rect 8102 11396 8126 11398
rect 7886 11376 8182 11396
rect 8220 11354 8248 11494
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8312 11014 8340 11494
rect 7932 11008 7984 11014
rect 7932 10950 7984 10956
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 7944 10606 7972 10950
rect 7932 10600 7984 10606
rect 7932 10542 7984 10548
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 7886 10364 8182 10384
rect 7942 10362 7966 10364
rect 8022 10362 8046 10364
rect 8102 10362 8126 10364
rect 7964 10310 7966 10362
rect 8028 10310 8040 10362
rect 8102 10310 8104 10362
rect 7942 10308 7966 10310
rect 8022 10308 8046 10310
rect 8102 10308 8126 10310
rect 7886 10288 8182 10308
rect 7656 10124 7708 10130
rect 7760 10118 7880 10146
rect 7656 10066 7708 10072
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 7760 9518 7788 9998
rect 7748 9512 7800 9518
rect 7748 9454 7800 9460
rect 7852 9364 7880 10118
rect 8220 10062 8248 10542
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8312 9994 8340 10202
rect 8404 10146 8432 13110
rect 8576 12980 8628 12986
rect 8576 12922 8628 12928
rect 8484 12776 8536 12782
rect 8482 12744 8484 12753
rect 8536 12744 8538 12753
rect 8482 12679 8538 12688
rect 8482 12472 8538 12481
rect 8482 12407 8484 12416
rect 8536 12407 8538 12416
rect 8484 12378 8536 12384
rect 8482 10704 8538 10713
rect 8482 10639 8538 10648
rect 8588 10656 8616 12922
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 8680 12442 8708 12786
rect 8772 12764 8800 13348
rect 9048 13326 9076 13874
rect 9036 13320 9088 13326
rect 8942 13288 8998 13297
rect 9036 13262 9088 13268
rect 8942 13223 8998 13232
rect 8772 12736 8892 12764
rect 8760 12640 8812 12646
rect 8760 12582 8812 12588
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 8680 11665 8708 12378
rect 8772 11898 8800 12582
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 8666 11656 8722 11665
rect 8666 11591 8722 11600
rect 8760 11620 8812 11626
rect 8680 11150 8708 11591
rect 8760 11562 8812 11568
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 8668 11008 8720 11014
rect 8668 10950 8720 10956
rect 8680 10849 8708 10950
rect 8666 10840 8722 10849
rect 8666 10775 8668 10784
rect 8720 10775 8722 10784
rect 8668 10746 8720 10752
rect 8680 10715 8708 10746
rect 8772 10713 8800 11562
rect 8864 10962 8892 12736
rect 8956 12374 8984 13223
rect 9036 13184 9088 13190
rect 9034 13152 9036 13161
rect 9088 13152 9090 13161
rect 9034 13087 9090 13096
rect 9048 12628 9076 13087
rect 9140 12986 9168 14334
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 9232 13870 9260 14214
rect 9220 13864 9272 13870
rect 9220 13806 9272 13812
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9126 12880 9182 12889
rect 9126 12815 9128 12824
rect 9180 12815 9182 12824
rect 9128 12786 9180 12792
rect 9128 12640 9180 12646
rect 9048 12600 9128 12628
rect 8944 12368 8996 12374
rect 8944 12310 8996 12316
rect 8944 12096 8996 12102
rect 8944 12038 8996 12044
rect 8956 11354 8984 12038
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 8864 10934 8984 10962
rect 8850 10840 8906 10849
rect 8850 10775 8906 10784
rect 8758 10704 8814 10713
rect 8496 10266 8524 10639
rect 8588 10628 8708 10656
rect 8758 10639 8814 10648
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8404 10118 8524 10146
rect 8300 9988 8352 9994
rect 8300 9930 8352 9936
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 7930 9480 7986 9489
rect 7930 9415 7932 9424
rect 7984 9415 7986 9424
rect 7932 9386 7984 9392
rect 7392 8486 7604 8514
rect 7760 9336 7880 9364
rect 7392 8430 7420 8486
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7288 8356 7340 8362
rect 7288 8298 7340 8304
rect 7472 8356 7524 8362
rect 7656 8356 7708 8362
rect 7472 8298 7524 8304
rect 7576 8316 7656 8344
rect 7196 8016 7248 8022
rect 7196 7958 7248 7964
rect 7300 7886 7328 8298
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7392 8090 7420 8230
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 7104 7336 7156 7342
rect 7104 7278 7156 7284
rect 7024 7002 7052 7278
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 7116 6905 7144 7278
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 7102 6896 7158 6905
rect 7102 6831 7158 6840
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6932 6322 6960 6598
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 6828 5704 6880 5710
rect 6932 5692 6960 6258
rect 7012 5908 7064 5914
rect 7064 5868 7144 5896
rect 7012 5850 7064 5856
rect 7012 5772 7064 5778
rect 7012 5714 7064 5720
rect 6880 5664 6960 5692
rect 6828 5646 6880 5652
rect 6736 5636 6788 5642
rect 6736 5578 6788 5584
rect 6644 5092 6696 5098
rect 6644 5034 6696 5040
rect 6656 4282 6684 5034
rect 6644 4276 6696 4282
rect 6644 4218 6696 4224
rect 6644 4004 6696 4010
rect 6644 3946 6696 3952
rect 6656 3534 6684 3946
rect 6748 3670 6776 5578
rect 7024 5545 7052 5714
rect 7010 5536 7066 5545
rect 7010 5471 7066 5480
rect 7024 5370 7052 5471
rect 7116 5370 7144 5868
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 7104 5364 7156 5370
rect 7104 5306 7156 5312
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 7116 4826 7144 5170
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 6736 3664 6788 3670
rect 6736 3606 6788 3612
rect 6920 3664 6972 3670
rect 6920 3606 6972 3612
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 6736 2916 6788 2922
rect 6736 2858 6788 2864
rect 6748 2378 6776 2858
rect 6736 2372 6788 2378
rect 6736 2314 6788 2320
rect 6840 800 6868 3130
rect 6932 3126 6960 3606
rect 7024 3398 7052 4014
rect 7116 3777 7144 4218
rect 7102 3768 7158 3777
rect 7102 3703 7158 3712
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 6920 3120 6972 3126
rect 6920 3062 6972 3068
rect 7024 2990 7052 3334
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 6920 2916 6972 2922
rect 6920 2858 6972 2864
rect 6932 2582 6960 2858
rect 6920 2576 6972 2582
rect 6920 2518 6972 2524
rect 6932 2106 6960 2518
rect 7208 2446 7236 6938
rect 7392 6730 7420 7346
rect 7380 6724 7432 6730
rect 7380 6666 7432 6672
rect 7392 6497 7420 6666
rect 7378 6488 7434 6497
rect 7378 6423 7434 6432
rect 7392 6322 7420 6423
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7378 6216 7434 6225
rect 7378 6151 7434 6160
rect 7288 5704 7340 5710
rect 7286 5672 7288 5681
rect 7340 5672 7342 5681
rect 7286 5607 7342 5616
rect 7286 5400 7342 5409
rect 7286 5335 7342 5344
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7208 2310 7236 2382
rect 7196 2304 7248 2310
rect 7196 2246 7248 2252
rect 6920 2100 6972 2106
rect 6920 2042 6972 2048
rect 7208 1902 7236 2246
rect 7196 1896 7248 1902
rect 7196 1838 7248 1844
rect 7300 800 7328 5335
rect 7392 5234 7420 6151
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7392 3738 7420 4966
rect 7484 4865 7512 8298
rect 7576 7449 7604 8316
rect 7656 8298 7708 8304
rect 7654 8256 7710 8265
rect 7654 8191 7710 8200
rect 7562 7440 7618 7449
rect 7562 7375 7618 7384
rect 7564 7268 7616 7274
rect 7564 7210 7616 7216
rect 7470 4856 7526 4865
rect 7470 4791 7526 4800
rect 7472 4684 7524 4690
rect 7472 4626 7524 4632
rect 7484 3942 7512 4626
rect 7576 4622 7604 7210
rect 7668 6866 7696 8191
rect 7760 7954 7788 9336
rect 7886 9276 8182 9296
rect 7942 9274 7966 9276
rect 8022 9274 8046 9276
rect 8102 9274 8126 9276
rect 7964 9222 7966 9274
rect 8028 9222 8040 9274
rect 8102 9222 8104 9274
rect 7942 9220 7966 9222
rect 8022 9220 8046 9222
rect 8102 9220 8126 9222
rect 7886 9200 8182 9220
rect 8220 9178 8248 9862
rect 8298 9752 8354 9761
rect 8298 9687 8354 9696
rect 8312 9353 8340 9687
rect 8392 9376 8444 9382
rect 8298 9344 8354 9353
rect 8392 9318 8444 9324
rect 8298 9279 8354 9288
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8024 9104 8076 9110
rect 8024 9046 8076 9052
rect 8206 9072 8262 9081
rect 7932 8832 7984 8838
rect 7932 8774 7984 8780
rect 7944 8401 7972 8774
rect 7930 8392 7986 8401
rect 8036 8362 8064 9046
rect 8206 9007 8208 9016
rect 8260 9007 8262 9016
rect 8300 9036 8352 9042
rect 8208 8978 8260 8984
rect 8300 8978 8352 8984
rect 8208 8900 8260 8906
rect 8208 8842 8260 8848
rect 7930 8327 7986 8336
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 7886 8188 8182 8208
rect 7942 8186 7966 8188
rect 8022 8186 8046 8188
rect 8102 8186 8126 8188
rect 7964 8134 7966 8186
rect 8028 8134 8040 8186
rect 8102 8134 8104 8186
rect 7942 8132 7966 8134
rect 8022 8132 8046 8134
rect 8102 8132 8126 8134
rect 7886 8112 8182 8132
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7748 7812 7800 7818
rect 7748 7754 7800 7760
rect 7760 7342 7788 7754
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 8036 7274 8064 7482
rect 8220 7426 8248 8842
rect 8312 8090 8340 8978
rect 8404 8498 8432 9318
rect 8496 9110 8524 10118
rect 8576 9716 8628 9722
rect 8576 9658 8628 9664
rect 8588 9382 8616 9658
rect 8576 9376 8628 9382
rect 8576 9318 8628 9324
rect 8484 9104 8536 9110
rect 8484 9046 8536 9052
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8390 8256 8446 8265
rect 8390 8191 8446 8200
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8312 7546 8340 7890
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8404 7426 8432 8191
rect 8496 7818 8524 8434
rect 8484 7812 8536 7818
rect 8484 7754 8536 7760
rect 8220 7398 8432 7426
rect 8024 7268 8076 7274
rect 8024 7210 8076 7216
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 7886 7100 8182 7120
rect 7942 7098 7966 7100
rect 8022 7098 8046 7100
rect 8102 7098 8126 7100
rect 7964 7046 7966 7098
rect 8028 7046 8040 7098
rect 8102 7046 8104 7098
rect 7942 7044 7966 7046
rect 8022 7044 8046 7046
rect 8102 7044 8126 7046
rect 7886 7024 8182 7044
rect 8022 6896 8078 6905
rect 7656 6860 7708 6866
rect 8022 6831 8078 6840
rect 7656 6802 7708 6808
rect 8036 6798 8064 6831
rect 7840 6792 7892 6798
rect 7838 6760 7840 6769
rect 8024 6792 8076 6798
rect 7892 6760 7894 6769
rect 8024 6734 8076 6740
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 7838 6695 7894 6704
rect 8116 6724 8168 6730
rect 8116 6666 8168 6672
rect 7838 6624 7894 6633
rect 7838 6559 7894 6568
rect 7852 6186 7880 6559
rect 8128 6361 8156 6666
rect 8220 6390 8248 6734
rect 8312 6730 8340 7142
rect 8300 6724 8352 6730
rect 8300 6666 8352 6672
rect 8404 6610 8432 7398
rect 8496 6746 8524 7754
rect 8588 7721 8616 9318
rect 8680 8022 8708 10628
rect 8758 10296 8814 10305
rect 8758 10231 8814 10240
rect 8772 10130 8800 10231
rect 8864 10198 8892 10775
rect 8956 10674 8984 10934
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 8956 10538 8984 10610
rect 8944 10532 8996 10538
rect 8944 10474 8996 10480
rect 8942 10432 8998 10441
rect 8942 10367 8998 10376
rect 8852 10192 8904 10198
rect 8852 10134 8904 10140
rect 8760 10124 8812 10130
rect 8760 10066 8812 10072
rect 8772 9722 8800 10066
rect 8956 9908 8984 10367
rect 8864 9880 8984 9908
rect 8760 9716 8812 9722
rect 8760 9658 8812 9664
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 8772 9382 8800 9522
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8772 8634 8800 9318
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8864 8378 8892 9880
rect 8942 9752 8998 9761
rect 8942 9687 8998 9696
rect 8956 9382 8984 9687
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 9048 9217 9076 12600
rect 9128 12582 9180 12588
rect 9128 12300 9180 12306
rect 9128 12242 9180 12248
rect 9034 9208 9090 9217
rect 9034 9143 9090 9152
rect 9036 9104 9088 9110
rect 9036 9046 9088 9052
rect 8772 8350 8892 8378
rect 8668 8016 8720 8022
rect 8668 7958 8720 7964
rect 8574 7712 8630 7721
rect 8574 7647 8630 7656
rect 8680 6866 8708 7958
rect 8772 7750 8800 8350
rect 9048 8294 9076 9046
rect 8852 8288 8904 8294
rect 8852 8230 8904 8236
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8496 6718 8708 6746
rect 8312 6582 8432 6610
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8208 6384 8260 6390
rect 8114 6352 8170 6361
rect 8208 6326 8260 6332
rect 8114 6287 8170 6296
rect 8128 6186 8156 6287
rect 7840 6180 7892 6186
rect 7840 6122 7892 6128
rect 8116 6180 8168 6186
rect 8116 6122 8168 6128
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7668 5098 7696 6054
rect 7760 5914 7788 6054
rect 7886 6012 8182 6032
rect 7942 6010 7966 6012
rect 8022 6010 8046 6012
rect 8102 6010 8126 6012
rect 7964 5958 7966 6010
rect 8028 5958 8040 6010
rect 8102 5958 8104 6010
rect 7942 5956 7966 5958
rect 8022 5956 8046 5958
rect 8102 5956 8126 5958
rect 7886 5936 8182 5956
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 7760 5234 7788 5510
rect 7852 5370 7880 5714
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 7656 5092 7708 5098
rect 7656 5034 7708 5040
rect 7944 5012 7972 5170
rect 8036 5098 8064 5510
rect 8024 5092 8076 5098
rect 8024 5034 8076 5040
rect 7760 4984 7972 5012
rect 7654 4856 7710 4865
rect 7654 4791 7710 4800
rect 7564 4616 7616 4622
rect 7564 4558 7616 4564
rect 7576 3942 7604 4558
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 7484 1630 7512 3538
rect 7564 2916 7616 2922
rect 7564 2858 7616 2864
rect 7576 2582 7604 2858
rect 7564 2576 7616 2582
rect 7564 2518 7616 2524
rect 7472 1624 7524 1630
rect 7472 1566 7524 1572
rect 7668 800 7696 4791
rect 7760 4078 7788 4984
rect 7886 4924 8182 4944
rect 7942 4922 7966 4924
rect 8022 4922 8046 4924
rect 8102 4922 8126 4924
rect 7964 4870 7966 4922
rect 8028 4870 8040 4922
rect 8102 4870 8104 4922
rect 7942 4868 7966 4870
rect 8022 4868 8046 4870
rect 8102 4868 8126 4870
rect 7886 4848 8182 4868
rect 8312 4706 8340 6582
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 8404 5710 8432 6258
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8392 5364 8444 5370
rect 8392 5306 8444 5312
rect 8404 4826 8432 5306
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8496 4729 8524 6598
rect 8574 5944 8630 5953
rect 8574 5879 8576 5888
rect 8628 5879 8630 5888
rect 8576 5850 8628 5856
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8482 4720 8538 4729
rect 8312 4678 8432 4706
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 7760 3194 7788 4014
rect 8220 4010 8248 4558
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8208 4004 8260 4010
rect 8208 3946 8260 3952
rect 7886 3836 8182 3856
rect 7942 3834 7966 3836
rect 8022 3834 8046 3836
rect 8102 3834 8126 3836
rect 7964 3782 7966 3834
rect 8028 3782 8040 3834
rect 8102 3782 8104 3834
rect 7942 3780 7966 3782
rect 8022 3780 8046 3782
rect 8102 3780 8126 3782
rect 7886 3760 8182 3780
rect 8220 3738 8248 3946
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8312 3505 8340 4082
rect 8298 3496 8354 3505
rect 7840 3460 7892 3466
rect 8298 3431 8354 3440
rect 7840 3402 7892 3408
rect 7748 3188 7800 3194
rect 7748 3130 7800 3136
rect 7746 3088 7802 3097
rect 7746 3023 7802 3032
rect 7760 2825 7788 3023
rect 7852 2990 7880 3402
rect 7840 2984 7892 2990
rect 7840 2926 7892 2932
rect 7746 2816 7802 2825
rect 7746 2751 7802 2760
rect 7760 2514 7788 2751
rect 7886 2748 8182 2768
rect 7942 2746 7966 2748
rect 8022 2746 8046 2748
rect 8102 2746 8126 2748
rect 7964 2694 7966 2746
rect 8028 2694 8040 2746
rect 8102 2694 8104 2746
rect 7942 2692 7966 2694
rect 8022 2692 8046 2694
rect 8102 2692 8126 2694
rect 7886 2672 8182 2692
rect 8404 2632 8432 4678
rect 8482 4655 8538 4664
rect 8588 4554 8616 5646
rect 8680 5302 8708 6718
rect 8760 6112 8812 6118
rect 8760 6054 8812 6060
rect 8772 5574 8800 6054
rect 8760 5568 8812 5574
rect 8760 5510 8812 5516
rect 8668 5296 8720 5302
rect 8668 5238 8720 5244
rect 8760 5092 8812 5098
rect 8760 5034 8812 5040
rect 8772 4826 8800 5034
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 8864 4706 8892 8230
rect 8942 8120 8998 8129
rect 8942 8055 8944 8064
rect 8996 8055 8998 8064
rect 8944 8026 8996 8032
rect 8944 7812 8996 7818
rect 8944 7754 8996 7760
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 8772 4678 8892 4706
rect 8576 4548 8628 4554
rect 8576 4490 8628 4496
rect 8484 4480 8536 4486
rect 8484 4422 8536 4428
rect 8496 2990 8524 4422
rect 8574 4312 8630 4321
rect 8574 4247 8630 4256
rect 8588 3913 8616 4247
rect 8574 3904 8630 3913
rect 8574 3839 8630 3848
rect 8680 3738 8708 4626
rect 8772 4282 8800 4678
rect 8852 4616 8904 4622
rect 8852 4558 8904 4564
rect 8760 4276 8812 4282
rect 8760 4218 8812 4224
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 8576 3664 8628 3670
rect 8574 3632 8576 3641
rect 8628 3632 8630 3641
rect 8574 3567 8630 3576
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 8482 2816 8538 2825
rect 8482 2751 8538 2760
rect 8128 2604 8432 2632
rect 7748 2508 7800 2514
rect 7748 2450 7800 2456
rect 8128 800 8156 2604
rect 8496 800 8524 2751
rect 8680 2446 8708 3334
rect 8772 2972 8800 4218
rect 8864 3942 8892 4558
rect 8956 4146 8984 7754
rect 9048 7274 9076 8230
rect 9140 8022 9168 12242
rect 9232 11014 9260 13806
rect 9324 13297 9352 14436
rect 9404 14340 9456 14346
rect 9404 14282 9456 14288
rect 9416 13938 9444 14282
rect 9404 13932 9456 13938
rect 9404 13874 9456 13880
rect 9508 13569 9536 16934
rect 9494 13560 9550 13569
rect 9494 13495 9496 13504
rect 9548 13495 9550 13504
rect 9496 13466 9548 13472
rect 9310 13288 9366 13297
rect 9310 13223 9366 13232
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 9324 12889 9352 13126
rect 9310 12880 9366 12889
rect 9310 12815 9366 12824
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 9324 12617 9352 12718
rect 9310 12608 9366 12617
rect 9310 12543 9366 12552
rect 9402 12336 9458 12345
rect 9402 12271 9458 12280
rect 9416 12238 9444 12271
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 9508 11762 9536 12786
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9600 11642 9628 17138
rect 9680 17128 9732 17134
rect 9678 17096 9680 17105
rect 9732 17096 9734 17105
rect 9678 17031 9734 17040
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9692 13530 9720 16594
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9784 12374 9812 22200
rect 9864 20528 9916 20534
rect 9864 20470 9916 20476
rect 9876 19310 9904 20470
rect 9956 19916 10008 19922
rect 9956 19858 10008 19864
rect 9864 19304 9916 19310
rect 9864 19246 9916 19252
rect 9862 19000 9918 19009
rect 9862 18935 9918 18944
rect 9876 18698 9904 18935
rect 9864 18692 9916 18698
rect 9864 18634 9916 18640
rect 9864 18216 9916 18222
rect 9864 18158 9916 18164
rect 9876 18057 9904 18158
rect 9862 18048 9918 18057
rect 9862 17983 9918 17992
rect 9968 17898 9996 19858
rect 10152 19446 10180 22200
rect 10140 19440 10192 19446
rect 10140 19382 10192 19388
rect 10140 19168 10192 19174
rect 10140 19110 10192 19116
rect 10152 18970 10180 19110
rect 10140 18964 10192 18970
rect 10140 18906 10192 18912
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 10140 18216 10192 18222
rect 10140 18158 10192 18164
rect 10152 18086 10180 18158
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 9959 17870 9996 17898
rect 10244 17882 10272 18702
rect 10416 18624 10468 18630
rect 10416 18566 10468 18572
rect 10324 18148 10376 18154
rect 10324 18090 10376 18096
rect 10232 17876 10284 17882
rect 9959 17796 9987 17870
rect 10232 17818 10284 17824
rect 9959 17768 9996 17796
rect 9864 17604 9916 17610
rect 9864 17546 9916 17552
rect 9876 17338 9904 17546
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9862 17232 9918 17241
rect 9862 17167 9864 17176
rect 9916 17167 9918 17176
rect 9864 17138 9916 17144
rect 9968 16794 9996 17768
rect 10140 17536 10192 17542
rect 10140 17478 10192 17484
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 9864 16516 9916 16522
rect 9864 16458 9916 16464
rect 9876 15978 9904 16458
rect 9864 15972 9916 15978
rect 9864 15914 9916 15920
rect 9876 15706 9904 15914
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 9968 15162 9996 15506
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9876 14618 9904 14894
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 9968 13954 9996 14350
rect 10060 14113 10088 15846
rect 10152 14929 10180 17478
rect 10230 15600 10286 15609
rect 10230 15535 10286 15544
rect 10138 14920 10194 14929
rect 10138 14855 10194 14864
rect 10140 14816 10192 14822
rect 10140 14758 10192 14764
rect 10046 14104 10102 14113
rect 10046 14039 10102 14048
rect 9864 13932 9916 13938
rect 9968 13926 10088 13954
rect 10152 13938 10180 14758
rect 10244 14618 10272 15535
rect 10336 14657 10364 18090
rect 10428 17882 10456 18566
rect 10416 17876 10468 17882
rect 10416 17818 10468 17824
rect 10520 16833 10548 22200
rect 10888 20058 10916 22200
rect 11256 20058 11284 22200
rect 11352 20700 11648 20720
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11430 20646 11432 20698
rect 11494 20646 11506 20698
rect 11568 20646 11570 20698
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11352 20624 11648 20644
rect 11716 20602 11744 22200
rect 11704 20596 11756 20602
rect 11704 20538 11756 20544
rect 12084 20058 12112 22200
rect 10876 20052 10928 20058
rect 10876 19994 10928 20000
rect 11244 20052 11296 20058
rect 11244 19994 11296 20000
rect 12072 20052 12124 20058
rect 12072 19994 12124 20000
rect 10876 19916 10928 19922
rect 10876 19858 10928 19864
rect 12164 19916 12216 19922
rect 12164 19858 12216 19864
rect 10600 19440 10652 19446
rect 10600 19382 10652 19388
rect 10612 17542 10640 19382
rect 10888 19378 10916 19858
rect 11352 19612 11648 19632
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11430 19558 11432 19610
rect 11494 19558 11506 19610
rect 11568 19558 11570 19610
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11352 19536 11648 19556
rect 10876 19372 10928 19378
rect 10876 19314 10928 19320
rect 10968 19372 11020 19378
rect 10968 19314 11020 19320
rect 11980 19372 12032 19378
rect 11980 19314 12032 19320
rect 10876 19168 10928 19174
rect 10876 19110 10928 19116
rect 10784 18216 10836 18222
rect 10784 18158 10836 18164
rect 10692 17808 10744 17814
rect 10692 17750 10744 17756
rect 10600 17536 10652 17542
rect 10600 17478 10652 17484
rect 10506 16824 10562 16833
rect 10506 16759 10562 16768
rect 10508 16720 10560 16726
rect 10508 16662 10560 16668
rect 10416 14816 10468 14822
rect 10414 14784 10416 14793
rect 10468 14784 10470 14793
rect 10414 14719 10470 14728
rect 10322 14648 10378 14657
rect 10232 14612 10284 14618
rect 10322 14583 10378 14592
rect 10232 14554 10284 14560
rect 10520 14396 10548 16662
rect 10704 16250 10732 17750
rect 10796 17678 10824 18158
rect 10888 17882 10916 19110
rect 10980 18222 11008 19314
rect 11704 19304 11756 19310
rect 11164 19242 11560 19258
rect 11704 19246 11756 19252
rect 11152 19236 11560 19242
rect 11204 19230 11560 19236
rect 11152 19178 11204 19184
rect 11336 19168 11388 19174
rect 11336 19110 11388 19116
rect 11348 19009 11376 19110
rect 11334 19000 11390 19009
rect 11072 18924 11284 18952
rect 11334 18935 11390 18944
rect 11532 18952 11560 19230
rect 11612 18964 11664 18970
rect 11532 18924 11612 18952
rect 11072 18601 11100 18924
rect 11256 18834 11284 18924
rect 11612 18906 11664 18912
rect 11152 18828 11204 18834
rect 11152 18770 11204 18776
rect 11244 18828 11296 18834
rect 11244 18770 11296 18776
rect 11058 18592 11114 18601
rect 11058 18527 11114 18536
rect 10968 18216 11020 18222
rect 10968 18158 11020 18164
rect 11164 18086 11192 18770
rect 11352 18524 11648 18544
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11430 18470 11432 18522
rect 11494 18470 11506 18522
rect 11568 18470 11570 18522
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11352 18448 11648 18468
rect 11336 18352 11388 18358
rect 11336 18294 11388 18300
rect 11152 18080 11204 18086
rect 11152 18022 11204 18028
rect 11348 17898 11376 18294
rect 11520 18216 11572 18222
rect 11520 18158 11572 18164
rect 10876 17876 10928 17882
rect 10876 17818 10928 17824
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 11164 17870 11376 17898
rect 11532 17882 11560 18158
rect 11716 17882 11744 19246
rect 11992 18630 12020 19314
rect 12072 19304 12124 19310
rect 12072 19246 12124 19252
rect 12084 18834 12112 19246
rect 12072 18828 12124 18834
rect 12072 18770 12124 18776
rect 12072 18692 12124 18698
rect 12072 18634 12124 18640
rect 11796 18624 11848 18630
rect 11796 18566 11848 18572
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11808 18290 11836 18566
rect 11796 18284 11848 18290
rect 11796 18226 11848 18232
rect 11992 18154 12020 18566
rect 11980 18148 12032 18154
rect 11980 18090 12032 18096
rect 10784 17672 10836 17678
rect 10784 17614 10836 17620
rect 10796 17202 10824 17614
rect 10966 17368 11022 17377
rect 10966 17303 11022 17312
rect 10784 17196 10836 17202
rect 10784 17138 10836 17144
rect 10980 16794 11008 17303
rect 11072 17134 11100 17818
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 10968 16788 11020 16794
rect 10968 16730 11020 16736
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 10692 16244 10744 16250
rect 10692 16186 10744 16192
rect 10600 15156 10652 15162
rect 10600 15098 10652 15104
rect 10428 14368 10548 14396
rect 9864 13874 9916 13880
rect 9876 13462 9904 13874
rect 10060 13870 10088 13926
rect 10140 13932 10192 13938
rect 10140 13874 10192 13880
rect 10048 13864 10100 13870
rect 9954 13832 10010 13841
rect 10048 13806 10100 13812
rect 9954 13767 10010 13776
rect 10324 13796 10376 13802
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 9864 13252 9916 13258
rect 9864 13194 9916 13200
rect 9772 12368 9824 12374
rect 9772 12310 9824 12316
rect 9784 11762 9812 12310
rect 9876 12238 9904 13194
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 9968 11812 9996 13767
rect 10324 13738 10376 13744
rect 10138 13560 10194 13569
rect 10138 13495 10194 13504
rect 10152 13326 10180 13495
rect 10336 13462 10364 13738
rect 10324 13456 10376 13462
rect 10324 13398 10376 13404
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10428 13258 10456 14368
rect 10612 14346 10640 15098
rect 10876 15020 10928 15026
rect 10876 14962 10928 14968
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 10600 14340 10652 14346
rect 10600 14282 10652 14288
rect 10508 14000 10560 14006
rect 10508 13942 10560 13948
rect 10520 13530 10548 13942
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 10612 13326 10640 14282
rect 10796 14278 10824 14554
rect 10888 14414 10916 14962
rect 11072 14618 11100 16594
rect 11164 16114 11192 17870
rect 11242 17776 11298 17785
rect 11242 17711 11244 17720
rect 11296 17711 11298 17720
rect 11244 17682 11296 17688
rect 11348 17678 11376 17870
rect 11520 17876 11572 17882
rect 11520 17818 11572 17824
rect 11704 17876 11756 17882
rect 11704 17818 11756 17824
rect 11980 17876 12032 17882
rect 11980 17818 12032 17824
rect 11796 17740 11848 17746
rect 11796 17682 11848 17688
rect 11336 17672 11388 17678
rect 11336 17614 11388 17620
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 11612 17196 11664 17202
rect 11612 17138 11664 17144
rect 11336 17128 11388 17134
rect 11336 17070 11388 17076
rect 11348 16561 11376 17070
rect 11624 16726 11652 17138
rect 11704 17060 11756 17066
rect 11704 17002 11756 17008
rect 11612 16720 11664 16726
rect 11612 16662 11664 16668
rect 11334 16552 11390 16561
rect 11334 16487 11336 16496
rect 11388 16487 11390 16496
rect 11336 16458 11388 16464
rect 11348 16427 11376 16458
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 11164 15910 11192 16050
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 11152 15428 11204 15434
rect 11152 15370 11204 15376
rect 11164 14618 11192 15370
rect 11244 15360 11296 15366
rect 11244 15302 11296 15308
rect 11256 15094 11284 15302
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 11244 15088 11296 15094
rect 11244 15030 11296 15036
rect 11060 14612 11112 14618
rect 11060 14554 11112 14560
rect 11152 14612 11204 14618
rect 11152 14554 11204 14560
rect 10876 14408 10928 14414
rect 10876 14350 10928 14356
rect 10968 14408 11020 14414
rect 10968 14350 11020 14356
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10600 13320 10652 13326
rect 10506 13288 10562 13297
rect 10416 13252 10468 13258
rect 10600 13262 10652 13268
rect 10506 13223 10562 13232
rect 10416 13194 10468 13200
rect 10140 12912 10192 12918
rect 10140 12854 10192 12860
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 10060 12442 10088 12718
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 10152 12345 10180 12854
rect 10520 12782 10548 13223
rect 10690 12880 10746 12889
rect 10690 12815 10746 12824
rect 10508 12776 10560 12782
rect 10508 12718 10560 12724
rect 10138 12336 10194 12345
rect 10138 12271 10194 12280
rect 10152 11898 10180 12271
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10048 11824 10100 11830
rect 9968 11784 10048 11812
rect 10048 11766 10100 11772
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9416 11614 9628 11642
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 9232 10169 9260 10950
rect 9312 10736 9364 10742
rect 9312 10678 9364 10684
rect 9218 10160 9274 10169
rect 9218 10095 9274 10104
rect 9232 10062 9260 10095
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9324 9994 9352 10678
rect 9312 9988 9364 9994
rect 9312 9930 9364 9936
rect 9218 9888 9274 9897
rect 9218 9823 9274 9832
rect 9128 8016 9180 8022
rect 9128 7958 9180 7964
rect 9036 7268 9088 7274
rect 9036 7210 9088 7216
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 9048 5710 9076 6598
rect 9232 6118 9260 9823
rect 9324 9761 9352 9930
rect 9310 9752 9366 9761
rect 9310 9687 9366 9696
rect 9416 9466 9444 11614
rect 10060 11558 10088 11766
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 9692 11150 9720 11494
rect 9770 11384 9826 11393
rect 10138 11384 10194 11393
rect 9770 11319 9826 11328
rect 9956 11348 10008 11354
rect 9784 11218 9812 11319
rect 10138 11319 10194 11328
rect 9956 11290 10008 11296
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9508 10674 9536 11086
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 9508 10130 9536 10610
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9600 10062 9628 10610
rect 9692 10470 9720 10746
rect 9784 10606 9812 11154
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9770 10432 9826 10441
rect 9770 10367 9826 10376
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 9496 9716 9548 9722
rect 9496 9658 9548 9664
rect 9324 9438 9444 9466
rect 9324 9364 9352 9438
rect 9324 9336 9444 9364
rect 9310 9208 9366 9217
rect 9310 9143 9366 9152
rect 9324 7818 9352 9143
rect 9312 7812 9364 7818
rect 9312 7754 9364 7760
rect 9312 7472 9364 7478
rect 9312 7414 9364 7420
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 9126 5808 9182 5817
rect 9126 5743 9182 5752
rect 9036 5704 9088 5710
rect 9034 5672 9036 5681
rect 9088 5672 9090 5681
rect 9034 5607 9090 5616
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8852 3936 8904 3942
rect 8852 3878 8904 3884
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8956 3670 8984 3878
rect 8944 3664 8996 3670
rect 8944 3606 8996 3612
rect 8942 3360 8998 3369
rect 8942 3295 8998 3304
rect 8956 3097 8984 3295
rect 8942 3088 8998 3097
rect 9048 3074 9076 5607
rect 9140 4826 9168 5743
rect 9220 5092 9272 5098
rect 9220 5034 9272 5040
rect 9232 4865 9260 5034
rect 9218 4856 9274 4865
rect 9128 4820 9180 4826
rect 9218 4791 9274 4800
rect 9128 4762 9180 4768
rect 9140 4690 9168 4762
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 9128 4548 9180 4554
rect 9128 4490 9180 4496
rect 9140 4321 9168 4490
rect 9126 4312 9182 4321
rect 9126 4247 9182 4256
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 9140 3194 9168 4082
rect 9220 3664 9272 3670
rect 9220 3606 9272 3612
rect 9232 3233 9260 3606
rect 9324 3398 9352 7414
rect 9416 6798 9444 9336
rect 9508 8838 9536 9658
rect 9600 9518 9628 9998
rect 9588 9512 9640 9518
rect 9588 9454 9640 9460
rect 9600 8838 9628 9454
rect 9784 9058 9812 10367
rect 9876 9926 9904 10542
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9876 9110 9904 9862
rect 9692 9030 9812 9058
rect 9864 9104 9916 9110
rect 9864 9046 9916 9052
rect 9692 8956 9720 9030
rect 9864 8968 9916 8974
rect 9692 8928 9812 8956
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9600 8566 9628 8774
rect 9588 8560 9640 8566
rect 9784 8514 9812 8928
rect 9864 8910 9916 8916
rect 9588 8502 9640 8508
rect 9496 8356 9548 8362
rect 9496 8298 9548 8304
rect 9508 7886 9536 8298
rect 9600 7954 9628 8502
rect 9692 8486 9812 8514
rect 9588 7948 9640 7954
rect 9588 7890 9640 7896
rect 9496 7880 9548 7886
rect 9494 7848 9496 7857
rect 9548 7848 9550 7857
rect 9494 7783 9550 7792
rect 9508 7410 9536 7783
rect 9586 7440 9642 7449
rect 9496 7404 9548 7410
rect 9586 7375 9642 7384
rect 9496 7346 9548 7352
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9416 6633 9444 6734
rect 9402 6624 9458 6633
rect 9402 6559 9458 6568
rect 9600 6458 9628 7375
rect 9588 6452 9640 6458
rect 9588 6394 9640 6400
rect 9692 5914 9720 8486
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9784 7750 9812 8366
rect 9876 7936 9904 8910
rect 9968 8072 9996 11290
rect 10152 11286 10180 11319
rect 10140 11280 10192 11286
rect 10140 11222 10192 11228
rect 10048 10532 10100 10538
rect 10048 10474 10100 10480
rect 10060 9586 10088 10474
rect 10140 10192 10192 10198
rect 10140 10134 10192 10140
rect 10152 9722 10180 10134
rect 10140 9716 10192 9722
rect 10140 9658 10192 9664
rect 10048 9580 10100 9586
rect 10048 9522 10100 9528
rect 10048 9444 10100 9450
rect 10048 9386 10100 9392
rect 10060 8498 10088 9386
rect 10152 9178 10180 9658
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10152 8634 10180 8910
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 10138 8392 10194 8401
rect 10138 8327 10194 8336
rect 9968 8044 10088 8072
rect 9956 7948 10008 7954
rect 9876 7908 9956 7936
rect 9956 7890 10008 7896
rect 9864 7812 9916 7818
rect 9864 7754 9916 7760
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9784 7410 9812 7686
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9680 5908 9732 5914
rect 9680 5850 9732 5856
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9416 5370 9444 5646
rect 9508 5574 9536 5714
rect 9496 5568 9548 5574
rect 9588 5568 9640 5574
rect 9496 5510 9548 5516
rect 9586 5536 9588 5545
rect 9640 5536 9642 5545
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9416 3754 9444 5306
rect 9508 4690 9536 5510
rect 9586 5471 9642 5480
rect 9680 5024 9732 5030
rect 9678 4992 9680 5001
rect 9732 4992 9734 5001
rect 9678 4927 9734 4936
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 9508 4214 9536 4626
rect 9680 4616 9732 4622
rect 9586 4584 9642 4593
rect 9680 4558 9732 4564
rect 9586 4519 9588 4528
rect 9640 4519 9642 4528
rect 9588 4490 9640 4496
rect 9496 4208 9548 4214
rect 9496 4150 9548 4156
rect 9692 4078 9720 4558
rect 9784 4214 9812 7346
rect 9876 6202 9904 7754
rect 9968 7206 9996 7890
rect 10060 7546 10088 8044
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 10060 7206 10088 7346
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 10048 7200 10100 7206
rect 10048 7142 10100 7148
rect 9968 7002 9996 7142
rect 9956 6996 10008 7002
rect 9956 6938 10008 6944
rect 9876 6174 9996 6202
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9772 4208 9824 4214
rect 9772 4150 9824 4156
rect 9876 4078 9904 6054
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 9508 3942 9536 4014
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9416 3726 9536 3754
rect 9692 3738 9720 4014
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9404 3664 9456 3670
rect 9404 3606 9456 3612
rect 9416 3505 9444 3606
rect 9508 3534 9536 3726
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9496 3528 9548 3534
rect 9402 3496 9458 3505
rect 9496 3470 9548 3476
rect 9402 3431 9458 3440
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9218 3224 9274 3233
rect 9128 3188 9180 3194
rect 9218 3159 9274 3168
rect 9128 3130 9180 3136
rect 9048 3046 9260 3074
rect 8942 3023 8998 3032
rect 9128 2984 9180 2990
rect 8772 2944 8984 2972
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 8680 1970 8708 2382
rect 8668 1964 8720 1970
rect 8668 1906 8720 1912
rect 8956 800 8984 2944
rect 9034 2952 9090 2961
rect 9128 2926 9180 2932
rect 9034 2887 9036 2896
rect 9088 2887 9090 2896
rect 9036 2858 9088 2864
rect 9048 2310 9076 2858
rect 9140 2417 9168 2926
rect 9126 2408 9182 2417
rect 9126 2343 9182 2352
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 9048 1698 9076 2246
rect 9232 2106 9260 3046
rect 9508 2904 9536 3470
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9600 3058 9628 3334
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9588 2916 9640 2922
rect 9508 2876 9588 2904
rect 9588 2858 9640 2864
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 9416 2689 9444 2790
rect 9402 2680 9458 2689
rect 9324 2624 9402 2632
rect 9324 2604 9404 2624
rect 9220 2100 9272 2106
rect 9220 2042 9272 2048
rect 9324 1766 9352 2604
rect 9456 2615 9458 2624
rect 9404 2586 9456 2592
rect 9416 2555 9444 2586
rect 9692 2582 9720 3674
rect 9784 2650 9812 3878
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 9680 2576 9732 2582
rect 9680 2518 9732 2524
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 9784 2378 9812 2450
rect 9772 2372 9824 2378
rect 9772 2314 9824 2320
rect 9404 2100 9456 2106
rect 9404 2042 9456 2048
rect 9312 1760 9364 1766
rect 9312 1702 9364 1708
rect 9036 1692 9088 1698
rect 9036 1634 9088 1640
rect 9416 800 9444 2042
rect 9876 1442 9904 3674
rect 9968 2582 9996 6174
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 10060 4826 10088 6054
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 10048 4208 10100 4214
rect 10048 4150 10100 4156
rect 10060 2961 10088 4150
rect 10046 2952 10102 2961
rect 10046 2887 10102 2896
rect 10152 2650 10180 8327
rect 10244 7410 10272 12174
rect 10520 11898 10548 12718
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 10506 11792 10562 11801
rect 10506 11727 10562 11736
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10336 10538 10364 11494
rect 10520 11286 10548 11727
rect 10612 11354 10640 12174
rect 10704 11898 10732 12815
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10508 11280 10560 11286
rect 10414 11248 10470 11257
rect 10508 11222 10560 11228
rect 10414 11183 10470 11192
rect 10324 10532 10376 10538
rect 10324 10474 10376 10480
rect 10428 9761 10456 11183
rect 10506 10704 10562 10713
rect 10506 10639 10562 10648
rect 10414 9752 10470 9761
rect 10414 9687 10470 9696
rect 10324 9104 10376 9110
rect 10324 9046 10376 9052
rect 10336 8888 10364 9046
rect 10428 9042 10456 9687
rect 10520 9450 10548 10639
rect 10690 9888 10746 9897
rect 10690 9823 10746 9832
rect 10508 9444 10560 9450
rect 10508 9386 10560 9392
rect 10520 9110 10548 9386
rect 10600 9172 10652 9178
rect 10600 9114 10652 9120
rect 10508 9104 10560 9110
rect 10508 9046 10560 9052
rect 10416 9036 10468 9042
rect 10416 8978 10468 8984
rect 10416 8900 10468 8906
rect 10336 8860 10416 8888
rect 10416 8842 10468 8848
rect 10612 8616 10640 9114
rect 10704 8906 10732 9823
rect 10692 8900 10744 8906
rect 10692 8842 10744 8848
rect 10336 8588 10640 8616
rect 10336 8090 10364 8588
rect 10508 8492 10560 8498
rect 10428 8452 10508 8480
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 10428 7857 10456 8452
rect 10508 8434 10560 8440
rect 10598 8392 10654 8401
rect 10598 8327 10654 8336
rect 10692 8356 10744 8362
rect 10414 7848 10470 7857
rect 10414 7783 10470 7792
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10336 7002 10364 7686
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 10416 7268 10468 7274
rect 10416 7210 10468 7216
rect 10428 7041 10456 7210
rect 10414 7032 10470 7041
rect 10324 6996 10376 7002
rect 10414 6967 10470 6976
rect 10324 6938 10376 6944
rect 10324 6792 10376 6798
rect 10244 6752 10324 6780
rect 10244 3738 10272 6752
rect 10324 6734 10376 6740
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 10336 6186 10364 6598
rect 10324 6180 10376 6186
rect 10324 6122 10376 6128
rect 10324 5772 10376 5778
rect 10324 5714 10376 5720
rect 10336 4622 10364 5714
rect 10520 5114 10548 7482
rect 10612 6730 10640 8327
rect 10692 8298 10744 8304
rect 10704 7954 10732 8298
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 10692 7812 10744 7818
rect 10692 7754 10744 7760
rect 10704 7546 10732 7754
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 10704 6769 10732 7346
rect 10796 7274 10824 14214
rect 10980 14074 11008 14350
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 11060 13796 11112 13802
rect 11060 13738 11112 13744
rect 10876 13252 10928 13258
rect 10876 13194 10928 13200
rect 10888 12714 10916 13194
rect 10876 12708 10928 12714
rect 10876 12650 10928 12656
rect 10888 12238 10916 12650
rect 11072 12288 11100 13738
rect 11256 12968 11284 15030
rect 11336 14884 11388 14890
rect 11336 14826 11388 14832
rect 11348 14521 11376 14826
rect 11334 14512 11390 14521
rect 11334 14447 11390 14456
rect 11716 14385 11744 17002
rect 11808 15042 11836 17682
rect 11992 17338 12020 17818
rect 11980 17332 12032 17338
rect 11980 17274 12032 17280
rect 12084 16046 12112 18634
rect 12176 18222 12204 19858
rect 12452 19786 12480 22200
rect 12440 19780 12492 19786
rect 12440 19722 12492 19728
rect 12256 19712 12308 19718
rect 12256 19654 12308 19660
rect 12164 18216 12216 18222
rect 12164 18158 12216 18164
rect 12164 18080 12216 18086
rect 12164 18022 12216 18028
rect 12176 17678 12204 18022
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 12268 17542 12296 19654
rect 12820 19174 12848 22200
rect 13084 19916 13136 19922
rect 13084 19858 13136 19864
rect 13096 19378 13124 19858
rect 13084 19372 13136 19378
rect 13084 19314 13136 19320
rect 12992 19304 13044 19310
rect 12992 19246 13044 19252
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 13004 18766 13032 19246
rect 13188 19156 13216 22200
rect 13452 20324 13504 20330
rect 13452 20266 13504 20272
rect 13360 19304 13412 19310
rect 13360 19246 13412 19252
rect 13268 19168 13320 19174
rect 13188 19128 13268 19156
rect 13268 19110 13320 19116
rect 12992 18760 13044 18766
rect 12992 18702 13044 18708
rect 13372 18698 13400 19246
rect 13360 18692 13412 18698
rect 13360 18634 13412 18640
rect 12440 18284 12492 18290
rect 12440 18226 12492 18232
rect 12256 17536 12308 17542
rect 12256 17478 12308 17484
rect 12452 17134 12480 18226
rect 12808 18080 12860 18086
rect 12622 18048 12678 18057
rect 12808 18022 12860 18028
rect 12622 17983 12678 17992
rect 12440 17128 12492 17134
rect 12360 17088 12440 17116
rect 12256 16516 12308 16522
rect 12256 16458 12308 16464
rect 12072 16040 12124 16046
rect 12072 15982 12124 15988
rect 11978 15872 12034 15881
rect 11978 15807 12034 15816
rect 11992 15638 12020 15807
rect 12164 15700 12216 15706
rect 12268 15688 12296 16458
rect 12360 16114 12388 17088
rect 12440 17070 12492 17076
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 12348 16108 12400 16114
rect 12348 16050 12400 16056
rect 12348 15972 12400 15978
rect 12348 15914 12400 15920
rect 12216 15660 12296 15688
rect 12164 15642 12216 15648
rect 11980 15632 12032 15638
rect 11980 15574 12032 15580
rect 12072 15632 12124 15638
rect 12072 15574 12124 15580
rect 12162 15600 12218 15609
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 11900 15162 11928 15438
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 12084 15094 12112 15574
rect 12162 15535 12218 15544
rect 12072 15088 12124 15094
rect 11808 15014 11928 15042
rect 12072 15030 12124 15036
rect 12176 15026 12204 15535
rect 11796 14612 11848 14618
rect 11796 14554 11848 14560
rect 11702 14376 11758 14385
rect 11702 14311 11758 14320
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11352 14096 11648 14116
rect 11808 13870 11836 14554
rect 11796 13864 11848 13870
rect 11610 13832 11666 13841
rect 11796 13806 11848 13812
rect 11610 13767 11612 13776
rect 11664 13767 11666 13776
rect 11612 13738 11664 13744
rect 11808 13512 11836 13806
rect 11900 13802 11928 15014
rect 12164 15020 12216 15026
rect 12164 14962 12216 14968
rect 12072 14952 12124 14958
rect 12072 14894 12124 14900
rect 11980 14816 12032 14822
rect 11980 14758 12032 14764
rect 11888 13796 11940 13802
rect 11888 13738 11940 13744
rect 11624 13484 11836 13512
rect 11624 13394 11652 13484
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 11624 13297 11652 13330
rect 11610 13288 11666 13297
rect 11610 13223 11666 13232
rect 11352 13084 11648 13104
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 11256 12940 11376 12968
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 10980 12260 11100 12288
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10888 11558 10916 12174
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10874 11248 10930 11257
rect 10874 11183 10930 11192
rect 10888 10849 10916 11183
rect 10874 10840 10930 10849
rect 10980 10810 11008 12260
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 11060 11892 11112 11898
rect 11060 11834 11112 11840
rect 10874 10775 10930 10784
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 11072 10606 11100 11834
rect 11164 11626 11192 12174
rect 11256 11898 11284 12582
rect 11348 12084 11376 12940
rect 11428 12708 11480 12714
rect 11428 12650 11480 12656
rect 11440 12617 11468 12650
rect 11426 12608 11482 12617
rect 11426 12543 11482 12552
rect 11440 12442 11468 12543
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11716 12306 11744 13484
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11808 12986 11836 13330
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 11900 12442 11928 12582
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 11886 12336 11942 12345
rect 11428 12300 11480 12306
rect 11428 12242 11480 12248
rect 11704 12300 11756 12306
rect 11886 12271 11942 12280
rect 11704 12242 11756 12248
rect 11440 12209 11468 12242
rect 11900 12238 11928 12271
rect 11888 12232 11940 12238
rect 11426 12200 11482 12209
rect 11888 12174 11940 12180
rect 11426 12135 11482 12144
rect 11348 12056 11744 12084
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11244 11892 11296 11898
rect 11716 11880 11744 12056
rect 11244 11834 11296 11840
rect 11624 11852 11744 11880
rect 11428 11824 11480 11830
rect 11428 11766 11480 11772
rect 11152 11620 11204 11626
rect 11152 11562 11204 11568
rect 11164 11150 11192 11562
rect 11440 11558 11468 11766
rect 11428 11552 11480 11558
rect 11428 11494 11480 11500
rect 11624 11370 11652 11852
rect 11900 11744 11928 12174
rect 11992 11937 12020 14758
rect 12084 14249 12112 14894
rect 12070 14240 12126 14249
rect 12070 14175 12126 14184
rect 11978 11928 12034 11937
rect 11978 11863 12034 11872
rect 12084 11812 12112 14175
rect 12254 14104 12310 14113
rect 12254 14039 12310 14048
rect 12268 14006 12296 14039
rect 12256 14000 12308 14006
rect 12256 13942 12308 13948
rect 12256 13796 12308 13802
rect 12256 13738 12308 13744
rect 12162 11928 12218 11937
rect 12162 11863 12218 11872
rect 11808 11716 11928 11744
rect 11992 11784 12112 11812
rect 11808 11626 11836 11716
rect 11992 11694 12020 11784
rect 11980 11688 12032 11694
rect 11900 11648 11980 11676
rect 11796 11620 11848 11626
rect 11256 11342 11652 11370
rect 11716 11580 11796 11608
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 11164 10810 11192 11086
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 11150 10432 11206 10441
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10888 7546 10916 8910
rect 10980 8401 11008 9114
rect 11072 8673 11100 10406
rect 11150 10367 11206 10376
rect 11058 8664 11114 8673
rect 11058 8599 11114 8608
rect 10966 8392 11022 8401
rect 10966 8327 10968 8336
rect 11020 8327 11022 8336
rect 10968 8298 11020 8304
rect 10980 7886 11008 8298
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 10874 7440 10930 7449
rect 10874 7375 10930 7384
rect 10784 7268 10836 7274
rect 10784 7210 10836 7216
rect 10690 6760 10746 6769
rect 10600 6724 10652 6730
rect 10690 6695 10746 6704
rect 10600 6666 10652 6672
rect 10692 6452 10744 6458
rect 10888 6440 10916 7375
rect 10980 6730 11008 7822
rect 11072 7410 11100 7890
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 11164 7290 11192 10367
rect 11256 8945 11284 11342
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 11336 10600 11388 10606
rect 11336 10542 11388 10548
rect 11348 10266 11376 10542
rect 11518 10432 11574 10441
rect 11518 10367 11574 10376
rect 11532 10266 11560 10367
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 11716 10198 11744 11580
rect 11796 11562 11848 11568
rect 11796 10736 11848 10742
rect 11796 10678 11848 10684
rect 11704 10192 11756 10198
rect 11704 10134 11756 10140
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11336 9444 11388 9450
rect 11336 9386 11388 9392
rect 11704 9444 11756 9450
rect 11704 9386 11756 9392
rect 11348 9178 11376 9386
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11428 9036 11480 9042
rect 11428 8978 11480 8984
rect 11440 8945 11468 8978
rect 11242 8936 11298 8945
rect 11242 8871 11298 8880
rect 11426 8936 11482 8945
rect 11426 8871 11482 8880
rect 11256 8242 11284 8871
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 11256 8214 11376 8242
rect 11348 8090 11376 8214
rect 11244 8084 11296 8090
rect 11244 8026 11296 8032
rect 11336 8084 11388 8090
rect 11336 8026 11388 8032
rect 11256 7857 11284 8026
rect 11242 7848 11298 7857
rect 11242 7783 11298 7792
rect 11256 7342 11284 7783
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 11072 7262 11192 7290
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 11520 7268 11572 7274
rect 10968 6724 11020 6730
rect 10968 6666 11020 6672
rect 10744 6412 10916 6440
rect 10692 6394 10744 6400
rect 10704 5914 10732 6394
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10690 5808 10746 5817
rect 10690 5743 10746 5752
rect 10704 5574 10732 5743
rect 10796 5574 10824 6258
rect 10968 6112 11020 6118
rect 10888 6072 10968 6100
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10796 5370 10824 5510
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10796 5234 10824 5306
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 10520 5086 10732 5114
rect 10888 5098 10916 6072
rect 10968 6054 11020 6060
rect 10968 5636 11020 5642
rect 10968 5578 11020 5584
rect 10980 5234 11008 5578
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10508 5024 10560 5030
rect 10508 4966 10560 4972
rect 10600 5024 10652 5030
rect 10600 4966 10652 4972
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10324 4616 10376 4622
rect 10324 4558 10376 4564
rect 10428 4486 10456 4762
rect 10520 4758 10548 4966
rect 10508 4752 10560 4758
rect 10508 4694 10560 4700
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 10414 4312 10470 4321
rect 10414 4247 10470 4256
rect 10322 3904 10378 3913
rect 10322 3839 10378 3848
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 10244 3641 10272 3674
rect 10230 3632 10286 3641
rect 10230 3567 10286 3576
rect 10230 3088 10286 3097
rect 10230 3023 10286 3032
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 9956 2576 10008 2582
rect 9956 2518 10008 2524
rect 9968 2310 9996 2518
rect 10140 2508 10192 2514
rect 10140 2450 10192 2456
rect 10152 2310 10180 2450
rect 9956 2304 10008 2310
rect 9956 2246 10008 2252
rect 10140 2304 10192 2310
rect 10140 2246 10192 2252
rect 9968 1834 9996 2246
rect 9956 1828 10008 1834
rect 9956 1770 10008 1776
rect 10152 1494 10180 2246
rect 9784 1414 9904 1442
rect 10140 1488 10192 1494
rect 10140 1430 10192 1436
rect 9784 800 9812 1414
rect 10244 800 10272 3023
rect 10336 2961 10364 3839
rect 10428 3398 10456 4247
rect 10520 4214 10548 4694
rect 10508 4208 10560 4214
rect 10508 4150 10560 4156
rect 10612 4078 10640 4966
rect 10704 4690 10732 5086
rect 10876 5092 10928 5098
rect 10876 5034 10928 5040
rect 10692 4684 10744 4690
rect 10692 4626 10744 4632
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 10796 4486 10824 4558
rect 10692 4480 10744 4486
rect 10692 4422 10744 4428
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 10600 4072 10652 4078
rect 10600 4014 10652 4020
rect 10704 3924 10732 4422
rect 10612 3896 10732 3924
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 10322 2952 10378 2961
rect 10322 2887 10378 2896
rect 10428 2446 10456 3334
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 10612 800 10640 3896
rect 10692 3528 10744 3534
rect 10690 3496 10692 3505
rect 10744 3496 10746 3505
rect 10690 3431 10746 3440
rect 10796 2310 10824 4422
rect 10888 3369 10916 4626
rect 10966 4176 11022 4185
rect 10966 4111 11022 4120
rect 10980 3738 11008 4111
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10874 3360 10930 3369
rect 10874 3295 10930 3304
rect 10980 3126 11008 3538
rect 10968 3120 11020 3126
rect 10968 3062 11020 3068
rect 10784 2304 10836 2310
rect 10784 2246 10836 2252
rect 11072 800 11100 7262
rect 11520 7210 11572 7216
rect 11428 7200 11480 7206
rect 11256 7148 11428 7154
rect 11256 7142 11480 7148
rect 11256 7126 11468 7142
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 11164 4622 11192 6190
rect 11256 5574 11284 7126
rect 11532 7002 11560 7210
rect 11716 7002 11744 9386
rect 11520 6996 11572 7002
rect 11520 6938 11572 6944
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11352 6480 11648 6500
rect 11428 6384 11480 6390
rect 11428 6326 11480 6332
rect 11440 6089 11468 6326
rect 11716 6322 11744 6938
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11426 6080 11482 6089
rect 11426 6015 11482 6024
rect 11716 5710 11744 6258
rect 11704 5704 11756 5710
rect 11704 5646 11756 5652
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 11256 5030 11284 5510
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 11336 5296 11388 5302
rect 11336 5238 11388 5244
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 11348 4826 11376 5238
rect 11716 5137 11744 5306
rect 11808 5166 11836 10678
rect 11900 10470 11928 11648
rect 12176 11642 12204 11863
rect 11980 11630 12032 11636
rect 12084 11614 12204 11642
rect 12084 11121 12112 11614
rect 12268 11218 12296 13738
rect 12256 11212 12308 11218
rect 12256 11154 12308 11160
rect 12070 11112 12126 11121
rect 12126 11070 12204 11098
rect 12070 11047 12126 11056
rect 12084 10987 12112 11047
rect 12070 10840 12126 10849
rect 12070 10775 12126 10784
rect 11888 10464 11940 10470
rect 11888 10406 11940 10412
rect 11980 10464 12032 10470
rect 12084 10441 12112 10775
rect 11980 10406 12032 10412
rect 12070 10432 12126 10441
rect 11992 10266 12020 10406
rect 12070 10367 12126 10376
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 11886 10160 11942 10169
rect 11886 10095 11888 10104
rect 11940 10095 11942 10104
rect 11888 10066 11940 10072
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 11888 9920 11940 9926
rect 11888 9862 11940 9868
rect 11900 9761 11928 9862
rect 11886 9752 11942 9761
rect 11886 9687 11942 9696
rect 11992 9518 12020 9998
rect 12084 9926 12112 10202
rect 12176 10010 12204 11070
rect 12360 10266 12388 15914
rect 12452 15706 12480 16594
rect 12532 16040 12584 16046
rect 12532 15982 12584 15988
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12544 14958 12572 15982
rect 12636 15570 12664 17983
rect 12716 16584 12768 16590
rect 12716 16526 12768 16532
rect 12728 16046 12756 16526
rect 12820 16454 12848 18022
rect 13268 17740 13320 17746
rect 13268 17682 13320 17688
rect 13174 17640 13230 17649
rect 13174 17575 13230 17584
rect 12808 16448 12860 16454
rect 12860 16408 12940 16436
rect 12808 16390 12860 16396
rect 12716 16040 12768 16046
rect 12716 15982 12768 15988
rect 12728 15609 12756 15982
rect 12808 15972 12860 15978
rect 12808 15914 12860 15920
rect 12714 15600 12770 15609
rect 12624 15564 12676 15570
rect 12714 15535 12770 15544
rect 12624 15506 12676 15512
rect 12636 15337 12664 15506
rect 12716 15496 12768 15502
rect 12714 15464 12716 15473
rect 12820 15484 12848 15914
rect 12912 15502 12940 16408
rect 13188 15586 13216 17575
rect 13280 17542 13308 17682
rect 13268 17536 13320 17542
rect 13268 17478 13320 17484
rect 13360 17060 13412 17066
rect 13360 17002 13412 17008
rect 13268 16652 13320 16658
rect 13268 16594 13320 16600
rect 13280 15706 13308 16594
rect 13372 16590 13400 17002
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 13372 15910 13400 16526
rect 13360 15904 13412 15910
rect 13360 15846 13412 15852
rect 13268 15700 13320 15706
rect 13268 15642 13320 15648
rect 13188 15558 13308 15586
rect 12768 15464 12848 15484
rect 12770 15456 12848 15464
rect 12900 15496 12952 15502
rect 12900 15438 12952 15444
rect 12714 15399 12770 15408
rect 12622 15328 12678 15337
rect 12622 15263 12678 15272
rect 12532 14952 12584 14958
rect 12912 14906 12940 15438
rect 13176 14952 13228 14958
rect 12532 14894 12584 14900
rect 12440 14612 12492 14618
rect 12544 14600 12572 14894
rect 12820 14890 13124 14906
rect 13176 14894 13228 14900
rect 12808 14884 13124 14890
rect 12860 14878 13124 14884
rect 12808 14826 12860 14832
rect 12492 14572 12572 14600
rect 12440 14554 12492 14560
rect 12532 14476 12584 14482
rect 12452 14436 12532 14464
rect 12452 13734 12480 14436
rect 12532 14418 12584 14424
rect 13096 14414 13124 14878
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 12624 14340 12676 14346
rect 12624 14282 12676 14288
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12452 13433 12480 13670
rect 12438 13424 12494 13433
rect 12438 13359 12494 13368
rect 12452 12986 12480 13359
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12532 12640 12584 12646
rect 12438 12608 12494 12617
rect 12532 12582 12584 12588
rect 12438 12543 12494 12552
rect 12452 12442 12480 12543
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12544 12374 12572 12582
rect 12532 12368 12584 12374
rect 12532 12310 12584 12316
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12452 11762 12480 12038
rect 12544 11830 12572 12174
rect 12532 11824 12584 11830
rect 12532 11766 12584 11772
rect 12440 11756 12492 11762
rect 12440 11698 12492 11704
rect 12440 11620 12492 11626
rect 12440 11562 12492 11568
rect 12452 11218 12480 11562
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12452 10742 12480 11154
rect 12544 10810 12572 11290
rect 12636 11257 12664 14282
rect 12716 13252 12768 13258
rect 12716 13194 12768 13200
rect 12728 12594 12756 13194
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 12820 12866 12848 13126
rect 12820 12838 12940 12866
rect 12912 12646 12940 12838
rect 12900 12640 12952 12646
rect 12728 12566 12848 12594
rect 12900 12582 12952 12588
rect 12820 12374 12848 12566
rect 12808 12368 12860 12374
rect 12808 12310 12860 12316
rect 13004 11665 13032 14350
rect 13188 14074 13216 14894
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13280 13954 13308 15558
rect 13096 13926 13308 13954
rect 12990 11656 13046 11665
rect 12912 11614 12990 11642
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 12820 11354 12848 11494
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 12622 11248 12678 11257
rect 12622 11183 12678 11192
rect 12806 11248 12862 11257
rect 12806 11183 12862 11192
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12440 10736 12492 10742
rect 12440 10678 12492 10684
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12348 10124 12400 10130
rect 12452 10112 12480 10542
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12400 10084 12480 10112
rect 12348 10066 12400 10072
rect 12176 9982 12296 10010
rect 12072 9920 12124 9926
rect 12072 9862 12124 9868
rect 11980 9512 12032 9518
rect 11980 9454 12032 9460
rect 11886 9344 11942 9353
rect 11886 9279 11942 9288
rect 11900 9042 11928 9279
rect 11978 9208 12034 9217
rect 11978 9143 12034 9152
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11888 8560 11940 8566
rect 11886 8528 11888 8537
rect 11940 8528 11942 8537
rect 11886 8463 11942 8472
rect 11888 8356 11940 8362
rect 11888 8298 11940 8304
rect 11900 7177 11928 8298
rect 11992 8265 12020 9143
rect 11978 8256 12034 8265
rect 11978 8191 12034 8200
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 11886 7168 11942 7177
rect 11886 7103 11942 7112
rect 11992 6746 12020 8026
rect 12084 7546 12112 9862
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 12176 9518 12204 9658
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 12268 9194 12296 9982
rect 12346 9888 12402 9897
rect 12346 9823 12402 9832
rect 12360 9654 12388 9823
rect 12348 9648 12400 9654
rect 12348 9590 12400 9596
rect 12176 9166 12296 9194
rect 12176 7970 12204 9166
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 12268 8294 12296 8910
rect 12346 8528 12402 8537
rect 12452 8498 12480 10084
rect 12544 9722 12572 10406
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 12820 9625 12848 11183
rect 12530 9616 12586 9625
rect 12806 9616 12862 9625
rect 12530 9551 12586 9560
rect 12624 9580 12676 9586
rect 12544 9217 12572 9551
rect 12806 9551 12862 9560
rect 12624 9522 12676 9528
rect 12530 9208 12586 9217
rect 12530 9143 12586 9152
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12346 8463 12402 8472
rect 12440 8492 12492 8498
rect 12360 8430 12388 8463
rect 12440 8434 12492 8440
rect 12348 8424 12400 8430
rect 12452 8401 12480 8434
rect 12348 8366 12400 8372
rect 12438 8392 12494 8401
rect 12438 8327 12494 8336
rect 12256 8288 12308 8294
rect 12308 8248 12388 8276
rect 12256 8230 12308 8236
rect 12176 7942 12296 7970
rect 12072 7540 12124 7546
rect 12072 7482 12124 7488
rect 12084 7206 12112 7237
rect 12072 7200 12124 7206
rect 12070 7168 12072 7177
rect 12124 7168 12126 7177
rect 12070 7103 12126 7112
rect 11900 6718 12020 6746
rect 11796 5160 11848 5166
rect 11702 5128 11758 5137
rect 11796 5102 11848 5108
rect 11702 5063 11758 5072
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 11164 4078 11192 4422
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 11716 4214 11744 4966
rect 11808 4826 11836 5102
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 11704 4208 11756 4214
rect 11704 4150 11756 4156
rect 11152 4072 11204 4078
rect 11152 4014 11204 4020
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 11164 2650 11192 3674
rect 11256 3398 11284 3878
rect 11244 3392 11296 3398
rect 11244 3334 11296 3340
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 11808 2938 11836 4762
rect 11624 2910 11836 2938
rect 11624 2689 11652 2910
rect 11796 2848 11848 2854
rect 11702 2816 11758 2825
rect 11796 2790 11848 2796
rect 11702 2751 11758 2760
rect 11610 2680 11666 2689
rect 11152 2644 11204 2650
rect 11610 2615 11666 2624
rect 11152 2586 11204 2592
rect 11164 2553 11192 2586
rect 11150 2544 11206 2553
rect 11150 2479 11206 2488
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 11716 1442 11744 2751
rect 11808 2514 11836 2790
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 11440 1414 11744 1442
rect 11440 800 11468 1414
rect 11900 800 11928 6718
rect 11978 6488 12034 6497
rect 11978 6423 12034 6432
rect 11992 5914 12020 6423
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 11992 5370 12020 5850
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 11980 5228 12032 5234
rect 11980 5170 12032 5176
rect 11992 5001 12020 5170
rect 11978 4992 12034 5001
rect 11978 4927 12034 4936
rect 11992 4622 12020 4927
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 11978 4448 12034 4457
rect 11978 4383 12034 4392
rect 11992 4146 12020 4383
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 12084 4049 12112 7103
rect 12268 5658 12296 7942
rect 12360 7886 12388 8248
rect 12452 8090 12480 8327
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 12360 6866 12388 7686
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 12452 6118 12480 8026
rect 12544 6458 12572 8910
rect 12636 7954 12664 9522
rect 12912 9466 12940 11614
rect 12990 11591 13046 11600
rect 12990 11248 13046 11257
rect 12990 11183 13046 11192
rect 12820 9438 12940 9466
rect 12716 9376 12768 9382
rect 12714 9344 12716 9353
rect 12768 9344 12770 9353
rect 12714 9279 12770 9288
rect 12820 8974 12848 9438
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12912 9178 12940 9318
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12624 7948 12676 7954
rect 12624 7890 12676 7896
rect 12624 7404 12676 7410
rect 12624 7346 12676 7352
rect 12636 7274 12664 7346
rect 12624 7268 12676 7274
rect 12624 7210 12676 7216
rect 12622 6760 12678 6769
rect 12622 6695 12678 6704
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 12636 6186 12664 6695
rect 12728 6322 12756 8570
rect 12820 8430 12848 8774
rect 13004 8616 13032 11183
rect 13096 9217 13124 13926
rect 13176 13728 13228 13734
rect 13176 13670 13228 13676
rect 13266 13696 13322 13705
rect 13188 13530 13216 13670
rect 13266 13631 13322 13640
rect 13176 13524 13228 13530
rect 13176 13466 13228 13472
rect 13280 13433 13308 13631
rect 13266 13424 13322 13433
rect 13266 13359 13322 13368
rect 13280 11257 13308 13359
rect 13360 11688 13412 11694
rect 13360 11630 13412 11636
rect 13266 11248 13322 11257
rect 13266 11183 13322 11192
rect 13372 11150 13400 11630
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 13464 10996 13492 20266
rect 13556 19156 13584 22200
rect 14016 20058 14044 22200
rect 14004 20052 14056 20058
rect 14004 19994 14056 20000
rect 13728 19304 13780 19310
rect 13728 19246 13780 19252
rect 14188 19304 14240 19310
rect 14188 19246 14240 19252
rect 13636 19168 13688 19174
rect 13556 19128 13636 19156
rect 13636 19110 13688 19116
rect 13544 18964 13596 18970
rect 13544 18906 13596 18912
rect 13556 17882 13584 18906
rect 13636 18624 13688 18630
rect 13740 18612 13768 19246
rect 14200 18630 14228 19246
rect 14384 19174 14412 22200
rect 14556 19916 14608 19922
rect 14556 19858 14608 19864
rect 14464 19304 14516 19310
rect 14464 19246 14516 19252
rect 14372 19168 14424 19174
rect 14372 19110 14424 19116
rect 14476 18630 14504 19246
rect 13688 18584 13768 18612
rect 14188 18624 14240 18630
rect 13636 18566 13688 18572
rect 14188 18566 14240 18572
rect 14464 18624 14516 18630
rect 14464 18566 14516 18572
rect 13544 17876 13596 17882
rect 13544 17818 13596 17824
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13556 14618 13584 15642
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13542 14512 13598 14521
rect 13648 14498 13676 18566
rect 13912 18216 13964 18222
rect 13912 18158 13964 18164
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 13832 16028 13860 17070
rect 13924 16658 13952 18158
rect 14200 17746 14228 18566
rect 14188 17740 14240 17746
rect 14188 17682 14240 17688
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 13912 16040 13964 16046
rect 13832 16000 13912 16028
rect 13912 15982 13964 15988
rect 13820 15904 13872 15910
rect 13726 15872 13782 15881
rect 13820 15846 13872 15852
rect 13726 15807 13782 15816
rect 13740 15706 13768 15807
rect 13728 15700 13780 15706
rect 13728 15642 13780 15648
rect 13726 15600 13782 15609
rect 13726 15535 13782 15544
rect 13740 15502 13768 15535
rect 13728 15496 13780 15502
rect 13728 15438 13780 15444
rect 13740 15094 13768 15438
rect 13832 15434 13860 15846
rect 13820 15428 13872 15434
rect 13820 15370 13872 15376
rect 13728 15088 13780 15094
rect 13924 15042 13952 15982
rect 14004 15904 14056 15910
rect 14056 15864 14136 15892
rect 14004 15846 14056 15852
rect 14108 15706 14136 15864
rect 14096 15700 14148 15706
rect 14096 15642 14148 15648
rect 14004 15564 14056 15570
rect 14004 15506 14056 15512
rect 14016 15434 14044 15506
rect 14004 15428 14056 15434
rect 14004 15370 14056 15376
rect 14108 15314 14136 15642
rect 13728 15030 13780 15036
rect 13832 15014 13952 15042
rect 14016 15286 14136 15314
rect 13832 14498 13860 15014
rect 13598 14470 13676 14498
rect 13740 14482 13860 14498
rect 13728 14476 13860 14482
rect 13542 14447 13598 14456
rect 13556 11880 13584 14447
rect 13780 14470 13860 14476
rect 13728 14418 13780 14424
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13832 14074 13860 14214
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 14016 13954 14044 15286
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 13832 13926 14044 13954
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 13740 13462 13768 13670
rect 13728 13456 13780 13462
rect 13728 13398 13780 13404
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13648 12850 13676 13126
rect 13636 12844 13688 12850
rect 13636 12786 13688 12792
rect 13636 11892 13688 11898
rect 13556 11852 13636 11880
rect 13636 11834 13688 11840
rect 13544 11620 13596 11626
rect 13544 11562 13596 11568
rect 13556 11286 13584 11562
rect 13740 11393 13768 13126
rect 13832 12646 13860 13926
rect 14108 13870 14136 14758
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 13912 13796 13964 13802
rect 13912 13738 13964 13744
rect 13924 13297 13952 13738
rect 14096 13728 14148 13734
rect 14016 13688 14096 13716
rect 14016 13462 14044 13688
rect 14096 13670 14148 13676
rect 14004 13456 14056 13462
rect 14004 13398 14056 13404
rect 14096 13456 14148 13462
rect 14096 13398 14148 13404
rect 13910 13288 13966 13297
rect 13910 13223 13966 13232
rect 13912 12912 13964 12918
rect 13910 12880 13912 12889
rect 13964 12880 13966 12889
rect 14108 12866 14136 13398
rect 14200 13190 14228 17682
rect 14476 17082 14504 18566
rect 14568 18290 14596 19858
rect 14752 19174 14780 22200
rect 15120 20346 15148 22200
rect 15120 20318 15240 20346
rect 14817 20156 15113 20176
rect 14873 20154 14897 20156
rect 14953 20154 14977 20156
rect 15033 20154 15057 20156
rect 14895 20102 14897 20154
rect 14959 20102 14971 20154
rect 15033 20102 15035 20154
rect 14873 20100 14897 20102
rect 14953 20100 14977 20102
rect 15033 20100 15057 20102
rect 14817 20080 15113 20100
rect 15212 20040 15240 20318
rect 15120 20012 15240 20040
rect 15384 20052 15436 20058
rect 15120 19514 15148 20012
rect 15488 20040 15516 22200
rect 15856 20058 15884 22200
rect 15436 20012 15516 20040
rect 15844 20052 15896 20058
rect 15384 19994 15436 20000
rect 15844 19994 15896 20000
rect 15200 19916 15252 19922
rect 15200 19858 15252 19864
rect 16120 19916 16172 19922
rect 16120 19858 16172 19864
rect 15108 19508 15160 19514
rect 15108 19450 15160 19456
rect 14740 19168 14792 19174
rect 14740 19110 14792 19116
rect 14817 19068 15113 19088
rect 14873 19066 14897 19068
rect 14953 19066 14977 19068
rect 15033 19066 15057 19068
rect 14895 19014 14897 19066
rect 14959 19014 14971 19066
rect 15033 19014 15035 19066
rect 14873 19012 14897 19014
rect 14953 19012 14977 19014
rect 15033 19012 15057 19014
rect 14817 18992 15113 19012
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14817 17980 15113 18000
rect 14873 17978 14897 17980
rect 14953 17978 14977 17980
rect 15033 17978 15057 17980
rect 14895 17926 14897 17978
rect 14959 17926 14971 17978
rect 15033 17926 15035 17978
rect 14873 17924 14897 17926
rect 14953 17924 14977 17926
rect 15033 17924 15057 17926
rect 14817 17904 15113 17924
rect 14280 17060 14332 17066
rect 14476 17054 14596 17082
rect 14280 17002 14332 17008
rect 14292 16590 14320 17002
rect 14464 16992 14516 16998
rect 14464 16934 14516 16940
rect 14476 16658 14504 16934
rect 14464 16652 14516 16658
rect 14464 16594 14516 16600
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14280 15564 14332 15570
rect 14280 15506 14332 15512
rect 14292 15026 14320 15506
rect 14280 15020 14332 15026
rect 14280 14962 14332 14968
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 14292 13462 14320 14554
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14280 13456 14332 13462
rect 14280 13398 14332 13404
rect 14384 13308 14412 14214
rect 14292 13280 14412 13308
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 14016 12850 14136 12866
rect 13910 12815 13966 12824
rect 14004 12844 14136 12850
rect 14056 12838 14136 12844
rect 14004 12786 14056 12792
rect 14096 12776 14148 12782
rect 14292 12730 14320 13280
rect 14370 12880 14426 12889
rect 14370 12815 14426 12824
rect 14096 12718 14148 12724
rect 13912 12708 13964 12714
rect 13912 12650 13964 12656
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 13924 12306 13952 12650
rect 14004 12640 14056 12646
rect 14004 12582 14056 12588
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 13924 11626 13952 12038
rect 13912 11620 13964 11626
rect 13912 11562 13964 11568
rect 13726 11384 13782 11393
rect 13726 11319 13782 11328
rect 13544 11280 13596 11286
rect 13544 11222 13596 11228
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 13832 11121 13860 11154
rect 13818 11112 13874 11121
rect 13818 11047 13874 11056
rect 13372 10968 13492 10996
rect 13176 10804 13228 10810
rect 13176 10746 13228 10752
rect 13188 10112 13216 10746
rect 13268 10124 13320 10130
rect 13188 10084 13268 10112
rect 13188 9586 13216 10084
rect 13268 10066 13320 10072
rect 13372 10010 13400 10968
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13556 10554 13584 10610
rect 13464 10538 13584 10554
rect 13452 10532 13584 10538
rect 13504 10526 13584 10532
rect 13452 10474 13504 10480
rect 13280 9982 13400 10010
rect 13176 9580 13228 9586
rect 13176 9522 13228 9528
rect 13174 9344 13230 9353
rect 13174 9279 13230 9288
rect 13082 9208 13138 9217
rect 13082 9143 13138 9152
rect 13084 9104 13136 9110
rect 13084 9046 13136 9052
rect 13096 8673 13124 9046
rect 12912 8588 13032 8616
rect 13082 8664 13138 8673
rect 13082 8599 13138 8608
rect 12808 8424 12860 8430
rect 12808 8366 12860 8372
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12820 8090 12848 8230
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 12912 7970 12940 8588
rect 13188 8537 13216 9279
rect 13280 8634 13308 9982
rect 13358 9888 13414 9897
rect 13358 9823 13414 9832
rect 13372 9722 13400 9823
rect 13360 9716 13412 9722
rect 13360 9658 13412 9664
rect 13358 9480 13414 9489
rect 13358 9415 13414 9424
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13174 8528 13230 8537
rect 13084 8492 13136 8498
rect 12820 7942 12940 7970
rect 13004 8452 13084 8480
rect 12820 7206 12848 7942
rect 13004 7750 13032 8452
rect 13174 8463 13230 8472
rect 13268 8492 13320 8498
rect 13084 8434 13136 8440
rect 13082 8392 13138 8401
rect 13082 8327 13138 8336
rect 12992 7744 13044 7750
rect 12898 7712 12954 7721
rect 12992 7686 13044 7692
rect 12898 7647 12954 7656
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12912 7002 12940 7647
rect 13004 7478 13032 7686
rect 13096 7546 13124 8327
rect 13084 7540 13136 7546
rect 13084 7482 13136 7488
rect 12992 7472 13044 7478
rect 12992 7414 13044 7420
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 12992 6656 13044 6662
rect 12992 6598 13044 6604
rect 13004 6322 13032 6598
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 12992 6316 13044 6322
rect 12992 6258 13044 6264
rect 12624 6180 12676 6186
rect 12624 6122 12676 6128
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12898 6080 12954 6089
rect 12452 5778 12480 6054
rect 12898 6015 12954 6024
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12624 5772 12676 5778
rect 12624 5714 12676 5720
rect 12176 5630 12296 5658
rect 12070 4040 12126 4049
rect 12070 3975 12126 3984
rect 12176 2825 12204 5630
rect 12254 5536 12310 5545
rect 12254 5471 12310 5480
rect 12268 5302 12296 5471
rect 12256 5296 12308 5302
rect 12256 5238 12308 5244
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12256 5092 12308 5098
rect 12256 5034 12308 5040
rect 12268 4826 12296 5034
rect 12452 4826 12480 5102
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12256 4820 12308 4826
rect 12256 4762 12308 4768
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12348 4752 12400 4758
rect 12348 4694 12400 4700
rect 12360 4298 12388 4694
rect 12268 4282 12388 4298
rect 12256 4276 12388 4282
rect 12308 4270 12388 4276
rect 12256 4218 12308 4224
rect 12544 4214 12572 4966
rect 12636 4622 12664 5714
rect 12912 5386 12940 6015
rect 13004 5846 13032 6258
rect 12992 5840 13044 5846
rect 12992 5782 13044 5788
rect 12716 5364 12768 5370
rect 12912 5358 13032 5386
rect 12716 5306 12768 5312
rect 12728 5098 12756 5306
rect 12900 5296 12952 5302
rect 12898 5264 12900 5273
rect 12952 5264 12954 5273
rect 12898 5199 12954 5208
rect 12716 5092 12768 5098
rect 12716 5034 12768 5040
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 12348 4208 12400 4214
rect 12348 4150 12400 4156
rect 12532 4208 12584 4214
rect 12532 4150 12584 4156
rect 12360 3602 12388 4150
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12452 3777 12480 3878
rect 12438 3768 12494 3777
rect 12438 3703 12494 3712
rect 12636 3670 12664 4558
rect 12912 4214 12940 5199
rect 13004 4486 13032 5358
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 13096 5001 13124 5170
rect 13188 5166 13216 8463
rect 13268 8434 13320 8440
rect 13280 7993 13308 8434
rect 13266 7984 13322 7993
rect 13266 7919 13322 7928
rect 13266 7712 13322 7721
rect 13266 7647 13322 7656
rect 13280 7313 13308 7647
rect 13372 7449 13400 9415
rect 13464 8974 13492 10474
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13556 9586 13584 9998
rect 13648 9994 13676 10406
rect 13832 10266 13860 11047
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13636 9988 13688 9994
rect 13636 9930 13688 9936
rect 13648 9710 13860 9738
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 13358 7440 13414 7449
rect 13358 7375 13414 7384
rect 13266 7304 13322 7313
rect 13266 7239 13322 7248
rect 13372 6798 13400 7375
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13372 6458 13400 6734
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13176 5160 13228 5166
rect 13176 5102 13228 5108
rect 13360 5024 13412 5030
rect 13082 4992 13138 5001
rect 13360 4966 13412 4972
rect 13082 4927 13138 4936
rect 13096 4758 13124 4927
rect 13084 4752 13136 4758
rect 13084 4694 13136 4700
rect 12992 4480 13044 4486
rect 12992 4422 13044 4428
rect 12716 4208 12768 4214
rect 12716 4150 12768 4156
rect 12900 4208 12952 4214
rect 12900 4150 12952 4156
rect 12728 3754 12756 4150
rect 13004 4026 13032 4422
rect 13268 4208 13320 4214
rect 13268 4150 13320 4156
rect 12808 4004 12860 4010
rect 12808 3946 12860 3952
rect 12912 3998 13032 4026
rect 12820 3913 12848 3946
rect 12912 3942 12940 3998
rect 12900 3936 12952 3942
rect 12806 3904 12862 3913
rect 12900 3878 12952 3884
rect 13084 3936 13136 3942
rect 13084 3878 13136 3884
rect 12806 3839 12862 3848
rect 12728 3738 13032 3754
rect 12728 3732 13044 3738
rect 12728 3726 12992 3732
rect 12992 3674 13044 3680
rect 12440 3664 12492 3670
rect 12440 3606 12492 3612
rect 12624 3664 12676 3670
rect 12624 3606 12676 3612
rect 12716 3664 12768 3670
rect 12716 3606 12768 3612
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12254 3360 12310 3369
rect 12254 3295 12310 3304
rect 12162 2816 12218 2825
rect 12162 2751 12218 2760
rect 12268 2038 12296 3295
rect 12348 3188 12400 3194
rect 12348 3130 12400 3136
rect 12360 2990 12388 3130
rect 12452 3126 12480 3606
rect 12440 3120 12492 3126
rect 12440 3062 12492 3068
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 12728 2922 12756 3606
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 12532 2916 12584 2922
rect 12532 2858 12584 2864
rect 12716 2916 12768 2922
rect 12716 2858 12768 2864
rect 12900 2916 12952 2922
rect 12900 2858 12952 2864
rect 12544 2650 12572 2858
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 12728 2446 12756 2858
rect 12912 2514 12940 2858
rect 13004 2650 13032 3334
rect 13096 2854 13124 3878
rect 13280 3584 13308 4150
rect 13372 4078 13400 4966
rect 13360 4072 13412 4078
rect 13360 4014 13412 4020
rect 13360 3596 13412 3602
rect 13280 3556 13360 3584
rect 13360 3538 13412 3544
rect 13464 3126 13492 8774
rect 13556 7954 13584 9522
rect 13648 9518 13676 9710
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13648 9042 13676 9318
rect 13740 9110 13768 9590
rect 13832 9466 13860 9710
rect 13924 9586 13952 11562
rect 14016 11286 14044 12582
rect 14108 11354 14136 12718
rect 14200 12702 14320 12730
rect 14200 12374 14228 12702
rect 14188 12368 14240 12374
rect 14188 12310 14240 12316
rect 14280 12300 14332 12306
rect 14280 12242 14332 12248
rect 14188 11552 14240 11558
rect 14188 11494 14240 11500
rect 14096 11348 14148 11354
rect 14096 11290 14148 11296
rect 14004 11280 14056 11286
rect 14004 11222 14056 11228
rect 14004 10464 14056 10470
rect 14004 10406 14056 10412
rect 13912 9580 13964 9586
rect 13912 9522 13964 9528
rect 14016 9466 14044 10406
rect 14108 9518 14136 11290
rect 14200 11150 14228 11494
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 14200 10674 14228 11086
rect 14188 10668 14240 10674
rect 14188 10610 14240 10616
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 14200 10266 14228 10406
rect 14188 10260 14240 10266
rect 14188 10202 14240 10208
rect 14188 10124 14240 10130
rect 14188 10066 14240 10072
rect 13832 9438 14044 9466
rect 14096 9512 14148 9518
rect 14096 9454 14148 9460
rect 14200 9110 14228 10066
rect 13728 9104 13780 9110
rect 14188 9104 14240 9110
rect 13728 9046 13780 9052
rect 13818 9072 13874 9081
rect 13636 9036 13688 9042
rect 13818 9007 13874 9016
rect 14186 9072 14188 9081
rect 14240 9072 14242 9081
rect 14186 9007 14242 9016
rect 13636 8978 13688 8984
rect 13544 7948 13596 7954
rect 13544 7890 13596 7896
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13648 7410 13676 7822
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13740 7410 13768 7482
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 13648 6798 13676 7346
rect 13726 7304 13782 7313
rect 13726 7239 13782 7248
rect 13740 7206 13768 7239
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 13726 6896 13782 6905
rect 13726 6831 13782 6840
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13544 6384 13596 6390
rect 13544 6326 13596 6332
rect 13452 3120 13504 3126
rect 13452 3062 13504 3068
rect 13556 3058 13584 6326
rect 13648 6118 13676 6598
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 13084 2848 13136 2854
rect 13084 2790 13136 2796
rect 12992 2644 13044 2650
rect 12992 2586 13044 2592
rect 13648 2553 13676 6054
rect 13740 5778 13768 6831
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 13740 5273 13768 5714
rect 13726 5264 13782 5273
rect 13726 5199 13782 5208
rect 13740 5166 13768 5199
rect 13728 5160 13780 5166
rect 13728 5102 13780 5108
rect 13832 5080 13860 9007
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13924 7954 13952 8230
rect 14002 7984 14058 7993
rect 13912 7948 13964 7954
rect 14200 7954 14228 8910
rect 14002 7919 14058 7928
rect 14188 7948 14240 7954
rect 13912 7890 13964 7896
rect 13924 7750 13952 7890
rect 14016 7886 14044 7919
rect 14188 7890 14240 7896
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 14016 6866 14044 7822
rect 14108 7410 14136 7822
rect 14200 7732 14228 7890
rect 14292 7857 14320 12242
rect 14278 7848 14334 7857
rect 14278 7783 14334 7792
rect 14200 7704 14320 7732
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 14016 6662 14044 6802
rect 14004 6656 14056 6662
rect 14004 6598 14056 6604
rect 14108 6458 14136 7142
rect 14188 6656 14240 6662
rect 14188 6598 14240 6604
rect 14200 6458 14228 6598
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 14004 6180 14056 6186
rect 14004 6122 14056 6128
rect 13912 6112 13964 6118
rect 13912 6054 13964 6060
rect 13924 5681 13952 6054
rect 13910 5672 13966 5681
rect 13910 5607 13966 5616
rect 13912 5568 13964 5574
rect 13912 5510 13964 5516
rect 13924 5234 13952 5510
rect 13912 5228 13964 5234
rect 13912 5170 13964 5176
rect 13912 5092 13964 5098
rect 13832 5052 13912 5080
rect 13912 5034 13964 5040
rect 14016 5030 14044 6122
rect 13728 5024 13780 5030
rect 13728 4966 13780 4972
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 13740 4570 13768 4966
rect 14016 4690 14044 4966
rect 14096 4752 14148 4758
rect 14094 4720 14096 4729
rect 14148 4720 14150 4729
rect 14004 4684 14056 4690
rect 14094 4655 14150 4664
rect 14004 4626 14056 4632
rect 13740 4554 13952 4570
rect 13740 4548 13964 4554
rect 13740 4542 13912 4548
rect 13912 4490 13964 4496
rect 13728 4480 13780 4486
rect 13728 4422 13780 4428
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 13740 2854 13768 4422
rect 13832 4214 13860 4422
rect 13820 4208 13872 4214
rect 13820 4150 13872 4156
rect 14094 4176 14150 4185
rect 13832 3534 13860 4150
rect 14094 4111 14150 4120
rect 14108 3738 14136 4111
rect 14200 4078 14228 4422
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 14188 3936 14240 3942
rect 14188 3878 14240 3884
rect 14200 3777 14228 3878
rect 14186 3768 14242 3777
rect 14096 3732 14148 3738
rect 14186 3703 14242 3712
rect 14096 3674 14148 3680
rect 14188 3596 14240 3602
rect 14188 3538 14240 3544
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 13912 3392 13964 3398
rect 13912 3334 13964 3340
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 13634 2544 13690 2553
rect 12900 2508 12952 2514
rect 13634 2479 13690 2488
rect 13820 2508 13872 2514
rect 12900 2450 12952 2456
rect 13820 2450 13872 2456
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 12716 2440 12768 2446
rect 13832 2417 13860 2450
rect 13924 2446 13952 3334
rect 14200 3058 14228 3538
rect 14292 3369 14320 7704
rect 14278 3360 14334 3369
rect 14278 3295 14334 3304
rect 14188 3052 14240 3058
rect 14188 2994 14240 3000
rect 14384 2990 14412 12815
rect 14476 10452 14504 16594
rect 14568 13530 14596 17054
rect 14817 16892 15113 16912
rect 14873 16890 14897 16892
rect 14953 16890 14977 16892
rect 15033 16890 15057 16892
rect 14895 16838 14897 16890
rect 14959 16838 14971 16890
rect 15033 16838 15035 16890
rect 14873 16836 14897 16838
rect 14953 16836 14977 16838
rect 15033 16836 15057 16838
rect 14817 16816 15113 16836
rect 14817 15804 15113 15824
rect 14873 15802 14897 15804
rect 14953 15802 14977 15804
rect 15033 15802 15057 15804
rect 14895 15750 14897 15802
rect 14959 15750 14971 15802
rect 15033 15750 15035 15802
rect 14873 15748 14897 15750
rect 14953 15748 14977 15750
rect 15033 15748 15057 15750
rect 14817 15728 15113 15748
rect 14817 14716 15113 14736
rect 14873 14714 14897 14716
rect 14953 14714 14977 14716
rect 15033 14714 15057 14716
rect 14895 14662 14897 14714
rect 14959 14662 14971 14714
rect 15033 14662 15035 14714
rect 14873 14660 14897 14662
rect 14953 14660 14977 14662
rect 15033 14660 15057 14662
rect 14817 14640 15113 14660
rect 14740 14000 14792 14006
rect 14740 13942 14792 13948
rect 14646 13560 14702 13569
rect 14556 13524 14608 13530
rect 14646 13495 14702 13504
rect 14556 13466 14608 13472
rect 14568 12918 14596 13466
rect 14660 13394 14688 13495
rect 14752 13444 14780 13942
rect 14817 13628 15113 13648
rect 14873 13626 14897 13628
rect 14953 13626 14977 13628
rect 15033 13626 15057 13628
rect 14895 13574 14897 13626
rect 14959 13574 14971 13626
rect 15033 13574 15035 13626
rect 14873 13572 14897 13574
rect 14953 13572 14977 13574
rect 15033 13572 15057 13574
rect 14817 13552 15113 13572
rect 14832 13456 14884 13462
rect 14752 13416 14832 13444
rect 14832 13398 14884 13404
rect 15106 13424 15162 13433
rect 14648 13388 14700 13394
rect 15106 13359 15108 13368
rect 14648 13330 14700 13336
rect 15160 13359 15162 13368
rect 15108 13330 15160 13336
rect 14660 12986 14688 13330
rect 14832 13320 14884 13326
rect 14924 13320 14976 13326
rect 14832 13262 14884 13268
rect 14922 13288 14924 13297
rect 14976 13288 14978 13297
rect 14844 12986 14872 13262
rect 14922 13223 14978 13232
rect 14648 12980 14700 12986
rect 14648 12922 14700 12928
rect 14832 12980 14884 12986
rect 14832 12922 14884 12928
rect 14556 12912 14608 12918
rect 14556 12854 14608 12860
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14568 11529 14596 12718
rect 14817 12540 15113 12560
rect 14873 12538 14897 12540
rect 14953 12538 14977 12540
rect 15033 12538 15057 12540
rect 14895 12486 14897 12538
rect 14959 12486 14971 12538
rect 15033 12486 15035 12538
rect 14873 12484 14897 12486
rect 14953 12484 14977 12486
rect 15033 12484 15057 12486
rect 14817 12464 15113 12484
rect 15212 12322 15240 19858
rect 15568 19304 15620 19310
rect 15568 19246 15620 19252
rect 16028 19304 16080 19310
rect 16028 19246 16080 19252
rect 15292 19168 15344 19174
rect 15292 19110 15344 19116
rect 15304 17814 15332 19110
rect 15580 18970 15608 19246
rect 15844 19236 15896 19242
rect 15844 19178 15896 19184
rect 15568 18964 15620 18970
rect 15568 18906 15620 18912
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 15292 17808 15344 17814
rect 15292 17750 15344 17756
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 15384 17672 15436 17678
rect 15384 17614 15436 17620
rect 15304 17270 15332 17614
rect 15396 17338 15424 17614
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 15292 17264 15344 17270
rect 15580 17241 15608 18566
rect 15856 18193 15884 19178
rect 16040 18630 16068 19246
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 15842 18184 15898 18193
rect 15842 18119 15898 18128
rect 15752 17808 15804 17814
rect 15752 17750 15804 17756
rect 15660 17740 15712 17746
rect 15660 17682 15712 17688
rect 15292 17206 15344 17212
rect 15566 17232 15622 17241
rect 15304 16046 15332 17206
rect 15566 17167 15622 17176
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 15580 16250 15608 16594
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15568 16244 15620 16250
rect 15568 16186 15620 16192
rect 15292 16040 15344 16046
rect 15292 15982 15344 15988
rect 15304 15434 15332 15982
rect 15488 15609 15516 16186
rect 15672 15706 15700 17682
rect 15764 17134 15792 17750
rect 15936 17672 15988 17678
rect 15936 17614 15988 17620
rect 15752 17128 15804 17134
rect 15752 17070 15804 17076
rect 15660 15700 15712 15706
rect 15660 15642 15712 15648
rect 15474 15600 15530 15609
rect 15764 15586 15792 17070
rect 15948 16658 15976 17614
rect 15936 16652 15988 16658
rect 15936 16594 15988 16600
rect 16132 16538 16160 19858
rect 16316 19174 16344 22200
rect 16684 19174 16712 22200
rect 16304 19168 16356 19174
rect 16304 19110 16356 19116
rect 16672 19168 16724 19174
rect 16672 19110 16724 19116
rect 16948 19168 17000 19174
rect 16948 19110 17000 19116
rect 16488 18216 16540 18222
rect 16488 18158 16540 18164
rect 16500 17814 16528 18158
rect 16488 17808 16540 17814
rect 16488 17750 16540 17756
rect 16212 17740 16264 17746
rect 16212 17682 16264 17688
rect 16224 17338 16252 17682
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 16592 17134 16620 17478
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16580 17128 16632 17134
rect 16580 17070 16632 17076
rect 15474 15535 15476 15544
rect 15528 15535 15530 15544
rect 15580 15558 15792 15586
rect 15856 16510 16160 16538
rect 16684 16522 16712 17138
rect 16764 16992 16816 16998
rect 16764 16934 16816 16940
rect 16776 16794 16804 16934
rect 16764 16788 16816 16794
rect 16764 16730 16816 16736
rect 16672 16516 16724 16522
rect 15476 15506 15528 15512
rect 15292 15428 15344 15434
rect 15292 15370 15344 15376
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 15304 14074 15332 14758
rect 15396 14550 15424 14962
rect 15384 14544 15436 14550
rect 15384 14486 15436 14492
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 15396 14006 15424 14486
rect 15384 14000 15436 14006
rect 15384 13942 15436 13948
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 15304 13326 15332 13874
rect 15488 13870 15516 15506
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 15384 13728 15436 13734
rect 15384 13670 15436 13676
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15396 12986 15424 13670
rect 15488 13530 15516 13670
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 15476 12708 15528 12714
rect 15476 12650 15528 12656
rect 15212 12294 15424 12322
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 14648 12164 14700 12170
rect 14648 12106 14700 12112
rect 14554 11520 14610 11529
rect 14554 11455 14610 11464
rect 14568 10588 14596 11455
rect 14660 11286 14688 12106
rect 14648 11280 14700 11286
rect 14648 11222 14700 11228
rect 14660 10742 14688 11222
rect 14752 11218 14780 12174
rect 14832 12096 14884 12102
rect 14832 12038 14884 12044
rect 14844 11762 14872 12038
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 15212 11558 15240 11834
rect 15304 11694 15332 12174
rect 15292 11688 15344 11694
rect 15292 11630 15344 11636
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 14817 11452 15113 11472
rect 14873 11450 14897 11452
rect 14953 11450 14977 11452
rect 15033 11450 15057 11452
rect 14895 11398 14897 11450
rect 14959 11398 14971 11450
rect 15033 11398 15035 11450
rect 14873 11396 14897 11398
rect 14953 11396 14977 11398
rect 15033 11396 15057 11398
rect 14817 11376 15113 11396
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 15120 11082 15148 11154
rect 15108 11076 15160 11082
rect 15108 11018 15160 11024
rect 14648 10736 14700 10742
rect 14648 10678 14700 10684
rect 15212 10606 15240 11494
rect 15292 11076 15344 11082
rect 15292 11018 15344 11024
rect 15304 10849 15332 11018
rect 15290 10840 15346 10849
rect 15290 10775 15346 10784
rect 15200 10600 15252 10606
rect 14568 10560 14688 10588
rect 14476 10424 14596 10452
rect 14568 10112 14596 10424
rect 14660 10266 14688 10560
rect 15200 10542 15252 10548
rect 15292 10532 15344 10538
rect 15292 10474 15344 10480
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14648 10260 14700 10266
rect 14648 10202 14700 10208
rect 14476 10084 14596 10112
rect 14476 7313 14504 10084
rect 14554 10024 14610 10033
rect 14554 9959 14610 9968
rect 14568 9110 14596 9959
rect 14556 9104 14608 9110
rect 14556 9046 14608 9052
rect 14660 8838 14688 10202
rect 14752 9654 14780 10406
rect 14817 10364 15113 10384
rect 14873 10362 14897 10364
rect 14953 10362 14977 10364
rect 15033 10362 15057 10364
rect 14895 10310 14897 10362
rect 14959 10310 14971 10362
rect 15033 10310 15035 10362
rect 14873 10308 14897 10310
rect 14953 10308 14977 10310
rect 15033 10308 15057 10310
rect 14817 10288 15113 10308
rect 15304 10266 15332 10474
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 14832 9988 14884 9994
rect 14832 9930 14884 9936
rect 15016 9988 15068 9994
rect 15016 9930 15068 9936
rect 14844 9897 14872 9930
rect 14830 9888 14886 9897
rect 14830 9823 14886 9832
rect 14740 9648 14792 9654
rect 14740 9590 14792 9596
rect 15028 9586 15056 9930
rect 15396 9874 15424 12294
rect 15488 11762 15516 12650
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15474 10160 15530 10169
rect 15474 10095 15476 10104
rect 15528 10095 15530 10104
rect 15476 10066 15528 10072
rect 15476 9988 15528 9994
rect 15476 9930 15528 9936
rect 15304 9846 15424 9874
rect 15198 9616 15254 9625
rect 15016 9580 15068 9586
rect 15198 9551 15200 9560
rect 15016 9522 15068 9528
rect 15252 9551 15254 9560
rect 15200 9522 15252 9528
rect 14817 9276 15113 9296
rect 14873 9274 14897 9276
rect 14953 9274 14977 9276
rect 15033 9274 15057 9276
rect 14895 9222 14897 9274
rect 14959 9222 14971 9274
rect 15033 9222 15035 9274
rect 14873 9220 14897 9222
rect 14953 9220 14977 9222
rect 15033 9220 15057 9222
rect 14817 9200 15113 9220
rect 14740 9172 14792 9178
rect 15200 9172 15252 9178
rect 14792 9132 14964 9160
rect 14740 9114 14792 9120
rect 14832 8900 14884 8906
rect 14832 8842 14884 8848
rect 14648 8832 14700 8838
rect 14844 8809 14872 8842
rect 14648 8774 14700 8780
rect 14830 8800 14886 8809
rect 14830 8735 14886 8744
rect 14936 8537 14964 9132
rect 15200 9114 15252 9120
rect 14922 8528 14978 8537
rect 15212 8498 15240 9114
rect 14922 8463 14978 8472
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 14646 8392 14702 8401
rect 14646 8327 14648 8336
rect 14700 8327 14702 8336
rect 14648 8298 14700 8304
rect 14554 8256 14610 8265
rect 14554 8191 14610 8200
rect 14568 8022 14596 8191
rect 14660 8090 14688 8298
rect 14740 8288 14792 8294
rect 14740 8230 14792 8236
rect 14648 8084 14700 8090
rect 14648 8026 14700 8032
rect 14556 8016 14608 8022
rect 14556 7958 14608 7964
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14462 7304 14518 7313
rect 14462 7239 14518 7248
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 14476 6730 14504 7142
rect 14568 7002 14596 7686
rect 14660 7546 14688 8026
rect 14752 7886 14780 8230
rect 14817 8188 15113 8208
rect 14873 8186 14897 8188
rect 14953 8186 14977 8188
rect 15033 8186 15057 8188
rect 14895 8134 14897 8186
rect 14959 8134 14971 8186
rect 15033 8134 15035 8186
rect 14873 8132 14897 8134
rect 14953 8132 14977 8134
rect 15033 8132 15057 8134
rect 14817 8112 15113 8132
rect 15200 8016 15252 8022
rect 15200 7958 15252 7964
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14648 7540 14700 7546
rect 14648 7482 14700 7488
rect 14648 7200 14700 7206
rect 14648 7142 14700 7148
rect 14556 6996 14608 7002
rect 14556 6938 14608 6944
rect 14464 6724 14516 6730
rect 14464 6666 14516 6672
rect 14568 6168 14596 6938
rect 14476 6140 14596 6168
rect 14476 5250 14504 6140
rect 14660 5914 14688 7142
rect 14817 7100 15113 7120
rect 14873 7098 14897 7100
rect 14953 7098 14977 7100
rect 15033 7098 15057 7100
rect 14895 7046 14897 7098
rect 14959 7046 14971 7098
rect 15033 7046 15035 7098
rect 14873 7044 14897 7046
rect 14953 7044 14977 7046
rect 15033 7044 15057 7046
rect 14817 7024 15113 7044
rect 15212 7002 15240 7958
rect 15200 6996 15252 7002
rect 15200 6938 15252 6944
rect 14832 6792 14884 6798
rect 14832 6734 14884 6740
rect 14844 6254 14872 6734
rect 15304 6610 15332 9846
rect 15382 9752 15438 9761
rect 15382 9687 15438 9696
rect 15212 6582 15332 6610
rect 14832 6248 14884 6254
rect 14752 6208 14832 6236
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 14556 5636 14608 5642
rect 14556 5578 14608 5584
rect 14568 5370 14596 5578
rect 14646 5536 14702 5545
rect 14646 5471 14702 5480
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14476 5222 14596 5250
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 14476 3670 14504 4082
rect 14568 4078 14596 5222
rect 14660 4758 14688 5471
rect 14752 5352 14780 6208
rect 14832 6190 14884 6196
rect 15212 6118 15240 6582
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 14817 6012 15113 6032
rect 14873 6010 14897 6012
rect 14953 6010 14977 6012
rect 15033 6010 15057 6012
rect 14895 5958 14897 6010
rect 14959 5958 14971 6010
rect 15033 5958 15035 6010
rect 14873 5956 14897 5958
rect 14953 5956 14977 5958
rect 15033 5956 15057 5958
rect 14817 5936 15113 5956
rect 15108 5568 15160 5574
rect 15106 5536 15108 5545
rect 15160 5536 15162 5545
rect 15106 5471 15162 5480
rect 14752 5324 14872 5352
rect 14844 5234 14872 5324
rect 15212 5250 15240 6054
rect 15304 5710 15332 6394
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 14832 5228 14884 5234
rect 14832 5170 14884 5176
rect 15120 5222 15240 5250
rect 14648 4752 14700 4758
rect 14648 4694 14700 4700
rect 14556 4072 14608 4078
rect 14556 4014 14608 4020
rect 14568 3913 14596 4014
rect 14554 3904 14610 3913
rect 14554 3839 14610 3848
rect 14464 3664 14516 3670
rect 14464 3606 14516 3612
rect 14660 3602 14688 4694
rect 14752 4622 14780 5170
rect 15016 5092 15068 5098
rect 15120 5080 15148 5222
rect 15200 5160 15252 5166
rect 15200 5102 15252 5108
rect 15068 5052 15148 5080
rect 15016 5034 15068 5040
rect 14817 4924 15113 4944
rect 14873 4922 14897 4924
rect 14953 4922 14977 4924
rect 15033 4922 15057 4924
rect 14895 4870 14897 4922
rect 14959 4870 14971 4922
rect 15033 4870 15035 4922
rect 14873 4868 14897 4870
rect 14953 4868 14977 4870
rect 15033 4868 15057 4870
rect 14817 4848 15113 4868
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 15120 4282 15148 4626
rect 15212 4622 15240 5102
rect 15304 5098 15332 5646
rect 15292 5092 15344 5098
rect 15292 5034 15344 5040
rect 15200 4616 15252 4622
rect 15200 4558 15252 4564
rect 15108 4276 15160 4282
rect 15108 4218 15160 4224
rect 15198 3904 15254 3913
rect 14817 3836 15113 3856
rect 15198 3839 15254 3848
rect 14873 3834 14897 3836
rect 14953 3834 14977 3836
rect 15033 3834 15057 3836
rect 14895 3782 14897 3834
rect 14959 3782 14971 3834
rect 15033 3782 15035 3834
rect 14873 3780 14897 3782
rect 14953 3780 14977 3782
rect 15033 3780 15057 3782
rect 14817 3760 15113 3780
rect 15212 3738 15240 3839
rect 15200 3732 15252 3738
rect 15200 3674 15252 3680
rect 15292 3664 15344 3670
rect 15292 3606 15344 3612
rect 14648 3596 14700 3602
rect 14648 3538 14700 3544
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 14740 3392 14792 3398
rect 14740 3334 14792 3340
rect 14646 3088 14702 3097
rect 14646 3023 14702 3032
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 14186 2544 14242 2553
rect 14660 2514 14688 3023
rect 14186 2479 14188 2488
rect 14240 2479 14242 2488
rect 14556 2508 14608 2514
rect 14188 2450 14240 2456
rect 14556 2450 14608 2456
rect 14648 2508 14700 2514
rect 14648 2450 14700 2456
rect 13912 2440 13964 2446
rect 12716 2382 12768 2388
rect 13818 2408 13874 2417
rect 12636 2038 12664 2382
rect 13544 2372 13596 2378
rect 13912 2382 13964 2388
rect 13818 2343 13874 2352
rect 13544 2314 13596 2320
rect 12716 2304 12768 2310
rect 12716 2246 12768 2252
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 12256 2032 12308 2038
rect 12256 1974 12308 1980
rect 12624 2032 12676 2038
rect 12624 1974 12676 1980
rect 12268 800 12296 1974
rect 12728 800 12756 2246
rect 13096 800 13124 2246
rect 13556 800 13584 2314
rect 14096 2304 14148 2310
rect 14096 2246 14148 2252
rect 14464 2304 14516 2310
rect 14464 2246 14516 2252
rect 14108 1170 14136 2246
rect 14476 1170 14504 2246
rect 14568 2038 14596 2450
rect 14556 2032 14608 2038
rect 14556 1974 14608 1980
rect 14752 1442 14780 3334
rect 15120 3194 15148 3538
rect 15304 3398 15332 3606
rect 15292 3392 15344 3398
rect 15292 3334 15344 3340
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 15396 2990 15424 9687
rect 15488 9586 15516 9930
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15474 9480 15530 9489
rect 15474 9415 15530 9424
rect 15488 8265 15516 9415
rect 15474 8256 15530 8265
rect 15474 8191 15530 8200
rect 15476 7880 15528 7886
rect 15580 7868 15608 15558
rect 15856 15502 15884 16510
rect 16672 16458 16724 16464
rect 15936 16448 15988 16454
rect 15936 16390 15988 16396
rect 15948 16046 15976 16390
rect 16684 16046 16712 16458
rect 15936 16040 15988 16046
rect 15936 15982 15988 15988
rect 16672 16040 16724 16046
rect 16672 15982 16724 15988
rect 15844 15496 15896 15502
rect 15764 15456 15844 15484
rect 15764 14006 15792 15456
rect 15844 15438 15896 15444
rect 15948 15162 15976 15982
rect 16304 15972 16356 15978
rect 16304 15914 16356 15920
rect 16316 15502 16344 15914
rect 16856 15564 16908 15570
rect 16856 15506 16908 15512
rect 16304 15496 16356 15502
rect 16304 15438 16356 15444
rect 15936 15156 15988 15162
rect 15936 15098 15988 15104
rect 16316 15094 16344 15438
rect 16868 15434 16896 15506
rect 16856 15428 16908 15434
rect 16856 15370 16908 15376
rect 16580 15156 16632 15162
rect 16580 15098 16632 15104
rect 16304 15088 16356 15094
rect 16304 15030 16356 15036
rect 15844 14952 15896 14958
rect 15844 14894 15896 14900
rect 15856 14618 15884 14894
rect 16120 14884 16172 14890
rect 16120 14826 16172 14832
rect 16028 14816 16080 14822
rect 16028 14758 16080 14764
rect 15844 14612 15896 14618
rect 15844 14554 15896 14560
rect 16040 14550 16068 14758
rect 16028 14544 16080 14550
rect 16028 14486 16080 14492
rect 15934 14240 15990 14249
rect 15934 14175 15990 14184
rect 15752 14000 15804 14006
rect 15752 13942 15804 13948
rect 15764 13734 15792 13942
rect 15948 13870 15976 14175
rect 15844 13864 15896 13870
rect 15844 13806 15896 13812
rect 15936 13864 15988 13870
rect 15936 13806 15988 13812
rect 15752 13728 15804 13734
rect 15752 13670 15804 13676
rect 15660 12368 15712 12374
rect 15660 12310 15712 12316
rect 15672 11898 15700 12310
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15672 8922 15700 11698
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 15764 11286 15792 11494
rect 15752 11280 15804 11286
rect 15752 11222 15804 11228
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 15764 10198 15792 10406
rect 15752 10192 15804 10198
rect 15752 10134 15804 10140
rect 15750 10024 15806 10033
rect 15750 9959 15806 9968
rect 15764 9926 15792 9959
rect 15752 9920 15804 9926
rect 15752 9862 15804 9868
rect 15856 9738 15884 13806
rect 15936 13456 15988 13462
rect 15936 13398 15988 13404
rect 15948 12646 15976 13398
rect 16040 13326 16068 14486
rect 16132 13530 16160 14826
rect 16120 13524 16172 13530
rect 16120 13466 16172 13472
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 16040 12850 16068 13262
rect 16212 13252 16264 13258
rect 16212 13194 16264 13200
rect 16028 12844 16080 12850
rect 16028 12786 16080 12792
rect 15936 12640 15988 12646
rect 15936 12582 15988 12588
rect 16224 12102 16252 13194
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 16212 12096 16264 12102
rect 16212 12038 16264 12044
rect 15936 11144 15988 11150
rect 15936 11086 15988 11092
rect 15948 10742 15976 11086
rect 15936 10736 15988 10742
rect 15936 10678 15988 10684
rect 15936 10600 15988 10606
rect 15936 10542 15988 10548
rect 15948 9926 15976 10542
rect 16040 10198 16068 12038
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 16132 10266 16160 11086
rect 16212 11076 16264 11082
rect 16212 11018 16264 11024
rect 16224 10606 16252 11018
rect 16212 10600 16264 10606
rect 16212 10542 16264 10548
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16028 10192 16080 10198
rect 16028 10134 16080 10140
rect 15936 9920 15988 9926
rect 15936 9862 15988 9868
rect 16212 9920 16264 9926
rect 16212 9862 16264 9868
rect 15856 9710 16068 9738
rect 15752 9580 15804 9586
rect 15752 9522 15804 9528
rect 15764 9178 15792 9522
rect 15934 9480 15990 9489
rect 15934 9415 15990 9424
rect 15844 9376 15896 9382
rect 15844 9318 15896 9324
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15764 9042 15792 9114
rect 15856 9110 15884 9318
rect 15844 9104 15896 9110
rect 15844 9046 15896 9052
rect 15752 9036 15804 9042
rect 15752 8978 15804 8984
rect 15672 8894 15884 8922
rect 15658 8256 15714 8265
rect 15658 8191 15714 8200
rect 15528 7840 15608 7868
rect 15476 7822 15528 7828
rect 15488 6662 15516 7822
rect 15568 7744 15620 7750
rect 15568 7686 15620 7692
rect 15580 7410 15608 7686
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15672 7018 15700 8191
rect 15580 6990 15700 7018
rect 15476 6656 15528 6662
rect 15476 6598 15528 6604
rect 15488 5953 15516 6598
rect 15474 5944 15530 5953
rect 15474 5879 15530 5888
rect 15476 5772 15528 5778
rect 15476 5714 15528 5720
rect 15488 5574 15516 5714
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 15488 5137 15516 5510
rect 15474 5128 15530 5137
rect 15474 5063 15530 5072
rect 15580 4978 15608 6990
rect 15658 6896 15714 6905
rect 15658 6831 15714 6840
rect 15672 6089 15700 6831
rect 15752 6792 15804 6798
rect 15752 6734 15804 6740
rect 15658 6080 15714 6089
rect 15658 6015 15714 6024
rect 15764 5930 15792 6734
rect 15856 6304 15884 8894
rect 15948 8838 15976 9415
rect 15936 8832 15988 8838
rect 15936 8774 15988 8780
rect 15936 8356 15988 8362
rect 15936 8298 15988 8304
rect 15948 7886 15976 8298
rect 15936 7880 15988 7886
rect 16040 7857 16068 9710
rect 16224 9586 16252 9862
rect 16212 9580 16264 9586
rect 16212 9522 16264 9528
rect 16212 9376 16264 9382
rect 16212 9318 16264 9324
rect 16118 9208 16174 9217
rect 16118 9143 16174 9152
rect 16132 7993 16160 9143
rect 16224 8809 16252 9318
rect 16210 8800 16266 8809
rect 16210 8735 16266 8744
rect 16118 7984 16174 7993
rect 16118 7919 16174 7928
rect 15936 7822 15988 7828
rect 16026 7848 16082 7857
rect 16026 7783 16082 7792
rect 16040 7206 16068 7783
rect 16028 7200 16080 7206
rect 16028 7142 16080 7148
rect 16028 6996 16080 7002
rect 16028 6938 16080 6944
rect 15856 6276 15976 6304
rect 15844 6180 15896 6186
rect 15844 6122 15896 6128
rect 15488 4950 15608 4978
rect 15672 5902 15792 5930
rect 15856 5914 15884 6122
rect 15948 5914 15976 6276
rect 15844 5908 15896 5914
rect 15488 4758 15516 4950
rect 15568 4820 15620 4826
rect 15568 4762 15620 4768
rect 15476 4752 15528 4758
rect 15476 4694 15528 4700
rect 15476 4616 15528 4622
rect 15476 4558 15528 4564
rect 15488 4214 15516 4558
rect 15476 4208 15528 4214
rect 15476 4150 15528 4156
rect 15580 4146 15608 4762
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 15476 3936 15528 3942
rect 15476 3878 15528 3884
rect 15488 3641 15516 3878
rect 15474 3632 15530 3641
rect 15474 3567 15530 3576
rect 15384 2984 15436 2990
rect 15384 2926 15436 2932
rect 15568 2916 15620 2922
rect 15568 2858 15620 2864
rect 15476 2848 15528 2854
rect 15476 2790 15528 2796
rect 14817 2748 15113 2768
rect 14873 2746 14897 2748
rect 14953 2746 14977 2748
rect 15033 2746 15057 2748
rect 14895 2694 14897 2746
rect 14959 2694 14971 2746
rect 15033 2694 15035 2746
rect 14873 2692 14897 2694
rect 14953 2692 14977 2694
rect 15033 2692 15057 2694
rect 14817 2672 15113 2692
rect 15488 2378 15516 2790
rect 15580 2514 15608 2858
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 15672 2446 15700 5902
rect 15844 5850 15896 5856
rect 15936 5908 15988 5914
rect 15936 5850 15988 5856
rect 16040 4593 16068 6938
rect 16132 6798 16160 7919
rect 16224 7585 16252 8735
rect 16316 8129 16344 15030
rect 16396 14952 16448 14958
rect 16592 14906 16620 15098
rect 16448 14900 16620 14906
rect 16396 14894 16620 14900
rect 16408 14878 16620 14894
rect 16592 14414 16620 14878
rect 16672 14476 16724 14482
rect 16672 14418 16724 14424
rect 16580 14408 16632 14414
rect 16580 14350 16632 14356
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16408 13938 16436 14214
rect 16396 13932 16448 13938
rect 16396 13874 16448 13880
rect 16408 13326 16436 13874
rect 16684 13818 16712 14418
rect 16592 13790 16712 13818
rect 16488 13728 16540 13734
rect 16488 13670 16540 13676
rect 16500 13530 16528 13670
rect 16488 13524 16540 13530
rect 16488 13466 16540 13472
rect 16396 13320 16448 13326
rect 16396 13262 16448 13268
rect 16592 13138 16620 13790
rect 16408 13110 16620 13138
rect 16408 11937 16436 13110
rect 16672 12708 16724 12714
rect 16672 12650 16724 12656
rect 16684 12238 16712 12650
rect 16764 12640 16816 12646
rect 16764 12582 16816 12588
rect 16776 12442 16804 12582
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16672 12232 16724 12238
rect 16672 12174 16724 12180
rect 16776 12102 16804 12378
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16764 12096 16816 12102
rect 16764 12038 16816 12044
rect 16394 11928 16450 11937
rect 16394 11863 16450 11872
rect 16394 10976 16450 10985
rect 16394 10911 16450 10920
rect 16408 10130 16436 10911
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 16396 10124 16448 10130
rect 16396 10066 16448 10072
rect 16408 9722 16436 10066
rect 16396 9716 16448 9722
rect 16396 9658 16448 9664
rect 16396 9444 16448 9450
rect 16396 9386 16448 9392
rect 16408 8634 16436 9386
rect 16500 9217 16528 10202
rect 16592 9586 16620 12038
rect 16764 11008 16816 11014
rect 16764 10950 16816 10956
rect 16776 10606 16804 10950
rect 16764 10600 16816 10606
rect 16764 10542 16816 10548
rect 16868 10470 16896 15370
rect 16960 14278 16988 19110
rect 17052 18426 17080 22200
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 17144 18902 17172 19246
rect 17420 19174 17448 22200
rect 17592 19304 17644 19310
rect 17592 19246 17644 19252
rect 17408 19168 17460 19174
rect 17408 19110 17460 19116
rect 17132 18896 17184 18902
rect 17132 18838 17184 18844
rect 17604 18834 17632 19246
rect 17788 19174 17816 22200
rect 18156 20058 18184 22200
rect 18282 20700 18578 20720
rect 18338 20698 18362 20700
rect 18418 20698 18442 20700
rect 18498 20698 18522 20700
rect 18360 20646 18362 20698
rect 18424 20646 18436 20698
rect 18498 20646 18500 20698
rect 18338 20644 18362 20646
rect 18418 20644 18442 20646
rect 18498 20644 18522 20646
rect 18282 20624 18578 20644
rect 18144 20052 18196 20058
rect 18144 19994 18196 20000
rect 18282 19612 18578 19632
rect 18338 19610 18362 19612
rect 18418 19610 18442 19612
rect 18498 19610 18522 19612
rect 18360 19558 18362 19610
rect 18424 19558 18436 19610
rect 18498 19558 18500 19610
rect 18338 19556 18362 19558
rect 18418 19556 18442 19558
rect 18498 19556 18522 19558
rect 18282 19536 18578 19556
rect 18512 19304 18564 19310
rect 18510 19272 18512 19281
rect 18564 19272 18566 19281
rect 18510 19207 18566 19216
rect 17776 19168 17828 19174
rect 17776 19110 17828 19116
rect 17868 18896 17920 18902
rect 17868 18838 17920 18844
rect 17592 18828 17644 18834
rect 17592 18770 17644 18776
rect 17040 18420 17092 18426
rect 17040 18362 17092 18368
rect 17224 17604 17276 17610
rect 17224 17546 17276 17552
rect 17236 16794 17264 17546
rect 17224 16788 17276 16794
rect 17224 16730 17276 16736
rect 17132 16652 17184 16658
rect 17132 16594 17184 16600
rect 17040 16108 17092 16114
rect 17040 16050 17092 16056
rect 17052 15910 17080 16050
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 17144 15638 17172 16594
rect 17500 16176 17552 16182
rect 17500 16118 17552 16124
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17420 15706 17448 15846
rect 17408 15700 17460 15706
rect 17408 15642 17460 15648
rect 17132 15632 17184 15638
rect 17224 15632 17276 15638
rect 17132 15574 17184 15580
rect 17222 15600 17224 15609
rect 17276 15600 17278 15609
rect 17222 15535 17278 15544
rect 17040 15496 17092 15502
rect 17040 15438 17092 15444
rect 16948 14272 17000 14278
rect 16948 14214 17000 14220
rect 17052 13530 17080 15438
rect 17316 15020 17368 15026
rect 17316 14962 17368 14968
rect 17328 14414 17356 14962
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 17328 12782 17356 14350
rect 17316 12776 17368 12782
rect 17316 12718 17368 12724
rect 16948 12708 17000 12714
rect 16948 12650 17000 12656
rect 16960 12442 16988 12650
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 17132 12436 17184 12442
rect 17132 12378 17184 12384
rect 16960 12345 16988 12378
rect 16946 12336 17002 12345
rect 16946 12271 17002 12280
rect 17144 12238 17172 12378
rect 17328 12306 17356 12718
rect 17512 12458 17540 16118
rect 17604 14482 17632 18770
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 17604 14074 17632 14418
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 17604 13734 17632 14010
rect 17592 13728 17644 13734
rect 17592 13670 17644 13676
rect 17684 13320 17736 13326
rect 17684 13262 17736 13268
rect 17696 12986 17724 13262
rect 17684 12980 17736 12986
rect 17684 12922 17736 12928
rect 17420 12430 17540 12458
rect 17684 12436 17736 12442
rect 17316 12300 17368 12306
rect 17316 12242 17368 12248
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16960 11082 16988 11494
rect 16948 11076 17000 11082
rect 16948 11018 17000 11024
rect 16856 10464 16908 10470
rect 16908 10424 16988 10452
rect 16856 10406 16908 10412
rect 16856 10056 16908 10062
rect 16776 10016 16856 10044
rect 16776 9926 16804 10016
rect 16856 9998 16908 10004
rect 16960 9926 16988 10424
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 16960 9761 16988 9862
rect 16946 9752 17002 9761
rect 16946 9687 17002 9696
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16580 9580 16632 9586
rect 16580 9522 16632 9528
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16486 9208 16542 9217
rect 16486 9143 16542 9152
rect 16488 9036 16540 9042
rect 16488 8978 16540 8984
rect 16500 8634 16528 8978
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 16488 8628 16540 8634
rect 16488 8570 16540 8576
rect 16302 8120 16358 8129
rect 16302 8055 16358 8064
rect 16316 7886 16344 8055
rect 16500 7954 16528 8570
rect 16488 7948 16540 7954
rect 16488 7890 16540 7896
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16210 7576 16266 7585
rect 16210 7511 16266 7520
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16120 6656 16172 6662
rect 16120 6598 16172 6604
rect 16132 6254 16160 6598
rect 16120 6248 16172 6254
rect 16120 6190 16172 6196
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 16026 4584 16082 4593
rect 16026 4519 16082 4528
rect 15844 4140 15896 4146
rect 15844 4082 15896 4088
rect 16028 4140 16080 4146
rect 16028 4082 16080 4088
rect 15856 3534 15884 4082
rect 15752 3528 15804 3534
rect 15752 3470 15804 3476
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 15764 3398 15792 3470
rect 16040 3466 16068 4082
rect 16132 3942 16160 4966
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 16132 3602 16160 3878
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 15936 3460 15988 3466
rect 15936 3402 15988 3408
rect 16028 3460 16080 3466
rect 16028 3402 16080 3408
rect 15752 3392 15804 3398
rect 15752 3334 15804 3340
rect 15764 2961 15792 3334
rect 15948 2990 15976 3402
rect 15936 2984 15988 2990
rect 15750 2952 15806 2961
rect 15936 2926 15988 2932
rect 15750 2887 15806 2896
rect 16224 2650 16252 7511
rect 16500 7410 16528 7890
rect 16592 7546 16620 9318
rect 16684 8022 16712 9590
rect 16764 9580 16816 9586
rect 16764 9522 16816 9528
rect 16856 9580 16908 9586
rect 16856 9522 16908 9528
rect 16776 8498 16804 9522
rect 16868 8838 16896 9522
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16868 8430 16896 8774
rect 16856 8424 16908 8430
rect 16856 8366 16908 8372
rect 16764 8288 16816 8294
rect 16764 8230 16816 8236
rect 16856 8288 16908 8294
rect 16856 8230 16908 8236
rect 16672 8016 16724 8022
rect 16672 7958 16724 7964
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 16672 7540 16724 7546
rect 16672 7482 16724 7488
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16396 7336 16448 7342
rect 16684 7290 16712 7482
rect 16396 7278 16448 7284
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16316 6934 16344 7142
rect 16304 6928 16356 6934
rect 16304 6870 16356 6876
rect 16408 4826 16436 7278
rect 16500 7262 16712 7290
rect 16776 7274 16804 8230
rect 16868 7546 16896 8230
rect 16960 7818 16988 9318
rect 16948 7812 17000 7818
rect 16948 7754 17000 7760
rect 17052 7698 17080 12038
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 17316 11212 17368 11218
rect 17316 11154 17368 11160
rect 17144 9178 17172 11154
rect 17328 10810 17356 11154
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17420 10282 17448 12430
rect 17684 12378 17736 12384
rect 17592 12300 17644 12306
rect 17592 12242 17644 12248
rect 17604 11898 17632 12242
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 17696 11778 17724 12378
rect 17604 11750 17724 11778
rect 17500 11620 17552 11626
rect 17500 11562 17552 11568
rect 17512 11082 17540 11562
rect 17500 11076 17552 11082
rect 17500 11018 17552 11024
rect 17512 10470 17540 11018
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17236 10254 17448 10282
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 17144 8129 17172 8366
rect 17130 8120 17186 8129
rect 17130 8055 17186 8064
rect 16960 7670 17080 7698
rect 16856 7540 16908 7546
rect 16856 7482 16908 7488
rect 16854 7440 16910 7449
rect 16854 7375 16856 7384
rect 16908 7375 16910 7384
rect 16856 7346 16908 7352
rect 16500 7002 16528 7262
rect 16684 7206 16712 7262
rect 16764 7268 16816 7274
rect 16764 7210 16816 7216
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 16672 7200 16724 7206
rect 16672 7142 16724 7148
rect 16488 6996 16540 7002
rect 16488 6938 16540 6944
rect 16486 6624 16542 6633
rect 16486 6559 16542 6568
rect 16500 4865 16528 6559
rect 16592 5370 16620 7142
rect 16764 6384 16816 6390
rect 16764 6326 16816 6332
rect 16672 5908 16724 5914
rect 16672 5850 16724 5856
rect 16684 5574 16712 5850
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 16580 5364 16632 5370
rect 16580 5306 16632 5312
rect 16672 5296 16724 5302
rect 16672 5238 16724 5244
rect 16580 5228 16632 5234
rect 16580 5170 16632 5176
rect 16486 4856 16542 4865
rect 16396 4820 16448 4826
rect 16486 4791 16542 4800
rect 16396 4762 16448 4768
rect 16408 4078 16436 4762
rect 16592 4554 16620 5170
rect 16684 4758 16712 5238
rect 16776 5234 16804 6326
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 16764 5228 16816 5234
rect 16764 5170 16816 5176
rect 16868 5166 16896 6054
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 16672 4752 16724 4758
rect 16672 4694 16724 4700
rect 16580 4548 16632 4554
rect 16580 4490 16632 4496
rect 16960 4486 16988 7670
rect 17132 7540 17184 7546
rect 17132 7482 17184 7488
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 17052 6798 17080 7346
rect 17144 7002 17172 7482
rect 17132 6996 17184 7002
rect 17132 6938 17184 6944
rect 17236 6866 17264 10254
rect 17314 9888 17370 9897
rect 17314 9823 17370 9832
rect 17328 7041 17356 9823
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 17420 9178 17448 9318
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 17420 8294 17448 9114
rect 17500 8968 17552 8974
rect 17500 8910 17552 8916
rect 17512 8634 17540 8910
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17406 7712 17462 7721
rect 17406 7647 17462 7656
rect 17420 7274 17448 7647
rect 17512 7546 17540 8570
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17604 7426 17632 11750
rect 17788 11642 17816 14214
rect 17880 13841 17908 18838
rect 18236 18760 18288 18766
rect 18234 18728 18236 18737
rect 18288 18728 18290 18737
rect 18234 18663 18290 18672
rect 18616 18630 18644 22200
rect 18984 20602 19012 22200
rect 19154 22199 19210 22208
rect 19338 22200 19394 23000
rect 19706 22200 19762 23000
rect 19982 22672 20038 22681
rect 19982 22607 20038 22616
rect 18972 20596 19024 20602
rect 18972 20538 19024 20544
rect 18984 19922 19012 20538
rect 19062 20224 19118 20233
rect 19062 20159 19118 20168
rect 18972 19916 19024 19922
rect 18972 19858 19024 19864
rect 18984 19378 19012 19858
rect 18972 19372 19024 19378
rect 18972 19314 19024 19320
rect 18694 19272 18750 19281
rect 18694 19207 18750 19216
rect 18972 19236 19024 19242
rect 18604 18624 18656 18630
rect 18604 18566 18656 18572
rect 18282 18524 18578 18544
rect 18338 18522 18362 18524
rect 18418 18522 18442 18524
rect 18498 18522 18522 18524
rect 18360 18470 18362 18522
rect 18424 18470 18436 18522
rect 18498 18470 18500 18522
rect 18338 18468 18362 18470
rect 18418 18468 18442 18470
rect 18498 18468 18522 18470
rect 18282 18448 18578 18468
rect 18708 18426 18736 19207
rect 18972 19178 19024 19184
rect 18984 18902 19012 19178
rect 18972 18896 19024 18902
rect 18972 18838 19024 18844
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18696 18420 18748 18426
rect 18696 18362 18748 18368
rect 18800 18329 18828 18702
rect 18786 18320 18842 18329
rect 18786 18255 18842 18264
rect 18052 18216 18104 18222
rect 18052 18158 18104 18164
rect 17960 15428 18012 15434
rect 17960 15370 18012 15376
rect 17972 15162 18000 15370
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 17972 14958 18000 15098
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 18064 14113 18092 18158
rect 18282 17436 18578 17456
rect 18338 17434 18362 17436
rect 18418 17434 18442 17436
rect 18498 17434 18522 17436
rect 18360 17382 18362 17434
rect 18424 17382 18436 17434
rect 18498 17382 18500 17434
rect 18338 17380 18362 17382
rect 18418 17380 18442 17382
rect 18498 17380 18522 17382
rect 18282 17360 18578 17380
rect 18282 16348 18578 16368
rect 18338 16346 18362 16348
rect 18418 16346 18442 16348
rect 18498 16346 18522 16348
rect 18360 16294 18362 16346
rect 18424 16294 18436 16346
rect 18498 16294 18500 16346
rect 18338 16292 18362 16294
rect 18418 16292 18442 16294
rect 18498 16292 18522 16294
rect 18282 16272 18578 16292
rect 19076 16250 19104 20159
rect 19168 18986 19196 22199
rect 19246 20632 19302 20641
rect 19352 20602 19380 22200
rect 19246 20567 19302 20576
rect 19340 20596 19392 20602
rect 19260 19990 19288 20567
rect 19340 20538 19392 20544
rect 19248 19984 19300 19990
rect 19248 19926 19300 19932
rect 19352 19854 19380 20538
rect 19616 20256 19668 20262
rect 19616 20198 19668 20204
rect 19432 19984 19484 19990
rect 19432 19926 19484 19932
rect 19340 19848 19392 19854
rect 19340 19790 19392 19796
rect 19168 18958 19288 18986
rect 19444 18970 19472 19926
rect 19628 19922 19656 20198
rect 19616 19916 19668 19922
rect 19616 19858 19668 19864
rect 19628 19360 19656 19858
rect 19720 19802 19748 22200
rect 19996 19990 20024 22607
rect 20074 22200 20130 23000
rect 20442 22200 20498 23000
rect 20902 22200 20958 23000
rect 21270 22200 21326 23000
rect 21638 22200 21694 23000
rect 22006 22200 22062 23000
rect 22374 22200 22430 23000
rect 22742 22200 22798 23000
rect 19984 19984 20036 19990
rect 19984 19926 20036 19932
rect 19720 19774 19840 19802
rect 19706 19680 19762 19689
rect 19706 19615 19762 19624
rect 19536 19332 19656 19360
rect 19536 19242 19564 19332
rect 19524 19236 19576 19242
rect 19524 19178 19576 19184
rect 19616 19236 19668 19242
rect 19616 19178 19668 19184
rect 19260 18902 19288 18958
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 19248 18896 19300 18902
rect 19248 18838 19300 18844
rect 19338 18864 19394 18873
rect 19338 18799 19394 18808
rect 19352 18766 19380 18799
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 19340 18080 19392 18086
rect 19340 18022 19392 18028
rect 19352 17066 19380 18022
rect 19536 17202 19564 19178
rect 19524 17196 19576 17202
rect 19524 17138 19576 17144
rect 19340 17060 19392 17066
rect 19392 17020 19472 17048
rect 19340 17002 19392 17008
rect 19064 16244 19116 16250
rect 19064 16186 19116 16192
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 18144 15564 18196 15570
rect 18144 15506 18196 15512
rect 18050 14104 18106 14113
rect 17960 14068 18012 14074
rect 18156 14074 18184 15506
rect 18696 15428 18748 15434
rect 18696 15370 18748 15376
rect 18282 15260 18578 15280
rect 18338 15258 18362 15260
rect 18418 15258 18442 15260
rect 18498 15258 18522 15260
rect 18360 15206 18362 15258
rect 18424 15206 18436 15258
rect 18498 15206 18500 15258
rect 18338 15204 18362 15206
rect 18418 15204 18442 15206
rect 18498 15204 18522 15206
rect 18282 15184 18578 15204
rect 18604 14476 18656 14482
rect 18604 14418 18656 14424
rect 18282 14172 18578 14192
rect 18338 14170 18362 14172
rect 18418 14170 18442 14172
rect 18498 14170 18522 14172
rect 18360 14118 18362 14170
rect 18424 14118 18436 14170
rect 18498 14118 18500 14170
rect 18338 14116 18362 14118
rect 18418 14116 18442 14118
rect 18498 14116 18522 14118
rect 18282 14096 18578 14116
rect 18050 14039 18106 14048
rect 18144 14068 18196 14074
rect 17960 14010 18012 14016
rect 17866 13832 17922 13841
rect 17972 13802 18000 14010
rect 17866 13767 17922 13776
rect 17960 13796 18012 13802
rect 17696 11614 17816 11642
rect 17696 10452 17724 11614
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 17788 10577 17816 11494
rect 17880 10674 17908 13767
rect 17960 13738 18012 13744
rect 18064 13512 18092 14039
rect 18144 14010 18196 14016
rect 18616 13938 18644 14418
rect 18604 13932 18656 13938
rect 18604 13874 18656 13880
rect 18064 13484 18184 13512
rect 18052 13388 18104 13394
rect 18052 13330 18104 13336
rect 18064 12986 18092 13330
rect 18052 12980 18104 12986
rect 18052 12922 18104 12928
rect 18156 11286 18184 13484
rect 18616 13326 18644 13874
rect 18708 13870 18736 15370
rect 19156 15360 19208 15366
rect 19156 15302 19208 15308
rect 18880 14884 18932 14890
rect 18880 14826 18932 14832
rect 18892 14346 18920 14826
rect 19168 14482 19196 15302
rect 19156 14476 19208 14482
rect 19156 14418 19208 14424
rect 19062 14376 19118 14385
rect 18880 14340 18932 14346
rect 19062 14311 19118 14320
rect 18880 14282 18932 14288
rect 18892 13938 18920 14282
rect 18972 14272 19024 14278
rect 18972 14214 19024 14220
rect 18880 13932 18932 13938
rect 18880 13874 18932 13880
rect 18696 13864 18748 13870
rect 18696 13806 18748 13812
rect 18788 13388 18840 13394
rect 18788 13330 18840 13336
rect 18604 13320 18656 13326
rect 18604 13262 18656 13268
rect 18282 13084 18578 13104
rect 18338 13082 18362 13084
rect 18418 13082 18442 13084
rect 18498 13082 18522 13084
rect 18360 13030 18362 13082
rect 18424 13030 18436 13082
rect 18498 13030 18500 13082
rect 18338 13028 18362 13030
rect 18418 13028 18442 13030
rect 18498 13028 18522 13030
rect 18282 13008 18578 13028
rect 18696 12708 18748 12714
rect 18696 12650 18748 12656
rect 18708 12170 18736 12650
rect 18800 12442 18828 13330
rect 18892 13258 18920 13874
rect 18984 13870 19012 14214
rect 19076 14074 19104 14311
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 18972 13864 19024 13870
rect 18972 13806 19024 13812
rect 18880 13252 18932 13258
rect 18880 13194 18932 13200
rect 18788 12436 18840 12442
rect 18788 12378 18840 12384
rect 18970 12200 19026 12209
rect 18696 12164 18748 12170
rect 18970 12135 19026 12144
rect 18696 12106 18748 12112
rect 18282 11996 18578 12016
rect 18338 11994 18362 11996
rect 18418 11994 18442 11996
rect 18498 11994 18522 11996
rect 18360 11942 18362 11994
rect 18424 11942 18436 11994
rect 18498 11942 18500 11994
rect 18338 11940 18362 11942
rect 18418 11940 18442 11942
rect 18498 11940 18522 11942
rect 18282 11920 18578 11940
rect 18708 11762 18736 12106
rect 18984 11830 19012 12135
rect 18972 11824 19024 11830
rect 18972 11766 19024 11772
rect 18696 11756 18748 11762
rect 18696 11698 18748 11704
rect 18144 11280 18196 11286
rect 18144 11222 18196 11228
rect 18156 10810 18184 11222
rect 18248 11218 18828 11234
rect 18236 11212 18828 11218
rect 18288 11206 18828 11212
rect 18236 11154 18288 11160
rect 18604 11144 18656 11150
rect 18656 11092 18736 11098
rect 18604 11086 18736 11092
rect 18616 11070 18736 11086
rect 18616 11014 18644 11070
rect 18604 11008 18656 11014
rect 18604 10950 18656 10956
rect 18282 10908 18578 10928
rect 18338 10906 18362 10908
rect 18418 10906 18442 10908
rect 18498 10906 18522 10908
rect 18360 10854 18362 10906
rect 18424 10854 18436 10906
rect 18498 10854 18500 10906
rect 18338 10852 18362 10854
rect 18418 10852 18442 10854
rect 18498 10852 18522 10854
rect 18282 10832 18578 10852
rect 18144 10804 18196 10810
rect 18144 10746 18196 10752
rect 18708 10674 18736 11070
rect 18800 10674 18828 11206
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18788 10668 18840 10674
rect 18788 10610 18840 10616
rect 17774 10568 17830 10577
rect 17774 10503 17830 10512
rect 18144 10532 18196 10538
rect 18144 10474 18196 10480
rect 17696 10424 17816 10452
rect 17684 10192 17736 10198
rect 17684 10134 17736 10140
rect 17696 8974 17724 10134
rect 17684 8968 17736 8974
rect 17788 8945 17816 10424
rect 17866 9752 17922 9761
rect 17866 9687 17922 9696
rect 17684 8910 17736 8916
rect 17774 8936 17830 8945
rect 17774 8871 17830 8880
rect 17684 8492 17736 8498
rect 17684 8434 17736 8440
rect 17696 7886 17724 8434
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 17788 7546 17816 8871
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 17512 7398 17632 7426
rect 17408 7268 17460 7274
rect 17408 7210 17460 7216
rect 17314 7032 17370 7041
rect 17314 6967 17370 6976
rect 17224 6860 17276 6866
rect 17144 6820 17224 6848
rect 17040 6792 17092 6798
rect 17040 6734 17092 6740
rect 17040 6112 17092 6118
rect 17040 6054 17092 6060
rect 17052 5914 17080 6054
rect 17040 5908 17092 5914
rect 17144 5896 17172 6820
rect 17224 6802 17276 6808
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17224 6724 17276 6730
rect 17224 6666 17276 6672
rect 17236 6322 17264 6666
rect 17420 6322 17448 6802
rect 17224 6316 17276 6322
rect 17224 6258 17276 6264
rect 17408 6316 17460 6322
rect 17408 6258 17460 6264
rect 17316 5908 17368 5914
rect 17144 5868 17264 5896
rect 17040 5850 17092 5856
rect 17132 5772 17184 5778
rect 17132 5714 17184 5720
rect 17144 5370 17172 5714
rect 17236 5710 17264 5868
rect 17512 5896 17540 7398
rect 17788 7342 17816 7482
rect 17776 7336 17828 7342
rect 17776 7278 17828 7284
rect 17592 6928 17644 6934
rect 17592 6870 17644 6876
rect 17604 5914 17632 6870
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17682 6216 17738 6225
rect 17682 6151 17684 6160
rect 17736 6151 17738 6160
rect 17684 6122 17736 6128
rect 17788 5914 17816 6598
rect 17368 5868 17540 5896
rect 17592 5908 17644 5914
rect 17316 5850 17368 5856
rect 17592 5850 17644 5856
rect 17776 5908 17828 5914
rect 17776 5850 17828 5856
rect 17224 5704 17276 5710
rect 17224 5646 17276 5652
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 17328 5166 17356 5850
rect 17880 5794 17908 9687
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 17972 7954 18000 8774
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 17972 6390 18000 7890
rect 18064 7546 18092 8910
rect 18156 8378 18184 10474
rect 18708 10266 18736 10610
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18432 10062 18460 10202
rect 18788 10124 18840 10130
rect 18788 10066 18840 10072
rect 18420 10056 18472 10062
rect 18420 9998 18472 10004
rect 18604 9920 18656 9926
rect 18604 9862 18656 9868
rect 18282 9820 18578 9840
rect 18338 9818 18362 9820
rect 18418 9818 18442 9820
rect 18498 9818 18522 9820
rect 18360 9766 18362 9818
rect 18424 9766 18436 9818
rect 18498 9766 18500 9818
rect 18338 9764 18362 9766
rect 18418 9764 18442 9766
rect 18498 9764 18522 9766
rect 18282 9744 18578 9764
rect 18616 9518 18644 9862
rect 18604 9512 18656 9518
rect 18604 9454 18656 9460
rect 18512 9376 18564 9382
rect 18512 9318 18564 9324
rect 18524 9178 18552 9318
rect 18512 9172 18564 9178
rect 18512 9114 18564 9120
rect 18616 8838 18644 9454
rect 18604 8832 18656 8838
rect 18604 8774 18656 8780
rect 18282 8732 18578 8752
rect 18338 8730 18362 8732
rect 18418 8730 18442 8732
rect 18498 8730 18522 8732
rect 18360 8678 18362 8730
rect 18424 8678 18436 8730
rect 18498 8678 18500 8730
rect 18338 8676 18362 8678
rect 18418 8676 18442 8678
rect 18498 8676 18522 8678
rect 18282 8656 18578 8676
rect 18510 8528 18566 8537
rect 18510 8463 18566 8472
rect 18604 8492 18656 8498
rect 18524 8430 18552 8463
rect 18604 8434 18656 8440
rect 18512 8424 18564 8430
rect 18156 8350 18276 8378
rect 18512 8366 18564 8372
rect 18144 8288 18196 8294
rect 18144 8230 18196 8236
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 18156 7002 18184 8230
rect 18248 8090 18276 8350
rect 18236 8084 18288 8090
rect 18236 8026 18288 8032
rect 18616 7954 18644 8434
rect 18696 8424 18748 8430
rect 18696 8366 18748 8372
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 18282 7644 18578 7664
rect 18338 7642 18362 7644
rect 18418 7642 18442 7644
rect 18498 7642 18522 7644
rect 18360 7590 18362 7642
rect 18424 7590 18436 7642
rect 18498 7590 18500 7642
rect 18338 7588 18362 7590
rect 18418 7588 18442 7590
rect 18498 7588 18522 7590
rect 18282 7568 18578 7588
rect 18616 7546 18644 7890
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 18616 7410 18644 7482
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18144 6996 18196 7002
rect 18144 6938 18196 6944
rect 18512 6928 18564 6934
rect 18512 6870 18564 6876
rect 18144 6792 18196 6798
rect 18144 6734 18196 6740
rect 18156 6458 18184 6734
rect 18524 6644 18552 6870
rect 18616 6798 18644 7346
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 18708 6662 18736 8366
rect 18800 7585 18828 10066
rect 18972 10056 19024 10062
rect 18972 9998 19024 10004
rect 18984 9518 19012 9998
rect 18972 9512 19024 9518
rect 18972 9454 19024 9460
rect 18880 9376 18932 9382
rect 18880 9318 18932 9324
rect 18972 9376 19024 9382
rect 18972 9318 19024 9324
rect 18786 7576 18842 7585
rect 18786 7511 18842 7520
rect 18892 6730 18920 9318
rect 18984 8634 19012 9318
rect 19076 9217 19104 14010
rect 19352 14006 19380 15642
rect 19444 14550 19472 17020
rect 19524 14816 19576 14822
rect 19524 14758 19576 14764
rect 19536 14618 19564 14758
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 19432 14544 19484 14550
rect 19432 14486 19484 14492
rect 19340 14000 19392 14006
rect 19340 13942 19392 13948
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19444 12918 19472 13262
rect 19432 12912 19484 12918
rect 19432 12854 19484 12860
rect 19340 12708 19392 12714
rect 19340 12650 19392 12656
rect 19352 11898 19380 12650
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 19444 11830 19472 12378
rect 19432 11824 19484 11830
rect 19628 11801 19656 19178
rect 19720 18426 19748 19615
rect 19812 18970 19840 19774
rect 20088 19174 20116 22200
rect 20456 21978 20484 22200
rect 20456 21950 20668 21978
rect 20534 21856 20590 21865
rect 20534 21791 20590 21800
rect 20442 21448 20498 21457
rect 20442 21383 20498 21392
rect 20456 19310 20484 21383
rect 20548 19990 20576 21791
rect 20640 20534 20668 21950
rect 20916 20602 20944 22200
rect 20994 21040 21050 21049
rect 20994 20975 21050 20984
rect 20904 20596 20956 20602
rect 20904 20538 20956 20544
rect 20628 20528 20680 20534
rect 20628 20470 20680 20476
rect 20640 19990 20668 20470
rect 20916 20398 20944 20538
rect 20720 20392 20772 20398
rect 20720 20334 20772 20340
rect 20904 20392 20956 20398
rect 20904 20334 20956 20340
rect 20536 19984 20588 19990
rect 20536 19926 20588 19932
rect 20628 19984 20680 19990
rect 20628 19926 20680 19932
rect 20628 19848 20680 19854
rect 20628 19790 20680 19796
rect 20640 19310 20668 19790
rect 20168 19304 20220 19310
rect 20168 19246 20220 19252
rect 20444 19304 20496 19310
rect 20444 19246 20496 19252
rect 20628 19304 20680 19310
rect 20628 19246 20680 19252
rect 20076 19168 20128 19174
rect 20076 19110 20128 19116
rect 20180 18970 20208 19246
rect 19800 18964 19852 18970
rect 19800 18906 19852 18912
rect 20168 18964 20220 18970
rect 20168 18906 20220 18912
rect 19812 18698 19840 18906
rect 19800 18692 19852 18698
rect 19800 18634 19852 18640
rect 19708 18420 19760 18426
rect 19708 18362 19760 18368
rect 20180 18358 20208 18906
rect 20732 18834 20760 20334
rect 21008 19310 21036 20975
rect 21284 20262 21312 22200
rect 21272 20256 21324 20262
rect 21272 20198 21324 20204
rect 21652 19990 21680 22200
rect 21640 19984 21692 19990
rect 21640 19926 21692 19932
rect 21272 19372 21324 19378
rect 21272 19314 21324 19320
rect 20996 19304 21048 19310
rect 20996 19246 21048 19252
rect 20720 18828 20772 18834
rect 20720 18770 20772 18776
rect 20536 18624 20588 18630
rect 20536 18566 20588 18572
rect 20168 18352 20220 18358
rect 20168 18294 20220 18300
rect 19984 18080 20036 18086
rect 19984 18022 20036 18028
rect 20074 18048 20130 18057
rect 19706 17640 19762 17649
rect 19706 17575 19708 17584
rect 19760 17575 19762 17584
rect 19708 17546 19760 17552
rect 19708 17128 19760 17134
rect 19708 17070 19760 17076
rect 19432 11766 19484 11772
rect 19614 11792 19670 11801
rect 19156 11144 19208 11150
rect 19156 11086 19208 11092
rect 19168 10742 19196 11086
rect 19156 10736 19208 10742
rect 19156 10678 19208 10684
rect 19444 10690 19472 11766
rect 19614 11727 19670 11736
rect 19444 10662 19564 10690
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 19156 9920 19208 9926
rect 19156 9862 19208 9868
rect 19168 9625 19196 9862
rect 19154 9616 19210 9625
rect 19154 9551 19210 9560
rect 19062 9208 19118 9217
rect 19062 9143 19118 9152
rect 19168 8786 19196 9551
rect 19248 9104 19300 9110
rect 19248 9046 19300 9052
rect 19076 8758 19196 8786
rect 18972 8628 19024 8634
rect 18972 8570 19024 8576
rect 18972 8084 19024 8090
rect 18972 8026 19024 8032
rect 18880 6724 18932 6730
rect 18880 6666 18932 6672
rect 18604 6656 18656 6662
rect 18524 6616 18604 6644
rect 18604 6598 18656 6604
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18282 6556 18578 6576
rect 18338 6554 18362 6556
rect 18418 6554 18442 6556
rect 18498 6554 18522 6556
rect 18360 6502 18362 6554
rect 18424 6502 18436 6554
rect 18498 6502 18500 6554
rect 18338 6500 18362 6502
rect 18418 6500 18442 6502
rect 18498 6500 18522 6502
rect 18282 6480 18578 6500
rect 18144 6452 18196 6458
rect 18144 6394 18196 6400
rect 17960 6384 18012 6390
rect 17960 6326 18012 6332
rect 18144 6112 18196 6118
rect 18144 6054 18196 6060
rect 18156 5914 18184 6054
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 17408 5772 17460 5778
rect 17408 5714 17460 5720
rect 17788 5766 17908 5794
rect 17420 5234 17448 5714
rect 17592 5296 17644 5302
rect 17592 5238 17644 5244
rect 17408 5228 17460 5234
rect 17408 5170 17460 5176
rect 17316 5160 17368 5166
rect 17316 5102 17368 5108
rect 17132 4684 17184 4690
rect 17132 4626 17184 4632
rect 16948 4480 17000 4486
rect 16948 4422 17000 4428
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16672 4072 16724 4078
rect 16672 4014 16724 4020
rect 16684 3534 16712 4014
rect 16764 3732 16816 3738
rect 16764 3674 16816 3680
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 16488 2848 16540 2854
rect 16488 2790 16540 2796
rect 16212 2644 16264 2650
rect 16212 2586 16264 2592
rect 16396 2576 16448 2582
rect 16396 2518 16448 2524
rect 16408 2446 16436 2518
rect 15660 2440 15712 2446
rect 15660 2382 15712 2388
rect 16396 2440 16448 2446
rect 16396 2382 16448 2388
rect 15476 2372 15528 2378
rect 15476 2314 15528 2320
rect 15200 2304 15252 2310
rect 15200 2246 15252 2252
rect 15660 2304 15712 2310
rect 15660 2246 15712 2252
rect 16028 2304 16080 2310
rect 16028 2246 16080 2252
rect 14752 1414 14872 1442
rect 14016 1142 14136 1170
rect 14384 1142 14504 1170
rect 14016 800 14044 1142
rect 14384 800 14412 1142
rect 14844 800 14872 1414
rect 15212 800 15240 2246
rect 15672 800 15700 2246
rect 16040 800 16068 2246
rect 16500 800 16528 2790
rect 16776 1442 16804 3674
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 16868 2514 16896 2994
rect 16960 2990 16988 4422
rect 17144 3194 17172 4626
rect 17500 4276 17552 4282
rect 17500 4218 17552 4224
rect 17512 3602 17540 4218
rect 17500 3596 17552 3602
rect 17500 3538 17552 3544
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 16948 2984 17000 2990
rect 16948 2926 17000 2932
rect 17224 2916 17276 2922
rect 17224 2858 17276 2864
rect 17236 2514 17264 2858
rect 16856 2508 16908 2514
rect 16856 2450 16908 2456
rect 17224 2508 17276 2514
rect 17224 2450 17276 2456
rect 17316 2372 17368 2378
rect 17316 2314 17368 2320
rect 16776 1414 16896 1442
rect 16868 800 16896 1414
rect 17328 800 17356 2314
rect 17604 2310 17632 5238
rect 17788 3641 17816 5766
rect 18156 5302 18184 5850
rect 18282 5468 18578 5488
rect 18338 5466 18362 5468
rect 18418 5466 18442 5468
rect 18498 5466 18522 5468
rect 18360 5414 18362 5466
rect 18424 5414 18436 5466
rect 18498 5414 18500 5466
rect 18338 5412 18362 5414
rect 18418 5412 18442 5414
rect 18498 5412 18522 5414
rect 18282 5392 18578 5412
rect 18144 5296 18196 5302
rect 18144 5238 18196 5244
rect 17868 5160 17920 5166
rect 17866 5128 17868 5137
rect 18052 5160 18104 5166
rect 17920 5128 17922 5137
rect 18052 5102 18104 5108
rect 17866 5063 17922 5072
rect 17868 5024 17920 5030
rect 17868 4966 17920 4972
rect 17880 4826 17908 4966
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 17960 4072 18012 4078
rect 17866 4040 17922 4049
rect 18064 4060 18092 5102
rect 18328 5092 18380 5098
rect 18328 5034 18380 5040
rect 18236 4684 18288 4690
rect 18236 4626 18288 4632
rect 18144 4616 18196 4622
rect 18144 4558 18196 4564
rect 18012 4032 18092 4060
rect 17960 4014 18012 4020
rect 17866 3975 17868 3984
rect 17920 3975 17922 3984
rect 17868 3946 17920 3952
rect 17774 3632 17830 3641
rect 17880 3602 17908 3946
rect 17960 3936 18012 3942
rect 17960 3878 18012 3884
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 17774 3567 17830 3576
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 17684 2644 17736 2650
rect 17684 2586 17736 2592
rect 17592 2304 17644 2310
rect 17592 2246 17644 2252
rect 17696 800 17724 2586
rect 17972 1986 18000 3878
rect 18064 3398 18092 3878
rect 18156 3738 18184 4558
rect 18248 4554 18276 4626
rect 18340 4622 18368 5034
rect 18616 5012 18644 6598
rect 18696 6384 18748 6390
rect 18696 6326 18748 6332
rect 18708 5778 18736 6326
rect 18696 5772 18748 5778
rect 18696 5714 18748 5720
rect 18708 5166 18736 5714
rect 18696 5160 18748 5166
rect 18696 5102 18748 5108
rect 18616 4984 18736 5012
rect 18328 4616 18380 4622
rect 18328 4558 18380 4564
rect 18236 4548 18288 4554
rect 18236 4490 18288 4496
rect 18282 4380 18578 4400
rect 18338 4378 18362 4380
rect 18418 4378 18442 4380
rect 18498 4378 18522 4380
rect 18360 4326 18362 4378
rect 18424 4326 18436 4378
rect 18498 4326 18500 4378
rect 18338 4324 18362 4326
rect 18418 4324 18442 4326
rect 18498 4324 18522 4326
rect 18282 4304 18578 4324
rect 18144 3732 18196 3738
rect 18144 3674 18196 3680
rect 18604 3528 18656 3534
rect 18708 3505 18736 4984
rect 18788 4276 18840 4282
rect 18788 4218 18840 4224
rect 18800 3534 18828 4218
rect 18984 4049 19012 8026
rect 19076 7886 19104 8758
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 19168 8498 19196 8570
rect 19156 8492 19208 8498
rect 19156 8434 19208 8440
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 19076 5370 19104 7822
rect 19168 7750 19196 8434
rect 19156 7744 19208 7750
rect 19156 7686 19208 7692
rect 19168 6798 19196 7686
rect 19156 6792 19208 6798
rect 19156 6734 19208 6740
rect 19260 6730 19288 9046
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19352 8634 19380 8978
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 19338 8528 19394 8537
rect 19338 8463 19394 8472
rect 19352 8090 19380 8463
rect 19340 8084 19392 8090
rect 19340 8026 19392 8032
rect 19340 7948 19392 7954
rect 19340 7890 19392 7896
rect 19352 7342 19380 7890
rect 19444 7478 19472 10542
rect 19536 9602 19564 10662
rect 19720 10554 19748 17070
rect 19892 13184 19944 13190
rect 19892 13126 19944 13132
rect 19904 12782 19932 13126
rect 19892 12776 19944 12782
rect 19892 12718 19944 12724
rect 19996 12594 20024 18022
rect 20074 17983 20130 17992
rect 20088 17882 20116 17983
rect 20076 17876 20128 17882
rect 20076 17818 20128 17824
rect 20444 17128 20496 17134
rect 20444 17070 20496 17076
rect 20456 16726 20484 17070
rect 20444 16720 20496 16726
rect 20444 16662 20496 16668
rect 20168 16176 20220 16182
rect 20168 16118 20220 16124
rect 20180 15026 20208 16118
rect 20168 15020 20220 15026
rect 20168 14962 20220 14968
rect 20352 14408 20404 14414
rect 20352 14350 20404 14356
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 19904 12566 20024 12594
rect 19904 12356 19932 12566
rect 20272 12374 20300 12718
rect 19628 10526 19748 10554
rect 19812 12328 19932 12356
rect 20260 12368 20312 12374
rect 19628 9722 19656 10526
rect 19708 10464 19760 10470
rect 19708 10406 19760 10412
rect 19616 9716 19668 9722
rect 19616 9658 19668 9664
rect 19527 9574 19564 9602
rect 19527 9500 19555 9574
rect 19527 9472 19564 9500
rect 19536 8922 19564 9472
rect 19720 9450 19748 10406
rect 19812 9636 19840 12328
rect 20260 12310 20312 12316
rect 20076 12096 20128 12102
rect 20076 12038 20128 12044
rect 19892 10668 19944 10674
rect 19892 10610 19944 10616
rect 19904 10130 19932 10610
rect 19892 10124 19944 10130
rect 19892 10066 19944 10072
rect 19812 9608 19932 9636
rect 19708 9444 19760 9450
rect 19708 9386 19760 9392
rect 19536 8894 19748 8922
rect 19524 8832 19576 8838
rect 19524 8774 19576 8780
rect 19536 8566 19564 8774
rect 19524 8560 19576 8566
rect 19524 8502 19576 8508
rect 19616 8560 19668 8566
rect 19616 8502 19668 8508
rect 19628 8294 19656 8502
rect 19616 8288 19668 8294
rect 19616 8230 19668 8236
rect 19616 7812 19668 7818
rect 19616 7754 19668 7760
rect 19432 7472 19484 7478
rect 19432 7414 19484 7420
rect 19340 7336 19392 7342
rect 19340 7278 19392 7284
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 19524 7200 19576 7206
rect 19524 7142 19576 7148
rect 19248 6724 19300 6730
rect 19248 6666 19300 6672
rect 19154 6624 19210 6633
rect 19154 6559 19210 6568
rect 19064 5364 19116 5370
rect 19064 5306 19116 5312
rect 18970 4040 19026 4049
rect 18970 3975 19026 3984
rect 18788 3528 18840 3534
rect 18604 3470 18656 3476
rect 18694 3496 18750 3505
rect 18616 3398 18644 3470
rect 18788 3470 18840 3476
rect 18694 3431 18750 3440
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 18144 3392 18196 3398
rect 18144 3334 18196 3340
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18064 3058 18092 3334
rect 18052 3052 18104 3058
rect 18052 2994 18104 3000
rect 18156 2990 18184 3334
rect 18282 3292 18578 3312
rect 18338 3290 18362 3292
rect 18418 3290 18442 3292
rect 18498 3290 18522 3292
rect 18360 3238 18362 3290
rect 18424 3238 18436 3290
rect 18498 3238 18500 3290
rect 18338 3236 18362 3238
rect 18418 3236 18442 3238
rect 18498 3236 18522 3238
rect 18282 3216 18578 3236
rect 18144 2984 18196 2990
rect 18144 2926 18196 2932
rect 18604 2848 18656 2854
rect 18604 2790 18656 2796
rect 18616 2514 18644 2790
rect 18708 2514 18736 3431
rect 18800 3058 18828 3470
rect 19076 3126 19104 5306
rect 19168 4758 19196 6559
rect 19156 4752 19208 4758
rect 19156 4694 19208 4700
rect 19352 3942 19380 7142
rect 19536 7002 19564 7142
rect 19524 6996 19576 7002
rect 19524 6938 19576 6944
rect 19432 6928 19484 6934
rect 19432 6870 19484 6876
rect 19444 6361 19472 6870
rect 19430 6352 19486 6361
rect 19430 6287 19486 6296
rect 19524 5772 19576 5778
rect 19524 5714 19576 5720
rect 19536 5370 19564 5714
rect 19524 5364 19576 5370
rect 19524 5306 19576 5312
rect 19524 4684 19576 4690
rect 19524 4626 19576 4632
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19444 4486 19472 4558
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19444 4282 19472 4422
rect 19432 4276 19484 4282
rect 19432 4218 19484 4224
rect 19536 4146 19564 4626
rect 19524 4140 19576 4146
rect 19524 4082 19576 4088
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 19340 3936 19392 3942
rect 19340 3878 19392 3884
rect 19340 3596 19392 3602
rect 19340 3538 19392 3544
rect 19352 3194 19380 3538
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 18972 3120 19024 3126
rect 18970 3088 18972 3097
rect 19064 3120 19116 3126
rect 19024 3088 19026 3097
rect 18788 3052 18840 3058
rect 19064 3062 19116 3068
rect 18970 3023 19026 3032
rect 18788 2994 18840 3000
rect 19340 2848 19392 2854
rect 19444 2836 19472 4014
rect 19536 3534 19564 4082
rect 19524 3528 19576 3534
rect 19524 3470 19576 3476
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 19392 2808 19472 2836
rect 19340 2790 19392 2796
rect 18604 2508 18656 2514
rect 18604 2450 18656 2456
rect 18696 2508 18748 2514
rect 18696 2450 18748 2456
rect 19340 2372 19392 2378
rect 19340 2314 19392 2320
rect 18604 2304 18656 2310
rect 18604 2246 18656 2252
rect 18972 2304 19024 2310
rect 18972 2246 19024 2252
rect 18282 2204 18578 2224
rect 18338 2202 18362 2204
rect 18418 2202 18442 2204
rect 18498 2202 18522 2204
rect 18360 2150 18362 2202
rect 18424 2150 18436 2202
rect 18498 2150 18500 2202
rect 18338 2148 18362 2150
rect 18418 2148 18442 2150
rect 18498 2148 18522 2150
rect 18282 2128 18578 2148
rect 17972 1958 18184 1986
rect 18156 800 18184 1958
rect 18616 800 18644 2246
rect 18984 800 19012 2246
rect 19352 1170 19380 2314
rect 19444 2292 19472 2808
rect 19536 2650 19564 3130
rect 19628 2922 19656 7754
rect 19720 5302 19748 8894
rect 19800 7540 19852 7546
rect 19800 7482 19852 7488
rect 19812 7410 19840 7482
rect 19800 7404 19852 7410
rect 19800 7346 19852 7352
rect 19800 6996 19852 7002
rect 19904 6984 19932 9608
rect 20088 8378 20116 12038
rect 20260 11620 20312 11626
rect 20260 11562 20312 11568
rect 20166 10296 20222 10305
rect 20166 10231 20222 10240
rect 20180 10033 20208 10231
rect 20166 10024 20222 10033
rect 20166 9959 20222 9968
rect 20168 9580 20220 9586
rect 20168 9522 20220 9528
rect 20180 9178 20208 9522
rect 20168 9172 20220 9178
rect 20168 9114 20220 9120
rect 19984 8356 20036 8362
rect 20088 8350 20208 8378
rect 19984 8298 20036 8304
rect 19996 8090 20024 8298
rect 20076 8288 20128 8294
rect 20076 8230 20128 8236
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 20088 7546 20116 8230
rect 20076 7540 20128 7546
rect 20076 7482 20128 7488
rect 20180 7274 20208 8350
rect 20272 8090 20300 11562
rect 20364 10538 20392 14350
rect 20548 13870 20576 18566
rect 20732 18426 20760 18770
rect 20720 18420 20772 18426
rect 20720 18362 20772 18368
rect 20732 17746 20760 18362
rect 20904 18148 20956 18154
rect 20904 18090 20956 18096
rect 20720 17740 20772 17746
rect 20720 17682 20772 17688
rect 20628 17672 20680 17678
rect 20628 17614 20680 17620
rect 20536 13864 20588 13870
rect 20536 13806 20588 13812
rect 20536 11688 20588 11694
rect 20536 11630 20588 11636
rect 20444 11212 20496 11218
rect 20444 11154 20496 11160
rect 20456 10674 20484 11154
rect 20444 10668 20496 10674
rect 20444 10610 20496 10616
rect 20352 10532 20404 10538
rect 20352 10474 20404 10480
rect 20444 10464 20496 10470
rect 20444 10406 20496 10412
rect 20352 10124 20404 10130
rect 20352 10066 20404 10072
rect 20364 9654 20392 10066
rect 20456 9722 20484 10406
rect 20444 9716 20496 9722
rect 20444 9658 20496 9664
rect 20352 9648 20404 9654
rect 20352 9590 20404 9596
rect 20444 8832 20496 8838
rect 20444 8774 20496 8780
rect 20260 8084 20312 8090
rect 20260 8026 20312 8032
rect 20076 7268 20128 7274
rect 20076 7210 20128 7216
rect 20168 7268 20220 7274
rect 20168 7210 20220 7216
rect 19984 7200 20036 7206
rect 19984 7142 20036 7148
rect 19852 6956 19932 6984
rect 19800 6938 19852 6944
rect 19996 6662 20024 7142
rect 20088 7002 20116 7210
rect 20076 6996 20128 7002
rect 20076 6938 20128 6944
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 19996 5846 20024 6598
rect 20076 6180 20128 6186
rect 20076 6122 20128 6128
rect 20088 5914 20116 6122
rect 20076 5908 20128 5914
rect 20076 5850 20128 5856
rect 19984 5840 20036 5846
rect 19984 5782 20036 5788
rect 20168 5772 20220 5778
rect 20168 5714 20220 5720
rect 20180 5370 20208 5714
rect 20168 5364 20220 5370
rect 20168 5306 20220 5312
rect 19708 5296 19760 5302
rect 19708 5238 19760 5244
rect 20076 5296 20128 5302
rect 20076 5238 20128 5244
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 19708 4684 19760 4690
rect 19708 4626 19760 4632
rect 19720 4282 19748 4626
rect 19996 4554 20024 4966
rect 19984 4548 20036 4554
rect 19984 4490 20036 4496
rect 19708 4276 19760 4282
rect 19708 4218 19760 4224
rect 19708 3936 19760 3942
rect 19708 3878 19760 3884
rect 19800 3936 19852 3942
rect 19984 3936 20036 3942
rect 19800 3878 19852 3884
rect 19982 3904 19984 3913
rect 20036 3904 20038 3913
rect 19720 3194 19748 3878
rect 19812 3738 19840 3878
rect 19982 3839 20038 3848
rect 19800 3732 19852 3738
rect 19800 3674 19852 3680
rect 19708 3188 19760 3194
rect 19708 3130 19760 3136
rect 19720 2972 19748 3130
rect 19982 3088 20038 3097
rect 19982 3023 20038 3032
rect 19996 2990 20024 3023
rect 20088 2990 20116 5238
rect 20272 3738 20300 8026
rect 20456 7342 20484 8774
rect 20352 7336 20404 7342
rect 20352 7278 20404 7284
rect 20444 7336 20496 7342
rect 20444 7278 20496 7284
rect 20364 6390 20392 7278
rect 20352 6384 20404 6390
rect 20352 6326 20404 6332
rect 20260 3732 20312 3738
rect 20260 3674 20312 3680
rect 20272 3058 20300 3674
rect 20364 3398 20392 6326
rect 20548 5846 20576 11630
rect 20536 5840 20588 5846
rect 20536 5782 20588 5788
rect 20640 4010 20668 17614
rect 20732 17338 20760 17682
rect 20720 17332 20772 17338
rect 20720 17274 20772 17280
rect 20812 16652 20864 16658
rect 20812 16594 20864 16600
rect 20824 15638 20852 16594
rect 20812 15632 20864 15638
rect 20812 15574 20864 15580
rect 20812 14952 20864 14958
rect 20812 14894 20864 14900
rect 20824 14550 20852 14894
rect 20812 14544 20864 14550
rect 20812 14486 20864 14492
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 20720 8288 20772 8294
rect 20720 8230 20772 8236
rect 20732 7818 20760 8230
rect 20720 7812 20772 7818
rect 20720 7754 20772 7760
rect 20824 7478 20852 9658
rect 20916 9518 20944 18090
rect 21284 17882 21312 19314
rect 22020 18902 22048 22200
rect 22388 20466 22416 22200
rect 22376 20460 22428 20466
rect 22376 20402 22428 20408
rect 22756 20330 22784 22200
rect 22744 20324 22796 20330
rect 22744 20266 22796 20272
rect 22008 18896 22060 18902
rect 21638 18864 21694 18873
rect 22008 18838 22060 18844
rect 21638 18799 21694 18808
rect 21454 18456 21510 18465
rect 21454 18391 21456 18400
rect 21508 18391 21510 18400
rect 21456 18362 21508 18368
rect 21272 17876 21324 17882
rect 21272 17818 21324 17824
rect 21548 17672 21600 17678
rect 21548 17614 21600 17620
rect 21362 17232 21418 17241
rect 21362 17167 21418 17176
rect 21272 16992 21324 16998
rect 21272 16934 21324 16940
rect 20994 16824 21050 16833
rect 20994 16759 21050 16768
rect 21008 16250 21036 16759
rect 20996 16244 21048 16250
rect 20996 16186 21048 16192
rect 21086 15872 21142 15881
rect 21086 15807 21142 15816
rect 21100 15706 21128 15807
rect 21088 15700 21140 15706
rect 21088 15642 21140 15648
rect 20994 15464 21050 15473
rect 20994 15399 21050 15408
rect 21008 15162 21036 15399
rect 20996 15156 21048 15162
rect 20996 15098 21048 15104
rect 21180 14816 21232 14822
rect 21180 14758 21232 14764
rect 21086 14648 21142 14657
rect 21086 14583 21088 14592
rect 21140 14583 21142 14592
rect 21088 14554 21140 14560
rect 21192 14550 21220 14758
rect 21180 14544 21232 14550
rect 21180 14486 21232 14492
rect 21284 14498 21312 16934
rect 21376 16250 21404 17167
rect 21454 16280 21510 16289
rect 21364 16244 21416 16250
rect 21454 16215 21510 16224
rect 21364 16186 21416 16192
rect 21468 15706 21496 16215
rect 21456 15700 21508 15706
rect 21456 15642 21508 15648
rect 21454 15056 21510 15065
rect 21560 15042 21588 17614
rect 21652 17338 21680 18799
rect 22006 17640 22062 17649
rect 22006 17575 22008 17584
rect 22060 17575 22062 17584
rect 22008 17546 22060 17552
rect 21640 17332 21692 17338
rect 21640 17274 21692 17280
rect 21560 15014 21680 15042
rect 21454 14991 21510 15000
rect 21468 14618 21496 14991
rect 21456 14612 21508 14618
rect 21456 14554 21508 14560
rect 21088 14476 21140 14482
rect 21284 14470 21588 14498
rect 21088 14418 21140 14424
rect 21100 14278 21128 14418
rect 21088 14272 21140 14278
rect 20994 14240 21050 14249
rect 21088 14214 21140 14220
rect 21456 14272 21508 14278
rect 21456 14214 21508 14220
rect 20994 14175 21050 14184
rect 21008 14074 21036 14175
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 21272 13864 21324 13870
rect 20994 13832 21050 13841
rect 21272 13806 21324 13812
rect 20994 13767 21050 13776
rect 21008 12986 21036 13767
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 21100 13433 21128 13466
rect 21086 13424 21142 13433
rect 21086 13359 21142 13368
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 20994 12472 21050 12481
rect 20994 12407 21050 12416
rect 21008 11898 21036 12407
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 21180 11688 21232 11694
rect 21180 11630 21232 11636
rect 21192 10674 21220 11630
rect 21180 10668 21232 10674
rect 21180 10610 21232 10616
rect 20904 9512 20956 9518
rect 20904 9454 20956 9460
rect 20904 9376 20956 9382
rect 20904 9318 20956 9324
rect 20916 8634 20944 9318
rect 20904 8628 20956 8634
rect 20904 8570 20956 8576
rect 21088 8492 21140 8498
rect 21088 8434 21140 8440
rect 21100 7886 21128 8434
rect 20904 7880 20956 7886
rect 20904 7822 20956 7828
rect 21088 7880 21140 7886
rect 21088 7822 21140 7828
rect 20812 7472 20864 7478
rect 20812 7414 20864 7420
rect 20916 7410 20944 7822
rect 21284 7562 21312 13806
rect 21362 12880 21418 12889
rect 21362 12815 21418 12824
rect 21376 11898 21404 12815
rect 21364 11892 21416 11898
rect 21364 11834 21416 11840
rect 21468 9722 21496 14214
rect 21456 9716 21508 9722
rect 21456 9658 21508 9664
rect 21456 8288 21508 8294
rect 21456 8230 21508 8236
rect 21008 7534 21312 7562
rect 20904 7404 20956 7410
rect 20904 7346 20956 7352
rect 20812 7336 20864 7342
rect 20812 7278 20864 7284
rect 20824 7206 20852 7278
rect 20720 7200 20772 7206
rect 20720 7142 20772 7148
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20732 4078 20760 7142
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 20628 4004 20680 4010
rect 20628 3946 20680 3952
rect 20352 3392 20404 3398
rect 20352 3334 20404 3340
rect 20364 3097 20392 3334
rect 20350 3088 20406 3097
rect 20260 3052 20312 3058
rect 20350 3023 20406 3032
rect 20260 2994 20312 3000
rect 19800 2984 19852 2990
rect 19720 2944 19800 2972
rect 19800 2926 19852 2932
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 20076 2984 20128 2990
rect 20272 2938 20300 2994
rect 20076 2926 20128 2932
rect 19616 2916 19668 2922
rect 19616 2858 19668 2864
rect 19892 2916 19944 2922
rect 19892 2858 19944 2864
rect 19800 2848 19852 2854
rect 19800 2790 19852 2796
rect 19524 2644 19576 2650
rect 19524 2586 19576 2592
rect 19524 2304 19576 2310
rect 19444 2264 19524 2292
rect 19524 2246 19576 2252
rect 19352 1142 19472 1170
rect 19444 800 19472 1142
rect 3790 232 3846 241
rect 3790 167 3846 176
rect 3882 0 3938 800
rect 4342 0 4398 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5630 0 5686 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7286 0 7342 800
rect 7654 0 7710 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8942 0 8998 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10230 0 10286 800
rect 10598 0 10654 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11886 0 11942 800
rect 12254 0 12310 800
rect 12714 0 12770 800
rect 13082 0 13138 800
rect 13542 0 13598 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14830 0 14886 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16026 0 16082 800
rect 16486 0 16542 800
rect 16854 0 16910 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18142 0 18198 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19430 0 19486 800
rect 19536 649 19564 2246
rect 19812 800 19840 2790
rect 19904 2310 19932 2858
rect 20088 2650 20116 2926
rect 20180 2910 20300 2938
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 19892 2304 19944 2310
rect 20180 2281 20208 2910
rect 20260 2848 20312 2854
rect 20260 2790 20312 2796
rect 20628 2848 20680 2854
rect 20628 2790 20680 2796
rect 19892 2246 19944 2252
rect 20166 2272 20222 2281
rect 19904 1465 19932 2246
rect 20166 2207 20222 2216
rect 19890 1456 19946 1465
rect 19890 1391 19946 1400
rect 20272 800 20300 2790
rect 20640 800 20668 2790
rect 19522 640 19578 649
rect 19522 575 19578 584
rect 19798 0 19854 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20824 241 20852 7142
rect 20916 6798 20944 7346
rect 20904 6792 20956 6798
rect 20904 6734 20956 6740
rect 20916 6458 20944 6734
rect 20904 6452 20956 6458
rect 20904 6394 20956 6400
rect 20904 3120 20956 3126
rect 20904 3062 20956 3068
rect 20916 1873 20944 3062
rect 20902 1864 20958 1873
rect 20902 1799 20958 1808
rect 21008 898 21036 7534
rect 21088 6724 21140 6730
rect 21088 6666 21140 6672
rect 21100 6390 21128 6666
rect 21088 6384 21140 6390
rect 21088 6326 21140 6332
rect 21468 5137 21496 8230
rect 21086 5128 21142 5137
rect 21086 5063 21142 5072
rect 21454 5128 21510 5137
rect 21454 5063 21510 5072
rect 21100 1057 21128 5063
rect 21560 4146 21588 14470
rect 21652 9654 21680 15014
rect 22006 12064 22062 12073
rect 22006 11999 22008 12008
rect 22060 11999 22062 12008
rect 22008 11970 22060 11976
rect 21640 9648 21692 9654
rect 21640 9590 21692 9596
rect 21824 9648 21876 9654
rect 21824 9590 21876 9596
rect 21548 4140 21600 4146
rect 21548 4082 21600 4088
rect 21086 1048 21142 1057
rect 21086 983 21142 992
rect 21836 921 21864 9590
rect 21916 9512 21968 9518
rect 21916 9454 21968 9460
rect 21454 912 21510 921
rect 21008 870 21128 898
rect 21100 800 21128 870
rect 21454 847 21510 856
rect 21822 912 21878 921
rect 21822 847 21878 856
rect 21468 800 21496 847
rect 21928 800 21956 9454
rect 22008 5568 22060 5574
rect 22008 5510 22060 5516
rect 22020 2689 22048 5510
rect 22744 4140 22796 4146
rect 22744 4082 22796 4088
rect 22284 4004 22336 4010
rect 22284 3946 22336 3952
rect 22006 2680 22062 2689
rect 22006 2615 22062 2624
rect 22296 800 22324 3946
rect 22756 800 22784 4082
rect 20810 232 20866 241
rect 20810 167 20866 176
rect 21086 0 21142 800
rect 21454 0 21510 800
rect 21914 0 21970 800
rect 22282 0 22338 800
rect 22742 0 22798 800
<< via2 >>
rect 3514 22616 3570 22672
rect 1950 20168 2006 20224
rect 1858 19624 1914 19680
rect 2134 18944 2190 19000
rect 1306 18536 1362 18592
rect 1582 18400 1638 18456
rect 1950 18028 1952 18048
rect 1952 18028 2004 18048
rect 2004 18028 2006 18048
rect 1950 17992 2006 18028
rect 2594 19216 2650 19272
rect 2502 18572 2504 18592
rect 2504 18572 2556 18592
rect 2556 18572 2558 18592
rect 2502 18536 2558 18572
rect 2962 19080 3018 19136
rect 2778 18808 2834 18864
rect 2410 17720 2466 17776
rect 1674 17584 1730 17640
rect 1582 17176 1638 17232
rect 1766 16088 1822 16144
rect 1950 15852 1952 15872
rect 1952 15852 2004 15872
rect 2004 15852 2006 15872
rect 1950 15816 2006 15852
rect 1766 15036 1768 15056
rect 1768 15036 1820 15056
rect 1820 15036 1822 15056
rect 1766 15000 1822 15036
rect 1858 14612 1914 14648
rect 1858 14592 1860 14612
rect 1860 14592 1912 14612
rect 1912 14592 1914 14612
rect 2042 14592 2098 14648
rect 1582 14320 1638 14376
rect 1766 14184 1822 14240
rect 1674 12824 1730 12880
rect 3146 18536 3202 18592
rect 2870 18028 2872 18048
rect 2872 18028 2924 18048
rect 2924 18028 2926 18048
rect 2870 17992 2926 18028
rect 2778 16904 2834 16960
rect 2778 16768 2834 16824
rect 2318 16244 2374 16280
rect 2318 16224 2320 16244
rect 2320 16224 2372 16244
rect 2372 16224 2374 16244
rect 3422 21800 3478 21856
rect 3790 22208 3846 22264
rect 3514 18672 3570 18728
rect 3422 18128 3478 18184
rect 3146 17448 3202 17504
rect 19154 22208 19210 22264
rect 3698 21392 3754 21448
rect 3882 20576 3938 20632
rect 3882 19216 3938 19272
rect 3790 18808 3846 18864
rect 3698 18264 3754 18320
rect 2410 13368 2466 13424
rect 1582 12008 1638 12064
rect 1398 9832 1454 9888
rect 1766 2216 1822 2272
rect 2778 13776 2834 13832
rect 3054 13252 3110 13288
rect 3054 13232 3056 13252
rect 3056 13232 3108 13252
rect 3108 13232 3110 13252
rect 3146 12416 3202 12472
rect 3790 16088 3846 16144
rect 3330 11464 3386 11520
rect 3698 15544 3754 15600
rect 3790 15408 3846 15464
rect 2870 7656 2926 7712
rect 2870 5616 2926 5672
rect 2962 3032 3018 3088
rect 2226 2760 2282 2816
rect 1306 1400 1362 1456
rect 2134 1808 2190 1864
rect 2778 2624 2834 2680
rect 3422 8880 3478 8936
rect 4066 20984 4122 21040
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4581 20698 4637 20700
rect 4661 20698 4717 20700
rect 4421 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4581 20646 4627 20698
rect 4627 20646 4637 20698
rect 4661 20646 4691 20698
rect 4691 20646 4717 20698
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4581 20644 4637 20646
rect 4661 20644 4717 20646
rect 4158 18944 4214 19000
rect 4158 18420 4214 18456
rect 4158 18400 4160 18420
rect 4160 18400 4212 18420
rect 4212 18400 4214 18420
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4581 19610 4637 19612
rect 4661 19610 4717 19612
rect 4421 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4581 19558 4627 19610
rect 4627 19558 4637 19610
rect 4661 19558 4691 19610
rect 4691 19558 4717 19610
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4581 19556 4637 19558
rect 4661 19556 4717 19558
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4581 18522 4637 18524
rect 4661 18522 4717 18524
rect 4421 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4581 18470 4627 18522
rect 4627 18470 4637 18522
rect 4661 18470 4691 18522
rect 4691 18470 4717 18522
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 4581 18468 4637 18470
rect 4661 18468 4717 18470
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4581 17434 4637 17436
rect 4661 17434 4717 17436
rect 4421 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4581 17382 4627 17434
rect 4627 17382 4637 17434
rect 4661 17382 4691 17434
rect 4691 17382 4717 17434
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 4581 17380 4637 17382
rect 4661 17380 4717 17382
rect 3974 14612 4030 14648
rect 3974 14592 3976 14612
rect 3976 14592 4028 14612
rect 4028 14592 4030 14612
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4581 16346 4637 16348
rect 4661 16346 4717 16348
rect 4421 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4581 16294 4627 16346
rect 4627 16294 4637 16346
rect 4661 16294 4691 16346
rect 4691 16294 4717 16346
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 4581 16292 4637 16294
rect 4661 16292 4717 16294
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4581 15258 4637 15260
rect 4661 15258 4717 15260
rect 4421 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4581 15206 4627 15258
rect 4627 15206 4637 15258
rect 4661 15206 4691 15258
rect 4691 15206 4717 15258
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 4581 15204 4637 15206
rect 4661 15204 4717 15206
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4581 14170 4637 14172
rect 4661 14170 4717 14172
rect 4421 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4581 14118 4627 14170
rect 4627 14118 4637 14170
rect 4661 14118 4691 14170
rect 4691 14118 4717 14170
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 4581 14116 4637 14118
rect 4661 14116 4717 14118
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4581 13082 4637 13084
rect 4661 13082 4717 13084
rect 4421 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4581 13030 4627 13082
rect 4627 13030 4637 13082
rect 4661 13030 4691 13082
rect 4691 13030 4717 13082
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4581 13028 4637 13030
rect 4661 13028 4717 13030
rect 3882 11872 3938 11928
rect 3882 11600 3938 11656
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4581 11994 4637 11996
rect 4661 11994 4717 11996
rect 4421 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4581 11942 4627 11994
rect 4627 11942 4637 11994
rect 4661 11942 4691 11994
rect 4691 11942 4717 11994
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 4581 11940 4637 11942
rect 4661 11940 4717 11942
rect 3606 9424 3662 9480
rect 4158 9968 4214 10024
rect 3790 7656 3846 7712
rect 4066 7792 4122 7848
rect 3974 7384 4030 7440
rect 5078 12008 5134 12064
rect 4710 11328 4766 11384
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4581 10906 4637 10908
rect 4661 10906 4717 10908
rect 4421 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4581 10854 4627 10906
rect 4627 10854 4637 10906
rect 4661 10854 4691 10906
rect 4691 10854 4717 10906
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 4581 10852 4637 10854
rect 4661 10852 4717 10854
rect 5078 11328 5134 11384
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4581 9818 4637 9820
rect 4661 9818 4717 9820
rect 4421 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4581 9766 4627 9818
rect 4627 9766 4637 9818
rect 4661 9766 4691 9818
rect 4691 9766 4717 9818
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 4581 9764 4637 9766
rect 4661 9764 4717 9766
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4581 8730 4637 8732
rect 4661 8730 4717 8732
rect 4421 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4581 8678 4627 8730
rect 4627 8678 4637 8730
rect 4661 8678 4691 8730
rect 4691 8678 4717 8730
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4581 8676 4637 8678
rect 4661 8676 4717 8678
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4581 7642 4637 7644
rect 4661 7642 4717 7644
rect 4421 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4581 7590 4627 7642
rect 4627 7590 4637 7642
rect 4661 7590 4691 7642
rect 4691 7590 4717 7642
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 4581 7588 4637 7590
rect 4661 7588 4717 7590
rect 4066 6432 4122 6488
rect 3974 6024 4030 6080
rect 3146 1808 3202 1864
rect 3606 992 3662 1048
rect 2962 584 3018 640
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4581 6554 4637 6556
rect 4661 6554 4717 6556
rect 4421 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4581 6502 4627 6554
rect 4627 6502 4637 6554
rect 4661 6502 4691 6554
rect 4691 6502 4717 6554
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 4581 6500 4637 6502
rect 4661 6500 4717 6502
rect 4250 5752 4306 5808
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4581 5466 4637 5468
rect 4661 5466 4717 5468
rect 4421 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4581 5414 4627 5466
rect 4627 5414 4637 5466
rect 4661 5414 4691 5466
rect 4691 5414 4717 5466
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4581 5412 4637 5414
rect 4661 5412 4717 5414
rect 4250 4276 4306 4312
rect 4250 4256 4252 4276
rect 4252 4256 4304 4276
rect 4304 4256 4306 4276
rect 5354 14900 5356 14920
rect 5356 14900 5408 14920
rect 5408 14900 5410 14920
rect 5354 14864 5410 14900
rect 5262 12280 5318 12336
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4581 4378 4637 4380
rect 4661 4378 4717 4380
rect 4421 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4581 4326 4627 4378
rect 4627 4326 4637 4378
rect 4661 4326 4691 4378
rect 4691 4326 4717 4378
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4581 4324 4637 4326
rect 4661 4324 4717 4326
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4581 3290 4637 3292
rect 4661 3290 4717 3292
rect 4421 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4581 3238 4627 3290
rect 4627 3238 4637 3290
rect 4661 3238 4691 3290
rect 4691 3238 4717 3290
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 4581 3236 4637 3238
rect 4661 3236 4717 3238
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4581 2202 4637 2204
rect 4661 2202 4717 2204
rect 4421 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4581 2150 4627 2202
rect 4627 2150 4637 2202
rect 4661 2150 4691 2202
rect 4691 2150 4717 2202
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 4581 2148 4637 2150
rect 4661 2148 4717 2150
rect 5170 6432 5226 6488
rect 5906 18964 5962 19000
rect 5906 18944 5908 18964
rect 5908 18944 5960 18964
rect 5960 18944 5962 18964
rect 5906 17176 5962 17232
rect 6274 18400 6330 18456
rect 6090 17040 6146 17096
rect 6274 14864 6330 14920
rect 5446 11328 5502 11384
rect 5722 12588 5724 12608
rect 5724 12588 5776 12608
rect 5776 12588 5778 12608
rect 5722 12552 5778 12588
rect 6090 11600 6146 11656
rect 5906 10784 5962 10840
rect 6366 12280 6422 12336
rect 7102 18964 7158 19000
rect 7102 18944 7104 18964
rect 7104 18944 7156 18964
rect 7156 18944 7158 18964
rect 7102 18400 7158 18456
rect 6550 17584 6606 17640
rect 6550 17196 6606 17232
rect 6550 17176 6552 17196
rect 6552 17176 6604 17196
rect 6604 17176 6606 17196
rect 6918 16904 6974 16960
rect 6550 13640 6606 13696
rect 6550 13268 6552 13288
rect 6552 13268 6604 13288
rect 6604 13268 6606 13288
rect 6550 13232 6606 13268
rect 6642 12824 6698 12880
rect 6458 11056 6514 11112
rect 6458 10920 6514 10976
rect 5906 10376 5962 10432
rect 5998 10240 6054 10296
rect 5722 9832 5778 9888
rect 5722 9696 5778 9752
rect 5354 7928 5410 7984
rect 5630 7792 5686 7848
rect 5262 4140 5318 4176
rect 5446 4256 5502 4312
rect 5262 4120 5264 4140
rect 5264 4120 5316 4140
rect 5316 4120 5318 4140
rect 6090 9696 6146 9752
rect 6366 9696 6422 9752
rect 6090 8608 6146 8664
rect 5722 4528 5778 4584
rect 6274 7384 6330 7440
rect 6458 6976 6514 7032
rect 6366 6296 6422 6352
rect 6274 3576 6330 3632
rect 5998 3304 6054 3360
rect 6458 3440 6514 3496
rect 6090 3168 6146 3224
rect 6642 11348 6698 11384
rect 6642 11328 6644 11348
rect 6644 11328 6696 11348
rect 6696 11328 6698 11348
rect 7886 20154 7942 20156
rect 7966 20154 8022 20156
rect 8046 20154 8102 20156
rect 8126 20154 8182 20156
rect 7886 20102 7912 20154
rect 7912 20102 7942 20154
rect 7966 20102 7976 20154
rect 7976 20102 8022 20154
rect 8046 20102 8092 20154
rect 8092 20102 8102 20154
rect 8126 20102 8156 20154
rect 8156 20102 8182 20154
rect 7886 20100 7942 20102
rect 7966 20100 8022 20102
rect 8046 20100 8102 20102
rect 8126 20100 8182 20102
rect 7562 19080 7618 19136
rect 8206 19352 8262 19408
rect 8574 19352 8630 19408
rect 7886 19066 7942 19068
rect 7966 19066 8022 19068
rect 8046 19066 8102 19068
rect 8126 19066 8182 19068
rect 7886 19014 7912 19066
rect 7912 19014 7942 19066
rect 7966 19014 7976 19066
rect 7976 19014 8022 19066
rect 8046 19014 8092 19066
rect 8092 19014 8102 19066
rect 8126 19014 8156 19066
rect 8156 19014 8182 19066
rect 7886 19012 7942 19014
rect 7966 19012 8022 19014
rect 8046 19012 8102 19014
rect 8126 19012 8182 19014
rect 7654 18536 7710 18592
rect 7562 17992 7618 18048
rect 7886 17978 7942 17980
rect 7966 17978 8022 17980
rect 8046 17978 8102 17980
rect 8126 17978 8182 17980
rect 7886 17926 7912 17978
rect 7912 17926 7942 17978
rect 7966 17926 7976 17978
rect 7976 17926 8022 17978
rect 8046 17926 8092 17978
rect 8092 17926 8102 17978
rect 8126 17926 8156 17978
rect 8156 17926 8182 17978
rect 7886 17924 7942 17926
rect 7966 17924 8022 17926
rect 8046 17924 8102 17926
rect 8126 17924 8182 17926
rect 8666 18400 8722 18456
rect 7654 17484 7656 17504
rect 7656 17484 7708 17504
rect 7708 17484 7710 17504
rect 7654 17448 7710 17484
rect 8206 17312 8262 17368
rect 7194 13504 7250 13560
rect 6918 11892 6974 11928
rect 6918 11872 6920 11892
rect 6920 11872 6972 11892
rect 6972 11872 6974 11892
rect 7102 11736 7158 11792
rect 6826 10512 6882 10568
rect 6642 8880 6698 8936
rect 6642 6704 6698 6760
rect 7286 11464 7342 11520
rect 7286 11328 7342 11384
rect 8206 17040 8262 17096
rect 7886 16890 7942 16892
rect 7966 16890 8022 16892
rect 8046 16890 8102 16892
rect 8126 16890 8182 16892
rect 7886 16838 7912 16890
rect 7912 16838 7942 16890
rect 7966 16838 7976 16890
rect 7976 16838 8022 16890
rect 8046 16838 8092 16890
rect 8092 16838 8102 16890
rect 8126 16838 8156 16890
rect 8156 16838 8182 16890
rect 7886 16836 7942 16838
rect 7966 16836 8022 16838
rect 8046 16836 8102 16838
rect 8126 16836 8182 16838
rect 7886 15802 7942 15804
rect 7966 15802 8022 15804
rect 8046 15802 8102 15804
rect 8126 15802 8182 15804
rect 7886 15750 7912 15802
rect 7912 15750 7942 15802
rect 7966 15750 7976 15802
rect 7976 15750 8022 15802
rect 8046 15750 8092 15802
rect 8092 15750 8102 15802
rect 8126 15750 8156 15802
rect 8156 15750 8182 15802
rect 7886 15748 7942 15750
rect 7966 15748 8022 15750
rect 8046 15748 8102 15750
rect 8126 15748 8182 15750
rect 8114 15564 8170 15600
rect 8114 15544 8116 15564
rect 8116 15544 8168 15564
rect 8168 15544 8170 15564
rect 7930 14864 7986 14920
rect 7886 14714 7942 14716
rect 7966 14714 8022 14716
rect 8046 14714 8102 14716
rect 8126 14714 8182 14716
rect 7886 14662 7912 14714
rect 7912 14662 7942 14714
rect 7966 14662 7976 14714
rect 7976 14662 8022 14714
rect 8046 14662 8092 14714
rect 8092 14662 8102 14714
rect 8126 14662 8156 14714
rect 8156 14662 8182 14714
rect 7886 14660 7942 14662
rect 7966 14660 8022 14662
rect 8046 14660 8102 14662
rect 8126 14660 8182 14662
rect 8114 14048 8170 14104
rect 8114 13812 8116 13832
rect 8116 13812 8168 13832
rect 8168 13812 8170 13832
rect 8114 13776 8170 13812
rect 7886 13626 7942 13628
rect 7966 13626 8022 13628
rect 8046 13626 8102 13628
rect 8126 13626 8182 13628
rect 7886 13574 7912 13626
rect 7912 13574 7942 13626
rect 7966 13574 7976 13626
rect 7976 13574 8022 13626
rect 8046 13574 8092 13626
rect 8092 13574 8102 13626
rect 8126 13574 8156 13626
rect 8156 13574 8182 13626
rect 7886 13572 7942 13574
rect 7966 13572 8022 13574
rect 8046 13572 8102 13574
rect 8126 13572 8182 13574
rect 7654 11328 7710 11384
rect 7470 11056 7526 11112
rect 7470 10376 7526 10432
rect 7470 8880 7526 8936
rect 8758 15444 8760 15464
rect 8760 15444 8812 15464
rect 8812 15444 8814 15464
rect 8758 15408 8814 15444
rect 8298 13368 8354 13424
rect 7886 12538 7942 12540
rect 7966 12538 8022 12540
rect 8046 12538 8102 12540
rect 8126 12538 8182 12540
rect 7886 12486 7912 12538
rect 7912 12486 7942 12538
rect 7966 12486 7976 12538
rect 7976 12486 8022 12538
rect 8046 12486 8092 12538
rect 8092 12486 8102 12538
rect 8126 12486 8156 12538
rect 8156 12486 8182 12538
rect 7886 12484 7942 12486
rect 7966 12484 8022 12486
rect 8046 12484 8102 12486
rect 8126 12484 8182 12486
rect 8666 14048 8722 14104
rect 8942 16360 8998 16416
rect 8942 16088 8998 16144
rect 8850 14864 8906 14920
rect 9126 16224 9182 16280
rect 9310 15580 9312 15600
rect 9312 15580 9364 15600
rect 9364 15580 9366 15600
rect 9310 15544 9366 15580
rect 9218 14864 9274 14920
rect 9494 17212 9496 17232
rect 9496 17212 9548 17232
rect 9548 17212 9550 17232
rect 9494 17176 9550 17212
rect 8758 13676 8760 13696
rect 8760 13676 8812 13696
rect 8812 13676 8814 13696
rect 8758 13640 8814 13676
rect 8850 13504 8906 13560
rect 8298 12824 8354 12880
rect 7886 11450 7942 11452
rect 7966 11450 8022 11452
rect 8046 11450 8102 11452
rect 8126 11450 8182 11452
rect 7886 11398 7912 11450
rect 7912 11398 7942 11450
rect 7966 11398 7976 11450
rect 7976 11398 8022 11450
rect 8046 11398 8092 11450
rect 8092 11398 8102 11450
rect 8126 11398 8156 11450
rect 8156 11398 8182 11450
rect 7886 11396 7942 11398
rect 7966 11396 8022 11398
rect 8046 11396 8102 11398
rect 8126 11396 8182 11398
rect 7886 10362 7942 10364
rect 7966 10362 8022 10364
rect 8046 10362 8102 10364
rect 8126 10362 8182 10364
rect 7886 10310 7912 10362
rect 7912 10310 7942 10362
rect 7966 10310 7976 10362
rect 7976 10310 8022 10362
rect 8046 10310 8092 10362
rect 8092 10310 8102 10362
rect 8126 10310 8156 10362
rect 8156 10310 8182 10362
rect 7886 10308 7942 10310
rect 7966 10308 8022 10310
rect 8046 10308 8102 10310
rect 8126 10308 8182 10310
rect 8482 12724 8484 12744
rect 8484 12724 8536 12744
rect 8536 12724 8538 12744
rect 8482 12688 8538 12724
rect 8482 12436 8538 12472
rect 8482 12416 8484 12436
rect 8484 12416 8536 12436
rect 8536 12416 8538 12436
rect 8482 10648 8538 10704
rect 8942 13232 8998 13288
rect 8666 11600 8722 11656
rect 8666 10804 8722 10840
rect 8666 10784 8668 10804
rect 8668 10784 8720 10804
rect 8720 10784 8722 10804
rect 9034 13132 9036 13152
rect 9036 13132 9088 13152
rect 9088 13132 9090 13152
rect 9034 13096 9090 13132
rect 9126 12844 9182 12880
rect 9126 12824 9128 12844
rect 9128 12824 9180 12844
rect 9180 12824 9182 12844
rect 8850 10784 8906 10840
rect 8758 10648 8814 10704
rect 7930 9444 7986 9480
rect 7930 9424 7932 9444
rect 7932 9424 7984 9444
rect 7984 9424 7986 9444
rect 7102 6840 7158 6896
rect 7010 5480 7066 5536
rect 7102 3712 7158 3768
rect 7378 6432 7434 6488
rect 7378 6160 7434 6216
rect 7286 5652 7288 5672
rect 7288 5652 7340 5672
rect 7340 5652 7342 5672
rect 7286 5616 7342 5652
rect 7286 5344 7342 5400
rect 7654 8200 7710 8256
rect 7562 7384 7618 7440
rect 7470 4800 7526 4856
rect 7886 9274 7942 9276
rect 7966 9274 8022 9276
rect 8046 9274 8102 9276
rect 8126 9274 8182 9276
rect 7886 9222 7912 9274
rect 7912 9222 7942 9274
rect 7966 9222 7976 9274
rect 7976 9222 8022 9274
rect 8046 9222 8092 9274
rect 8092 9222 8102 9274
rect 8126 9222 8156 9274
rect 8156 9222 8182 9274
rect 7886 9220 7942 9222
rect 7966 9220 8022 9222
rect 8046 9220 8102 9222
rect 8126 9220 8182 9222
rect 8298 9696 8354 9752
rect 8298 9288 8354 9344
rect 7930 8336 7986 8392
rect 8206 9036 8262 9072
rect 8206 9016 8208 9036
rect 8208 9016 8260 9036
rect 8260 9016 8262 9036
rect 7886 8186 7942 8188
rect 7966 8186 8022 8188
rect 8046 8186 8102 8188
rect 8126 8186 8182 8188
rect 7886 8134 7912 8186
rect 7912 8134 7942 8186
rect 7966 8134 7976 8186
rect 7976 8134 8022 8186
rect 8046 8134 8092 8186
rect 8092 8134 8102 8186
rect 8126 8134 8156 8186
rect 8156 8134 8182 8186
rect 7886 8132 7942 8134
rect 7966 8132 8022 8134
rect 8046 8132 8102 8134
rect 8126 8132 8182 8134
rect 8390 8200 8446 8256
rect 7886 7098 7942 7100
rect 7966 7098 8022 7100
rect 8046 7098 8102 7100
rect 8126 7098 8182 7100
rect 7886 7046 7912 7098
rect 7912 7046 7942 7098
rect 7966 7046 7976 7098
rect 7976 7046 8022 7098
rect 8046 7046 8092 7098
rect 8092 7046 8102 7098
rect 8126 7046 8156 7098
rect 8156 7046 8182 7098
rect 7886 7044 7942 7046
rect 7966 7044 8022 7046
rect 8046 7044 8102 7046
rect 8126 7044 8182 7046
rect 8022 6840 8078 6896
rect 7838 6740 7840 6760
rect 7840 6740 7892 6760
rect 7892 6740 7894 6760
rect 7838 6704 7894 6740
rect 7838 6568 7894 6624
rect 8758 10240 8814 10296
rect 8942 10376 8998 10432
rect 8942 9696 8998 9752
rect 9034 9152 9090 9208
rect 8574 7656 8630 7712
rect 8114 6296 8170 6352
rect 7886 6010 7942 6012
rect 7966 6010 8022 6012
rect 8046 6010 8102 6012
rect 8126 6010 8182 6012
rect 7886 5958 7912 6010
rect 7912 5958 7942 6010
rect 7966 5958 7976 6010
rect 7976 5958 8022 6010
rect 8046 5958 8092 6010
rect 8092 5958 8102 6010
rect 8126 5958 8156 6010
rect 8156 5958 8182 6010
rect 7886 5956 7942 5958
rect 7966 5956 8022 5958
rect 8046 5956 8102 5958
rect 8126 5956 8182 5958
rect 7654 4800 7710 4856
rect 7886 4922 7942 4924
rect 7966 4922 8022 4924
rect 8046 4922 8102 4924
rect 8126 4922 8182 4924
rect 7886 4870 7912 4922
rect 7912 4870 7942 4922
rect 7966 4870 7976 4922
rect 7976 4870 8022 4922
rect 8046 4870 8092 4922
rect 8092 4870 8102 4922
rect 8126 4870 8156 4922
rect 8156 4870 8182 4922
rect 7886 4868 7942 4870
rect 7966 4868 8022 4870
rect 8046 4868 8102 4870
rect 8126 4868 8182 4870
rect 8574 5908 8630 5944
rect 8574 5888 8576 5908
rect 8576 5888 8628 5908
rect 8628 5888 8630 5908
rect 7886 3834 7942 3836
rect 7966 3834 8022 3836
rect 8046 3834 8102 3836
rect 8126 3834 8182 3836
rect 7886 3782 7912 3834
rect 7912 3782 7942 3834
rect 7966 3782 7976 3834
rect 7976 3782 8022 3834
rect 8046 3782 8092 3834
rect 8092 3782 8102 3834
rect 8126 3782 8156 3834
rect 8156 3782 8182 3834
rect 7886 3780 7942 3782
rect 7966 3780 8022 3782
rect 8046 3780 8102 3782
rect 8126 3780 8182 3782
rect 8298 3440 8354 3496
rect 7746 3032 7802 3088
rect 7746 2760 7802 2816
rect 7886 2746 7942 2748
rect 7966 2746 8022 2748
rect 8046 2746 8102 2748
rect 8126 2746 8182 2748
rect 7886 2694 7912 2746
rect 7912 2694 7942 2746
rect 7966 2694 7976 2746
rect 7976 2694 8022 2746
rect 8046 2694 8092 2746
rect 8092 2694 8102 2746
rect 8126 2694 8156 2746
rect 8156 2694 8182 2746
rect 7886 2692 7942 2694
rect 7966 2692 8022 2694
rect 8046 2692 8102 2694
rect 8126 2692 8182 2694
rect 8482 4664 8538 4720
rect 8942 8084 8998 8120
rect 8942 8064 8944 8084
rect 8944 8064 8996 8084
rect 8996 8064 8998 8084
rect 8574 4256 8630 4312
rect 8574 3848 8630 3904
rect 8574 3612 8576 3632
rect 8576 3612 8628 3632
rect 8628 3612 8630 3632
rect 8574 3576 8630 3612
rect 8482 2760 8538 2816
rect 9494 13524 9550 13560
rect 9494 13504 9496 13524
rect 9496 13504 9548 13524
rect 9548 13504 9550 13524
rect 9310 13232 9366 13288
rect 9310 12824 9366 12880
rect 9310 12552 9366 12608
rect 9402 12280 9458 12336
rect 9678 17076 9680 17096
rect 9680 17076 9732 17096
rect 9732 17076 9734 17096
rect 9678 17040 9734 17076
rect 9862 18944 9918 19000
rect 9862 17992 9918 18048
rect 9862 17196 9918 17232
rect 9862 17176 9864 17196
rect 9864 17176 9916 17196
rect 9916 17176 9918 17196
rect 10230 15544 10286 15600
rect 10138 14864 10194 14920
rect 10046 14048 10102 14104
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11378 20698
rect 11378 20646 11408 20698
rect 11432 20646 11442 20698
rect 11442 20646 11488 20698
rect 11512 20646 11558 20698
rect 11558 20646 11568 20698
rect 11592 20646 11622 20698
rect 11622 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11378 19610
rect 11378 19558 11408 19610
rect 11432 19558 11442 19610
rect 11442 19558 11488 19610
rect 11512 19558 11558 19610
rect 11558 19558 11568 19610
rect 11592 19558 11622 19610
rect 11622 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 10506 16768 10562 16824
rect 10414 14764 10416 14784
rect 10416 14764 10468 14784
rect 10468 14764 10470 14784
rect 10414 14728 10470 14764
rect 10322 14592 10378 14648
rect 11334 18944 11390 19000
rect 11058 18536 11114 18592
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11378 18522
rect 11378 18470 11408 18522
rect 11432 18470 11442 18522
rect 11442 18470 11488 18522
rect 11512 18470 11558 18522
rect 11558 18470 11568 18522
rect 11592 18470 11622 18522
rect 11622 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 10966 17312 11022 17368
rect 9954 13776 10010 13832
rect 10138 13504 10194 13560
rect 11242 17740 11298 17776
rect 11242 17720 11244 17740
rect 11244 17720 11296 17740
rect 11296 17720 11298 17740
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11334 16516 11390 16552
rect 11334 16496 11336 16516
rect 11336 16496 11388 16516
rect 11388 16496 11390 16516
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 10506 13232 10562 13288
rect 10690 12824 10746 12880
rect 10138 12280 10194 12336
rect 9218 10104 9274 10160
rect 9218 9832 9274 9888
rect 9310 9696 9366 9752
rect 9770 11328 9826 11384
rect 10138 11328 10194 11384
rect 9770 10376 9826 10432
rect 9310 9152 9366 9208
rect 9126 5752 9182 5808
rect 9034 5652 9036 5672
rect 9036 5652 9088 5672
rect 9088 5652 9090 5672
rect 9034 5616 9090 5652
rect 8942 3304 8998 3360
rect 8942 3032 8998 3088
rect 9218 4800 9274 4856
rect 9126 4256 9182 4312
rect 9494 7828 9496 7848
rect 9496 7828 9548 7848
rect 9548 7828 9550 7848
rect 9494 7792 9550 7828
rect 9586 7384 9642 7440
rect 9402 6568 9458 6624
rect 10138 8336 10194 8392
rect 9586 5516 9588 5536
rect 9588 5516 9640 5536
rect 9640 5516 9642 5536
rect 9586 5480 9642 5516
rect 9678 4972 9680 4992
rect 9680 4972 9732 4992
rect 9732 4972 9734 4992
rect 9678 4936 9734 4972
rect 9586 4548 9642 4584
rect 9586 4528 9588 4548
rect 9588 4528 9640 4548
rect 9640 4528 9642 4548
rect 9402 3440 9458 3496
rect 9218 3168 9274 3224
rect 9034 2916 9090 2952
rect 9034 2896 9036 2916
rect 9036 2896 9088 2916
rect 9088 2896 9090 2916
rect 9126 2352 9182 2408
rect 9402 2644 9458 2680
rect 9402 2624 9404 2644
rect 9404 2624 9456 2644
rect 9456 2624 9458 2644
rect 10046 2896 10102 2952
rect 10506 11736 10562 11792
rect 10414 11192 10470 11248
rect 10506 10648 10562 10704
rect 10414 9696 10470 9752
rect 10690 9832 10746 9888
rect 10598 8336 10654 8392
rect 10414 7792 10470 7848
rect 10414 6976 10470 7032
rect 11334 14456 11390 14512
rect 12622 17992 12678 18048
rect 11978 15816 12034 15872
rect 12162 15544 12218 15600
rect 11702 14320 11758 14376
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11610 13796 11666 13832
rect 11610 13776 11612 13796
rect 11612 13776 11664 13796
rect 11664 13776 11666 13796
rect 11610 13232 11666 13288
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 10874 11192 10930 11248
rect 10874 10784 10930 10840
rect 11426 12552 11482 12608
rect 11886 12280 11942 12336
rect 11426 12144 11482 12200
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 12070 14184 12126 14240
rect 11978 11872 12034 11928
rect 12254 14048 12310 14104
rect 12162 11872 12218 11928
rect 11150 10376 11206 10432
rect 11058 8608 11114 8664
rect 10966 8356 11022 8392
rect 10966 8336 10968 8356
rect 10968 8336 11020 8356
rect 11020 8336 11022 8356
rect 10874 7384 10930 7440
rect 10690 6704 10746 6760
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11518 10376 11574 10432
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11242 8880 11298 8936
rect 11426 8880 11482 8936
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11242 7792 11298 7848
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 10690 5752 10746 5808
rect 10414 4256 10470 4312
rect 10322 3848 10378 3904
rect 10230 3576 10286 3632
rect 10230 3032 10286 3088
rect 10322 2896 10378 2952
rect 10690 3476 10692 3496
rect 10692 3476 10744 3496
rect 10744 3476 10746 3496
rect 10690 3440 10746 3476
rect 10966 4120 11022 4176
rect 10874 3304 10930 3360
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11426 6024 11482 6080
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 12070 11056 12126 11112
rect 12070 10784 12126 10840
rect 12070 10376 12126 10432
rect 11886 10124 11942 10160
rect 11886 10104 11888 10124
rect 11888 10104 11940 10124
rect 11940 10104 11942 10124
rect 11886 9696 11942 9752
rect 13174 17584 13230 17640
rect 12714 15544 12770 15600
rect 12714 15444 12716 15464
rect 12716 15444 12768 15464
rect 12768 15444 12770 15464
rect 12714 15408 12770 15444
rect 12622 15272 12678 15328
rect 12438 13368 12494 13424
rect 12438 12552 12494 12608
rect 12622 11192 12678 11248
rect 12806 11192 12862 11248
rect 11886 9288 11942 9344
rect 11978 9152 12034 9208
rect 11886 8508 11888 8528
rect 11888 8508 11940 8528
rect 11940 8508 11942 8528
rect 11886 8472 11942 8508
rect 11978 8200 12034 8256
rect 11886 7112 11942 7168
rect 12346 9832 12402 9888
rect 12346 8472 12402 8528
rect 12530 9560 12586 9616
rect 12806 9560 12862 9616
rect 12530 9152 12586 9208
rect 12438 8336 12494 8392
rect 12070 7148 12072 7168
rect 12072 7148 12124 7168
rect 12124 7148 12126 7168
rect 12070 7112 12126 7148
rect 11702 5072 11758 5128
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11702 2760 11758 2816
rect 11610 2624 11666 2680
rect 11150 2488 11206 2544
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 11978 6432 12034 6488
rect 11978 4936 12034 4992
rect 11978 4392 12034 4448
rect 12990 11600 13046 11656
rect 12990 11192 13046 11248
rect 12714 9324 12716 9344
rect 12716 9324 12768 9344
rect 12768 9324 12770 9344
rect 12714 9288 12770 9324
rect 12622 6704 12678 6760
rect 13266 13640 13322 13696
rect 13266 13368 13322 13424
rect 13266 11192 13322 11248
rect 13542 14456 13598 14512
rect 13726 15816 13782 15872
rect 13726 15544 13782 15600
rect 13910 13232 13966 13288
rect 13910 12860 13912 12880
rect 13912 12860 13964 12880
rect 13964 12860 13966 12880
rect 14817 20154 14873 20156
rect 14897 20154 14953 20156
rect 14977 20154 15033 20156
rect 15057 20154 15113 20156
rect 14817 20102 14843 20154
rect 14843 20102 14873 20154
rect 14897 20102 14907 20154
rect 14907 20102 14953 20154
rect 14977 20102 15023 20154
rect 15023 20102 15033 20154
rect 15057 20102 15087 20154
rect 15087 20102 15113 20154
rect 14817 20100 14873 20102
rect 14897 20100 14953 20102
rect 14977 20100 15033 20102
rect 15057 20100 15113 20102
rect 14817 19066 14873 19068
rect 14897 19066 14953 19068
rect 14977 19066 15033 19068
rect 15057 19066 15113 19068
rect 14817 19014 14843 19066
rect 14843 19014 14873 19066
rect 14897 19014 14907 19066
rect 14907 19014 14953 19066
rect 14977 19014 15023 19066
rect 15023 19014 15033 19066
rect 15057 19014 15087 19066
rect 15087 19014 15113 19066
rect 14817 19012 14873 19014
rect 14897 19012 14953 19014
rect 14977 19012 15033 19014
rect 15057 19012 15113 19014
rect 14817 17978 14873 17980
rect 14897 17978 14953 17980
rect 14977 17978 15033 17980
rect 15057 17978 15113 17980
rect 14817 17926 14843 17978
rect 14843 17926 14873 17978
rect 14897 17926 14907 17978
rect 14907 17926 14953 17978
rect 14977 17926 15023 17978
rect 15023 17926 15033 17978
rect 15057 17926 15087 17978
rect 15087 17926 15113 17978
rect 14817 17924 14873 17926
rect 14897 17924 14953 17926
rect 14977 17924 15033 17926
rect 15057 17924 15113 17926
rect 13910 12824 13966 12860
rect 14370 12824 14426 12880
rect 13726 11328 13782 11384
rect 13818 11056 13874 11112
rect 13174 9288 13230 9344
rect 13082 9152 13138 9208
rect 13082 8608 13138 8664
rect 13358 9832 13414 9888
rect 13358 9424 13414 9480
rect 13174 8472 13230 8528
rect 13082 8336 13138 8392
rect 12898 7656 12954 7712
rect 12898 6024 12954 6080
rect 12070 3984 12126 4040
rect 12254 5480 12310 5536
rect 12898 5244 12900 5264
rect 12900 5244 12952 5264
rect 12952 5244 12954 5264
rect 12898 5208 12954 5244
rect 12438 3712 12494 3768
rect 13266 7928 13322 7984
rect 13266 7656 13322 7712
rect 13358 7384 13414 7440
rect 13266 7248 13322 7304
rect 13082 4936 13138 4992
rect 12806 3848 12862 3904
rect 12254 3304 12310 3360
rect 12162 2760 12218 2816
rect 13818 9016 13874 9072
rect 14186 9052 14188 9072
rect 14188 9052 14240 9072
rect 14240 9052 14242 9072
rect 14186 9016 14242 9052
rect 13726 7248 13782 7304
rect 13726 6840 13782 6896
rect 13726 5208 13782 5264
rect 14002 7928 14058 7984
rect 14278 7792 14334 7848
rect 13910 5616 13966 5672
rect 14094 4700 14096 4720
rect 14096 4700 14148 4720
rect 14148 4700 14150 4720
rect 14094 4664 14150 4700
rect 14094 4120 14150 4176
rect 14186 3712 14242 3768
rect 13634 2488 13690 2544
rect 14278 3304 14334 3360
rect 14817 16890 14873 16892
rect 14897 16890 14953 16892
rect 14977 16890 15033 16892
rect 15057 16890 15113 16892
rect 14817 16838 14843 16890
rect 14843 16838 14873 16890
rect 14897 16838 14907 16890
rect 14907 16838 14953 16890
rect 14977 16838 15023 16890
rect 15023 16838 15033 16890
rect 15057 16838 15087 16890
rect 15087 16838 15113 16890
rect 14817 16836 14873 16838
rect 14897 16836 14953 16838
rect 14977 16836 15033 16838
rect 15057 16836 15113 16838
rect 14817 15802 14873 15804
rect 14897 15802 14953 15804
rect 14977 15802 15033 15804
rect 15057 15802 15113 15804
rect 14817 15750 14843 15802
rect 14843 15750 14873 15802
rect 14897 15750 14907 15802
rect 14907 15750 14953 15802
rect 14977 15750 15023 15802
rect 15023 15750 15033 15802
rect 15057 15750 15087 15802
rect 15087 15750 15113 15802
rect 14817 15748 14873 15750
rect 14897 15748 14953 15750
rect 14977 15748 15033 15750
rect 15057 15748 15113 15750
rect 14817 14714 14873 14716
rect 14897 14714 14953 14716
rect 14977 14714 15033 14716
rect 15057 14714 15113 14716
rect 14817 14662 14843 14714
rect 14843 14662 14873 14714
rect 14897 14662 14907 14714
rect 14907 14662 14953 14714
rect 14977 14662 15023 14714
rect 15023 14662 15033 14714
rect 15057 14662 15087 14714
rect 15087 14662 15113 14714
rect 14817 14660 14873 14662
rect 14897 14660 14953 14662
rect 14977 14660 15033 14662
rect 15057 14660 15113 14662
rect 14646 13504 14702 13560
rect 14817 13626 14873 13628
rect 14897 13626 14953 13628
rect 14977 13626 15033 13628
rect 15057 13626 15113 13628
rect 14817 13574 14843 13626
rect 14843 13574 14873 13626
rect 14897 13574 14907 13626
rect 14907 13574 14953 13626
rect 14977 13574 15023 13626
rect 15023 13574 15033 13626
rect 15057 13574 15087 13626
rect 15087 13574 15113 13626
rect 14817 13572 14873 13574
rect 14897 13572 14953 13574
rect 14977 13572 15033 13574
rect 15057 13572 15113 13574
rect 15106 13388 15162 13424
rect 15106 13368 15108 13388
rect 15108 13368 15160 13388
rect 15160 13368 15162 13388
rect 14922 13268 14924 13288
rect 14924 13268 14976 13288
rect 14976 13268 14978 13288
rect 14922 13232 14978 13268
rect 14817 12538 14873 12540
rect 14897 12538 14953 12540
rect 14977 12538 15033 12540
rect 15057 12538 15113 12540
rect 14817 12486 14843 12538
rect 14843 12486 14873 12538
rect 14897 12486 14907 12538
rect 14907 12486 14953 12538
rect 14977 12486 15023 12538
rect 15023 12486 15033 12538
rect 15057 12486 15087 12538
rect 15087 12486 15113 12538
rect 14817 12484 14873 12486
rect 14897 12484 14953 12486
rect 14977 12484 15033 12486
rect 15057 12484 15113 12486
rect 15842 18128 15898 18184
rect 15566 17176 15622 17232
rect 15474 15564 15530 15600
rect 15474 15544 15476 15564
rect 15476 15544 15528 15564
rect 15528 15544 15530 15564
rect 14554 11464 14610 11520
rect 14817 11450 14873 11452
rect 14897 11450 14953 11452
rect 14977 11450 15033 11452
rect 15057 11450 15113 11452
rect 14817 11398 14843 11450
rect 14843 11398 14873 11450
rect 14897 11398 14907 11450
rect 14907 11398 14953 11450
rect 14977 11398 15023 11450
rect 15023 11398 15033 11450
rect 15057 11398 15087 11450
rect 15087 11398 15113 11450
rect 14817 11396 14873 11398
rect 14897 11396 14953 11398
rect 14977 11396 15033 11398
rect 15057 11396 15113 11398
rect 15290 10784 15346 10840
rect 14554 9968 14610 10024
rect 14817 10362 14873 10364
rect 14897 10362 14953 10364
rect 14977 10362 15033 10364
rect 15057 10362 15113 10364
rect 14817 10310 14843 10362
rect 14843 10310 14873 10362
rect 14897 10310 14907 10362
rect 14907 10310 14953 10362
rect 14977 10310 15023 10362
rect 15023 10310 15033 10362
rect 15057 10310 15087 10362
rect 15087 10310 15113 10362
rect 14817 10308 14873 10310
rect 14897 10308 14953 10310
rect 14977 10308 15033 10310
rect 15057 10308 15113 10310
rect 14830 9832 14886 9888
rect 15474 10124 15530 10160
rect 15474 10104 15476 10124
rect 15476 10104 15528 10124
rect 15528 10104 15530 10124
rect 15198 9580 15254 9616
rect 15198 9560 15200 9580
rect 15200 9560 15252 9580
rect 15252 9560 15254 9580
rect 14817 9274 14873 9276
rect 14897 9274 14953 9276
rect 14977 9274 15033 9276
rect 15057 9274 15113 9276
rect 14817 9222 14843 9274
rect 14843 9222 14873 9274
rect 14897 9222 14907 9274
rect 14907 9222 14953 9274
rect 14977 9222 15023 9274
rect 15023 9222 15033 9274
rect 15057 9222 15087 9274
rect 15087 9222 15113 9274
rect 14817 9220 14873 9222
rect 14897 9220 14953 9222
rect 14977 9220 15033 9222
rect 15057 9220 15113 9222
rect 14830 8744 14886 8800
rect 14922 8472 14978 8528
rect 14646 8356 14702 8392
rect 14646 8336 14648 8356
rect 14648 8336 14700 8356
rect 14700 8336 14702 8356
rect 14554 8200 14610 8256
rect 14462 7248 14518 7304
rect 14817 8186 14873 8188
rect 14897 8186 14953 8188
rect 14977 8186 15033 8188
rect 15057 8186 15113 8188
rect 14817 8134 14843 8186
rect 14843 8134 14873 8186
rect 14897 8134 14907 8186
rect 14907 8134 14953 8186
rect 14977 8134 15023 8186
rect 15023 8134 15033 8186
rect 15057 8134 15087 8186
rect 15087 8134 15113 8186
rect 14817 8132 14873 8134
rect 14897 8132 14953 8134
rect 14977 8132 15033 8134
rect 15057 8132 15113 8134
rect 14817 7098 14873 7100
rect 14897 7098 14953 7100
rect 14977 7098 15033 7100
rect 15057 7098 15113 7100
rect 14817 7046 14843 7098
rect 14843 7046 14873 7098
rect 14897 7046 14907 7098
rect 14907 7046 14953 7098
rect 14977 7046 15023 7098
rect 15023 7046 15033 7098
rect 15057 7046 15087 7098
rect 15087 7046 15113 7098
rect 14817 7044 14873 7046
rect 14897 7044 14953 7046
rect 14977 7044 15033 7046
rect 15057 7044 15113 7046
rect 15382 9696 15438 9752
rect 14646 5480 14702 5536
rect 14817 6010 14873 6012
rect 14897 6010 14953 6012
rect 14977 6010 15033 6012
rect 15057 6010 15113 6012
rect 14817 5958 14843 6010
rect 14843 5958 14873 6010
rect 14897 5958 14907 6010
rect 14907 5958 14953 6010
rect 14977 5958 15023 6010
rect 15023 5958 15033 6010
rect 15057 5958 15087 6010
rect 15087 5958 15113 6010
rect 14817 5956 14873 5958
rect 14897 5956 14953 5958
rect 14977 5956 15033 5958
rect 15057 5956 15113 5958
rect 15106 5516 15108 5536
rect 15108 5516 15160 5536
rect 15160 5516 15162 5536
rect 15106 5480 15162 5516
rect 14554 3848 14610 3904
rect 14817 4922 14873 4924
rect 14897 4922 14953 4924
rect 14977 4922 15033 4924
rect 15057 4922 15113 4924
rect 14817 4870 14843 4922
rect 14843 4870 14873 4922
rect 14897 4870 14907 4922
rect 14907 4870 14953 4922
rect 14977 4870 15023 4922
rect 15023 4870 15033 4922
rect 15057 4870 15087 4922
rect 15087 4870 15113 4922
rect 14817 4868 14873 4870
rect 14897 4868 14953 4870
rect 14977 4868 15033 4870
rect 15057 4868 15113 4870
rect 15198 3848 15254 3904
rect 14817 3834 14873 3836
rect 14897 3834 14953 3836
rect 14977 3834 15033 3836
rect 15057 3834 15113 3836
rect 14817 3782 14843 3834
rect 14843 3782 14873 3834
rect 14897 3782 14907 3834
rect 14907 3782 14953 3834
rect 14977 3782 15023 3834
rect 15023 3782 15033 3834
rect 15057 3782 15087 3834
rect 15087 3782 15113 3834
rect 14817 3780 14873 3782
rect 14897 3780 14953 3782
rect 14977 3780 15033 3782
rect 15057 3780 15113 3782
rect 14646 3032 14702 3088
rect 14186 2508 14242 2544
rect 14186 2488 14188 2508
rect 14188 2488 14240 2508
rect 14240 2488 14242 2508
rect 13818 2352 13874 2408
rect 15474 9424 15530 9480
rect 15474 8200 15530 8256
rect 15934 14184 15990 14240
rect 15750 9968 15806 10024
rect 15934 9424 15990 9480
rect 15658 8200 15714 8256
rect 15474 5888 15530 5944
rect 15474 5072 15530 5128
rect 15658 6840 15714 6896
rect 15658 6024 15714 6080
rect 16118 9152 16174 9208
rect 16210 8744 16266 8800
rect 16118 7928 16174 7984
rect 16026 7792 16082 7848
rect 15474 3576 15530 3632
rect 14817 2746 14873 2748
rect 14897 2746 14953 2748
rect 14977 2746 15033 2748
rect 15057 2746 15113 2748
rect 14817 2694 14843 2746
rect 14843 2694 14873 2746
rect 14897 2694 14907 2746
rect 14907 2694 14953 2746
rect 14977 2694 15023 2746
rect 15023 2694 15033 2746
rect 15057 2694 15087 2746
rect 15087 2694 15113 2746
rect 14817 2692 14873 2694
rect 14897 2692 14953 2694
rect 14977 2692 15033 2694
rect 15057 2692 15113 2694
rect 16394 11872 16450 11928
rect 16394 10920 16450 10976
rect 18282 20698 18338 20700
rect 18362 20698 18418 20700
rect 18442 20698 18498 20700
rect 18522 20698 18578 20700
rect 18282 20646 18308 20698
rect 18308 20646 18338 20698
rect 18362 20646 18372 20698
rect 18372 20646 18418 20698
rect 18442 20646 18488 20698
rect 18488 20646 18498 20698
rect 18522 20646 18552 20698
rect 18552 20646 18578 20698
rect 18282 20644 18338 20646
rect 18362 20644 18418 20646
rect 18442 20644 18498 20646
rect 18522 20644 18578 20646
rect 18282 19610 18338 19612
rect 18362 19610 18418 19612
rect 18442 19610 18498 19612
rect 18522 19610 18578 19612
rect 18282 19558 18308 19610
rect 18308 19558 18338 19610
rect 18362 19558 18372 19610
rect 18372 19558 18418 19610
rect 18442 19558 18488 19610
rect 18488 19558 18498 19610
rect 18522 19558 18552 19610
rect 18552 19558 18578 19610
rect 18282 19556 18338 19558
rect 18362 19556 18418 19558
rect 18442 19556 18498 19558
rect 18522 19556 18578 19558
rect 18510 19252 18512 19272
rect 18512 19252 18564 19272
rect 18564 19252 18566 19272
rect 18510 19216 18566 19252
rect 17222 15580 17224 15600
rect 17224 15580 17276 15600
rect 17276 15580 17278 15600
rect 17222 15544 17278 15580
rect 16946 12280 17002 12336
rect 16946 9696 17002 9752
rect 16486 9152 16542 9208
rect 16302 8064 16358 8120
rect 16210 7520 16266 7576
rect 16026 4528 16082 4584
rect 15750 2896 15806 2952
rect 17130 8064 17186 8120
rect 16854 7404 16910 7440
rect 16854 7384 16856 7404
rect 16856 7384 16908 7404
rect 16908 7384 16910 7404
rect 16486 6568 16542 6624
rect 16486 4800 16542 4856
rect 17314 9832 17370 9888
rect 17406 7656 17462 7712
rect 18234 18708 18236 18728
rect 18236 18708 18288 18728
rect 18288 18708 18290 18728
rect 18234 18672 18290 18708
rect 19982 22616 20038 22672
rect 19062 20168 19118 20224
rect 18694 19216 18750 19272
rect 18282 18522 18338 18524
rect 18362 18522 18418 18524
rect 18442 18522 18498 18524
rect 18522 18522 18578 18524
rect 18282 18470 18308 18522
rect 18308 18470 18338 18522
rect 18362 18470 18372 18522
rect 18372 18470 18418 18522
rect 18442 18470 18488 18522
rect 18488 18470 18498 18522
rect 18522 18470 18552 18522
rect 18552 18470 18578 18522
rect 18282 18468 18338 18470
rect 18362 18468 18418 18470
rect 18442 18468 18498 18470
rect 18522 18468 18578 18470
rect 18786 18264 18842 18320
rect 18282 17434 18338 17436
rect 18362 17434 18418 17436
rect 18442 17434 18498 17436
rect 18522 17434 18578 17436
rect 18282 17382 18308 17434
rect 18308 17382 18338 17434
rect 18362 17382 18372 17434
rect 18372 17382 18418 17434
rect 18442 17382 18488 17434
rect 18488 17382 18498 17434
rect 18522 17382 18552 17434
rect 18552 17382 18578 17434
rect 18282 17380 18338 17382
rect 18362 17380 18418 17382
rect 18442 17380 18498 17382
rect 18522 17380 18578 17382
rect 18282 16346 18338 16348
rect 18362 16346 18418 16348
rect 18442 16346 18498 16348
rect 18522 16346 18578 16348
rect 18282 16294 18308 16346
rect 18308 16294 18338 16346
rect 18362 16294 18372 16346
rect 18372 16294 18418 16346
rect 18442 16294 18488 16346
rect 18488 16294 18498 16346
rect 18522 16294 18552 16346
rect 18552 16294 18578 16346
rect 18282 16292 18338 16294
rect 18362 16292 18418 16294
rect 18442 16292 18498 16294
rect 18522 16292 18578 16294
rect 19246 20576 19302 20632
rect 19706 19624 19762 19680
rect 19338 18808 19394 18864
rect 18050 14048 18106 14104
rect 18282 15258 18338 15260
rect 18362 15258 18418 15260
rect 18442 15258 18498 15260
rect 18522 15258 18578 15260
rect 18282 15206 18308 15258
rect 18308 15206 18338 15258
rect 18362 15206 18372 15258
rect 18372 15206 18418 15258
rect 18442 15206 18488 15258
rect 18488 15206 18498 15258
rect 18522 15206 18552 15258
rect 18552 15206 18578 15258
rect 18282 15204 18338 15206
rect 18362 15204 18418 15206
rect 18442 15204 18498 15206
rect 18522 15204 18578 15206
rect 18282 14170 18338 14172
rect 18362 14170 18418 14172
rect 18442 14170 18498 14172
rect 18522 14170 18578 14172
rect 18282 14118 18308 14170
rect 18308 14118 18338 14170
rect 18362 14118 18372 14170
rect 18372 14118 18418 14170
rect 18442 14118 18488 14170
rect 18488 14118 18498 14170
rect 18522 14118 18552 14170
rect 18552 14118 18578 14170
rect 18282 14116 18338 14118
rect 18362 14116 18418 14118
rect 18442 14116 18498 14118
rect 18522 14116 18578 14118
rect 17866 13776 17922 13832
rect 19062 14320 19118 14376
rect 18282 13082 18338 13084
rect 18362 13082 18418 13084
rect 18442 13082 18498 13084
rect 18522 13082 18578 13084
rect 18282 13030 18308 13082
rect 18308 13030 18338 13082
rect 18362 13030 18372 13082
rect 18372 13030 18418 13082
rect 18442 13030 18488 13082
rect 18488 13030 18498 13082
rect 18522 13030 18552 13082
rect 18552 13030 18578 13082
rect 18282 13028 18338 13030
rect 18362 13028 18418 13030
rect 18442 13028 18498 13030
rect 18522 13028 18578 13030
rect 18970 12144 19026 12200
rect 18282 11994 18338 11996
rect 18362 11994 18418 11996
rect 18442 11994 18498 11996
rect 18522 11994 18578 11996
rect 18282 11942 18308 11994
rect 18308 11942 18338 11994
rect 18362 11942 18372 11994
rect 18372 11942 18418 11994
rect 18442 11942 18488 11994
rect 18488 11942 18498 11994
rect 18522 11942 18552 11994
rect 18552 11942 18578 11994
rect 18282 11940 18338 11942
rect 18362 11940 18418 11942
rect 18442 11940 18498 11942
rect 18522 11940 18578 11942
rect 18282 10906 18338 10908
rect 18362 10906 18418 10908
rect 18442 10906 18498 10908
rect 18522 10906 18578 10908
rect 18282 10854 18308 10906
rect 18308 10854 18338 10906
rect 18362 10854 18372 10906
rect 18372 10854 18418 10906
rect 18442 10854 18488 10906
rect 18488 10854 18498 10906
rect 18522 10854 18552 10906
rect 18552 10854 18578 10906
rect 18282 10852 18338 10854
rect 18362 10852 18418 10854
rect 18442 10852 18498 10854
rect 18522 10852 18578 10854
rect 17774 10512 17830 10568
rect 17866 9696 17922 9752
rect 17774 8880 17830 8936
rect 17314 6976 17370 7032
rect 17682 6180 17738 6216
rect 17682 6160 17684 6180
rect 17684 6160 17736 6180
rect 17736 6160 17738 6180
rect 18282 9818 18338 9820
rect 18362 9818 18418 9820
rect 18442 9818 18498 9820
rect 18522 9818 18578 9820
rect 18282 9766 18308 9818
rect 18308 9766 18338 9818
rect 18362 9766 18372 9818
rect 18372 9766 18418 9818
rect 18442 9766 18488 9818
rect 18488 9766 18498 9818
rect 18522 9766 18552 9818
rect 18552 9766 18578 9818
rect 18282 9764 18338 9766
rect 18362 9764 18418 9766
rect 18442 9764 18498 9766
rect 18522 9764 18578 9766
rect 18282 8730 18338 8732
rect 18362 8730 18418 8732
rect 18442 8730 18498 8732
rect 18522 8730 18578 8732
rect 18282 8678 18308 8730
rect 18308 8678 18338 8730
rect 18362 8678 18372 8730
rect 18372 8678 18418 8730
rect 18442 8678 18488 8730
rect 18488 8678 18498 8730
rect 18522 8678 18552 8730
rect 18552 8678 18578 8730
rect 18282 8676 18338 8678
rect 18362 8676 18418 8678
rect 18442 8676 18498 8678
rect 18522 8676 18578 8678
rect 18510 8472 18566 8528
rect 18282 7642 18338 7644
rect 18362 7642 18418 7644
rect 18442 7642 18498 7644
rect 18522 7642 18578 7644
rect 18282 7590 18308 7642
rect 18308 7590 18338 7642
rect 18362 7590 18372 7642
rect 18372 7590 18418 7642
rect 18442 7590 18488 7642
rect 18488 7590 18498 7642
rect 18522 7590 18552 7642
rect 18552 7590 18578 7642
rect 18282 7588 18338 7590
rect 18362 7588 18418 7590
rect 18442 7588 18498 7590
rect 18522 7588 18578 7590
rect 18786 7520 18842 7576
rect 20534 21800 20590 21856
rect 20442 21392 20498 21448
rect 20994 20984 21050 21040
rect 19706 17604 19762 17640
rect 19706 17584 19708 17604
rect 19708 17584 19760 17604
rect 19760 17584 19762 17604
rect 19614 11736 19670 11792
rect 19154 9560 19210 9616
rect 19062 9152 19118 9208
rect 18282 6554 18338 6556
rect 18362 6554 18418 6556
rect 18442 6554 18498 6556
rect 18522 6554 18578 6556
rect 18282 6502 18308 6554
rect 18308 6502 18338 6554
rect 18362 6502 18372 6554
rect 18372 6502 18418 6554
rect 18442 6502 18488 6554
rect 18488 6502 18498 6554
rect 18522 6502 18552 6554
rect 18552 6502 18578 6554
rect 18282 6500 18338 6502
rect 18362 6500 18418 6502
rect 18442 6500 18498 6502
rect 18522 6500 18578 6502
rect 18282 5466 18338 5468
rect 18362 5466 18418 5468
rect 18442 5466 18498 5468
rect 18522 5466 18578 5468
rect 18282 5414 18308 5466
rect 18308 5414 18338 5466
rect 18362 5414 18372 5466
rect 18372 5414 18418 5466
rect 18442 5414 18488 5466
rect 18488 5414 18498 5466
rect 18522 5414 18552 5466
rect 18552 5414 18578 5466
rect 18282 5412 18338 5414
rect 18362 5412 18418 5414
rect 18442 5412 18498 5414
rect 18522 5412 18578 5414
rect 17866 5108 17868 5128
rect 17868 5108 17920 5128
rect 17920 5108 17922 5128
rect 17866 5072 17922 5108
rect 17866 4004 17922 4040
rect 17866 3984 17868 4004
rect 17868 3984 17920 4004
rect 17920 3984 17922 4004
rect 17774 3576 17830 3632
rect 18282 4378 18338 4380
rect 18362 4378 18418 4380
rect 18442 4378 18498 4380
rect 18522 4378 18578 4380
rect 18282 4326 18308 4378
rect 18308 4326 18338 4378
rect 18362 4326 18372 4378
rect 18372 4326 18418 4378
rect 18442 4326 18488 4378
rect 18488 4326 18498 4378
rect 18522 4326 18552 4378
rect 18552 4326 18578 4378
rect 18282 4324 18338 4326
rect 18362 4324 18418 4326
rect 18442 4324 18498 4326
rect 18522 4324 18578 4326
rect 19338 8472 19394 8528
rect 20074 17992 20130 18048
rect 19154 6568 19210 6624
rect 18970 3984 19026 4040
rect 18694 3440 18750 3496
rect 18282 3290 18338 3292
rect 18362 3290 18418 3292
rect 18442 3290 18498 3292
rect 18522 3290 18578 3292
rect 18282 3238 18308 3290
rect 18308 3238 18338 3290
rect 18362 3238 18372 3290
rect 18372 3238 18418 3290
rect 18442 3238 18488 3290
rect 18488 3238 18498 3290
rect 18522 3238 18552 3290
rect 18552 3238 18578 3290
rect 18282 3236 18338 3238
rect 18362 3236 18418 3238
rect 18442 3236 18498 3238
rect 18522 3236 18578 3238
rect 19430 6296 19486 6352
rect 18970 3068 18972 3088
rect 18972 3068 19024 3088
rect 19024 3068 19026 3088
rect 18970 3032 19026 3068
rect 18282 2202 18338 2204
rect 18362 2202 18418 2204
rect 18442 2202 18498 2204
rect 18522 2202 18578 2204
rect 18282 2150 18308 2202
rect 18308 2150 18338 2202
rect 18362 2150 18372 2202
rect 18372 2150 18418 2202
rect 18442 2150 18488 2202
rect 18488 2150 18498 2202
rect 18522 2150 18552 2202
rect 18552 2150 18578 2202
rect 18282 2148 18338 2150
rect 18362 2148 18418 2150
rect 18442 2148 18498 2150
rect 18522 2148 18578 2150
rect 20166 10240 20222 10296
rect 20166 9968 20222 10024
rect 19982 3884 19984 3904
rect 19984 3884 20036 3904
rect 20036 3884 20038 3904
rect 19982 3848 20038 3884
rect 19982 3032 20038 3088
rect 21638 18808 21694 18864
rect 21454 18420 21510 18456
rect 21454 18400 21456 18420
rect 21456 18400 21508 18420
rect 21508 18400 21510 18420
rect 21362 17176 21418 17232
rect 20994 16768 21050 16824
rect 21086 15816 21142 15872
rect 20994 15408 21050 15464
rect 21086 14612 21142 14648
rect 21086 14592 21088 14612
rect 21088 14592 21140 14612
rect 21140 14592 21142 14612
rect 21454 16224 21510 16280
rect 21454 15000 21510 15056
rect 22006 17604 22062 17640
rect 22006 17584 22008 17604
rect 22008 17584 22060 17604
rect 22060 17584 22062 17604
rect 20994 14184 21050 14240
rect 20994 13776 21050 13832
rect 21086 13368 21142 13424
rect 20994 12416 21050 12472
rect 21362 12824 21418 12880
rect 20350 3032 20406 3088
rect 3790 176 3846 232
rect 20166 2216 20222 2272
rect 19890 1400 19946 1456
rect 19522 584 19578 640
rect 20902 1808 20958 1864
rect 21086 5072 21142 5128
rect 21454 5072 21510 5128
rect 22006 12028 22062 12064
rect 22006 12008 22008 12028
rect 22008 12008 22060 12028
rect 22060 12008 22062 12028
rect 21086 992 21142 1048
rect 21454 856 21510 912
rect 21822 856 21878 912
rect 22006 2624 22062 2680
rect 20810 176 20866 232
<< metal3 >>
rect 0 22674 800 22704
rect 3509 22674 3575 22677
rect 0 22672 3575 22674
rect 0 22616 3514 22672
rect 3570 22616 3575 22672
rect 0 22614 3575 22616
rect 0 22584 800 22614
rect 3509 22611 3575 22614
rect 19977 22674 20043 22677
rect 22200 22674 23000 22704
rect 19977 22672 23000 22674
rect 19977 22616 19982 22672
rect 20038 22616 23000 22672
rect 19977 22614 23000 22616
rect 19977 22611 20043 22614
rect 22200 22584 23000 22614
rect 0 22266 800 22296
rect 3785 22266 3851 22269
rect 0 22264 3851 22266
rect 0 22208 3790 22264
rect 3846 22208 3851 22264
rect 0 22206 3851 22208
rect 0 22176 800 22206
rect 3785 22203 3851 22206
rect 19149 22266 19215 22269
rect 22200 22266 23000 22296
rect 19149 22264 23000 22266
rect 19149 22208 19154 22264
rect 19210 22208 23000 22264
rect 19149 22206 23000 22208
rect 19149 22203 19215 22206
rect 22200 22176 23000 22206
rect 0 21858 800 21888
rect 3417 21858 3483 21861
rect 0 21856 3483 21858
rect 0 21800 3422 21856
rect 3478 21800 3483 21856
rect 0 21798 3483 21800
rect 0 21768 800 21798
rect 3417 21795 3483 21798
rect 20529 21858 20595 21861
rect 22200 21858 23000 21888
rect 20529 21856 23000 21858
rect 20529 21800 20534 21856
rect 20590 21800 23000 21856
rect 20529 21798 23000 21800
rect 20529 21795 20595 21798
rect 22200 21768 23000 21798
rect 0 21450 800 21480
rect 3693 21450 3759 21453
rect 0 21448 3759 21450
rect 0 21392 3698 21448
rect 3754 21392 3759 21448
rect 0 21390 3759 21392
rect 0 21360 800 21390
rect 3693 21387 3759 21390
rect 20437 21450 20503 21453
rect 22200 21450 23000 21480
rect 20437 21448 23000 21450
rect 20437 21392 20442 21448
rect 20498 21392 23000 21448
rect 20437 21390 23000 21392
rect 20437 21387 20503 21390
rect 22200 21360 23000 21390
rect 0 21042 800 21072
rect 4061 21042 4127 21045
rect 0 21040 4127 21042
rect 0 20984 4066 21040
rect 4122 20984 4127 21040
rect 0 20982 4127 20984
rect 0 20952 800 20982
rect 4061 20979 4127 20982
rect 20989 21042 21055 21045
rect 22200 21042 23000 21072
rect 20989 21040 23000 21042
rect 20989 20984 20994 21040
rect 21050 20984 23000 21040
rect 20989 20982 23000 20984
rect 20989 20979 21055 20982
rect 22200 20952 23000 20982
rect 4409 20704 4729 20705
rect 0 20634 800 20664
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 20639 4729 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 18270 20704 18590 20705
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 18270 20639 18590 20640
rect 3877 20634 3943 20637
rect 0 20632 3943 20634
rect 0 20576 3882 20632
rect 3938 20576 3943 20632
rect 0 20574 3943 20576
rect 0 20544 800 20574
rect 3877 20571 3943 20574
rect 19241 20634 19307 20637
rect 22200 20634 23000 20664
rect 19241 20632 23000 20634
rect 19241 20576 19246 20632
rect 19302 20576 23000 20632
rect 19241 20574 23000 20576
rect 19241 20571 19307 20574
rect 22200 20544 23000 20574
rect 0 20226 800 20256
rect 1945 20226 2011 20229
rect 0 20224 2011 20226
rect 0 20168 1950 20224
rect 2006 20168 2011 20224
rect 0 20166 2011 20168
rect 0 20136 800 20166
rect 1945 20163 2011 20166
rect 19057 20226 19123 20229
rect 22200 20226 23000 20256
rect 19057 20224 23000 20226
rect 19057 20168 19062 20224
rect 19118 20168 23000 20224
rect 19057 20166 23000 20168
rect 19057 20163 19123 20166
rect 7874 20160 8194 20161
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8194 20160
rect 7874 20095 8194 20096
rect 14805 20160 15125 20161
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 22200 20136 23000 20166
rect 14805 20095 15125 20096
rect 0 19682 800 19712
rect 1853 19682 1919 19685
rect 0 19680 1919 19682
rect 0 19624 1858 19680
rect 1914 19624 1919 19680
rect 0 19622 1919 19624
rect 0 19592 800 19622
rect 1853 19619 1919 19622
rect 19701 19682 19767 19685
rect 22200 19682 23000 19712
rect 19701 19680 23000 19682
rect 19701 19624 19706 19680
rect 19762 19624 23000 19680
rect 19701 19622 23000 19624
rect 19701 19619 19767 19622
rect 4409 19616 4729 19617
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 19551 4729 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 18270 19616 18590 19617
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 22200 19592 23000 19622
rect 18270 19551 18590 19552
rect 7598 19348 7604 19412
rect 7668 19410 7674 19412
rect 8201 19410 8267 19413
rect 8569 19412 8635 19413
rect 8518 19410 8524 19412
rect 7668 19408 8267 19410
rect 7668 19352 8206 19408
rect 8262 19352 8267 19408
rect 7668 19350 8267 19352
rect 8478 19350 8524 19410
rect 8588 19408 8635 19412
rect 8630 19352 8635 19408
rect 7668 19348 7674 19350
rect 8201 19347 8267 19350
rect 8518 19348 8524 19350
rect 8588 19348 8635 19352
rect 8569 19347 8635 19348
rect 0 19274 800 19304
rect 2589 19274 2655 19277
rect 0 19272 2655 19274
rect 0 19216 2594 19272
rect 2650 19216 2655 19272
rect 0 19214 2655 19216
rect 0 19184 800 19214
rect 2589 19211 2655 19214
rect 3877 19274 3943 19277
rect 18505 19274 18571 19277
rect 3877 19272 18571 19274
rect 3877 19216 3882 19272
rect 3938 19216 18510 19272
rect 18566 19216 18571 19272
rect 3877 19214 18571 19216
rect 3877 19211 3943 19214
rect 18505 19211 18571 19214
rect 18689 19274 18755 19277
rect 22200 19274 23000 19304
rect 18689 19272 23000 19274
rect 18689 19216 18694 19272
rect 18750 19216 23000 19272
rect 18689 19214 23000 19216
rect 18689 19211 18755 19214
rect 22200 19184 23000 19214
rect 2957 19138 3023 19141
rect 7557 19138 7623 19141
rect 2957 19136 7623 19138
rect 2957 19080 2962 19136
rect 3018 19080 7562 19136
rect 7618 19080 7623 19136
rect 2957 19078 7623 19080
rect 2957 19075 3023 19078
rect 7557 19075 7623 19078
rect 7874 19072 8194 19073
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8194 19072
rect 7874 19007 8194 19008
rect 14805 19072 15125 19073
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 19007 15125 19008
rect 2129 19002 2195 19005
rect 4153 19002 4219 19005
rect 2129 19000 4219 19002
rect 2129 18944 2134 19000
rect 2190 18944 4158 19000
rect 4214 18944 4219 19000
rect 2129 18942 4219 18944
rect 2129 18939 2195 18942
rect 4153 18939 4219 18942
rect 5901 19002 5967 19005
rect 7097 19002 7163 19005
rect 5901 19000 7163 19002
rect 5901 18944 5906 19000
rect 5962 18944 7102 19000
rect 7158 18944 7163 19000
rect 5901 18942 7163 18944
rect 5901 18939 5967 18942
rect 7097 18939 7163 18942
rect 9857 19002 9923 19005
rect 11329 19002 11395 19005
rect 9857 19000 11395 19002
rect 9857 18944 9862 19000
rect 9918 18944 11334 19000
rect 11390 18944 11395 19000
rect 9857 18942 11395 18944
rect 9857 18939 9923 18942
rect 11329 18939 11395 18942
rect 0 18866 800 18896
rect 2773 18866 2839 18869
rect 0 18864 2839 18866
rect 0 18808 2778 18864
rect 2834 18808 2839 18864
rect 0 18806 2839 18808
rect 0 18776 800 18806
rect 2773 18803 2839 18806
rect 3785 18866 3851 18869
rect 19333 18866 19399 18869
rect 3785 18864 19399 18866
rect 3785 18808 3790 18864
rect 3846 18808 19338 18864
rect 19394 18808 19399 18864
rect 3785 18806 19399 18808
rect 3785 18803 3851 18806
rect 19333 18803 19399 18806
rect 21633 18866 21699 18869
rect 22200 18866 23000 18896
rect 21633 18864 23000 18866
rect 21633 18808 21638 18864
rect 21694 18808 23000 18864
rect 21633 18806 23000 18808
rect 21633 18803 21699 18806
rect 22200 18776 23000 18806
rect 3509 18730 3575 18733
rect 18229 18730 18295 18733
rect 3509 18728 18295 18730
rect 3509 18672 3514 18728
rect 3570 18672 18234 18728
rect 18290 18672 18295 18728
rect 3509 18670 18295 18672
rect 3509 18667 3575 18670
rect 18229 18667 18295 18670
rect 1301 18594 1367 18597
rect 2497 18594 2563 18597
rect 3141 18594 3207 18597
rect 1301 18592 2376 18594
rect 1301 18536 1306 18592
rect 1362 18536 2376 18592
rect 1301 18534 2376 18536
rect 1301 18531 1367 18534
rect 0 18458 800 18488
rect 1577 18458 1643 18461
rect 0 18456 1643 18458
rect 0 18400 1582 18456
rect 1638 18400 1643 18456
rect 0 18398 1643 18400
rect 2316 18458 2376 18534
rect 2497 18592 3207 18594
rect 2497 18536 2502 18592
rect 2558 18536 3146 18592
rect 3202 18536 3207 18592
rect 2497 18534 3207 18536
rect 2497 18531 2563 18534
rect 3141 18531 3207 18534
rect 7649 18594 7715 18597
rect 11053 18594 11119 18597
rect 7649 18592 11119 18594
rect 7649 18536 7654 18592
rect 7710 18536 11058 18592
rect 11114 18536 11119 18592
rect 7649 18534 11119 18536
rect 7649 18531 7715 18534
rect 11053 18531 11119 18534
rect 4409 18528 4729 18529
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 18463 4729 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 18270 18528 18590 18529
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 18463 18590 18464
rect 4153 18458 4219 18461
rect 2316 18456 4219 18458
rect 2316 18400 4158 18456
rect 4214 18400 4219 18456
rect 2316 18398 4219 18400
rect 0 18368 800 18398
rect 1577 18395 1643 18398
rect 4153 18395 4219 18398
rect 6269 18458 6335 18461
rect 6862 18458 6868 18460
rect 6269 18456 6868 18458
rect 6269 18400 6274 18456
rect 6330 18400 6868 18456
rect 6269 18398 6868 18400
rect 6269 18395 6335 18398
rect 6862 18396 6868 18398
rect 6932 18396 6938 18460
rect 7097 18458 7163 18461
rect 8661 18458 8727 18461
rect 7097 18456 8727 18458
rect 7097 18400 7102 18456
rect 7158 18400 8666 18456
rect 8722 18400 8727 18456
rect 7097 18398 8727 18400
rect 7097 18395 7163 18398
rect 8661 18395 8727 18398
rect 21449 18458 21515 18461
rect 22200 18458 23000 18488
rect 21449 18456 23000 18458
rect 21449 18400 21454 18456
rect 21510 18400 23000 18456
rect 21449 18398 23000 18400
rect 21449 18395 21515 18398
rect 22200 18368 23000 18398
rect 3693 18322 3759 18325
rect 18781 18322 18847 18325
rect 3693 18320 18847 18322
rect 3693 18264 3698 18320
rect 3754 18264 18786 18320
rect 18842 18264 18847 18320
rect 3693 18262 18847 18264
rect 3693 18259 3759 18262
rect 18781 18259 18847 18262
rect 3417 18186 3483 18189
rect 15837 18186 15903 18189
rect 3417 18184 15903 18186
rect 3417 18128 3422 18184
rect 3478 18128 15842 18184
rect 15898 18128 15903 18184
rect 3417 18126 15903 18128
rect 3417 18123 3483 18126
rect 15837 18123 15903 18126
rect 0 18050 800 18080
rect 1945 18050 2011 18053
rect 0 18048 2011 18050
rect 0 17992 1950 18048
rect 2006 17992 2011 18048
rect 0 17990 2011 17992
rect 0 17960 800 17990
rect 1945 17987 2011 17990
rect 2865 18050 2931 18053
rect 7557 18050 7623 18053
rect 2865 18048 7623 18050
rect 2865 17992 2870 18048
rect 2926 17992 7562 18048
rect 7618 17992 7623 18048
rect 2865 17990 7623 17992
rect 2865 17987 2931 17990
rect 7557 17987 7623 17990
rect 9857 18050 9923 18053
rect 12617 18050 12683 18053
rect 9857 18048 12683 18050
rect 9857 17992 9862 18048
rect 9918 17992 12622 18048
rect 12678 17992 12683 18048
rect 9857 17990 12683 17992
rect 9857 17987 9923 17990
rect 12617 17987 12683 17990
rect 20069 18050 20135 18053
rect 22200 18050 23000 18080
rect 20069 18048 23000 18050
rect 20069 17992 20074 18048
rect 20130 17992 23000 18048
rect 20069 17990 23000 17992
rect 20069 17987 20135 17990
rect 7874 17984 8194 17985
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8194 17984
rect 7874 17919 8194 17920
rect 14805 17984 15125 17985
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 22200 17960 23000 17990
rect 14805 17919 15125 17920
rect 2405 17778 2471 17781
rect 11237 17778 11303 17781
rect 2405 17776 11303 17778
rect 2405 17720 2410 17776
rect 2466 17720 11242 17776
rect 11298 17720 11303 17776
rect 2405 17718 11303 17720
rect 2405 17715 2471 17718
rect 11237 17715 11303 17718
rect 0 17642 800 17672
rect 1669 17642 1735 17645
rect 0 17640 1735 17642
rect 0 17584 1674 17640
rect 1730 17584 1735 17640
rect 0 17582 1735 17584
rect 0 17552 800 17582
rect 1669 17579 1735 17582
rect 6545 17642 6611 17645
rect 13169 17642 13235 17645
rect 19701 17642 19767 17645
rect 6545 17640 19767 17642
rect 6545 17584 6550 17640
rect 6606 17584 13174 17640
rect 13230 17584 19706 17640
rect 19762 17584 19767 17640
rect 6545 17582 19767 17584
rect 6545 17579 6611 17582
rect 13169 17579 13235 17582
rect 19701 17579 19767 17582
rect 22001 17642 22067 17645
rect 22200 17642 23000 17672
rect 22001 17640 23000 17642
rect 22001 17584 22006 17640
rect 22062 17584 23000 17640
rect 22001 17582 23000 17584
rect 22001 17579 22067 17582
rect 22200 17552 23000 17582
rect 3141 17504 3207 17509
rect 3141 17448 3146 17504
rect 3202 17448 3207 17504
rect 3141 17443 3207 17448
rect 7046 17444 7052 17508
rect 7116 17506 7122 17508
rect 7649 17506 7715 17509
rect 7116 17504 7715 17506
rect 7116 17448 7654 17504
rect 7710 17448 7715 17504
rect 7116 17446 7715 17448
rect 7116 17444 7122 17446
rect 7649 17443 7715 17446
rect 0 17234 800 17264
rect 1577 17234 1643 17237
rect 0 17232 1643 17234
rect 0 17176 1582 17232
rect 1638 17176 1643 17232
rect 0 17174 1643 17176
rect 3144 17234 3204 17443
rect 4409 17440 4729 17441
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 17375 4729 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 18270 17440 18590 17441
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 18270 17375 18590 17376
rect 8201 17370 8267 17373
rect 10961 17370 11027 17373
rect 8201 17368 11027 17370
rect 8201 17312 8206 17368
rect 8262 17312 10966 17368
rect 11022 17312 11027 17368
rect 8201 17310 11027 17312
rect 8201 17307 8267 17310
rect 10961 17307 11027 17310
rect 5901 17234 5967 17237
rect 6545 17234 6611 17237
rect 9489 17234 9555 17237
rect 3144 17232 9555 17234
rect 3144 17176 5906 17232
rect 5962 17176 6550 17232
rect 6606 17176 9494 17232
rect 9550 17176 9555 17232
rect 3144 17174 9555 17176
rect 0 17144 800 17174
rect 1577 17171 1643 17174
rect 5901 17171 5967 17174
rect 6545 17171 6611 17174
rect 9489 17171 9555 17174
rect 9857 17234 9923 17237
rect 15561 17234 15627 17237
rect 9857 17232 15627 17234
rect 9857 17176 9862 17232
rect 9918 17176 15566 17232
rect 15622 17176 15627 17232
rect 9857 17174 15627 17176
rect 9857 17171 9923 17174
rect 15561 17171 15627 17174
rect 21357 17234 21423 17237
rect 22200 17234 23000 17264
rect 21357 17232 23000 17234
rect 21357 17176 21362 17232
rect 21418 17176 23000 17232
rect 21357 17174 23000 17176
rect 21357 17171 21423 17174
rect 22200 17144 23000 17174
rect 6085 17098 6151 17101
rect 8201 17098 8267 17101
rect 6085 17096 8267 17098
rect 6085 17040 6090 17096
rect 6146 17040 8206 17096
rect 8262 17040 8267 17096
rect 6085 17038 8267 17040
rect 6085 17035 6151 17038
rect 8201 17035 8267 17038
rect 9673 17098 9739 17101
rect 9806 17098 9812 17100
rect 9673 17096 9812 17098
rect 9673 17040 9678 17096
rect 9734 17040 9812 17096
rect 9673 17038 9812 17040
rect 9673 17035 9739 17038
rect 9806 17036 9812 17038
rect 9876 17036 9882 17100
rect 2773 16962 2839 16965
rect 6913 16962 6979 16965
rect 2773 16960 6979 16962
rect 2773 16904 2778 16960
rect 2834 16904 6918 16960
rect 6974 16904 6979 16960
rect 2773 16902 6979 16904
rect 2773 16899 2839 16902
rect 6913 16899 6979 16902
rect 7874 16896 8194 16897
rect 0 16826 800 16856
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8194 16896
rect 7874 16831 8194 16832
rect 14805 16896 15125 16897
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 16831 15125 16832
rect 2773 16826 2839 16829
rect 10501 16828 10567 16829
rect 10501 16826 10548 16828
rect 0 16824 2839 16826
rect 0 16768 2778 16824
rect 2834 16768 2839 16824
rect 0 16766 2839 16768
rect 10456 16824 10548 16826
rect 10456 16768 10506 16824
rect 10456 16766 10548 16768
rect 0 16736 800 16766
rect 2773 16763 2839 16766
rect 10501 16764 10548 16766
rect 10612 16764 10618 16828
rect 20989 16826 21055 16829
rect 22200 16826 23000 16856
rect 20989 16824 23000 16826
rect 20989 16768 20994 16824
rect 21050 16768 23000 16824
rect 20989 16766 23000 16768
rect 10501 16763 10567 16764
rect 20989 16763 21055 16766
rect 22200 16736 23000 16766
rect 11329 16554 11395 16557
rect 11830 16554 11836 16556
rect 11329 16552 11836 16554
rect 11329 16496 11334 16552
rect 11390 16496 11836 16552
rect 11329 16494 11836 16496
rect 11329 16491 11395 16494
rect 11830 16492 11836 16494
rect 11900 16492 11906 16556
rect 8937 16418 9003 16421
rect 9254 16418 9260 16420
rect 8937 16416 9260 16418
rect 8937 16360 8942 16416
rect 8998 16360 9260 16416
rect 8937 16358 9260 16360
rect 8937 16355 9003 16358
rect 9254 16356 9260 16358
rect 9324 16356 9330 16420
rect 4409 16352 4729 16353
rect 0 16282 800 16312
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 16287 4729 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 18270 16352 18590 16353
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 16287 18590 16288
rect 2313 16282 2379 16285
rect 0 16280 2379 16282
rect 0 16224 2318 16280
rect 2374 16224 2379 16280
rect 0 16222 2379 16224
rect 0 16192 800 16222
rect 2313 16219 2379 16222
rect 7414 16220 7420 16284
rect 7484 16282 7490 16284
rect 9121 16282 9187 16285
rect 7484 16280 9187 16282
rect 7484 16224 9126 16280
rect 9182 16224 9187 16280
rect 7484 16222 9187 16224
rect 7484 16220 7490 16222
rect 9121 16219 9187 16222
rect 21449 16282 21515 16285
rect 22200 16282 23000 16312
rect 21449 16280 23000 16282
rect 21449 16224 21454 16280
rect 21510 16224 23000 16280
rect 21449 16222 23000 16224
rect 21449 16219 21515 16222
rect 22200 16192 23000 16222
rect 1761 16146 1827 16149
rect 3785 16146 3851 16149
rect 8937 16146 9003 16149
rect 1761 16144 9003 16146
rect 1761 16088 1766 16144
rect 1822 16088 3790 16144
rect 3846 16088 8942 16144
rect 8998 16088 9003 16144
rect 1761 16086 9003 16088
rect 1761 16083 1827 16086
rect 3785 16083 3851 16086
rect 8937 16083 9003 16086
rect 0 15874 800 15904
rect 1945 15874 2011 15877
rect 0 15872 2011 15874
rect 0 15816 1950 15872
rect 2006 15816 2011 15872
rect 0 15814 2011 15816
rect 0 15784 800 15814
rect 1945 15811 2011 15814
rect 11973 15874 12039 15877
rect 13721 15874 13787 15877
rect 11973 15872 13787 15874
rect 11973 15816 11978 15872
rect 12034 15816 13726 15872
rect 13782 15816 13787 15872
rect 11973 15814 13787 15816
rect 11973 15811 12039 15814
rect 13721 15811 13787 15814
rect 21081 15874 21147 15877
rect 22200 15874 23000 15904
rect 21081 15872 23000 15874
rect 21081 15816 21086 15872
rect 21142 15816 23000 15872
rect 21081 15814 23000 15816
rect 21081 15811 21147 15814
rect 7874 15808 8194 15809
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8194 15808
rect 7874 15743 8194 15744
rect 14805 15808 15125 15809
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 22200 15784 23000 15814
rect 14805 15743 15125 15744
rect 3693 15602 3759 15605
rect 7230 15602 7236 15604
rect 3693 15600 7236 15602
rect 3693 15544 3698 15600
rect 3754 15544 7236 15600
rect 3693 15542 7236 15544
rect 3693 15539 3759 15542
rect 7230 15540 7236 15542
rect 7300 15602 7306 15604
rect 8109 15602 8175 15605
rect 7300 15600 8175 15602
rect 7300 15544 8114 15600
rect 8170 15544 8175 15600
rect 7300 15542 8175 15544
rect 7300 15540 7306 15542
rect 8109 15539 8175 15542
rect 9305 15602 9371 15605
rect 10225 15602 10291 15605
rect 9305 15600 10291 15602
rect 9305 15544 9310 15600
rect 9366 15544 10230 15600
rect 10286 15544 10291 15600
rect 9305 15542 10291 15544
rect 9305 15539 9371 15542
rect 10225 15539 10291 15542
rect 12157 15602 12223 15605
rect 12709 15602 12775 15605
rect 13721 15602 13787 15605
rect 12157 15600 13787 15602
rect 12157 15544 12162 15600
rect 12218 15544 12714 15600
rect 12770 15544 13726 15600
rect 13782 15544 13787 15600
rect 12157 15542 13787 15544
rect 12157 15539 12223 15542
rect 12709 15539 12775 15542
rect 13721 15539 13787 15542
rect 15469 15602 15535 15605
rect 17217 15602 17283 15605
rect 15469 15600 17283 15602
rect 15469 15544 15474 15600
rect 15530 15544 17222 15600
rect 17278 15544 17283 15600
rect 15469 15542 17283 15544
rect 15469 15539 15535 15542
rect 17217 15539 17283 15542
rect 0 15466 800 15496
rect 3785 15466 3851 15469
rect 0 15464 3851 15466
rect 0 15408 3790 15464
rect 3846 15408 3851 15464
rect 0 15406 3851 15408
rect 0 15376 800 15406
rect 3785 15403 3851 15406
rect 8753 15466 8819 15469
rect 12709 15466 12775 15469
rect 8753 15464 12775 15466
rect 8753 15408 8758 15464
rect 8814 15408 12714 15464
rect 12770 15408 12775 15464
rect 8753 15406 12775 15408
rect 8753 15403 8819 15406
rect 12709 15403 12775 15406
rect 20989 15466 21055 15469
rect 22200 15466 23000 15496
rect 20989 15464 23000 15466
rect 20989 15408 20994 15464
rect 21050 15408 23000 15464
rect 20989 15406 23000 15408
rect 20989 15403 21055 15406
rect 22200 15376 23000 15406
rect 12617 15332 12683 15333
rect 12566 15268 12572 15332
rect 12636 15330 12683 15332
rect 12636 15328 12728 15330
rect 12678 15272 12728 15328
rect 12636 15270 12728 15272
rect 12636 15268 12683 15270
rect 12617 15267 12683 15268
rect 4409 15264 4729 15265
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 15199 4729 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 18270 15264 18590 15265
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 15199 18590 15200
rect 0 15058 800 15088
rect 1761 15058 1827 15061
rect 0 15056 1827 15058
rect 0 15000 1766 15056
rect 1822 15000 1827 15056
rect 0 14998 1827 15000
rect 0 14968 800 14998
rect 1761 14995 1827 14998
rect 21449 15058 21515 15061
rect 22200 15058 23000 15088
rect 21449 15056 23000 15058
rect 21449 15000 21454 15056
rect 21510 15000 23000 15056
rect 21449 14998 23000 15000
rect 21449 14995 21515 14998
rect 22200 14968 23000 14998
rect 5349 14922 5415 14925
rect 6269 14922 6335 14925
rect 7925 14922 7991 14925
rect 5349 14920 7991 14922
rect 5349 14864 5354 14920
rect 5410 14864 6274 14920
rect 6330 14864 7930 14920
rect 7986 14864 7991 14920
rect 5349 14862 7991 14864
rect 5349 14859 5415 14862
rect 6269 14859 6335 14862
rect 7925 14859 7991 14862
rect 8845 14922 8911 14925
rect 9213 14922 9279 14925
rect 8845 14920 9279 14922
rect 8845 14864 8850 14920
rect 8906 14864 9218 14920
rect 9274 14864 9279 14920
rect 8845 14862 9279 14864
rect 8845 14859 8911 14862
rect 9213 14859 9279 14862
rect 9990 14860 9996 14924
rect 10060 14922 10066 14924
rect 10133 14922 10199 14925
rect 10060 14920 10199 14922
rect 10060 14864 10138 14920
rect 10194 14864 10199 14920
rect 10060 14862 10199 14864
rect 10060 14860 10066 14862
rect 10133 14859 10199 14862
rect 10409 14788 10475 14789
rect 10358 14724 10364 14788
rect 10428 14786 10475 14788
rect 10428 14784 10520 14786
rect 10470 14728 10520 14784
rect 10428 14726 10520 14728
rect 10428 14724 10475 14726
rect 10409 14723 10475 14724
rect 7874 14720 8194 14721
rect 0 14650 800 14680
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8194 14720
rect 7874 14655 8194 14656
rect 14805 14720 15125 14721
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 14655 15125 14656
rect 1853 14650 1919 14653
rect 0 14648 1919 14650
rect 0 14592 1858 14648
rect 1914 14592 1919 14648
rect 0 14590 1919 14592
rect 0 14560 800 14590
rect 1853 14587 1919 14590
rect 2037 14650 2103 14653
rect 3969 14650 4035 14653
rect 2037 14648 4035 14650
rect 2037 14592 2042 14648
rect 2098 14592 3974 14648
rect 4030 14592 4035 14648
rect 2037 14590 4035 14592
rect 2037 14587 2103 14590
rect 3969 14587 4035 14590
rect 9622 14588 9628 14652
rect 9692 14650 9698 14652
rect 10317 14650 10383 14653
rect 9692 14648 10383 14650
rect 9692 14592 10322 14648
rect 10378 14592 10383 14648
rect 9692 14590 10383 14592
rect 9692 14588 9698 14590
rect 10317 14587 10383 14590
rect 21081 14650 21147 14653
rect 22200 14650 23000 14680
rect 21081 14648 23000 14650
rect 21081 14592 21086 14648
rect 21142 14592 23000 14648
rect 21081 14590 23000 14592
rect 21081 14587 21147 14590
rect 22200 14560 23000 14590
rect 11329 14514 11395 14517
rect 13537 14514 13603 14517
rect 11329 14512 13603 14514
rect 11329 14456 11334 14512
rect 11390 14456 13542 14512
rect 13598 14456 13603 14512
rect 11329 14454 13603 14456
rect 11329 14451 11395 14454
rect 13537 14451 13603 14454
rect 1577 14378 1643 14381
rect 7414 14378 7420 14380
rect 1577 14376 7420 14378
rect 1577 14320 1582 14376
rect 1638 14320 7420 14376
rect 1577 14318 7420 14320
rect 1577 14315 1643 14318
rect 7414 14316 7420 14318
rect 7484 14316 7490 14380
rect 11697 14378 11763 14381
rect 19057 14378 19123 14381
rect 11697 14376 19123 14378
rect 11697 14320 11702 14376
rect 11758 14320 19062 14376
rect 19118 14320 19123 14376
rect 11697 14318 19123 14320
rect 11697 14315 11763 14318
rect 19057 14315 19123 14318
rect 0 14242 800 14272
rect 1761 14242 1827 14245
rect 0 14240 1827 14242
rect 0 14184 1766 14240
rect 1822 14184 1827 14240
rect 0 14182 1827 14184
rect 0 14152 800 14182
rect 1761 14179 1827 14182
rect 12065 14242 12131 14245
rect 15929 14242 15995 14245
rect 12065 14240 15995 14242
rect 12065 14184 12070 14240
rect 12126 14184 15934 14240
rect 15990 14184 15995 14240
rect 12065 14182 15995 14184
rect 12065 14179 12131 14182
rect 15929 14179 15995 14182
rect 20989 14242 21055 14245
rect 22200 14242 23000 14272
rect 20989 14240 23000 14242
rect 20989 14184 20994 14240
rect 21050 14184 23000 14240
rect 20989 14182 23000 14184
rect 20989 14179 21055 14182
rect 4409 14176 4729 14177
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 14111 4729 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 18270 14176 18590 14177
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 22200 14152 23000 14182
rect 18270 14111 18590 14112
rect 8109 14106 8175 14109
rect 6548 14104 8175 14106
rect 6548 14048 8114 14104
rect 8170 14048 8175 14104
rect 6548 14046 8175 14048
rect 0 13834 800 13864
rect 2773 13834 2839 13837
rect 0 13832 2839 13834
rect 0 13776 2778 13832
rect 2834 13776 2839 13832
rect 0 13774 2839 13776
rect 0 13744 800 13774
rect 2773 13771 2839 13774
rect 6548 13701 6608 14046
rect 8109 14043 8175 14046
rect 8661 14106 8727 14109
rect 9622 14106 9628 14108
rect 8661 14104 9628 14106
rect 8661 14048 8666 14104
rect 8722 14048 9628 14104
rect 8661 14046 9628 14048
rect 8661 14043 8727 14046
rect 9622 14044 9628 14046
rect 9692 14044 9698 14108
rect 10041 14106 10107 14109
rect 9998 14104 10107 14106
rect 9998 14048 10046 14104
rect 10102 14048 10107 14104
rect 9998 14043 10107 14048
rect 12249 14106 12315 14109
rect 18045 14106 18111 14109
rect 12249 14104 18111 14106
rect 12249 14048 12254 14104
rect 12310 14048 18050 14104
rect 18106 14048 18111 14104
rect 12249 14046 18111 14048
rect 12249 14043 12315 14046
rect 18045 14043 18111 14046
rect 9998 13837 10058 14043
rect 8109 13834 8175 13837
rect 8702 13834 8708 13836
rect 8109 13832 8708 13834
rect 8109 13776 8114 13832
rect 8170 13776 8708 13832
rect 8109 13774 8708 13776
rect 8109 13771 8175 13774
rect 8702 13772 8708 13774
rect 8772 13772 8778 13836
rect 9949 13832 10058 13837
rect 9949 13776 9954 13832
rect 10010 13776 10058 13832
rect 9949 13774 10058 13776
rect 9949 13771 10015 13774
rect 11094 13772 11100 13836
rect 11164 13834 11170 13836
rect 11605 13834 11671 13837
rect 17861 13834 17927 13837
rect 11164 13832 17927 13834
rect 11164 13776 11610 13832
rect 11666 13776 17866 13832
rect 17922 13776 17927 13832
rect 11164 13774 17927 13776
rect 11164 13772 11170 13774
rect 11605 13771 11671 13774
rect 17861 13771 17927 13774
rect 20989 13834 21055 13837
rect 22200 13834 23000 13864
rect 20989 13832 23000 13834
rect 20989 13776 20994 13832
rect 21050 13776 23000 13832
rect 20989 13774 23000 13776
rect 20989 13771 21055 13774
rect 22200 13744 23000 13774
rect 6545 13696 6611 13701
rect 6545 13640 6550 13696
rect 6606 13640 6611 13696
rect 6545 13635 6611 13640
rect 8753 13698 8819 13701
rect 13261 13698 13327 13701
rect 8753 13696 13327 13698
rect 8753 13640 8758 13696
rect 8814 13640 13266 13696
rect 13322 13640 13327 13696
rect 8753 13638 13327 13640
rect 8753 13635 8819 13638
rect 13261 13635 13327 13638
rect 7874 13632 8194 13633
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8194 13632
rect 7874 13567 8194 13568
rect 14805 13632 15125 13633
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 13567 15125 13568
rect 7189 13562 7255 13565
rect 8845 13564 8911 13565
rect 9489 13564 9555 13565
rect 8845 13562 8892 13564
rect 7189 13560 7666 13562
rect 7189 13504 7194 13560
rect 7250 13504 7666 13560
rect 7189 13502 7666 13504
rect 8800 13560 8892 13562
rect 8800 13504 8850 13560
rect 8800 13502 8892 13504
rect 7189 13499 7255 13502
rect 0 13426 800 13456
rect 2405 13426 2471 13429
rect 0 13424 2471 13426
rect 0 13368 2410 13424
rect 2466 13368 2471 13424
rect 0 13366 2471 13368
rect 7606 13426 7666 13502
rect 8845 13500 8892 13502
rect 8956 13500 8962 13564
rect 9438 13500 9444 13564
rect 9508 13562 9555 13564
rect 10133 13562 10199 13565
rect 14641 13562 14707 13565
rect 9508 13560 9600 13562
rect 9550 13504 9600 13560
rect 9508 13502 9600 13504
rect 10133 13560 14707 13562
rect 10133 13504 10138 13560
rect 10194 13504 14646 13560
rect 14702 13504 14707 13560
rect 10133 13502 14707 13504
rect 9508 13500 9555 13502
rect 8845 13499 8911 13500
rect 9489 13499 9555 13500
rect 10133 13499 10199 13502
rect 14641 13499 14707 13502
rect 8293 13426 8359 13429
rect 7606 13424 8359 13426
rect 7606 13368 8298 13424
rect 8354 13368 8359 13424
rect 7606 13366 8359 13368
rect 0 13336 800 13366
rect 2405 13363 2471 13366
rect 8293 13363 8359 13366
rect 10910 13364 10916 13428
rect 10980 13426 10986 13428
rect 12433 13426 12499 13429
rect 10980 13424 12499 13426
rect 10980 13368 12438 13424
rect 12494 13368 12499 13424
rect 10980 13366 12499 13368
rect 10980 13364 10986 13366
rect 12433 13363 12499 13366
rect 13261 13426 13327 13429
rect 15101 13426 15167 13429
rect 13261 13424 15167 13426
rect 13261 13368 13266 13424
rect 13322 13368 15106 13424
rect 15162 13368 15167 13424
rect 13261 13366 15167 13368
rect 13261 13363 13327 13366
rect 15101 13363 15167 13366
rect 21081 13426 21147 13429
rect 22200 13426 23000 13456
rect 21081 13424 23000 13426
rect 21081 13368 21086 13424
rect 21142 13368 23000 13424
rect 21081 13366 23000 13368
rect 21081 13363 21147 13366
rect 22200 13336 23000 13366
rect 3049 13290 3115 13293
rect 6545 13290 6611 13293
rect 8937 13290 9003 13293
rect 9305 13290 9371 13293
rect 3049 13288 6424 13290
rect 3049 13232 3054 13288
rect 3110 13232 6424 13288
rect 3049 13230 6424 13232
rect 3049 13227 3115 13230
rect 6364 13154 6424 13230
rect 6545 13288 9371 13290
rect 6545 13232 6550 13288
rect 6606 13232 8942 13288
rect 8998 13232 9310 13288
rect 9366 13232 9371 13288
rect 6545 13230 9371 13232
rect 6545 13227 6611 13230
rect 8937 13227 9003 13230
rect 9305 13227 9371 13230
rect 10501 13290 10567 13293
rect 11605 13290 11671 13293
rect 10501 13288 11671 13290
rect 10501 13232 10506 13288
rect 10562 13232 11610 13288
rect 11666 13232 11671 13288
rect 10501 13230 11671 13232
rect 10501 13227 10567 13230
rect 11605 13227 11671 13230
rect 13905 13290 13971 13293
rect 14917 13290 14983 13293
rect 13905 13288 14983 13290
rect 13905 13232 13910 13288
rect 13966 13232 14922 13288
rect 14978 13232 14983 13288
rect 13905 13230 14983 13232
rect 13905 13227 13971 13230
rect 14917 13227 14983 13230
rect 9029 13154 9095 13157
rect 6364 13152 9095 13154
rect 6364 13096 9034 13152
rect 9090 13096 9095 13152
rect 6364 13094 9095 13096
rect 9029 13091 9095 13094
rect 4409 13088 4729 13089
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 13023 4729 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 18270 13088 18590 13089
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 13023 18590 13024
rect 0 12882 800 12912
rect 1669 12882 1735 12885
rect 0 12880 1735 12882
rect 0 12824 1674 12880
rect 1730 12824 1735 12880
rect 0 12822 1735 12824
rect 0 12792 800 12822
rect 1669 12819 1735 12822
rect 6637 12882 6703 12885
rect 8293 12882 8359 12885
rect 9121 12882 9187 12885
rect 6637 12880 6746 12882
rect 6637 12824 6642 12880
rect 6698 12824 6746 12880
rect 6637 12819 6746 12824
rect 8293 12880 9187 12882
rect 8293 12824 8298 12880
rect 8354 12824 9126 12880
rect 9182 12824 9187 12880
rect 8293 12822 9187 12824
rect 8293 12819 8359 12822
rect 9121 12819 9187 12822
rect 9305 12882 9371 12885
rect 10685 12882 10751 12885
rect 9305 12880 10751 12882
rect 9305 12824 9310 12880
rect 9366 12824 10690 12880
rect 10746 12824 10751 12880
rect 9305 12822 10751 12824
rect 9305 12819 9371 12822
rect 10685 12819 10751 12822
rect 13905 12882 13971 12885
rect 14365 12882 14431 12885
rect 13905 12880 14431 12882
rect 13905 12824 13910 12880
rect 13966 12824 14370 12880
rect 14426 12824 14431 12880
rect 13905 12822 14431 12824
rect 13905 12819 13971 12822
rect 14365 12819 14431 12822
rect 21357 12882 21423 12885
rect 22200 12882 23000 12912
rect 21357 12880 23000 12882
rect 21357 12824 21362 12880
rect 21418 12824 23000 12880
rect 21357 12822 23000 12824
rect 21357 12819 21423 12822
rect 5717 12612 5783 12613
rect 5717 12610 5764 12612
rect 5672 12608 5764 12610
rect 5672 12552 5722 12608
rect 5672 12550 5764 12552
rect 5717 12548 5764 12550
rect 5828 12548 5834 12612
rect 5717 12547 5783 12548
rect 0 12474 800 12504
rect 3141 12474 3207 12477
rect 0 12472 3207 12474
rect 0 12416 3146 12472
rect 3202 12416 3207 12472
rect 0 12414 3207 12416
rect 0 12384 800 12414
rect 3141 12411 3207 12414
rect 5257 12338 5323 12341
rect 5214 12336 5323 12338
rect 5214 12280 5262 12336
rect 5318 12280 5323 12336
rect 5214 12275 5323 12280
rect 6361 12338 6427 12341
rect 6686 12338 6746 12819
rect 22200 12792 23000 12822
rect 6862 12684 6868 12748
rect 6932 12746 6938 12748
rect 8477 12746 8543 12749
rect 6932 12744 8543 12746
rect 6932 12688 8482 12744
rect 8538 12688 8543 12744
rect 6932 12686 8543 12688
rect 6932 12684 6938 12686
rect 8477 12683 8543 12686
rect 9305 12610 9371 12613
rect 11421 12610 11487 12613
rect 12433 12610 12499 12613
rect 9305 12608 12499 12610
rect 9305 12552 9310 12608
rect 9366 12552 11426 12608
rect 11482 12552 12438 12608
rect 12494 12552 12499 12608
rect 9305 12550 12499 12552
rect 9305 12547 9371 12550
rect 11421 12547 11487 12550
rect 12433 12547 12499 12550
rect 7874 12544 8194 12545
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8194 12544
rect 7874 12479 8194 12480
rect 14805 12544 15125 12545
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 12479 15125 12480
rect 8477 12474 8543 12477
rect 11094 12474 11100 12476
rect 8477 12472 11100 12474
rect 8477 12416 8482 12472
rect 8538 12416 11100 12472
rect 8477 12414 11100 12416
rect 8477 12411 8543 12414
rect 11094 12412 11100 12414
rect 11164 12412 11170 12476
rect 20989 12474 21055 12477
rect 22200 12474 23000 12504
rect 11700 12414 12496 12474
rect 9397 12338 9463 12341
rect 6361 12336 9463 12338
rect 6361 12280 6366 12336
rect 6422 12280 9402 12336
rect 9458 12280 9463 12336
rect 6361 12278 9463 12280
rect 6361 12275 6427 12278
rect 9397 12275 9463 12278
rect 10133 12338 10199 12341
rect 11700 12338 11760 12414
rect 11881 12340 11947 12341
rect 10133 12336 11760 12338
rect 10133 12280 10138 12336
rect 10194 12280 11760 12336
rect 10133 12278 11760 12280
rect 10133 12275 10199 12278
rect 11830 12276 11836 12340
rect 11900 12338 11947 12340
rect 12436 12338 12496 12414
rect 20989 12472 23000 12474
rect 20989 12416 20994 12472
rect 21050 12416 23000 12472
rect 20989 12414 23000 12416
rect 20989 12411 21055 12414
rect 22200 12384 23000 12414
rect 16941 12338 17007 12341
rect 11900 12336 11992 12338
rect 11942 12280 11992 12336
rect 11900 12278 11992 12280
rect 12436 12336 17007 12338
rect 12436 12280 16946 12336
rect 17002 12280 17007 12336
rect 12436 12278 17007 12280
rect 11900 12276 11947 12278
rect 11881 12275 11947 12276
rect 16941 12275 17007 12278
rect 0 12066 800 12096
rect 1577 12066 1643 12069
rect 0 12064 1643 12066
rect 0 12008 1582 12064
rect 1638 12008 1643 12064
rect 0 12006 1643 12008
rect 0 11976 800 12006
rect 1577 12003 1643 12006
rect 5073 12066 5139 12069
rect 5214 12066 5274 12275
rect 11421 12202 11487 12205
rect 18965 12202 19031 12205
rect 11421 12200 19031 12202
rect 11421 12144 11426 12200
rect 11482 12144 18970 12200
rect 19026 12144 19031 12200
rect 11421 12142 19031 12144
rect 11421 12139 11487 12142
rect 18965 12139 19031 12142
rect 5073 12064 5274 12066
rect 5073 12008 5078 12064
rect 5134 12008 5274 12064
rect 5073 12006 5274 12008
rect 22001 12066 22067 12069
rect 22200 12066 23000 12096
rect 22001 12064 23000 12066
rect 22001 12008 22006 12064
rect 22062 12008 23000 12064
rect 22001 12006 23000 12008
rect 5073 12003 5139 12006
rect 22001 12003 22067 12006
rect 4409 12000 4729 12001
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 11935 4729 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 18270 12000 18590 12001
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 22200 11976 23000 12006
rect 18270 11935 18590 11936
rect 3877 11932 3943 11933
rect 6913 11932 6979 11933
rect 3877 11928 3924 11932
rect 3988 11930 3994 11932
rect 3877 11872 3882 11928
rect 3877 11868 3924 11872
rect 3988 11870 4034 11930
rect 3988 11868 3994 11870
rect 6862 11868 6868 11932
rect 6932 11930 6979 11932
rect 11973 11932 12039 11933
rect 11973 11930 12020 11932
rect 6932 11928 7024 11930
rect 6974 11872 7024 11928
rect 6932 11870 7024 11872
rect 11928 11928 12020 11930
rect 11928 11872 11978 11928
rect 11928 11870 12020 11872
rect 6932 11868 6979 11870
rect 3877 11867 3943 11868
rect 6913 11867 6979 11868
rect 11973 11868 12020 11870
rect 12084 11868 12090 11932
rect 12157 11930 12223 11933
rect 16389 11930 16455 11933
rect 12157 11928 16455 11930
rect 12157 11872 12162 11928
rect 12218 11872 16394 11928
rect 16450 11872 16455 11928
rect 12157 11870 16455 11872
rect 11973 11867 12039 11868
rect 12157 11867 12223 11870
rect 16389 11867 16455 11870
rect 7097 11794 7163 11797
rect 7414 11794 7420 11796
rect 7097 11792 7420 11794
rect 7097 11736 7102 11792
rect 7158 11736 7420 11792
rect 7097 11734 7420 11736
rect 7097 11731 7163 11734
rect 7414 11732 7420 11734
rect 7484 11732 7490 11796
rect 10501 11794 10567 11797
rect 19609 11794 19675 11797
rect 10501 11792 19675 11794
rect 10501 11736 10506 11792
rect 10562 11736 19614 11792
rect 19670 11736 19675 11792
rect 10501 11734 19675 11736
rect 10501 11731 10567 11734
rect 19609 11731 19675 11734
rect 0 11658 800 11688
rect 3877 11658 3943 11661
rect 0 11656 3943 11658
rect 0 11600 3882 11656
rect 3938 11600 3943 11656
rect 0 11598 3943 11600
rect 0 11568 800 11598
rect 3877 11595 3943 11598
rect 6085 11658 6151 11661
rect 8661 11658 8727 11661
rect 6085 11656 8727 11658
rect 6085 11600 6090 11656
rect 6146 11600 8666 11656
rect 8722 11600 8727 11656
rect 6085 11598 8727 11600
rect 6085 11595 6151 11598
rect 8661 11595 8727 11598
rect 12985 11658 13051 11661
rect 22200 11658 23000 11688
rect 12985 11656 23000 11658
rect 12985 11600 12990 11656
rect 13046 11600 23000 11656
rect 12985 11598 23000 11600
rect 12985 11595 13051 11598
rect 22200 11568 23000 11598
rect 3325 11524 3391 11525
rect 3325 11520 3372 11524
rect 3436 11522 3442 11524
rect 7281 11522 7347 11525
rect 14549 11522 14615 11525
rect 3325 11464 3330 11520
rect 3325 11460 3372 11464
rect 3436 11462 3482 11522
rect 4478 11520 7347 11522
rect 4478 11464 7286 11520
rect 7342 11464 7347 11520
rect 4478 11462 7347 11464
rect 3436 11460 3442 11462
rect 3325 11459 3391 11460
rect 0 11250 800 11280
rect 4478 11250 4538 11462
rect 7281 11459 7347 11462
rect 9998 11520 14615 11522
rect 9998 11464 14554 11520
rect 14610 11464 14615 11520
rect 9998 11462 14615 11464
rect 7874 11456 8194 11457
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8194 11456
rect 7874 11391 8194 11392
rect 4705 11386 4771 11389
rect 5073 11386 5139 11389
rect 5441 11386 5507 11389
rect 6637 11386 6703 11389
rect 4705 11384 5274 11386
rect 4705 11328 4710 11384
rect 4766 11328 5078 11384
rect 5134 11328 5274 11384
rect 4705 11326 5274 11328
rect 4705 11323 4771 11326
rect 5073 11323 5139 11326
rect 0 11190 4538 11250
rect 5214 11250 5274 11326
rect 5441 11384 6703 11386
rect 5441 11328 5446 11384
rect 5502 11328 6642 11384
rect 6698 11328 6703 11384
rect 5441 11326 6703 11328
rect 5441 11323 5507 11326
rect 6637 11323 6703 11326
rect 7281 11386 7347 11389
rect 7649 11386 7715 11389
rect 7281 11384 7715 11386
rect 7281 11328 7286 11384
rect 7342 11328 7654 11384
rect 7710 11328 7715 11384
rect 7281 11326 7715 11328
rect 7281 11323 7347 11326
rect 7649 11323 7715 11326
rect 9765 11386 9831 11389
rect 9998 11388 10058 11462
rect 14549 11459 14615 11462
rect 14805 11456 15125 11457
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 11391 15125 11392
rect 9990 11386 9996 11388
rect 9765 11384 9996 11386
rect 9765 11328 9770 11384
rect 9826 11328 9996 11384
rect 9765 11326 9996 11328
rect 9765 11323 9831 11326
rect 9990 11324 9996 11326
rect 10060 11324 10066 11388
rect 10133 11386 10199 11389
rect 13721 11386 13787 11389
rect 10133 11384 13787 11386
rect 10133 11328 10138 11384
rect 10194 11328 13726 11384
rect 13782 11328 13787 11384
rect 10133 11326 13787 11328
rect 10133 11323 10199 11326
rect 13721 11323 13787 11326
rect 10409 11250 10475 11253
rect 5214 11248 10475 11250
rect 5214 11192 10414 11248
rect 10470 11192 10475 11248
rect 5214 11190 10475 11192
rect 0 11160 800 11190
rect 10409 11187 10475 11190
rect 10869 11250 10935 11253
rect 12617 11250 12683 11253
rect 12801 11250 12867 11253
rect 10869 11248 12496 11250
rect 10869 11192 10874 11248
rect 10930 11192 12496 11248
rect 10869 11190 12496 11192
rect 10869 11187 10935 11190
rect 6453 11114 6519 11117
rect 7465 11114 7531 11117
rect 12065 11114 12131 11117
rect 6453 11112 12131 11114
rect 6453 11056 6458 11112
rect 6514 11056 7470 11112
rect 7526 11056 12070 11112
rect 12126 11056 12131 11112
rect 6453 11054 12131 11056
rect 6453 11051 6519 11054
rect 7465 11051 7531 11054
rect 12065 11051 12131 11054
rect 6453 10978 6519 10981
rect 9254 10978 9260 10980
rect 6453 10976 9260 10978
rect 6453 10920 6458 10976
rect 6514 10920 9260 10976
rect 6453 10918 9260 10920
rect 6453 10915 6519 10918
rect 9254 10916 9260 10918
rect 9324 10916 9330 10980
rect 12436 10978 12496 11190
rect 12617 11248 12867 11250
rect 12617 11192 12622 11248
rect 12678 11192 12806 11248
rect 12862 11192 12867 11248
rect 12617 11190 12867 11192
rect 12617 11187 12683 11190
rect 12801 11187 12867 11190
rect 12985 11250 13051 11253
rect 13261 11250 13327 11253
rect 22200 11250 23000 11280
rect 12985 11248 13327 11250
rect 12985 11192 12990 11248
rect 13046 11192 13266 11248
rect 13322 11192 13327 11248
rect 12985 11190 13327 11192
rect 12985 11187 13051 11190
rect 13261 11187 13327 11190
rect 13494 11190 23000 11250
rect 12566 11052 12572 11116
rect 12636 11114 12642 11116
rect 13494 11114 13554 11190
rect 22200 11160 23000 11190
rect 12636 11054 13554 11114
rect 13813 11114 13879 11117
rect 17902 11114 17908 11116
rect 13813 11112 17908 11114
rect 13813 11056 13818 11112
rect 13874 11056 17908 11112
rect 13813 11054 17908 11056
rect 12636 11052 12642 11054
rect 13813 11051 13879 11054
rect 17902 11052 17908 11054
rect 17972 11052 17978 11116
rect 16389 10978 16455 10981
rect 12436 10976 16455 10978
rect 12436 10920 16394 10976
rect 16450 10920 16455 10976
rect 12436 10918 16455 10920
rect 16389 10915 16455 10918
rect 4409 10912 4729 10913
rect 0 10842 800 10872
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 10847 4729 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 18270 10912 18590 10913
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 18270 10847 18590 10848
rect 5901 10842 5967 10845
rect 8661 10842 8727 10845
rect 0 10782 4216 10842
rect 0 10752 800 10782
rect 4156 10706 4216 10782
rect 5901 10840 8727 10842
rect 5901 10784 5906 10840
rect 5962 10784 8666 10840
rect 8722 10784 8727 10840
rect 5901 10782 8727 10784
rect 5901 10779 5967 10782
rect 8661 10779 8727 10782
rect 8845 10842 8911 10845
rect 10869 10842 10935 10845
rect 8845 10840 10935 10842
rect 8845 10784 8850 10840
rect 8906 10784 10874 10840
rect 10930 10784 10935 10840
rect 8845 10782 10935 10784
rect 8845 10779 8911 10782
rect 10869 10779 10935 10782
rect 12065 10842 12131 10845
rect 15285 10842 15351 10845
rect 12065 10840 15351 10842
rect 12065 10784 12070 10840
rect 12126 10784 15290 10840
rect 15346 10784 15351 10840
rect 12065 10782 15351 10784
rect 12065 10779 12131 10782
rect 15285 10779 15351 10782
rect 17902 10780 17908 10844
rect 17972 10842 17978 10844
rect 22200 10842 23000 10872
rect 17972 10782 18108 10842
rect 17972 10780 17978 10782
rect 8477 10706 8543 10709
rect 4156 10704 8543 10706
rect 4156 10648 8482 10704
rect 8538 10648 8543 10704
rect 4156 10646 8543 10648
rect 8477 10643 8543 10646
rect 8753 10706 8819 10709
rect 10358 10706 10364 10708
rect 8753 10704 10364 10706
rect 8753 10648 8758 10704
rect 8814 10648 10364 10704
rect 8753 10646 10364 10648
rect 8753 10643 8819 10646
rect 10358 10644 10364 10646
rect 10428 10706 10434 10708
rect 10501 10706 10567 10709
rect 18048 10706 18108 10782
rect 22142 10752 23000 10842
rect 22142 10706 22202 10752
rect 10428 10704 17970 10706
rect 10428 10648 10506 10704
rect 10562 10648 17970 10704
rect 10428 10646 17970 10648
rect 18048 10646 22202 10706
rect 10428 10644 10434 10646
rect 10501 10643 10567 10646
rect 6821 10570 6887 10573
rect 17769 10570 17835 10573
rect 6821 10568 17835 10570
rect 6821 10512 6826 10568
rect 6882 10512 17774 10568
rect 17830 10512 17835 10568
rect 6821 10510 17835 10512
rect 6821 10507 6887 10510
rect 17769 10507 17835 10510
rect 0 10434 800 10464
rect 5901 10434 5967 10437
rect 0 10432 5967 10434
rect 0 10376 5906 10432
rect 5962 10376 5967 10432
rect 0 10374 5967 10376
rect 0 10344 800 10374
rect 5901 10371 5967 10374
rect 7465 10434 7531 10437
rect 7598 10434 7604 10436
rect 7465 10432 7604 10434
rect 7465 10376 7470 10432
rect 7526 10376 7604 10432
rect 7465 10374 7604 10376
rect 7465 10371 7531 10374
rect 7598 10372 7604 10374
rect 7668 10372 7674 10436
rect 8937 10434 9003 10437
rect 9765 10436 9831 10437
rect 11145 10436 11211 10437
rect 9438 10434 9444 10436
rect 8937 10432 9444 10434
rect 8937 10376 8942 10432
rect 8998 10376 9444 10432
rect 8937 10374 9444 10376
rect 8937 10371 9003 10374
rect 9438 10372 9444 10374
rect 9508 10372 9514 10436
rect 9765 10432 9812 10436
rect 9876 10434 9882 10436
rect 9765 10376 9770 10432
rect 9765 10372 9812 10376
rect 9876 10374 9922 10434
rect 9876 10372 9882 10374
rect 11094 10372 11100 10436
rect 11164 10434 11211 10436
rect 11513 10434 11579 10437
rect 12065 10434 12131 10437
rect 11164 10432 11256 10434
rect 11206 10376 11256 10432
rect 11164 10374 11256 10376
rect 11513 10432 12131 10434
rect 11513 10376 11518 10432
rect 11574 10376 12070 10432
rect 12126 10376 12131 10432
rect 11513 10374 12131 10376
rect 17910 10434 17970 10646
rect 22200 10434 23000 10464
rect 17910 10374 23000 10434
rect 11164 10372 11211 10374
rect 9765 10371 9831 10372
rect 11145 10371 11211 10372
rect 11513 10371 11579 10374
rect 12065 10371 12131 10374
rect 7874 10368 8194 10369
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8194 10368
rect 7874 10303 8194 10304
rect 14805 10368 15125 10369
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 22200 10344 23000 10374
rect 14805 10303 15125 10304
rect 5993 10298 6059 10301
rect 7046 10298 7052 10300
rect 5993 10296 7052 10298
rect 5993 10240 5998 10296
rect 6054 10240 7052 10296
rect 5993 10238 7052 10240
rect 5993 10235 6059 10238
rect 7046 10236 7052 10238
rect 7116 10236 7122 10300
rect 8753 10298 8819 10301
rect 8886 10298 8892 10300
rect 8753 10296 8892 10298
rect 8753 10240 8758 10296
rect 8814 10240 8892 10296
rect 8753 10238 8892 10240
rect 8753 10235 8819 10238
rect 8886 10236 8892 10238
rect 8956 10236 8962 10300
rect 9622 10236 9628 10300
rect 9692 10298 9698 10300
rect 11830 10298 11836 10300
rect 9692 10238 11836 10298
rect 9692 10236 9698 10238
rect 11830 10236 11836 10238
rect 11900 10236 11906 10300
rect 17902 10236 17908 10300
rect 17972 10298 17978 10300
rect 20161 10298 20227 10301
rect 17972 10296 20227 10298
rect 17972 10240 20166 10296
rect 20222 10240 20227 10296
rect 17972 10238 20227 10240
rect 17972 10236 17978 10238
rect 20161 10235 20227 10238
rect 9213 10162 9279 10165
rect 9032 10160 9279 10162
rect 9032 10104 9218 10160
rect 9274 10104 9279 10160
rect 9032 10102 9279 10104
rect 4153 10026 4219 10029
rect 9032 10026 9092 10102
rect 9213 10099 9279 10102
rect 11881 10162 11947 10165
rect 15469 10162 15535 10165
rect 11881 10160 15535 10162
rect 11881 10104 11886 10160
rect 11942 10104 15474 10160
rect 15530 10104 15535 10160
rect 11881 10102 15535 10104
rect 11881 10099 11947 10102
rect 15469 10099 15535 10102
rect 4153 10024 9092 10026
rect 4153 9968 4158 10024
rect 4214 9968 9092 10024
rect 4153 9966 9092 9968
rect 4153 9963 4219 9966
rect 9254 9964 9260 10028
rect 9324 10026 9330 10028
rect 14549 10026 14615 10029
rect 9324 10024 14615 10026
rect 9324 9968 14554 10024
rect 14610 9968 14615 10024
rect 9324 9966 14615 9968
rect 9324 9964 9330 9966
rect 14549 9963 14615 9966
rect 15745 10026 15811 10029
rect 17902 10026 17908 10028
rect 15745 10024 17908 10026
rect 15745 9968 15750 10024
rect 15806 9968 17908 10024
rect 15745 9966 17908 9968
rect 15745 9963 15811 9966
rect 17902 9964 17908 9966
rect 17972 9964 17978 10028
rect 20161 10026 20227 10029
rect 20161 10024 22202 10026
rect 20161 9968 20166 10024
rect 20222 9968 22202 10024
rect 20161 9966 22202 9968
rect 20161 9963 20227 9966
rect 22142 9920 22202 9966
rect 0 9890 800 9920
rect 1393 9890 1459 9893
rect 0 9888 1459 9890
rect 0 9832 1398 9888
rect 1454 9832 1459 9888
rect 0 9830 1459 9832
rect 0 9800 800 9830
rect 1393 9827 1459 9830
rect 5717 9890 5783 9893
rect 9213 9890 9279 9893
rect 10685 9890 10751 9893
rect 5717 9888 10751 9890
rect 5717 9832 5722 9888
rect 5778 9832 9218 9888
rect 9274 9832 10690 9888
rect 10746 9832 10751 9888
rect 5717 9830 10751 9832
rect 5717 9827 5783 9830
rect 9213 9827 9279 9830
rect 10685 9827 10751 9830
rect 12341 9890 12407 9893
rect 13353 9890 13419 9893
rect 12341 9888 13419 9890
rect 12341 9832 12346 9888
rect 12402 9832 13358 9888
rect 13414 9832 13419 9888
rect 12341 9830 13419 9832
rect 12341 9827 12407 9830
rect 13353 9827 13419 9830
rect 14825 9890 14891 9893
rect 17309 9890 17375 9893
rect 14825 9888 17375 9890
rect 14825 9832 14830 9888
rect 14886 9832 17314 9888
rect 17370 9832 17375 9888
rect 14825 9830 17375 9832
rect 22142 9830 23000 9920
rect 14825 9827 14891 9830
rect 17309 9827 17375 9830
rect 4409 9824 4729 9825
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 9759 4729 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 18270 9824 18590 9825
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 22200 9800 23000 9830
rect 18270 9759 18590 9760
rect 5717 9756 5783 9757
rect 5717 9752 5764 9756
rect 5828 9754 5834 9756
rect 6085 9754 6151 9757
rect 6361 9754 6427 9757
rect 8293 9754 8359 9757
rect 5717 9696 5722 9752
rect 5717 9692 5764 9696
rect 5828 9694 5874 9754
rect 6085 9752 8359 9754
rect 6085 9696 6090 9752
rect 6146 9696 6366 9752
rect 6422 9696 8298 9752
rect 8354 9696 8359 9752
rect 6085 9694 8359 9696
rect 5828 9692 5834 9694
rect 5717 9691 5783 9692
rect 6085 9691 6151 9694
rect 6361 9691 6427 9694
rect 8293 9691 8359 9694
rect 8937 9754 9003 9757
rect 9305 9754 9371 9757
rect 10409 9756 10475 9757
rect 10358 9754 10364 9756
rect 8937 9752 9371 9754
rect 8937 9696 8942 9752
rect 8998 9696 9310 9752
rect 9366 9696 9371 9752
rect 8937 9694 9371 9696
rect 10318 9694 10364 9754
rect 10428 9752 10475 9756
rect 10470 9696 10475 9752
rect 8937 9691 9003 9694
rect 9305 9691 9371 9694
rect 10358 9692 10364 9694
rect 10428 9692 10475 9696
rect 10409 9691 10475 9692
rect 11881 9754 11947 9757
rect 15377 9754 15443 9757
rect 11881 9752 15443 9754
rect 11881 9696 11886 9752
rect 11942 9696 15382 9752
rect 15438 9696 15443 9752
rect 11881 9694 15443 9696
rect 11881 9691 11947 9694
rect 15377 9691 15443 9694
rect 16941 9754 17007 9757
rect 17861 9754 17927 9757
rect 16941 9752 17927 9754
rect 16941 9696 16946 9752
rect 17002 9696 17866 9752
rect 17922 9696 17927 9752
rect 16941 9694 17927 9696
rect 16941 9691 17007 9694
rect 17861 9691 17927 9694
rect 12525 9618 12591 9621
rect 7606 9616 12591 9618
rect 7606 9560 12530 9616
rect 12586 9560 12591 9616
rect 7606 9558 12591 9560
rect 0 9482 800 9512
rect 3601 9482 3667 9485
rect 0 9480 3667 9482
rect 0 9424 3606 9480
rect 3662 9424 3667 9480
rect 0 9422 3667 9424
rect 0 9392 800 9422
rect 3601 9419 3667 9422
rect 0 9074 800 9104
rect 7606 9074 7666 9558
rect 12525 9555 12591 9558
rect 12801 9618 12867 9621
rect 15193 9618 15259 9621
rect 19149 9618 19215 9621
rect 12801 9616 13738 9618
rect 12801 9560 12806 9616
rect 12862 9560 13738 9616
rect 12801 9558 13738 9560
rect 12801 9555 12867 9558
rect 7925 9482 7991 9485
rect 13353 9482 13419 9485
rect 7925 9480 13419 9482
rect 7925 9424 7930 9480
rect 7986 9424 13358 9480
rect 13414 9424 13419 9480
rect 7925 9422 13419 9424
rect 13678 9482 13738 9558
rect 15193 9616 19215 9618
rect 15193 9560 15198 9616
rect 15254 9560 19154 9616
rect 19210 9560 19215 9616
rect 15193 9558 19215 9560
rect 15193 9555 15259 9558
rect 19149 9555 19215 9558
rect 15469 9482 15535 9485
rect 13678 9480 15535 9482
rect 13678 9424 15474 9480
rect 15530 9424 15535 9480
rect 13678 9422 15535 9424
rect 7925 9419 7991 9422
rect 13353 9419 13419 9422
rect 15469 9419 15535 9422
rect 15929 9482 15995 9485
rect 22200 9482 23000 9512
rect 15929 9480 23000 9482
rect 15929 9424 15934 9480
rect 15990 9424 23000 9480
rect 15929 9422 23000 9424
rect 15929 9419 15995 9422
rect 22200 9392 23000 9422
rect 8293 9346 8359 9349
rect 11881 9346 11947 9349
rect 8293 9344 11947 9346
rect 8293 9288 8298 9344
rect 8354 9288 11886 9344
rect 11942 9288 11947 9344
rect 8293 9286 11947 9288
rect 8293 9283 8359 9286
rect 11881 9283 11947 9286
rect 12566 9284 12572 9348
rect 12636 9346 12642 9348
rect 12709 9346 12775 9349
rect 12636 9344 12775 9346
rect 12636 9288 12714 9344
rect 12770 9288 12775 9344
rect 12636 9286 12775 9288
rect 12636 9284 12642 9286
rect 12709 9283 12775 9286
rect 13169 9346 13235 9349
rect 13169 9344 14428 9346
rect 13169 9288 13174 9344
rect 13230 9288 14428 9344
rect 13169 9286 14428 9288
rect 13169 9283 13235 9286
rect 7874 9280 8194 9281
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8194 9280
rect 7874 9215 8194 9216
rect 9029 9210 9095 9213
rect 9305 9210 9371 9213
rect 11973 9210 12039 9213
rect 9029 9208 12039 9210
rect 9029 9152 9034 9208
rect 9090 9152 9310 9208
rect 9366 9152 11978 9208
rect 12034 9152 12039 9208
rect 9029 9150 12039 9152
rect 9029 9147 9095 9150
rect 9305 9147 9371 9150
rect 11973 9147 12039 9150
rect 12525 9210 12591 9213
rect 13077 9210 13143 9213
rect 14038 9210 14044 9212
rect 12525 9208 14044 9210
rect 12525 9152 12530 9208
rect 12586 9152 13082 9208
rect 13138 9152 14044 9208
rect 12525 9150 14044 9152
rect 12525 9147 12591 9150
rect 13077 9147 13143 9150
rect 14038 9148 14044 9150
rect 14108 9148 14114 9212
rect 0 9014 7666 9074
rect 8201 9074 8267 9077
rect 13813 9074 13879 9077
rect 14181 9074 14247 9077
rect 8201 9072 14247 9074
rect 8201 9016 8206 9072
rect 8262 9016 13818 9072
rect 13874 9016 14186 9072
rect 14242 9016 14247 9072
rect 8201 9014 14247 9016
rect 14368 9074 14428 9286
rect 14805 9280 15125 9281
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 9215 15125 9216
rect 16113 9210 16179 9213
rect 16481 9210 16547 9213
rect 16113 9208 16547 9210
rect 16113 9152 16118 9208
rect 16174 9152 16486 9208
rect 16542 9152 16547 9208
rect 16113 9150 16547 9152
rect 16113 9147 16179 9150
rect 16481 9147 16547 9150
rect 19057 9210 19123 9213
rect 19190 9210 19196 9212
rect 19057 9208 19196 9210
rect 19057 9152 19062 9208
rect 19118 9152 19196 9208
rect 19057 9150 19196 9152
rect 19057 9147 19123 9150
rect 19190 9148 19196 9150
rect 19260 9148 19266 9212
rect 22200 9074 23000 9104
rect 14368 9014 23000 9074
rect 0 8984 800 9014
rect 8201 9011 8267 9014
rect 13813 9011 13879 9014
rect 14181 9011 14247 9014
rect 22200 8984 23000 9014
rect 3417 8940 3483 8941
rect 3366 8876 3372 8940
rect 3436 8938 3483 8940
rect 6637 8938 6703 8941
rect 3436 8936 3528 8938
rect 3478 8880 3528 8936
rect 3436 8878 3528 8880
rect 4156 8936 6703 8938
rect 4156 8880 6642 8936
rect 6698 8880 6703 8936
rect 4156 8878 6703 8880
rect 3436 8876 3483 8878
rect 3417 8875 3483 8876
rect 0 8666 800 8696
rect 4156 8666 4216 8878
rect 6637 8875 6703 8878
rect 7465 8938 7531 8941
rect 11237 8938 11303 8941
rect 7465 8936 11303 8938
rect 7465 8880 7470 8936
rect 7526 8880 11242 8936
rect 11298 8880 11303 8936
rect 7465 8878 11303 8880
rect 7465 8875 7531 8878
rect 11237 8875 11303 8878
rect 11421 8938 11487 8941
rect 17769 8938 17835 8941
rect 11421 8936 17835 8938
rect 11421 8880 11426 8936
rect 11482 8880 17774 8936
rect 17830 8880 17835 8936
rect 11421 8878 17835 8880
rect 11421 8875 11487 8878
rect 17769 8875 17835 8878
rect 7230 8740 7236 8804
rect 7300 8802 7306 8804
rect 11094 8802 11100 8804
rect 7300 8742 11100 8802
rect 7300 8740 7306 8742
rect 11094 8740 11100 8742
rect 11164 8740 11170 8804
rect 14825 8802 14891 8805
rect 16205 8802 16271 8805
rect 14825 8800 16271 8802
rect 14825 8744 14830 8800
rect 14886 8744 16210 8800
rect 16266 8744 16271 8800
rect 14825 8742 16271 8744
rect 14825 8739 14891 8742
rect 16205 8739 16271 8742
rect 4409 8736 4729 8737
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 8671 4729 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 18270 8736 18590 8737
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 8671 18590 8672
rect 0 8606 4216 8666
rect 6085 8666 6151 8669
rect 11053 8666 11119 8669
rect 6085 8664 11119 8666
rect 6085 8608 6090 8664
rect 6146 8608 11058 8664
rect 11114 8608 11119 8664
rect 6085 8606 11119 8608
rect 0 8576 800 8606
rect 6085 8603 6151 8606
rect 11053 8603 11119 8606
rect 13077 8668 13143 8669
rect 13077 8664 13124 8668
rect 13188 8666 13194 8668
rect 13077 8608 13082 8664
rect 13077 8604 13124 8608
rect 13188 8606 13234 8666
rect 13188 8604 13194 8606
rect 18822 8604 18828 8668
rect 18892 8666 18898 8668
rect 22200 8666 23000 8696
rect 18892 8606 23000 8666
rect 18892 8604 18898 8606
rect 13077 8603 13143 8604
rect 22200 8576 23000 8606
rect 7598 8468 7604 8532
rect 7668 8530 7674 8532
rect 11881 8530 11947 8533
rect 7668 8528 11947 8530
rect 7668 8472 11886 8528
rect 11942 8472 11947 8528
rect 7668 8470 11947 8472
rect 7668 8468 7674 8470
rect 11881 8467 11947 8470
rect 12341 8530 12407 8533
rect 13169 8530 13235 8533
rect 12341 8528 13235 8530
rect 12341 8472 12346 8528
rect 12402 8472 13174 8528
rect 13230 8472 13235 8528
rect 12341 8470 13235 8472
rect 12341 8467 12407 8470
rect 13169 8467 13235 8470
rect 14917 8530 14983 8533
rect 18505 8530 18571 8533
rect 19333 8530 19399 8533
rect 14917 8528 19399 8530
rect 14917 8472 14922 8528
rect 14978 8472 18510 8528
rect 18566 8472 19338 8528
rect 19394 8472 19399 8528
rect 14917 8470 19399 8472
rect 14917 8467 14983 8470
rect 18505 8467 18571 8470
rect 19333 8467 19399 8470
rect 7414 8332 7420 8396
rect 7484 8394 7490 8396
rect 7925 8394 7991 8397
rect 10133 8394 10199 8397
rect 10593 8396 10659 8397
rect 10542 8394 10548 8396
rect 7484 8334 7712 8394
rect 7484 8332 7490 8334
rect 0 8258 800 8288
rect 7652 8261 7712 8334
rect 7925 8392 10199 8394
rect 7925 8336 7930 8392
rect 7986 8336 10138 8392
rect 10194 8336 10199 8392
rect 7925 8334 10199 8336
rect 10502 8334 10548 8394
rect 10612 8392 10659 8396
rect 10654 8336 10659 8392
rect 7925 8331 7991 8334
rect 10133 8331 10199 8334
rect 10542 8332 10548 8334
rect 10612 8332 10659 8336
rect 10593 8331 10659 8332
rect 10961 8394 11027 8397
rect 12433 8394 12499 8397
rect 13077 8396 13143 8397
rect 13077 8394 13124 8396
rect 10961 8392 12499 8394
rect 10961 8336 10966 8392
rect 11022 8336 12438 8392
rect 12494 8336 12499 8392
rect 10961 8334 12499 8336
rect 13032 8392 13124 8394
rect 13032 8336 13082 8392
rect 13032 8334 13124 8336
rect 10961 8331 11027 8334
rect 12433 8331 12499 8334
rect 13077 8332 13124 8334
rect 13188 8332 13194 8396
rect 14641 8394 14707 8397
rect 18822 8394 18828 8396
rect 14641 8392 18828 8394
rect 14641 8336 14646 8392
rect 14702 8336 18828 8392
rect 14641 8334 18828 8336
rect 13077 8331 13143 8332
rect 14641 8331 14707 8334
rect 18822 8332 18828 8334
rect 18892 8332 18898 8396
rect 0 8198 5274 8258
rect 0 8168 800 8198
rect 0 7850 800 7880
rect 4061 7850 4127 7853
rect 0 7848 4127 7850
rect 0 7792 4066 7848
rect 4122 7792 4127 7848
rect 0 7790 4127 7792
rect 0 7760 800 7790
rect 4061 7787 4127 7790
rect 2865 7714 2931 7717
rect 3785 7714 3851 7717
rect 5214 7714 5274 8198
rect 7649 8256 7715 8261
rect 7649 8200 7654 8256
rect 7710 8200 7715 8256
rect 7649 8195 7715 8200
rect 8385 8258 8451 8261
rect 10910 8258 10916 8260
rect 8385 8256 10916 8258
rect 8385 8200 8390 8256
rect 8446 8200 10916 8256
rect 8385 8198 10916 8200
rect 8385 8195 8451 8198
rect 10910 8196 10916 8198
rect 10980 8196 10986 8260
rect 11973 8258 12039 8261
rect 14549 8258 14615 8261
rect 11973 8256 14615 8258
rect 11973 8200 11978 8256
rect 12034 8200 14554 8256
rect 14610 8200 14615 8256
rect 11973 8198 14615 8200
rect 11973 8195 12039 8198
rect 14549 8195 14615 8198
rect 15469 8258 15535 8261
rect 15653 8258 15719 8261
rect 22200 8258 23000 8288
rect 15469 8256 23000 8258
rect 15469 8200 15474 8256
rect 15530 8200 15658 8256
rect 15714 8200 23000 8256
rect 15469 8198 23000 8200
rect 15469 8195 15535 8198
rect 15653 8195 15719 8198
rect 7874 8192 8194 8193
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8194 8192
rect 7874 8127 8194 8128
rect 14805 8192 15125 8193
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 22200 8168 23000 8198
rect 14805 8127 15125 8128
rect 8937 8122 9003 8125
rect 16297 8122 16363 8125
rect 17125 8122 17191 8125
rect 8937 8120 14244 8122
rect 8937 8064 8942 8120
rect 8998 8064 14244 8120
rect 8937 8062 14244 8064
rect 8937 8059 9003 8062
rect 5349 7986 5415 7989
rect 13261 7986 13327 7989
rect 13997 7986 14063 7989
rect 5349 7984 12220 7986
rect 5349 7928 5354 7984
rect 5410 7928 12220 7984
rect 5349 7926 12220 7928
rect 5349 7923 5415 7926
rect 5625 7850 5691 7853
rect 8518 7850 8524 7852
rect 5625 7848 8524 7850
rect 5625 7792 5630 7848
rect 5686 7792 8524 7848
rect 5625 7790 8524 7792
rect 5625 7787 5691 7790
rect 8518 7788 8524 7790
rect 8588 7788 8594 7852
rect 9489 7850 9555 7853
rect 10409 7850 10475 7853
rect 9489 7848 10475 7850
rect 9489 7792 9494 7848
rect 9550 7792 10414 7848
rect 10470 7792 10475 7848
rect 9489 7790 10475 7792
rect 9489 7787 9555 7790
rect 10409 7787 10475 7790
rect 11237 7850 11303 7853
rect 12160 7850 12220 7926
rect 13261 7984 14063 7986
rect 13261 7928 13266 7984
rect 13322 7928 14002 7984
rect 14058 7928 14063 7984
rect 13261 7926 14063 7928
rect 14184 7986 14244 8062
rect 16297 8120 17191 8122
rect 16297 8064 16302 8120
rect 16358 8064 17130 8120
rect 17186 8064 17191 8120
rect 16297 8062 17191 8064
rect 16297 8059 16363 8062
rect 17125 8059 17191 8062
rect 16113 7986 16179 7989
rect 14184 7984 16179 7986
rect 14184 7928 16118 7984
rect 16174 7928 16179 7984
rect 14184 7926 16179 7928
rect 13261 7923 13327 7926
rect 13997 7923 14063 7926
rect 16113 7923 16179 7926
rect 14273 7850 14339 7853
rect 11237 7848 12082 7850
rect 11237 7792 11242 7848
rect 11298 7792 12082 7848
rect 11237 7790 12082 7792
rect 12160 7848 14339 7850
rect 12160 7792 14278 7848
rect 14334 7792 14339 7848
rect 12160 7790 14339 7792
rect 11237 7787 11303 7790
rect 8569 7714 8635 7717
rect 2865 7712 4170 7714
rect 2865 7656 2870 7712
rect 2926 7656 3790 7712
rect 3846 7656 4170 7712
rect 2865 7654 4170 7656
rect 5214 7712 8635 7714
rect 5214 7656 8574 7712
rect 8630 7656 8635 7712
rect 5214 7654 8635 7656
rect 12022 7714 12082 7790
rect 14273 7787 14339 7790
rect 16021 7850 16087 7853
rect 22200 7850 23000 7880
rect 16021 7848 23000 7850
rect 16021 7792 16026 7848
rect 16082 7792 23000 7848
rect 16021 7790 23000 7792
rect 16021 7787 16087 7790
rect 22200 7760 23000 7790
rect 12893 7714 12959 7717
rect 12022 7712 12959 7714
rect 12022 7656 12898 7712
rect 12954 7656 12959 7712
rect 12022 7654 12959 7656
rect 2865 7651 2931 7654
rect 3785 7651 3851 7654
rect 0 7442 800 7472
rect 3969 7442 4035 7445
rect 0 7440 4035 7442
rect 0 7384 3974 7440
rect 4030 7384 4035 7440
rect 0 7382 4035 7384
rect 0 7352 800 7382
rect 3969 7379 4035 7382
rect 4110 7306 4170 7654
rect 8569 7651 8635 7654
rect 12893 7651 12959 7654
rect 13261 7714 13327 7717
rect 17401 7714 17467 7717
rect 13261 7712 17467 7714
rect 13261 7656 13266 7712
rect 13322 7656 17406 7712
rect 17462 7656 17467 7712
rect 13261 7654 17467 7656
rect 13261 7651 13327 7654
rect 17401 7651 17467 7654
rect 4409 7648 4729 7649
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 7583 4729 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 18270 7648 18590 7649
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 18270 7583 18590 7584
rect 16205 7578 16271 7581
rect 13126 7576 16271 7578
rect 13126 7520 16210 7576
rect 16266 7520 16271 7576
rect 13126 7518 16271 7520
rect 6269 7442 6335 7445
rect 7557 7442 7623 7445
rect 9581 7442 9647 7445
rect 6269 7440 9647 7442
rect 6269 7384 6274 7440
rect 6330 7384 7562 7440
rect 7618 7384 9586 7440
rect 9642 7384 9647 7440
rect 6269 7382 9647 7384
rect 6269 7379 6335 7382
rect 7557 7379 7623 7382
rect 9581 7379 9647 7382
rect 10869 7442 10935 7445
rect 13126 7442 13186 7518
rect 16205 7515 16271 7518
rect 18781 7578 18847 7581
rect 18781 7576 19074 7578
rect 18781 7520 18786 7576
rect 18842 7520 19074 7576
rect 18781 7518 19074 7520
rect 18781 7515 18847 7518
rect 10869 7440 13186 7442
rect 10869 7384 10874 7440
rect 10930 7384 13186 7440
rect 10869 7382 13186 7384
rect 13353 7442 13419 7445
rect 16849 7442 16915 7445
rect 13353 7440 16915 7442
rect 13353 7384 13358 7440
rect 13414 7384 16854 7440
rect 16910 7384 16915 7440
rect 13353 7382 16915 7384
rect 19014 7442 19074 7518
rect 22200 7442 23000 7472
rect 19014 7382 23000 7442
rect 10869 7379 10935 7382
rect 13353 7379 13419 7382
rect 16849 7379 16915 7382
rect 22200 7352 23000 7382
rect 13261 7306 13327 7309
rect 13721 7306 13787 7309
rect 14457 7306 14523 7309
rect 4110 7304 13327 7306
rect 4110 7248 13266 7304
rect 13322 7248 13327 7304
rect 4110 7246 13327 7248
rect 13261 7243 13327 7246
rect 13494 7304 14523 7306
rect 13494 7248 13726 7304
rect 13782 7248 14462 7304
rect 14518 7248 14523 7304
rect 13494 7246 14523 7248
rect 11094 7108 11100 7172
rect 11164 7170 11170 7172
rect 11881 7170 11947 7173
rect 11164 7168 11947 7170
rect 11164 7112 11886 7168
rect 11942 7112 11947 7168
rect 11164 7110 11947 7112
rect 11164 7108 11170 7110
rect 11881 7107 11947 7110
rect 12065 7170 12131 7173
rect 13494 7170 13554 7246
rect 13721 7243 13787 7246
rect 14457 7243 14523 7246
rect 12065 7168 13554 7170
rect 12065 7112 12070 7168
rect 12126 7112 13554 7168
rect 12065 7110 13554 7112
rect 12065 7107 12131 7110
rect 7874 7104 8194 7105
rect 0 7034 800 7064
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8194 7104
rect 7874 7039 8194 7040
rect 14805 7104 15125 7105
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 7039 15125 7040
rect 6453 7034 6519 7037
rect 0 7032 6519 7034
rect 0 6976 6458 7032
rect 6514 6976 6519 7032
rect 0 6974 6519 6976
rect 0 6944 800 6974
rect 6453 6971 6519 6974
rect 10409 7034 10475 7037
rect 17309 7034 17375 7037
rect 22200 7034 23000 7064
rect 10409 7032 13922 7034
rect 10409 6976 10414 7032
rect 10470 6976 13922 7032
rect 10409 6974 13922 6976
rect 10409 6971 10475 6974
rect 7097 6898 7163 6901
rect 8017 6898 8083 6901
rect 13721 6898 13787 6901
rect 7097 6896 13787 6898
rect 7097 6840 7102 6896
rect 7158 6840 8022 6896
rect 8078 6840 13726 6896
rect 13782 6840 13787 6896
rect 7097 6838 13787 6840
rect 13862 6898 13922 6974
rect 17309 7032 23000 7034
rect 17309 6976 17314 7032
rect 17370 6976 23000 7032
rect 17309 6974 23000 6976
rect 17309 6971 17375 6974
rect 22200 6944 23000 6974
rect 15653 6898 15719 6901
rect 13862 6896 15719 6898
rect 13862 6840 15658 6896
rect 15714 6840 15719 6896
rect 13862 6838 15719 6840
rect 7097 6835 7163 6838
rect 8017 6835 8083 6838
rect 13721 6835 13787 6838
rect 15653 6835 15719 6838
rect 6637 6762 6703 6765
rect 7833 6762 7899 6765
rect 6637 6760 7899 6762
rect 6637 6704 6642 6760
rect 6698 6704 7838 6760
rect 7894 6704 7899 6760
rect 6637 6702 7899 6704
rect 6637 6699 6703 6702
rect 7833 6699 7899 6702
rect 10685 6762 10751 6765
rect 12617 6762 12683 6765
rect 10685 6760 11898 6762
rect 10685 6704 10690 6760
rect 10746 6704 11898 6760
rect 10685 6702 11898 6704
rect 10685 6699 10751 6702
rect 7833 6626 7899 6629
rect 9397 6626 9463 6629
rect 7833 6624 9463 6626
rect 7833 6568 7838 6624
rect 7894 6568 9402 6624
rect 9458 6568 9463 6624
rect 7833 6566 9463 6568
rect 11838 6626 11898 6702
rect 12617 6760 18752 6762
rect 12617 6704 12622 6760
rect 12678 6704 18752 6760
rect 12617 6702 18752 6704
rect 12617 6699 12683 6702
rect 16481 6626 16547 6629
rect 11838 6624 16547 6626
rect 11838 6568 16486 6624
rect 16542 6568 16547 6624
rect 11838 6566 16547 6568
rect 7833 6563 7899 6566
rect 9397 6563 9463 6566
rect 16481 6563 16547 6566
rect 4409 6560 4729 6561
rect 0 6490 800 6520
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 6495 4729 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 18270 6560 18590 6561
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 6495 18590 6496
rect 4061 6490 4127 6493
rect 0 6488 4127 6490
rect 0 6432 4066 6488
rect 4122 6432 4127 6488
rect 0 6430 4127 6432
rect 0 6400 800 6430
rect 4061 6427 4127 6430
rect 5165 6490 5231 6493
rect 7373 6490 7439 6493
rect 11973 6492 12039 6493
rect 11973 6490 12020 6492
rect 5165 6488 7439 6490
rect 5165 6432 5170 6488
rect 5226 6432 7378 6488
rect 7434 6432 7439 6488
rect 5165 6430 7439 6432
rect 11928 6488 12020 6490
rect 11928 6432 11978 6488
rect 11928 6430 12020 6432
rect 5165 6427 5231 6430
rect 7373 6427 7439 6430
rect 11973 6428 12020 6430
rect 12084 6428 12090 6492
rect 18692 6490 18752 6702
rect 19149 6628 19215 6629
rect 19149 6626 19196 6628
rect 19104 6624 19196 6626
rect 19104 6568 19154 6624
rect 19104 6566 19196 6568
rect 19149 6564 19196 6566
rect 19260 6564 19266 6628
rect 19149 6563 19215 6564
rect 22200 6490 23000 6520
rect 18692 6430 23000 6490
rect 11973 6427 12039 6428
rect 22200 6400 23000 6430
rect 6361 6354 6427 6357
rect 8109 6354 8175 6357
rect 19425 6354 19491 6357
rect 6361 6352 7666 6354
rect 6361 6296 6366 6352
rect 6422 6296 7666 6352
rect 6361 6294 7666 6296
rect 6361 6291 6427 6294
rect 7230 6156 7236 6220
rect 7300 6218 7306 6220
rect 7373 6218 7439 6221
rect 7300 6216 7439 6218
rect 7300 6160 7378 6216
rect 7434 6160 7439 6216
rect 7300 6158 7439 6160
rect 7606 6218 7666 6294
rect 8109 6352 19491 6354
rect 8109 6296 8114 6352
rect 8170 6296 19430 6352
rect 19486 6296 19491 6352
rect 8109 6294 19491 6296
rect 8109 6291 8175 6294
rect 19425 6291 19491 6294
rect 17677 6218 17743 6221
rect 7606 6216 17743 6218
rect 7606 6160 17682 6216
rect 17738 6160 17743 6216
rect 7606 6158 17743 6160
rect 7300 6156 7306 6158
rect 7373 6155 7439 6158
rect 17677 6155 17743 6158
rect 0 6082 800 6112
rect 3969 6082 4035 6085
rect 0 6080 4035 6082
rect 0 6024 3974 6080
rect 4030 6024 4035 6080
rect 0 6022 4035 6024
rect 0 5992 800 6022
rect 3969 6019 4035 6022
rect 11421 6082 11487 6085
rect 12893 6082 12959 6085
rect 11421 6080 12959 6082
rect 11421 6024 11426 6080
rect 11482 6024 12898 6080
rect 12954 6024 12959 6080
rect 11421 6022 12959 6024
rect 11421 6019 11487 6022
rect 12893 6019 12959 6022
rect 15653 6082 15719 6085
rect 22200 6082 23000 6112
rect 15653 6080 23000 6082
rect 15653 6024 15658 6080
rect 15714 6024 23000 6080
rect 15653 6022 23000 6024
rect 15653 6019 15719 6022
rect 7874 6016 8194 6017
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8194 6016
rect 7874 5951 8194 5952
rect 14805 6016 15125 6017
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 22200 5992 23000 6022
rect 14805 5951 15125 5952
rect 8569 5946 8635 5949
rect 8702 5946 8708 5948
rect 8569 5944 8708 5946
rect 8569 5888 8574 5944
rect 8630 5888 8708 5944
rect 8569 5886 8708 5888
rect 8569 5883 8635 5886
rect 8702 5884 8708 5886
rect 8772 5884 8778 5948
rect 15469 5944 15535 5949
rect 15469 5888 15474 5944
rect 15530 5888 15535 5944
rect 15469 5883 15535 5888
rect 4245 5810 4311 5813
rect 9121 5810 9187 5813
rect 4245 5808 9187 5810
rect 4245 5752 4250 5808
rect 4306 5752 9126 5808
rect 9182 5752 9187 5808
rect 4245 5750 9187 5752
rect 4245 5747 4311 5750
rect 9121 5747 9187 5750
rect 10685 5810 10751 5813
rect 15472 5810 15532 5883
rect 10685 5808 15532 5810
rect 10685 5752 10690 5808
rect 10746 5752 15532 5808
rect 10685 5750 15532 5752
rect 10685 5747 10751 5750
rect 0 5674 800 5704
rect 2865 5674 2931 5677
rect 7281 5674 7347 5677
rect 0 5672 7347 5674
rect 0 5616 2870 5672
rect 2926 5616 7286 5672
rect 7342 5616 7347 5672
rect 0 5614 7347 5616
rect 0 5584 800 5614
rect 2865 5611 2931 5614
rect 7281 5611 7347 5614
rect 9029 5674 9095 5677
rect 13905 5674 13971 5677
rect 22200 5674 23000 5704
rect 9029 5672 13971 5674
rect 9029 5616 9034 5672
rect 9090 5616 13910 5672
rect 13966 5616 13971 5672
rect 9029 5614 13971 5616
rect 9029 5611 9095 5614
rect 13905 5611 13971 5614
rect 14046 5614 23000 5674
rect 7005 5538 7071 5541
rect 9438 5538 9444 5540
rect 7005 5536 9444 5538
rect 7005 5480 7010 5536
rect 7066 5480 9444 5536
rect 7005 5478 9444 5480
rect 7005 5475 7071 5478
rect 9438 5476 9444 5478
rect 9508 5538 9514 5540
rect 9581 5538 9647 5541
rect 9508 5536 9647 5538
rect 9508 5480 9586 5536
rect 9642 5480 9647 5536
rect 9508 5478 9647 5480
rect 9508 5476 9514 5478
rect 9581 5475 9647 5478
rect 12249 5538 12315 5541
rect 14046 5538 14106 5614
rect 22200 5584 23000 5614
rect 12249 5536 14106 5538
rect 12249 5480 12254 5536
rect 12310 5480 14106 5536
rect 12249 5478 14106 5480
rect 14641 5538 14707 5541
rect 15101 5538 15167 5541
rect 14641 5536 15167 5538
rect 14641 5480 14646 5536
rect 14702 5480 15106 5536
rect 15162 5480 15167 5536
rect 14641 5478 15167 5480
rect 12249 5475 12315 5478
rect 14641 5475 14707 5478
rect 15101 5475 15167 5478
rect 4409 5472 4729 5473
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 5407 4729 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 18270 5472 18590 5473
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 5407 18590 5408
rect 7281 5402 7347 5405
rect 7598 5402 7604 5404
rect 7281 5400 7604 5402
rect 7281 5344 7286 5400
rect 7342 5344 7604 5400
rect 7281 5342 7604 5344
rect 7281 5339 7347 5342
rect 7598 5340 7604 5342
rect 7668 5340 7674 5404
rect 0 5266 800 5296
rect 12893 5266 12959 5269
rect 0 5264 12959 5266
rect 0 5208 12898 5264
rect 12954 5208 12959 5264
rect 0 5206 12959 5208
rect 0 5176 800 5206
rect 12893 5203 12959 5206
rect 13721 5266 13787 5269
rect 22200 5266 23000 5296
rect 13721 5264 23000 5266
rect 13721 5208 13726 5264
rect 13782 5208 23000 5264
rect 13721 5206 23000 5208
rect 13721 5203 13787 5206
rect 22200 5176 23000 5206
rect 11697 5130 11763 5133
rect 4846 5128 11763 5130
rect 4846 5072 11702 5128
rect 11758 5072 11763 5128
rect 4846 5070 11763 5072
rect 0 4858 800 4888
rect 4846 4858 4906 5070
rect 11697 5067 11763 5070
rect 11830 5068 11836 5132
rect 11900 5130 11906 5132
rect 15469 5130 15535 5133
rect 11900 5128 15535 5130
rect 11900 5072 15474 5128
rect 15530 5072 15535 5128
rect 11900 5070 15535 5072
rect 11900 5068 11906 5070
rect 9673 4994 9739 4997
rect 11838 4994 11898 5068
rect 15469 5067 15535 5070
rect 17861 5130 17927 5133
rect 21081 5130 21147 5133
rect 21449 5130 21515 5133
rect 17861 5128 21515 5130
rect 17861 5072 17866 5128
rect 17922 5072 21086 5128
rect 21142 5072 21454 5128
rect 21510 5072 21515 5128
rect 17861 5070 21515 5072
rect 17861 5067 17927 5070
rect 21081 5067 21147 5070
rect 21449 5067 21515 5070
rect 9673 4992 11898 4994
rect 9673 4936 9678 4992
rect 9734 4936 11898 4992
rect 9673 4934 11898 4936
rect 11973 4994 12039 4997
rect 13077 4994 13143 4997
rect 11973 4992 13143 4994
rect 11973 4936 11978 4992
rect 12034 4936 13082 4992
rect 13138 4936 13143 4992
rect 11973 4934 13143 4936
rect 9673 4931 9739 4934
rect 11973 4931 12039 4934
rect 13077 4931 13143 4934
rect 7874 4928 8194 4929
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8194 4928
rect 7874 4863 8194 4864
rect 14805 4928 15125 4929
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 4863 15125 4864
rect 0 4798 4906 4858
rect 7465 4858 7531 4861
rect 7649 4858 7715 4861
rect 9213 4858 9279 4861
rect 7465 4856 7715 4858
rect 7465 4800 7470 4856
rect 7526 4800 7654 4856
rect 7710 4800 7715 4856
rect 7465 4798 7715 4800
rect 0 4768 800 4798
rect 7465 4795 7531 4798
rect 7649 4795 7715 4798
rect 8296 4856 9279 4858
rect 8296 4800 9218 4856
rect 9274 4800 9279 4856
rect 8296 4798 9279 4800
rect 8296 4722 8356 4798
rect 9213 4795 9279 4798
rect 16481 4858 16547 4861
rect 22200 4858 23000 4888
rect 16481 4856 23000 4858
rect 16481 4800 16486 4856
rect 16542 4800 23000 4856
rect 16481 4798 23000 4800
rect 16481 4795 16547 4798
rect 22200 4768 23000 4798
rect 4156 4662 8356 4722
rect 8477 4722 8543 4725
rect 14089 4722 14155 4725
rect 8477 4720 14155 4722
rect 8477 4664 8482 4720
rect 8538 4664 14094 4720
rect 14150 4664 14155 4720
rect 8477 4662 14155 4664
rect 0 4450 800 4480
rect 4156 4450 4216 4662
rect 8477 4659 8543 4662
rect 5717 4586 5783 4589
rect 9581 4586 9647 4589
rect 5717 4584 9647 4586
rect 5717 4528 5722 4584
rect 5778 4528 9586 4584
rect 9642 4528 9647 4584
rect 5717 4526 9647 4528
rect 5717 4523 5783 4526
rect 9581 4523 9647 4526
rect 12022 4453 12082 4662
rect 14089 4659 14155 4662
rect 16021 4586 16087 4589
rect 17902 4586 17908 4588
rect 16021 4584 17908 4586
rect 16021 4528 16026 4584
rect 16082 4528 17908 4584
rect 16021 4526 17908 4528
rect 16021 4523 16087 4526
rect 17902 4524 17908 4526
rect 17972 4524 17978 4588
rect 0 4390 4216 4450
rect 11973 4448 12082 4453
rect 22200 4450 23000 4480
rect 11973 4392 11978 4448
rect 12034 4392 12082 4448
rect 11973 4390 12082 4392
rect 0 4360 800 4390
rect 11973 4387 12039 4390
rect 4409 4384 4729 4385
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 4319 4729 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 18270 4384 18590 4385
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 18270 4319 18590 4320
rect 22142 4360 23000 4450
rect 3918 4252 3924 4316
rect 3988 4314 3994 4316
rect 4245 4314 4311 4317
rect 3988 4312 4311 4314
rect 3988 4256 4250 4312
rect 4306 4256 4311 4312
rect 3988 4254 4311 4256
rect 3988 4252 3994 4254
rect 4245 4251 4311 4254
rect 5441 4314 5507 4317
rect 8569 4314 8635 4317
rect 5441 4312 8635 4314
rect 5441 4256 5446 4312
rect 5502 4256 8574 4312
rect 8630 4256 8635 4312
rect 5441 4254 8635 4256
rect 5441 4251 5507 4254
rect 8569 4251 8635 4254
rect 9121 4314 9187 4317
rect 10409 4314 10475 4317
rect 22142 4314 22202 4360
rect 9121 4312 10475 4314
rect 9121 4256 9126 4312
rect 9182 4256 10414 4312
rect 10470 4256 10475 4312
rect 9121 4254 10475 4256
rect 9121 4251 9187 4254
rect 10409 4251 10475 4254
rect 18692 4254 22202 4314
rect 5257 4178 5323 4181
rect 10961 4178 11027 4181
rect 14089 4180 14155 4181
rect 5257 4176 11027 4178
rect 5257 4120 5262 4176
rect 5318 4120 10966 4176
rect 11022 4120 11027 4176
rect 5257 4118 11027 4120
rect 5257 4115 5323 4118
rect 10961 4115 11027 4118
rect 14038 4116 14044 4180
rect 14108 4178 14155 4180
rect 14108 4176 14200 4178
rect 14150 4120 14200 4176
rect 14108 4118 14200 4120
rect 14108 4116 14155 4118
rect 17902 4116 17908 4180
rect 17972 4178 17978 4180
rect 18692 4178 18752 4254
rect 17972 4118 18752 4178
rect 17972 4116 17978 4118
rect 14089 4115 14155 4116
rect 0 4042 800 4072
rect 12065 4042 12131 4045
rect 17861 4042 17927 4045
rect 0 4040 12131 4042
rect 0 3984 12070 4040
rect 12126 3984 12131 4040
rect 0 3982 12131 3984
rect 0 3952 800 3982
rect 12065 3979 12131 3982
rect 12206 4040 17927 4042
rect 12206 3984 17866 4040
rect 17922 3984 17927 4040
rect 12206 3982 17927 3984
rect 8569 3906 8635 3909
rect 10317 3906 10383 3909
rect 8569 3904 10383 3906
rect 8569 3848 8574 3904
rect 8630 3848 10322 3904
rect 10378 3848 10383 3904
rect 8569 3846 10383 3848
rect 8569 3843 8635 3846
rect 10317 3843 10383 3846
rect 7874 3840 8194 3841
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8194 3840
rect 7874 3775 8194 3776
rect 7097 3770 7163 3773
rect 12206 3770 12266 3982
rect 17861 3979 17927 3982
rect 18965 4042 19031 4045
rect 22200 4042 23000 4072
rect 18965 4040 23000 4042
rect 18965 3984 18970 4040
rect 19026 3984 23000 4040
rect 18965 3982 23000 3984
rect 18965 3979 19031 3982
rect 22200 3952 23000 3982
rect 12801 3906 12867 3909
rect 14549 3906 14615 3909
rect 12801 3904 14615 3906
rect 12801 3848 12806 3904
rect 12862 3848 14554 3904
rect 14610 3848 14615 3904
rect 12801 3846 14615 3848
rect 12801 3843 12867 3846
rect 14549 3843 14615 3846
rect 15193 3906 15259 3909
rect 19977 3906 20043 3909
rect 15193 3904 20043 3906
rect 15193 3848 15198 3904
rect 15254 3848 19982 3904
rect 20038 3848 20043 3904
rect 15193 3846 20043 3848
rect 15193 3843 15259 3846
rect 19977 3843 20043 3846
rect 14805 3840 15125 3841
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 3775 15125 3776
rect 6134 3768 7163 3770
rect 6134 3712 7102 3768
rect 7158 3712 7163 3768
rect 6134 3710 7163 3712
rect 0 3634 800 3664
rect 6134 3634 6194 3710
rect 7097 3707 7163 3710
rect 8710 3710 12266 3770
rect 12433 3770 12499 3773
rect 14181 3770 14247 3773
rect 12433 3768 14247 3770
rect 12433 3712 12438 3768
rect 12494 3712 14186 3768
rect 14242 3712 14247 3768
rect 12433 3710 14247 3712
rect 0 3574 6194 3634
rect 6269 3634 6335 3637
rect 8569 3634 8635 3637
rect 6269 3632 8635 3634
rect 6269 3576 6274 3632
rect 6330 3576 8574 3632
rect 8630 3576 8635 3632
rect 6269 3574 8635 3576
rect 0 3544 800 3574
rect 6269 3571 6335 3574
rect 8569 3571 8635 3574
rect 6453 3498 6519 3501
rect 8293 3498 8359 3501
rect 6453 3496 8359 3498
rect 6453 3440 6458 3496
rect 6514 3440 8298 3496
rect 8354 3440 8359 3496
rect 6453 3438 8359 3440
rect 6453 3435 6519 3438
rect 8293 3435 8359 3438
rect 5993 3362 6059 3365
rect 8710 3362 8770 3710
rect 12433 3707 12499 3710
rect 14181 3707 14247 3710
rect 10225 3634 10291 3637
rect 15469 3634 15535 3637
rect 10225 3632 15535 3634
rect 10225 3576 10230 3632
rect 10286 3576 15474 3632
rect 15530 3576 15535 3632
rect 10225 3574 15535 3576
rect 10225 3571 10291 3574
rect 15469 3571 15535 3574
rect 17769 3634 17835 3637
rect 22200 3634 23000 3664
rect 17769 3632 23000 3634
rect 17769 3576 17774 3632
rect 17830 3576 23000 3632
rect 17769 3574 23000 3576
rect 17769 3571 17835 3574
rect 22200 3544 23000 3574
rect 8886 3436 8892 3500
rect 8956 3498 8962 3500
rect 9397 3498 9463 3501
rect 10685 3498 10751 3501
rect 18689 3498 18755 3501
rect 8956 3496 18755 3498
rect 8956 3440 9402 3496
rect 9458 3440 10690 3496
rect 10746 3440 18694 3496
rect 18750 3440 18755 3496
rect 8956 3438 18755 3440
rect 8956 3436 8962 3438
rect 9397 3435 9463 3438
rect 10685 3435 10751 3438
rect 18689 3435 18755 3438
rect 5993 3360 8770 3362
rect 5993 3304 5998 3360
rect 6054 3304 8770 3360
rect 5993 3302 8770 3304
rect 8937 3362 9003 3365
rect 10869 3362 10935 3365
rect 8937 3360 10935 3362
rect 8937 3304 8942 3360
rect 8998 3304 10874 3360
rect 10930 3304 10935 3360
rect 8937 3302 10935 3304
rect 5993 3299 6059 3302
rect 8937 3299 9003 3302
rect 10869 3299 10935 3302
rect 12249 3362 12315 3365
rect 14273 3362 14339 3365
rect 12249 3360 14339 3362
rect 12249 3304 12254 3360
rect 12310 3304 14278 3360
rect 14334 3304 14339 3360
rect 12249 3302 14339 3304
rect 12249 3299 12315 3302
rect 14273 3299 14339 3302
rect 4409 3296 4729 3297
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 3231 4729 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 18270 3296 18590 3297
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18270 3231 18590 3232
rect 6085 3226 6151 3229
rect 9213 3226 9279 3229
rect 6085 3224 11208 3226
rect 6085 3168 6090 3224
rect 6146 3168 9218 3224
rect 9274 3168 11208 3224
rect 6085 3166 11208 3168
rect 6085 3163 6151 3166
rect 9213 3163 9279 3166
rect 0 3090 800 3120
rect 2957 3090 3023 3093
rect 0 3088 3023 3090
rect 0 3032 2962 3088
rect 3018 3032 3023 3088
rect 0 3030 3023 3032
rect 0 3000 800 3030
rect 2957 3027 3023 3030
rect 7741 3090 7807 3093
rect 8937 3090 9003 3093
rect 7741 3088 9003 3090
rect 7741 3032 7746 3088
rect 7802 3032 8942 3088
rect 8998 3032 9003 3088
rect 7741 3030 9003 3032
rect 7741 3027 7807 3030
rect 8937 3027 9003 3030
rect 10225 3090 10291 3093
rect 10358 3090 10364 3092
rect 10225 3088 10364 3090
rect 10225 3032 10230 3088
rect 10286 3032 10364 3088
rect 10225 3030 10364 3032
rect 10225 3027 10291 3030
rect 10358 3028 10364 3030
rect 10428 3028 10434 3092
rect 11148 3090 11208 3166
rect 14641 3090 14707 3093
rect 11148 3088 14707 3090
rect 11148 3032 14646 3088
rect 14702 3032 14707 3088
rect 11148 3030 14707 3032
rect 14641 3027 14707 3030
rect 18965 3090 19031 3093
rect 19977 3090 20043 3093
rect 18965 3088 20043 3090
rect 18965 3032 18970 3088
rect 19026 3032 19982 3088
rect 20038 3032 20043 3088
rect 18965 3030 20043 3032
rect 18965 3027 19031 3030
rect 19977 3027 20043 3030
rect 20345 3090 20411 3093
rect 22200 3090 23000 3120
rect 20345 3088 23000 3090
rect 20345 3032 20350 3088
rect 20406 3032 23000 3088
rect 20345 3030 23000 3032
rect 20345 3027 20411 3030
rect 22200 3000 23000 3030
rect 9029 2954 9095 2957
rect 10041 2954 10107 2957
rect 9029 2952 10107 2954
rect 9029 2896 9034 2952
rect 9090 2896 10046 2952
rect 10102 2896 10107 2952
rect 9029 2894 10107 2896
rect 9029 2891 9095 2894
rect 10041 2891 10107 2894
rect 10317 2954 10383 2957
rect 15745 2954 15811 2957
rect 10317 2952 15811 2954
rect 10317 2896 10322 2952
rect 10378 2896 15750 2952
rect 15806 2896 15811 2952
rect 10317 2894 15811 2896
rect 10317 2891 10383 2894
rect 15745 2891 15811 2894
rect 2221 2818 2287 2821
rect 7741 2818 7807 2821
rect 2221 2816 7807 2818
rect 2221 2760 2226 2816
rect 2282 2760 7746 2816
rect 7802 2760 7807 2816
rect 2221 2758 7807 2760
rect 2221 2755 2287 2758
rect 7741 2755 7807 2758
rect 8477 2818 8543 2821
rect 9438 2818 9444 2820
rect 8477 2816 9444 2818
rect 8477 2760 8482 2816
rect 8538 2760 9444 2816
rect 8477 2758 9444 2760
rect 8477 2755 8543 2758
rect 9438 2756 9444 2758
rect 9508 2756 9514 2820
rect 11697 2818 11763 2821
rect 12157 2818 12223 2821
rect 11697 2816 12223 2818
rect 11697 2760 11702 2816
rect 11758 2760 12162 2816
rect 12218 2760 12223 2816
rect 11697 2758 12223 2760
rect 11697 2755 11763 2758
rect 12157 2755 12223 2758
rect 7874 2752 8194 2753
rect 0 2682 800 2712
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8194 2752
rect 7874 2687 8194 2688
rect 14805 2752 15125 2753
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2687 15125 2688
rect 2773 2682 2839 2685
rect 0 2680 2839 2682
rect 0 2624 2778 2680
rect 2834 2624 2839 2680
rect 0 2622 2839 2624
rect 0 2592 800 2622
rect 2773 2619 2839 2622
rect 9397 2682 9463 2685
rect 11605 2682 11671 2685
rect 9397 2680 11671 2682
rect 9397 2624 9402 2680
rect 9458 2624 11610 2680
rect 11666 2624 11671 2680
rect 9397 2622 11671 2624
rect 9397 2619 9463 2622
rect 11605 2619 11671 2622
rect 22001 2682 22067 2685
rect 22200 2682 23000 2712
rect 22001 2680 23000 2682
rect 22001 2624 22006 2680
rect 22062 2624 23000 2680
rect 22001 2622 23000 2624
rect 22001 2619 22067 2622
rect 22200 2592 23000 2622
rect 11145 2546 11211 2549
rect 13629 2546 13695 2549
rect 14181 2546 14247 2549
rect 11145 2544 14247 2546
rect 11145 2488 11150 2544
rect 11206 2488 13634 2544
rect 13690 2488 14186 2544
rect 14242 2488 14247 2544
rect 11145 2486 14247 2488
rect 11145 2483 11211 2486
rect 13629 2483 13695 2486
rect 14181 2483 14247 2486
rect 9121 2410 9187 2413
rect 13813 2410 13879 2413
rect 9121 2408 13879 2410
rect 9121 2352 9126 2408
rect 9182 2352 13818 2408
rect 13874 2352 13879 2408
rect 9121 2350 13879 2352
rect 9121 2347 9187 2350
rect 13813 2347 13879 2350
rect 0 2274 800 2304
rect 1761 2274 1827 2277
rect 0 2272 1827 2274
rect 0 2216 1766 2272
rect 1822 2216 1827 2272
rect 0 2214 1827 2216
rect 0 2184 800 2214
rect 1761 2211 1827 2214
rect 20161 2274 20227 2277
rect 22200 2274 23000 2304
rect 20161 2272 23000 2274
rect 20161 2216 20166 2272
rect 20222 2216 23000 2272
rect 20161 2214 23000 2216
rect 20161 2211 20227 2214
rect 4409 2208 4729 2209
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2143 4729 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 18270 2208 18590 2209
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 22200 2184 23000 2214
rect 18270 2143 18590 2144
rect 0 1866 800 1896
rect 2129 1866 2195 1869
rect 3141 1866 3207 1869
rect 0 1864 3207 1866
rect 0 1808 2134 1864
rect 2190 1808 3146 1864
rect 3202 1808 3207 1864
rect 0 1806 3207 1808
rect 0 1776 800 1806
rect 2129 1803 2195 1806
rect 3141 1803 3207 1806
rect 20897 1866 20963 1869
rect 22200 1866 23000 1896
rect 20897 1864 23000 1866
rect 20897 1808 20902 1864
rect 20958 1808 23000 1864
rect 20897 1806 23000 1808
rect 20897 1803 20963 1806
rect 22200 1776 23000 1806
rect 0 1458 800 1488
rect 1301 1458 1367 1461
rect 0 1456 1367 1458
rect 0 1400 1306 1456
rect 1362 1400 1367 1456
rect 0 1398 1367 1400
rect 0 1368 800 1398
rect 1301 1395 1367 1398
rect 19885 1458 19951 1461
rect 22200 1458 23000 1488
rect 19885 1456 23000 1458
rect 19885 1400 19890 1456
rect 19946 1400 23000 1456
rect 19885 1398 23000 1400
rect 19885 1395 19951 1398
rect 22200 1368 23000 1398
rect 0 1050 800 1080
rect 3601 1050 3667 1053
rect 0 1048 3667 1050
rect 0 992 3606 1048
rect 3662 992 3667 1048
rect 0 990 3667 992
rect 0 960 800 990
rect 3601 987 3667 990
rect 21081 1050 21147 1053
rect 22200 1050 23000 1080
rect 21081 1048 23000 1050
rect 21081 992 21086 1048
rect 21142 992 23000 1048
rect 21081 990 23000 992
rect 21081 987 21147 990
rect 22200 960 23000 990
rect 21449 914 21515 917
rect 21817 914 21883 917
rect 21449 912 21883 914
rect 21449 856 21454 912
rect 21510 856 21822 912
rect 21878 856 21883 912
rect 21449 854 21883 856
rect 21449 851 21515 854
rect 21817 851 21883 854
rect 0 642 800 672
rect 2957 642 3023 645
rect 0 640 3023 642
rect 0 584 2962 640
rect 3018 584 3023 640
rect 0 582 3023 584
rect 0 552 800 582
rect 2957 579 3023 582
rect 19517 642 19583 645
rect 22200 642 23000 672
rect 19517 640 23000 642
rect 19517 584 19522 640
rect 19578 584 23000 640
rect 19517 582 23000 584
rect 19517 579 19583 582
rect 22200 552 23000 582
rect 0 234 800 264
rect 3785 234 3851 237
rect 0 232 3851 234
rect 0 176 3790 232
rect 3846 176 3851 232
rect 0 174 3851 176
rect 0 144 800 174
rect 3785 171 3851 174
rect 20805 234 20871 237
rect 22200 234 23000 264
rect 20805 232 23000 234
rect 20805 176 20810 232
rect 20866 176 23000 232
rect 20805 174 23000 176
rect 20805 171 20871 174
rect 22200 144 23000 174
<< via3 >>
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 4577 20700 4641 20704
rect 4577 20644 4581 20700
rect 4581 20644 4637 20700
rect 4637 20644 4641 20700
rect 4577 20640 4641 20644
rect 4657 20700 4721 20704
rect 4657 20644 4661 20700
rect 4661 20644 4717 20700
rect 4717 20644 4721 20700
rect 4657 20640 4721 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 18278 20700 18342 20704
rect 18278 20644 18282 20700
rect 18282 20644 18338 20700
rect 18338 20644 18342 20700
rect 18278 20640 18342 20644
rect 18358 20700 18422 20704
rect 18358 20644 18362 20700
rect 18362 20644 18418 20700
rect 18418 20644 18422 20700
rect 18358 20640 18422 20644
rect 18438 20700 18502 20704
rect 18438 20644 18442 20700
rect 18442 20644 18498 20700
rect 18498 20644 18502 20700
rect 18438 20640 18502 20644
rect 18518 20700 18582 20704
rect 18518 20644 18522 20700
rect 18522 20644 18578 20700
rect 18578 20644 18582 20700
rect 18518 20640 18582 20644
rect 7882 20156 7946 20160
rect 7882 20100 7886 20156
rect 7886 20100 7942 20156
rect 7942 20100 7946 20156
rect 7882 20096 7946 20100
rect 7962 20156 8026 20160
rect 7962 20100 7966 20156
rect 7966 20100 8022 20156
rect 8022 20100 8026 20156
rect 7962 20096 8026 20100
rect 8042 20156 8106 20160
rect 8042 20100 8046 20156
rect 8046 20100 8102 20156
rect 8102 20100 8106 20156
rect 8042 20096 8106 20100
rect 8122 20156 8186 20160
rect 8122 20100 8126 20156
rect 8126 20100 8182 20156
rect 8182 20100 8186 20156
rect 8122 20096 8186 20100
rect 14813 20156 14877 20160
rect 14813 20100 14817 20156
rect 14817 20100 14873 20156
rect 14873 20100 14877 20156
rect 14813 20096 14877 20100
rect 14893 20156 14957 20160
rect 14893 20100 14897 20156
rect 14897 20100 14953 20156
rect 14953 20100 14957 20156
rect 14893 20096 14957 20100
rect 14973 20156 15037 20160
rect 14973 20100 14977 20156
rect 14977 20100 15033 20156
rect 15033 20100 15037 20156
rect 14973 20096 15037 20100
rect 15053 20156 15117 20160
rect 15053 20100 15057 20156
rect 15057 20100 15113 20156
rect 15113 20100 15117 20156
rect 15053 20096 15117 20100
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 4577 19612 4641 19616
rect 4577 19556 4581 19612
rect 4581 19556 4637 19612
rect 4637 19556 4641 19612
rect 4577 19552 4641 19556
rect 4657 19612 4721 19616
rect 4657 19556 4661 19612
rect 4661 19556 4717 19612
rect 4717 19556 4721 19612
rect 4657 19552 4721 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 18278 19612 18342 19616
rect 18278 19556 18282 19612
rect 18282 19556 18338 19612
rect 18338 19556 18342 19612
rect 18278 19552 18342 19556
rect 18358 19612 18422 19616
rect 18358 19556 18362 19612
rect 18362 19556 18418 19612
rect 18418 19556 18422 19612
rect 18358 19552 18422 19556
rect 18438 19612 18502 19616
rect 18438 19556 18442 19612
rect 18442 19556 18498 19612
rect 18498 19556 18502 19612
rect 18438 19552 18502 19556
rect 18518 19612 18582 19616
rect 18518 19556 18522 19612
rect 18522 19556 18578 19612
rect 18578 19556 18582 19612
rect 18518 19552 18582 19556
rect 7604 19348 7668 19412
rect 8524 19408 8588 19412
rect 8524 19352 8574 19408
rect 8574 19352 8588 19408
rect 8524 19348 8588 19352
rect 7882 19068 7946 19072
rect 7882 19012 7886 19068
rect 7886 19012 7942 19068
rect 7942 19012 7946 19068
rect 7882 19008 7946 19012
rect 7962 19068 8026 19072
rect 7962 19012 7966 19068
rect 7966 19012 8022 19068
rect 8022 19012 8026 19068
rect 7962 19008 8026 19012
rect 8042 19068 8106 19072
rect 8042 19012 8046 19068
rect 8046 19012 8102 19068
rect 8102 19012 8106 19068
rect 8042 19008 8106 19012
rect 8122 19068 8186 19072
rect 8122 19012 8126 19068
rect 8126 19012 8182 19068
rect 8182 19012 8186 19068
rect 8122 19008 8186 19012
rect 14813 19068 14877 19072
rect 14813 19012 14817 19068
rect 14817 19012 14873 19068
rect 14873 19012 14877 19068
rect 14813 19008 14877 19012
rect 14893 19068 14957 19072
rect 14893 19012 14897 19068
rect 14897 19012 14953 19068
rect 14953 19012 14957 19068
rect 14893 19008 14957 19012
rect 14973 19068 15037 19072
rect 14973 19012 14977 19068
rect 14977 19012 15033 19068
rect 15033 19012 15037 19068
rect 14973 19008 15037 19012
rect 15053 19068 15117 19072
rect 15053 19012 15057 19068
rect 15057 19012 15113 19068
rect 15113 19012 15117 19068
rect 15053 19008 15117 19012
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 4577 18524 4641 18528
rect 4577 18468 4581 18524
rect 4581 18468 4637 18524
rect 4637 18468 4641 18524
rect 4577 18464 4641 18468
rect 4657 18524 4721 18528
rect 4657 18468 4661 18524
rect 4661 18468 4717 18524
rect 4717 18468 4721 18524
rect 4657 18464 4721 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 18278 18524 18342 18528
rect 18278 18468 18282 18524
rect 18282 18468 18338 18524
rect 18338 18468 18342 18524
rect 18278 18464 18342 18468
rect 18358 18524 18422 18528
rect 18358 18468 18362 18524
rect 18362 18468 18418 18524
rect 18418 18468 18422 18524
rect 18358 18464 18422 18468
rect 18438 18524 18502 18528
rect 18438 18468 18442 18524
rect 18442 18468 18498 18524
rect 18498 18468 18502 18524
rect 18438 18464 18502 18468
rect 18518 18524 18582 18528
rect 18518 18468 18522 18524
rect 18522 18468 18578 18524
rect 18578 18468 18582 18524
rect 18518 18464 18582 18468
rect 6868 18396 6932 18460
rect 7882 17980 7946 17984
rect 7882 17924 7886 17980
rect 7886 17924 7942 17980
rect 7942 17924 7946 17980
rect 7882 17920 7946 17924
rect 7962 17980 8026 17984
rect 7962 17924 7966 17980
rect 7966 17924 8022 17980
rect 8022 17924 8026 17980
rect 7962 17920 8026 17924
rect 8042 17980 8106 17984
rect 8042 17924 8046 17980
rect 8046 17924 8102 17980
rect 8102 17924 8106 17980
rect 8042 17920 8106 17924
rect 8122 17980 8186 17984
rect 8122 17924 8126 17980
rect 8126 17924 8182 17980
rect 8182 17924 8186 17980
rect 8122 17920 8186 17924
rect 14813 17980 14877 17984
rect 14813 17924 14817 17980
rect 14817 17924 14873 17980
rect 14873 17924 14877 17980
rect 14813 17920 14877 17924
rect 14893 17980 14957 17984
rect 14893 17924 14897 17980
rect 14897 17924 14953 17980
rect 14953 17924 14957 17980
rect 14893 17920 14957 17924
rect 14973 17980 15037 17984
rect 14973 17924 14977 17980
rect 14977 17924 15033 17980
rect 15033 17924 15037 17980
rect 14973 17920 15037 17924
rect 15053 17980 15117 17984
rect 15053 17924 15057 17980
rect 15057 17924 15113 17980
rect 15113 17924 15117 17980
rect 15053 17920 15117 17924
rect 7052 17444 7116 17508
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 4577 17436 4641 17440
rect 4577 17380 4581 17436
rect 4581 17380 4637 17436
rect 4637 17380 4641 17436
rect 4577 17376 4641 17380
rect 4657 17436 4721 17440
rect 4657 17380 4661 17436
rect 4661 17380 4717 17436
rect 4717 17380 4721 17436
rect 4657 17376 4721 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 18278 17436 18342 17440
rect 18278 17380 18282 17436
rect 18282 17380 18338 17436
rect 18338 17380 18342 17436
rect 18278 17376 18342 17380
rect 18358 17436 18422 17440
rect 18358 17380 18362 17436
rect 18362 17380 18418 17436
rect 18418 17380 18422 17436
rect 18358 17376 18422 17380
rect 18438 17436 18502 17440
rect 18438 17380 18442 17436
rect 18442 17380 18498 17436
rect 18498 17380 18502 17436
rect 18438 17376 18502 17380
rect 18518 17436 18582 17440
rect 18518 17380 18522 17436
rect 18522 17380 18578 17436
rect 18578 17380 18582 17436
rect 18518 17376 18582 17380
rect 9812 17036 9876 17100
rect 7882 16892 7946 16896
rect 7882 16836 7886 16892
rect 7886 16836 7942 16892
rect 7942 16836 7946 16892
rect 7882 16832 7946 16836
rect 7962 16892 8026 16896
rect 7962 16836 7966 16892
rect 7966 16836 8022 16892
rect 8022 16836 8026 16892
rect 7962 16832 8026 16836
rect 8042 16892 8106 16896
rect 8042 16836 8046 16892
rect 8046 16836 8102 16892
rect 8102 16836 8106 16892
rect 8042 16832 8106 16836
rect 8122 16892 8186 16896
rect 8122 16836 8126 16892
rect 8126 16836 8182 16892
rect 8182 16836 8186 16892
rect 8122 16832 8186 16836
rect 14813 16892 14877 16896
rect 14813 16836 14817 16892
rect 14817 16836 14873 16892
rect 14873 16836 14877 16892
rect 14813 16832 14877 16836
rect 14893 16892 14957 16896
rect 14893 16836 14897 16892
rect 14897 16836 14953 16892
rect 14953 16836 14957 16892
rect 14893 16832 14957 16836
rect 14973 16892 15037 16896
rect 14973 16836 14977 16892
rect 14977 16836 15033 16892
rect 15033 16836 15037 16892
rect 14973 16832 15037 16836
rect 15053 16892 15117 16896
rect 15053 16836 15057 16892
rect 15057 16836 15113 16892
rect 15113 16836 15117 16892
rect 15053 16832 15117 16836
rect 10548 16824 10612 16828
rect 10548 16768 10562 16824
rect 10562 16768 10612 16824
rect 10548 16764 10612 16768
rect 11836 16492 11900 16556
rect 9260 16356 9324 16420
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 4577 16348 4641 16352
rect 4577 16292 4581 16348
rect 4581 16292 4637 16348
rect 4637 16292 4641 16348
rect 4577 16288 4641 16292
rect 4657 16348 4721 16352
rect 4657 16292 4661 16348
rect 4661 16292 4717 16348
rect 4717 16292 4721 16348
rect 4657 16288 4721 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 18278 16348 18342 16352
rect 18278 16292 18282 16348
rect 18282 16292 18338 16348
rect 18338 16292 18342 16348
rect 18278 16288 18342 16292
rect 18358 16348 18422 16352
rect 18358 16292 18362 16348
rect 18362 16292 18418 16348
rect 18418 16292 18422 16348
rect 18358 16288 18422 16292
rect 18438 16348 18502 16352
rect 18438 16292 18442 16348
rect 18442 16292 18498 16348
rect 18498 16292 18502 16348
rect 18438 16288 18502 16292
rect 18518 16348 18582 16352
rect 18518 16292 18522 16348
rect 18522 16292 18578 16348
rect 18578 16292 18582 16348
rect 18518 16288 18582 16292
rect 7420 16220 7484 16284
rect 7882 15804 7946 15808
rect 7882 15748 7886 15804
rect 7886 15748 7942 15804
rect 7942 15748 7946 15804
rect 7882 15744 7946 15748
rect 7962 15804 8026 15808
rect 7962 15748 7966 15804
rect 7966 15748 8022 15804
rect 8022 15748 8026 15804
rect 7962 15744 8026 15748
rect 8042 15804 8106 15808
rect 8042 15748 8046 15804
rect 8046 15748 8102 15804
rect 8102 15748 8106 15804
rect 8042 15744 8106 15748
rect 8122 15804 8186 15808
rect 8122 15748 8126 15804
rect 8126 15748 8182 15804
rect 8182 15748 8186 15804
rect 8122 15744 8186 15748
rect 14813 15804 14877 15808
rect 14813 15748 14817 15804
rect 14817 15748 14873 15804
rect 14873 15748 14877 15804
rect 14813 15744 14877 15748
rect 14893 15804 14957 15808
rect 14893 15748 14897 15804
rect 14897 15748 14953 15804
rect 14953 15748 14957 15804
rect 14893 15744 14957 15748
rect 14973 15804 15037 15808
rect 14973 15748 14977 15804
rect 14977 15748 15033 15804
rect 15033 15748 15037 15804
rect 14973 15744 15037 15748
rect 15053 15804 15117 15808
rect 15053 15748 15057 15804
rect 15057 15748 15113 15804
rect 15113 15748 15117 15804
rect 15053 15744 15117 15748
rect 7236 15540 7300 15604
rect 12572 15328 12636 15332
rect 12572 15272 12622 15328
rect 12622 15272 12636 15328
rect 12572 15268 12636 15272
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 4577 15260 4641 15264
rect 4577 15204 4581 15260
rect 4581 15204 4637 15260
rect 4637 15204 4641 15260
rect 4577 15200 4641 15204
rect 4657 15260 4721 15264
rect 4657 15204 4661 15260
rect 4661 15204 4717 15260
rect 4717 15204 4721 15260
rect 4657 15200 4721 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 18278 15260 18342 15264
rect 18278 15204 18282 15260
rect 18282 15204 18338 15260
rect 18338 15204 18342 15260
rect 18278 15200 18342 15204
rect 18358 15260 18422 15264
rect 18358 15204 18362 15260
rect 18362 15204 18418 15260
rect 18418 15204 18422 15260
rect 18358 15200 18422 15204
rect 18438 15260 18502 15264
rect 18438 15204 18442 15260
rect 18442 15204 18498 15260
rect 18498 15204 18502 15260
rect 18438 15200 18502 15204
rect 18518 15260 18582 15264
rect 18518 15204 18522 15260
rect 18522 15204 18578 15260
rect 18578 15204 18582 15260
rect 18518 15200 18582 15204
rect 9996 14860 10060 14924
rect 10364 14784 10428 14788
rect 10364 14728 10414 14784
rect 10414 14728 10428 14784
rect 10364 14724 10428 14728
rect 7882 14716 7946 14720
rect 7882 14660 7886 14716
rect 7886 14660 7942 14716
rect 7942 14660 7946 14716
rect 7882 14656 7946 14660
rect 7962 14716 8026 14720
rect 7962 14660 7966 14716
rect 7966 14660 8022 14716
rect 8022 14660 8026 14716
rect 7962 14656 8026 14660
rect 8042 14716 8106 14720
rect 8042 14660 8046 14716
rect 8046 14660 8102 14716
rect 8102 14660 8106 14716
rect 8042 14656 8106 14660
rect 8122 14716 8186 14720
rect 8122 14660 8126 14716
rect 8126 14660 8182 14716
rect 8182 14660 8186 14716
rect 8122 14656 8186 14660
rect 14813 14716 14877 14720
rect 14813 14660 14817 14716
rect 14817 14660 14873 14716
rect 14873 14660 14877 14716
rect 14813 14656 14877 14660
rect 14893 14716 14957 14720
rect 14893 14660 14897 14716
rect 14897 14660 14953 14716
rect 14953 14660 14957 14716
rect 14893 14656 14957 14660
rect 14973 14716 15037 14720
rect 14973 14660 14977 14716
rect 14977 14660 15033 14716
rect 15033 14660 15037 14716
rect 14973 14656 15037 14660
rect 15053 14716 15117 14720
rect 15053 14660 15057 14716
rect 15057 14660 15113 14716
rect 15113 14660 15117 14716
rect 15053 14656 15117 14660
rect 9628 14588 9692 14652
rect 7420 14316 7484 14380
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 4577 14172 4641 14176
rect 4577 14116 4581 14172
rect 4581 14116 4637 14172
rect 4637 14116 4641 14172
rect 4577 14112 4641 14116
rect 4657 14172 4721 14176
rect 4657 14116 4661 14172
rect 4661 14116 4717 14172
rect 4717 14116 4721 14172
rect 4657 14112 4721 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 18278 14172 18342 14176
rect 18278 14116 18282 14172
rect 18282 14116 18338 14172
rect 18338 14116 18342 14172
rect 18278 14112 18342 14116
rect 18358 14172 18422 14176
rect 18358 14116 18362 14172
rect 18362 14116 18418 14172
rect 18418 14116 18422 14172
rect 18358 14112 18422 14116
rect 18438 14172 18502 14176
rect 18438 14116 18442 14172
rect 18442 14116 18498 14172
rect 18498 14116 18502 14172
rect 18438 14112 18502 14116
rect 18518 14172 18582 14176
rect 18518 14116 18522 14172
rect 18522 14116 18578 14172
rect 18578 14116 18582 14172
rect 18518 14112 18582 14116
rect 9628 14044 9692 14108
rect 8708 13772 8772 13836
rect 11100 13772 11164 13836
rect 7882 13628 7946 13632
rect 7882 13572 7886 13628
rect 7886 13572 7942 13628
rect 7942 13572 7946 13628
rect 7882 13568 7946 13572
rect 7962 13628 8026 13632
rect 7962 13572 7966 13628
rect 7966 13572 8022 13628
rect 8022 13572 8026 13628
rect 7962 13568 8026 13572
rect 8042 13628 8106 13632
rect 8042 13572 8046 13628
rect 8046 13572 8102 13628
rect 8102 13572 8106 13628
rect 8042 13568 8106 13572
rect 8122 13628 8186 13632
rect 8122 13572 8126 13628
rect 8126 13572 8182 13628
rect 8182 13572 8186 13628
rect 8122 13568 8186 13572
rect 14813 13628 14877 13632
rect 14813 13572 14817 13628
rect 14817 13572 14873 13628
rect 14873 13572 14877 13628
rect 14813 13568 14877 13572
rect 14893 13628 14957 13632
rect 14893 13572 14897 13628
rect 14897 13572 14953 13628
rect 14953 13572 14957 13628
rect 14893 13568 14957 13572
rect 14973 13628 15037 13632
rect 14973 13572 14977 13628
rect 14977 13572 15033 13628
rect 15033 13572 15037 13628
rect 14973 13568 15037 13572
rect 15053 13628 15117 13632
rect 15053 13572 15057 13628
rect 15057 13572 15113 13628
rect 15113 13572 15117 13628
rect 15053 13568 15117 13572
rect 8892 13560 8956 13564
rect 8892 13504 8906 13560
rect 8906 13504 8956 13560
rect 8892 13500 8956 13504
rect 9444 13560 9508 13564
rect 9444 13504 9494 13560
rect 9494 13504 9508 13560
rect 9444 13500 9508 13504
rect 10916 13364 10980 13428
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 4577 13084 4641 13088
rect 4577 13028 4581 13084
rect 4581 13028 4637 13084
rect 4637 13028 4641 13084
rect 4577 13024 4641 13028
rect 4657 13084 4721 13088
rect 4657 13028 4661 13084
rect 4661 13028 4717 13084
rect 4717 13028 4721 13084
rect 4657 13024 4721 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 18278 13084 18342 13088
rect 18278 13028 18282 13084
rect 18282 13028 18338 13084
rect 18338 13028 18342 13084
rect 18278 13024 18342 13028
rect 18358 13084 18422 13088
rect 18358 13028 18362 13084
rect 18362 13028 18418 13084
rect 18418 13028 18422 13084
rect 18358 13024 18422 13028
rect 18438 13084 18502 13088
rect 18438 13028 18442 13084
rect 18442 13028 18498 13084
rect 18498 13028 18502 13084
rect 18438 13024 18502 13028
rect 18518 13084 18582 13088
rect 18518 13028 18522 13084
rect 18522 13028 18578 13084
rect 18578 13028 18582 13084
rect 18518 13024 18582 13028
rect 5764 12608 5828 12612
rect 5764 12552 5778 12608
rect 5778 12552 5828 12608
rect 5764 12548 5828 12552
rect 6868 12684 6932 12748
rect 7882 12540 7946 12544
rect 7882 12484 7886 12540
rect 7886 12484 7942 12540
rect 7942 12484 7946 12540
rect 7882 12480 7946 12484
rect 7962 12540 8026 12544
rect 7962 12484 7966 12540
rect 7966 12484 8022 12540
rect 8022 12484 8026 12540
rect 7962 12480 8026 12484
rect 8042 12540 8106 12544
rect 8042 12484 8046 12540
rect 8046 12484 8102 12540
rect 8102 12484 8106 12540
rect 8042 12480 8106 12484
rect 8122 12540 8186 12544
rect 8122 12484 8126 12540
rect 8126 12484 8182 12540
rect 8182 12484 8186 12540
rect 8122 12480 8186 12484
rect 14813 12540 14877 12544
rect 14813 12484 14817 12540
rect 14817 12484 14873 12540
rect 14873 12484 14877 12540
rect 14813 12480 14877 12484
rect 14893 12540 14957 12544
rect 14893 12484 14897 12540
rect 14897 12484 14953 12540
rect 14953 12484 14957 12540
rect 14893 12480 14957 12484
rect 14973 12540 15037 12544
rect 14973 12484 14977 12540
rect 14977 12484 15033 12540
rect 15033 12484 15037 12540
rect 14973 12480 15037 12484
rect 15053 12540 15117 12544
rect 15053 12484 15057 12540
rect 15057 12484 15113 12540
rect 15113 12484 15117 12540
rect 15053 12480 15117 12484
rect 11100 12412 11164 12476
rect 11836 12336 11900 12340
rect 11836 12280 11886 12336
rect 11886 12280 11900 12336
rect 11836 12276 11900 12280
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 4577 11996 4641 12000
rect 4577 11940 4581 11996
rect 4581 11940 4637 11996
rect 4637 11940 4641 11996
rect 4577 11936 4641 11940
rect 4657 11996 4721 12000
rect 4657 11940 4661 11996
rect 4661 11940 4717 11996
rect 4717 11940 4721 11996
rect 4657 11936 4721 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 18278 11996 18342 12000
rect 18278 11940 18282 11996
rect 18282 11940 18338 11996
rect 18338 11940 18342 11996
rect 18278 11936 18342 11940
rect 18358 11996 18422 12000
rect 18358 11940 18362 11996
rect 18362 11940 18418 11996
rect 18418 11940 18422 11996
rect 18358 11936 18422 11940
rect 18438 11996 18502 12000
rect 18438 11940 18442 11996
rect 18442 11940 18498 11996
rect 18498 11940 18502 11996
rect 18438 11936 18502 11940
rect 18518 11996 18582 12000
rect 18518 11940 18522 11996
rect 18522 11940 18578 11996
rect 18578 11940 18582 11996
rect 18518 11936 18582 11940
rect 3924 11928 3988 11932
rect 3924 11872 3938 11928
rect 3938 11872 3988 11928
rect 3924 11868 3988 11872
rect 6868 11928 6932 11932
rect 6868 11872 6918 11928
rect 6918 11872 6932 11928
rect 6868 11868 6932 11872
rect 12020 11928 12084 11932
rect 12020 11872 12034 11928
rect 12034 11872 12084 11928
rect 12020 11868 12084 11872
rect 7420 11732 7484 11796
rect 3372 11520 3436 11524
rect 3372 11464 3386 11520
rect 3386 11464 3436 11520
rect 3372 11460 3436 11464
rect 7882 11452 7946 11456
rect 7882 11396 7886 11452
rect 7886 11396 7942 11452
rect 7942 11396 7946 11452
rect 7882 11392 7946 11396
rect 7962 11452 8026 11456
rect 7962 11396 7966 11452
rect 7966 11396 8022 11452
rect 8022 11396 8026 11452
rect 7962 11392 8026 11396
rect 8042 11452 8106 11456
rect 8042 11396 8046 11452
rect 8046 11396 8102 11452
rect 8102 11396 8106 11452
rect 8042 11392 8106 11396
rect 8122 11452 8186 11456
rect 8122 11396 8126 11452
rect 8126 11396 8182 11452
rect 8182 11396 8186 11452
rect 8122 11392 8186 11396
rect 14813 11452 14877 11456
rect 14813 11396 14817 11452
rect 14817 11396 14873 11452
rect 14873 11396 14877 11452
rect 14813 11392 14877 11396
rect 14893 11452 14957 11456
rect 14893 11396 14897 11452
rect 14897 11396 14953 11452
rect 14953 11396 14957 11452
rect 14893 11392 14957 11396
rect 14973 11452 15037 11456
rect 14973 11396 14977 11452
rect 14977 11396 15033 11452
rect 15033 11396 15037 11452
rect 14973 11392 15037 11396
rect 15053 11452 15117 11456
rect 15053 11396 15057 11452
rect 15057 11396 15113 11452
rect 15113 11396 15117 11452
rect 15053 11392 15117 11396
rect 9996 11324 10060 11388
rect 9260 10916 9324 10980
rect 12572 11052 12636 11116
rect 17908 11052 17972 11116
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 4577 10908 4641 10912
rect 4577 10852 4581 10908
rect 4581 10852 4637 10908
rect 4637 10852 4641 10908
rect 4577 10848 4641 10852
rect 4657 10908 4721 10912
rect 4657 10852 4661 10908
rect 4661 10852 4717 10908
rect 4717 10852 4721 10908
rect 4657 10848 4721 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 18278 10908 18342 10912
rect 18278 10852 18282 10908
rect 18282 10852 18338 10908
rect 18338 10852 18342 10908
rect 18278 10848 18342 10852
rect 18358 10908 18422 10912
rect 18358 10852 18362 10908
rect 18362 10852 18418 10908
rect 18418 10852 18422 10908
rect 18358 10848 18422 10852
rect 18438 10908 18502 10912
rect 18438 10852 18442 10908
rect 18442 10852 18498 10908
rect 18498 10852 18502 10908
rect 18438 10848 18502 10852
rect 18518 10908 18582 10912
rect 18518 10852 18522 10908
rect 18522 10852 18578 10908
rect 18578 10852 18582 10908
rect 18518 10848 18582 10852
rect 17908 10780 17972 10844
rect 10364 10644 10428 10708
rect 7604 10372 7668 10436
rect 9444 10372 9508 10436
rect 9812 10432 9876 10436
rect 9812 10376 9826 10432
rect 9826 10376 9876 10432
rect 9812 10372 9876 10376
rect 11100 10432 11164 10436
rect 11100 10376 11150 10432
rect 11150 10376 11164 10432
rect 11100 10372 11164 10376
rect 7882 10364 7946 10368
rect 7882 10308 7886 10364
rect 7886 10308 7942 10364
rect 7942 10308 7946 10364
rect 7882 10304 7946 10308
rect 7962 10364 8026 10368
rect 7962 10308 7966 10364
rect 7966 10308 8022 10364
rect 8022 10308 8026 10364
rect 7962 10304 8026 10308
rect 8042 10364 8106 10368
rect 8042 10308 8046 10364
rect 8046 10308 8102 10364
rect 8102 10308 8106 10364
rect 8042 10304 8106 10308
rect 8122 10364 8186 10368
rect 8122 10308 8126 10364
rect 8126 10308 8182 10364
rect 8182 10308 8186 10364
rect 8122 10304 8186 10308
rect 14813 10364 14877 10368
rect 14813 10308 14817 10364
rect 14817 10308 14873 10364
rect 14873 10308 14877 10364
rect 14813 10304 14877 10308
rect 14893 10364 14957 10368
rect 14893 10308 14897 10364
rect 14897 10308 14953 10364
rect 14953 10308 14957 10364
rect 14893 10304 14957 10308
rect 14973 10364 15037 10368
rect 14973 10308 14977 10364
rect 14977 10308 15033 10364
rect 15033 10308 15037 10364
rect 14973 10304 15037 10308
rect 15053 10364 15117 10368
rect 15053 10308 15057 10364
rect 15057 10308 15113 10364
rect 15113 10308 15117 10364
rect 15053 10304 15117 10308
rect 7052 10236 7116 10300
rect 8892 10236 8956 10300
rect 9628 10236 9692 10300
rect 11836 10236 11900 10300
rect 17908 10236 17972 10300
rect 9260 9964 9324 10028
rect 17908 9964 17972 10028
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 4577 9820 4641 9824
rect 4577 9764 4581 9820
rect 4581 9764 4637 9820
rect 4637 9764 4641 9820
rect 4577 9760 4641 9764
rect 4657 9820 4721 9824
rect 4657 9764 4661 9820
rect 4661 9764 4717 9820
rect 4717 9764 4721 9820
rect 4657 9760 4721 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 18278 9820 18342 9824
rect 18278 9764 18282 9820
rect 18282 9764 18338 9820
rect 18338 9764 18342 9820
rect 18278 9760 18342 9764
rect 18358 9820 18422 9824
rect 18358 9764 18362 9820
rect 18362 9764 18418 9820
rect 18418 9764 18422 9820
rect 18358 9760 18422 9764
rect 18438 9820 18502 9824
rect 18438 9764 18442 9820
rect 18442 9764 18498 9820
rect 18498 9764 18502 9820
rect 18438 9760 18502 9764
rect 18518 9820 18582 9824
rect 18518 9764 18522 9820
rect 18522 9764 18578 9820
rect 18578 9764 18582 9820
rect 18518 9760 18582 9764
rect 5764 9752 5828 9756
rect 5764 9696 5778 9752
rect 5778 9696 5828 9752
rect 5764 9692 5828 9696
rect 10364 9752 10428 9756
rect 10364 9696 10414 9752
rect 10414 9696 10428 9752
rect 10364 9692 10428 9696
rect 12572 9284 12636 9348
rect 7882 9276 7946 9280
rect 7882 9220 7886 9276
rect 7886 9220 7942 9276
rect 7942 9220 7946 9276
rect 7882 9216 7946 9220
rect 7962 9276 8026 9280
rect 7962 9220 7966 9276
rect 7966 9220 8022 9276
rect 8022 9220 8026 9276
rect 7962 9216 8026 9220
rect 8042 9276 8106 9280
rect 8042 9220 8046 9276
rect 8046 9220 8102 9276
rect 8102 9220 8106 9276
rect 8042 9216 8106 9220
rect 8122 9276 8186 9280
rect 8122 9220 8126 9276
rect 8126 9220 8182 9276
rect 8182 9220 8186 9276
rect 8122 9216 8186 9220
rect 14044 9148 14108 9212
rect 14813 9276 14877 9280
rect 14813 9220 14817 9276
rect 14817 9220 14873 9276
rect 14873 9220 14877 9276
rect 14813 9216 14877 9220
rect 14893 9276 14957 9280
rect 14893 9220 14897 9276
rect 14897 9220 14953 9276
rect 14953 9220 14957 9276
rect 14893 9216 14957 9220
rect 14973 9276 15037 9280
rect 14973 9220 14977 9276
rect 14977 9220 15033 9276
rect 15033 9220 15037 9276
rect 14973 9216 15037 9220
rect 15053 9276 15117 9280
rect 15053 9220 15057 9276
rect 15057 9220 15113 9276
rect 15113 9220 15117 9276
rect 15053 9216 15117 9220
rect 19196 9148 19260 9212
rect 3372 8936 3436 8940
rect 3372 8880 3422 8936
rect 3422 8880 3436 8936
rect 3372 8876 3436 8880
rect 7236 8740 7300 8804
rect 11100 8740 11164 8804
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 4577 8732 4641 8736
rect 4577 8676 4581 8732
rect 4581 8676 4637 8732
rect 4637 8676 4641 8732
rect 4577 8672 4641 8676
rect 4657 8732 4721 8736
rect 4657 8676 4661 8732
rect 4661 8676 4717 8732
rect 4717 8676 4721 8732
rect 4657 8672 4721 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 18278 8732 18342 8736
rect 18278 8676 18282 8732
rect 18282 8676 18338 8732
rect 18338 8676 18342 8732
rect 18278 8672 18342 8676
rect 18358 8732 18422 8736
rect 18358 8676 18362 8732
rect 18362 8676 18418 8732
rect 18418 8676 18422 8732
rect 18358 8672 18422 8676
rect 18438 8732 18502 8736
rect 18438 8676 18442 8732
rect 18442 8676 18498 8732
rect 18498 8676 18502 8732
rect 18438 8672 18502 8676
rect 18518 8732 18582 8736
rect 18518 8676 18522 8732
rect 18522 8676 18578 8732
rect 18578 8676 18582 8732
rect 18518 8672 18582 8676
rect 13124 8664 13188 8668
rect 13124 8608 13138 8664
rect 13138 8608 13188 8664
rect 13124 8604 13188 8608
rect 18828 8604 18892 8668
rect 7604 8468 7668 8532
rect 7420 8332 7484 8396
rect 10548 8392 10612 8396
rect 10548 8336 10598 8392
rect 10598 8336 10612 8392
rect 10548 8332 10612 8336
rect 13124 8392 13188 8396
rect 13124 8336 13138 8392
rect 13138 8336 13188 8392
rect 13124 8332 13188 8336
rect 18828 8332 18892 8396
rect 10916 8196 10980 8260
rect 7882 8188 7946 8192
rect 7882 8132 7886 8188
rect 7886 8132 7942 8188
rect 7942 8132 7946 8188
rect 7882 8128 7946 8132
rect 7962 8188 8026 8192
rect 7962 8132 7966 8188
rect 7966 8132 8022 8188
rect 8022 8132 8026 8188
rect 7962 8128 8026 8132
rect 8042 8188 8106 8192
rect 8042 8132 8046 8188
rect 8046 8132 8102 8188
rect 8102 8132 8106 8188
rect 8042 8128 8106 8132
rect 8122 8188 8186 8192
rect 8122 8132 8126 8188
rect 8126 8132 8182 8188
rect 8182 8132 8186 8188
rect 8122 8128 8186 8132
rect 14813 8188 14877 8192
rect 14813 8132 14817 8188
rect 14817 8132 14873 8188
rect 14873 8132 14877 8188
rect 14813 8128 14877 8132
rect 14893 8188 14957 8192
rect 14893 8132 14897 8188
rect 14897 8132 14953 8188
rect 14953 8132 14957 8188
rect 14893 8128 14957 8132
rect 14973 8188 15037 8192
rect 14973 8132 14977 8188
rect 14977 8132 15033 8188
rect 15033 8132 15037 8188
rect 14973 8128 15037 8132
rect 15053 8188 15117 8192
rect 15053 8132 15057 8188
rect 15057 8132 15113 8188
rect 15113 8132 15117 8188
rect 15053 8128 15117 8132
rect 8524 7788 8588 7852
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 4577 7644 4641 7648
rect 4577 7588 4581 7644
rect 4581 7588 4637 7644
rect 4637 7588 4641 7644
rect 4577 7584 4641 7588
rect 4657 7644 4721 7648
rect 4657 7588 4661 7644
rect 4661 7588 4717 7644
rect 4717 7588 4721 7644
rect 4657 7584 4721 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 18278 7644 18342 7648
rect 18278 7588 18282 7644
rect 18282 7588 18338 7644
rect 18338 7588 18342 7644
rect 18278 7584 18342 7588
rect 18358 7644 18422 7648
rect 18358 7588 18362 7644
rect 18362 7588 18418 7644
rect 18418 7588 18422 7644
rect 18358 7584 18422 7588
rect 18438 7644 18502 7648
rect 18438 7588 18442 7644
rect 18442 7588 18498 7644
rect 18498 7588 18502 7644
rect 18438 7584 18502 7588
rect 18518 7644 18582 7648
rect 18518 7588 18522 7644
rect 18522 7588 18578 7644
rect 18578 7588 18582 7644
rect 18518 7584 18582 7588
rect 11100 7108 11164 7172
rect 7882 7100 7946 7104
rect 7882 7044 7886 7100
rect 7886 7044 7942 7100
rect 7942 7044 7946 7100
rect 7882 7040 7946 7044
rect 7962 7100 8026 7104
rect 7962 7044 7966 7100
rect 7966 7044 8022 7100
rect 8022 7044 8026 7100
rect 7962 7040 8026 7044
rect 8042 7100 8106 7104
rect 8042 7044 8046 7100
rect 8046 7044 8102 7100
rect 8102 7044 8106 7100
rect 8042 7040 8106 7044
rect 8122 7100 8186 7104
rect 8122 7044 8126 7100
rect 8126 7044 8182 7100
rect 8182 7044 8186 7100
rect 8122 7040 8186 7044
rect 14813 7100 14877 7104
rect 14813 7044 14817 7100
rect 14817 7044 14873 7100
rect 14873 7044 14877 7100
rect 14813 7040 14877 7044
rect 14893 7100 14957 7104
rect 14893 7044 14897 7100
rect 14897 7044 14953 7100
rect 14953 7044 14957 7100
rect 14893 7040 14957 7044
rect 14973 7100 15037 7104
rect 14973 7044 14977 7100
rect 14977 7044 15033 7100
rect 15033 7044 15037 7100
rect 14973 7040 15037 7044
rect 15053 7100 15117 7104
rect 15053 7044 15057 7100
rect 15057 7044 15113 7100
rect 15113 7044 15117 7100
rect 15053 7040 15117 7044
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 4577 6556 4641 6560
rect 4577 6500 4581 6556
rect 4581 6500 4637 6556
rect 4637 6500 4641 6556
rect 4577 6496 4641 6500
rect 4657 6556 4721 6560
rect 4657 6500 4661 6556
rect 4661 6500 4717 6556
rect 4717 6500 4721 6556
rect 4657 6496 4721 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 18278 6556 18342 6560
rect 18278 6500 18282 6556
rect 18282 6500 18338 6556
rect 18338 6500 18342 6556
rect 18278 6496 18342 6500
rect 18358 6556 18422 6560
rect 18358 6500 18362 6556
rect 18362 6500 18418 6556
rect 18418 6500 18422 6556
rect 18358 6496 18422 6500
rect 18438 6556 18502 6560
rect 18438 6500 18442 6556
rect 18442 6500 18498 6556
rect 18498 6500 18502 6556
rect 18438 6496 18502 6500
rect 18518 6556 18582 6560
rect 18518 6500 18522 6556
rect 18522 6500 18578 6556
rect 18578 6500 18582 6556
rect 18518 6496 18582 6500
rect 12020 6488 12084 6492
rect 12020 6432 12034 6488
rect 12034 6432 12084 6488
rect 12020 6428 12084 6432
rect 19196 6624 19260 6628
rect 19196 6568 19210 6624
rect 19210 6568 19260 6624
rect 19196 6564 19260 6568
rect 7236 6156 7300 6220
rect 7882 6012 7946 6016
rect 7882 5956 7886 6012
rect 7886 5956 7942 6012
rect 7942 5956 7946 6012
rect 7882 5952 7946 5956
rect 7962 6012 8026 6016
rect 7962 5956 7966 6012
rect 7966 5956 8022 6012
rect 8022 5956 8026 6012
rect 7962 5952 8026 5956
rect 8042 6012 8106 6016
rect 8042 5956 8046 6012
rect 8046 5956 8102 6012
rect 8102 5956 8106 6012
rect 8042 5952 8106 5956
rect 8122 6012 8186 6016
rect 8122 5956 8126 6012
rect 8126 5956 8182 6012
rect 8182 5956 8186 6012
rect 8122 5952 8186 5956
rect 14813 6012 14877 6016
rect 14813 5956 14817 6012
rect 14817 5956 14873 6012
rect 14873 5956 14877 6012
rect 14813 5952 14877 5956
rect 14893 6012 14957 6016
rect 14893 5956 14897 6012
rect 14897 5956 14953 6012
rect 14953 5956 14957 6012
rect 14893 5952 14957 5956
rect 14973 6012 15037 6016
rect 14973 5956 14977 6012
rect 14977 5956 15033 6012
rect 15033 5956 15037 6012
rect 14973 5952 15037 5956
rect 15053 6012 15117 6016
rect 15053 5956 15057 6012
rect 15057 5956 15113 6012
rect 15113 5956 15117 6012
rect 15053 5952 15117 5956
rect 8708 5884 8772 5948
rect 9444 5476 9508 5540
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 4577 5468 4641 5472
rect 4577 5412 4581 5468
rect 4581 5412 4637 5468
rect 4637 5412 4641 5468
rect 4577 5408 4641 5412
rect 4657 5468 4721 5472
rect 4657 5412 4661 5468
rect 4661 5412 4717 5468
rect 4717 5412 4721 5468
rect 4657 5408 4721 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 18278 5468 18342 5472
rect 18278 5412 18282 5468
rect 18282 5412 18338 5468
rect 18338 5412 18342 5468
rect 18278 5408 18342 5412
rect 18358 5468 18422 5472
rect 18358 5412 18362 5468
rect 18362 5412 18418 5468
rect 18418 5412 18422 5468
rect 18358 5408 18422 5412
rect 18438 5468 18502 5472
rect 18438 5412 18442 5468
rect 18442 5412 18498 5468
rect 18498 5412 18502 5468
rect 18438 5408 18502 5412
rect 18518 5468 18582 5472
rect 18518 5412 18522 5468
rect 18522 5412 18578 5468
rect 18578 5412 18582 5468
rect 18518 5408 18582 5412
rect 7604 5340 7668 5404
rect 11836 5068 11900 5132
rect 7882 4924 7946 4928
rect 7882 4868 7886 4924
rect 7886 4868 7942 4924
rect 7942 4868 7946 4924
rect 7882 4864 7946 4868
rect 7962 4924 8026 4928
rect 7962 4868 7966 4924
rect 7966 4868 8022 4924
rect 8022 4868 8026 4924
rect 7962 4864 8026 4868
rect 8042 4924 8106 4928
rect 8042 4868 8046 4924
rect 8046 4868 8102 4924
rect 8102 4868 8106 4924
rect 8042 4864 8106 4868
rect 8122 4924 8186 4928
rect 8122 4868 8126 4924
rect 8126 4868 8182 4924
rect 8182 4868 8186 4924
rect 8122 4864 8186 4868
rect 14813 4924 14877 4928
rect 14813 4868 14817 4924
rect 14817 4868 14873 4924
rect 14873 4868 14877 4924
rect 14813 4864 14877 4868
rect 14893 4924 14957 4928
rect 14893 4868 14897 4924
rect 14897 4868 14953 4924
rect 14953 4868 14957 4924
rect 14893 4864 14957 4868
rect 14973 4924 15037 4928
rect 14973 4868 14977 4924
rect 14977 4868 15033 4924
rect 15033 4868 15037 4924
rect 14973 4864 15037 4868
rect 15053 4924 15117 4928
rect 15053 4868 15057 4924
rect 15057 4868 15113 4924
rect 15113 4868 15117 4924
rect 15053 4864 15117 4868
rect 17908 4524 17972 4588
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 4577 4380 4641 4384
rect 4577 4324 4581 4380
rect 4581 4324 4637 4380
rect 4637 4324 4641 4380
rect 4577 4320 4641 4324
rect 4657 4380 4721 4384
rect 4657 4324 4661 4380
rect 4661 4324 4717 4380
rect 4717 4324 4721 4380
rect 4657 4320 4721 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 18278 4380 18342 4384
rect 18278 4324 18282 4380
rect 18282 4324 18338 4380
rect 18338 4324 18342 4380
rect 18278 4320 18342 4324
rect 18358 4380 18422 4384
rect 18358 4324 18362 4380
rect 18362 4324 18418 4380
rect 18418 4324 18422 4380
rect 18358 4320 18422 4324
rect 18438 4380 18502 4384
rect 18438 4324 18442 4380
rect 18442 4324 18498 4380
rect 18498 4324 18502 4380
rect 18438 4320 18502 4324
rect 18518 4380 18582 4384
rect 18518 4324 18522 4380
rect 18522 4324 18578 4380
rect 18578 4324 18582 4380
rect 18518 4320 18582 4324
rect 3924 4252 3988 4316
rect 14044 4176 14108 4180
rect 14044 4120 14094 4176
rect 14094 4120 14108 4176
rect 14044 4116 14108 4120
rect 17908 4116 17972 4180
rect 7882 3836 7946 3840
rect 7882 3780 7886 3836
rect 7886 3780 7942 3836
rect 7942 3780 7946 3836
rect 7882 3776 7946 3780
rect 7962 3836 8026 3840
rect 7962 3780 7966 3836
rect 7966 3780 8022 3836
rect 8022 3780 8026 3836
rect 7962 3776 8026 3780
rect 8042 3836 8106 3840
rect 8042 3780 8046 3836
rect 8046 3780 8102 3836
rect 8102 3780 8106 3836
rect 8042 3776 8106 3780
rect 8122 3836 8186 3840
rect 8122 3780 8126 3836
rect 8126 3780 8182 3836
rect 8182 3780 8186 3836
rect 8122 3776 8186 3780
rect 14813 3836 14877 3840
rect 14813 3780 14817 3836
rect 14817 3780 14873 3836
rect 14873 3780 14877 3836
rect 14813 3776 14877 3780
rect 14893 3836 14957 3840
rect 14893 3780 14897 3836
rect 14897 3780 14953 3836
rect 14953 3780 14957 3836
rect 14893 3776 14957 3780
rect 14973 3836 15037 3840
rect 14973 3780 14977 3836
rect 14977 3780 15033 3836
rect 15033 3780 15037 3836
rect 14973 3776 15037 3780
rect 15053 3836 15117 3840
rect 15053 3780 15057 3836
rect 15057 3780 15113 3836
rect 15113 3780 15117 3836
rect 15053 3776 15117 3780
rect 8892 3436 8956 3500
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 4577 3292 4641 3296
rect 4577 3236 4581 3292
rect 4581 3236 4637 3292
rect 4637 3236 4641 3292
rect 4577 3232 4641 3236
rect 4657 3292 4721 3296
rect 4657 3236 4661 3292
rect 4661 3236 4717 3292
rect 4717 3236 4721 3292
rect 4657 3232 4721 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 18278 3292 18342 3296
rect 18278 3236 18282 3292
rect 18282 3236 18338 3292
rect 18338 3236 18342 3292
rect 18278 3232 18342 3236
rect 18358 3292 18422 3296
rect 18358 3236 18362 3292
rect 18362 3236 18418 3292
rect 18418 3236 18422 3292
rect 18358 3232 18422 3236
rect 18438 3292 18502 3296
rect 18438 3236 18442 3292
rect 18442 3236 18498 3292
rect 18498 3236 18502 3292
rect 18438 3232 18502 3236
rect 18518 3292 18582 3296
rect 18518 3236 18522 3292
rect 18522 3236 18578 3292
rect 18578 3236 18582 3292
rect 18518 3232 18582 3236
rect 10364 3028 10428 3092
rect 9444 2756 9508 2820
rect 7882 2748 7946 2752
rect 7882 2692 7886 2748
rect 7886 2692 7942 2748
rect 7942 2692 7946 2748
rect 7882 2688 7946 2692
rect 7962 2748 8026 2752
rect 7962 2692 7966 2748
rect 7966 2692 8022 2748
rect 8022 2692 8026 2748
rect 7962 2688 8026 2692
rect 8042 2748 8106 2752
rect 8042 2692 8046 2748
rect 8046 2692 8102 2748
rect 8102 2692 8106 2748
rect 8042 2688 8106 2692
rect 8122 2748 8186 2752
rect 8122 2692 8126 2748
rect 8126 2692 8182 2748
rect 8182 2692 8186 2748
rect 8122 2688 8186 2692
rect 14813 2748 14877 2752
rect 14813 2692 14817 2748
rect 14817 2692 14873 2748
rect 14873 2692 14877 2748
rect 14813 2688 14877 2692
rect 14893 2748 14957 2752
rect 14893 2692 14897 2748
rect 14897 2692 14953 2748
rect 14953 2692 14957 2748
rect 14893 2688 14957 2692
rect 14973 2748 15037 2752
rect 14973 2692 14977 2748
rect 14977 2692 15033 2748
rect 15033 2692 15037 2748
rect 14973 2688 15037 2692
rect 15053 2748 15117 2752
rect 15053 2692 15057 2748
rect 15057 2692 15113 2748
rect 15113 2692 15117 2748
rect 15053 2688 15117 2692
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 4577 2204 4641 2208
rect 4577 2148 4581 2204
rect 4581 2148 4637 2204
rect 4637 2148 4641 2204
rect 4577 2144 4641 2148
rect 4657 2204 4721 2208
rect 4657 2148 4661 2204
rect 4661 2148 4717 2204
rect 4717 2148 4721 2204
rect 4657 2144 4721 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 18278 2204 18342 2208
rect 18278 2148 18282 2204
rect 18282 2148 18338 2204
rect 18338 2148 18342 2204
rect 18278 2144 18342 2148
rect 18358 2204 18422 2208
rect 18358 2148 18362 2204
rect 18362 2148 18418 2204
rect 18418 2148 18422 2204
rect 18358 2144 18422 2148
rect 18438 2204 18502 2208
rect 18438 2148 18442 2204
rect 18442 2148 18498 2204
rect 18498 2148 18502 2204
rect 18438 2144 18502 2148
rect 18518 2204 18582 2208
rect 18518 2148 18522 2204
rect 18522 2148 18578 2204
rect 18578 2148 18582 2204
rect 18518 2144 18582 2148
<< metal4 >>
rect 4409 20704 4729 20720
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 19616 4729 20640
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 18528 4729 19552
rect 7874 20160 8195 20720
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8195 20160
rect 7603 19412 7669 19413
rect 7603 19348 7604 19412
rect 7668 19348 7669 19412
rect 7603 19347 7669 19348
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 17440 4729 18464
rect 6867 18460 6933 18461
rect 6867 18396 6868 18460
rect 6932 18396 6933 18460
rect 6867 18395 6933 18396
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 16352 4729 17376
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 15264 4729 16288
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 14176 4729 15200
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 13088 4729 14112
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 12000 4729 13024
rect 6870 12749 6930 18395
rect 7051 17508 7117 17509
rect 7051 17444 7052 17508
rect 7116 17444 7117 17508
rect 7051 17443 7117 17444
rect 6867 12748 6933 12749
rect 6867 12684 6868 12748
rect 6932 12684 6933 12748
rect 6867 12683 6933 12684
rect 5763 12612 5829 12613
rect 5763 12548 5764 12612
rect 5828 12548 5829 12612
rect 5763 12547 5829 12548
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 3923 11932 3989 11933
rect 3923 11868 3924 11932
rect 3988 11868 3989 11932
rect 3923 11867 3989 11868
rect 3371 11524 3437 11525
rect 3371 11460 3372 11524
rect 3436 11460 3437 11524
rect 3371 11459 3437 11460
rect 3374 8941 3434 11459
rect 3371 8940 3437 8941
rect 3371 8876 3372 8940
rect 3436 8876 3437 8940
rect 3371 8875 3437 8876
rect 3926 4317 3986 11867
rect 4409 10912 4729 11936
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 9824 4729 10848
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 8736 4729 9760
rect 5766 9757 5826 12547
rect 6870 11933 6930 12683
rect 6867 11932 6933 11933
rect 6867 11868 6868 11932
rect 6932 11868 6933 11932
rect 6867 11867 6933 11868
rect 7054 10301 7114 17443
rect 7419 16284 7485 16285
rect 7419 16220 7420 16284
rect 7484 16220 7485 16284
rect 7419 16219 7485 16220
rect 7235 15604 7301 15605
rect 7235 15540 7236 15604
rect 7300 15540 7301 15604
rect 7235 15539 7301 15540
rect 7051 10300 7117 10301
rect 7051 10236 7052 10300
rect 7116 10236 7117 10300
rect 7051 10235 7117 10236
rect 5763 9756 5829 9757
rect 5763 9692 5764 9756
rect 5828 9692 5829 9756
rect 5763 9691 5829 9692
rect 7238 8805 7298 15539
rect 7422 14381 7482 16219
rect 7419 14380 7485 14381
rect 7419 14316 7420 14380
rect 7484 14316 7485 14380
rect 7419 14315 7485 14316
rect 7422 11797 7482 14315
rect 7419 11796 7485 11797
rect 7419 11732 7420 11796
rect 7484 11732 7485 11796
rect 7419 11731 7485 11732
rect 7606 10570 7666 19347
rect 7422 10510 7666 10570
rect 7874 19072 8195 20096
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 8523 19412 8589 19413
rect 8523 19348 8524 19412
rect 8588 19348 8589 19412
rect 8523 19347 8589 19348
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8195 19072
rect 7874 17984 8195 19008
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8195 17984
rect 7874 16896 8195 17920
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8195 16896
rect 7874 15808 8195 16832
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8195 15808
rect 7874 14720 8195 15744
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8195 14720
rect 7874 13632 8195 14656
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8195 13632
rect 7874 12544 8195 13568
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8195 12544
rect 7874 11456 8195 12480
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8195 11456
rect 7235 8804 7301 8805
rect 7235 8740 7236 8804
rect 7300 8740 7301 8804
rect 7235 8739 7301 8740
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 7648 4729 8672
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 6560 4729 7584
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 5472 4729 6496
rect 7238 6221 7298 8739
rect 7422 8397 7482 10510
rect 7603 10436 7669 10437
rect 7603 10372 7604 10436
rect 7668 10372 7669 10436
rect 7603 10371 7669 10372
rect 7606 8533 7666 10371
rect 7874 10368 8195 11392
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8195 10368
rect 7874 9280 8195 10304
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8195 9280
rect 7603 8532 7669 8533
rect 7603 8468 7604 8532
rect 7668 8468 7669 8532
rect 7603 8467 7669 8468
rect 7419 8396 7485 8397
rect 7419 8332 7420 8396
rect 7484 8332 7485 8396
rect 7419 8331 7485 8332
rect 7235 6220 7301 6221
rect 7235 6156 7236 6220
rect 7300 6156 7301 6220
rect 7235 6155 7301 6156
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 4384 4729 5408
rect 7606 5405 7666 8467
rect 7874 8192 8195 9216
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8195 8192
rect 7874 7104 8195 8128
rect 8526 7853 8586 19347
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 9811 17100 9877 17101
rect 9811 17036 9812 17100
rect 9876 17036 9877 17100
rect 9811 17035 9877 17036
rect 9259 16420 9325 16421
rect 9259 16356 9260 16420
rect 9324 16356 9325 16420
rect 9259 16355 9325 16356
rect 8707 13836 8773 13837
rect 8707 13772 8708 13836
rect 8772 13772 8773 13836
rect 8707 13771 8773 13772
rect 8523 7852 8589 7853
rect 8523 7788 8524 7852
rect 8588 7788 8589 7852
rect 8523 7787 8589 7788
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8195 7104
rect 7874 6016 8195 7040
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8195 6016
rect 7603 5404 7669 5405
rect 7603 5340 7604 5404
rect 7668 5340 7669 5404
rect 7603 5339 7669 5340
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 3923 4316 3989 4317
rect 3923 4252 3924 4316
rect 3988 4252 3989 4316
rect 3923 4251 3989 4252
rect 4409 3296 4729 4320
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 2208 4729 3232
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2128 4729 2144
rect 7874 4928 8195 5952
rect 8526 5810 8586 7787
rect 8710 5949 8770 13771
rect 8891 13564 8957 13565
rect 8891 13500 8892 13564
rect 8956 13500 8957 13564
rect 8891 13499 8957 13500
rect 8894 10301 8954 13499
rect 9262 10981 9322 16355
rect 9627 14652 9693 14653
rect 9627 14588 9628 14652
rect 9692 14588 9693 14652
rect 9627 14587 9693 14588
rect 9630 14109 9690 14587
rect 9627 14108 9693 14109
rect 9627 14044 9628 14108
rect 9692 14044 9693 14108
rect 9627 14043 9693 14044
rect 9443 13564 9509 13565
rect 9443 13500 9444 13564
rect 9508 13500 9509 13564
rect 9443 13499 9509 13500
rect 9259 10980 9325 10981
rect 9259 10916 9260 10980
rect 9324 10916 9325 10980
rect 9259 10915 9325 10916
rect 8891 10300 8957 10301
rect 8891 10236 8892 10300
rect 8956 10236 8957 10300
rect 8891 10235 8957 10236
rect 9262 10029 9322 10915
rect 9446 10437 9506 13499
rect 9443 10436 9509 10437
rect 9443 10372 9444 10436
rect 9508 10372 9509 10436
rect 9443 10371 9509 10372
rect 9630 10301 9690 14043
rect 9814 10437 9874 17035
rect 10547 16828 10613 16829
rect 10547 16764 10548 16828
rect 10612 16764 10613 16828
rect 10547 16763 10613 16764
rect 9995 14924 10061 14925
rect 9995 14860 9996 14924
rect 10060 14860 10061 14924
rect 9995 14859 10061 14860
rect 9998 11389 10058 14859
rect 10363 14788 10429 14789
rect 10363 14724 10364 14788
rect 10428 14724 10429 14788
rect 10363 14723 10429 14724
rect 9995 11388 10061 11389
rect 9995 11324 9996 11388
rect 10060 11324 10061 11388
rect 9995 11323 10061 11324
rect 10366 10709 10426 14723
rect 10363 10708 10429 10709
rect 10363 10644 10364 10708
rect 10428 10644 10429 10708
rect 10363 10643 10429 10644
rect 9811 10436 9877 10437
rect 9811 10372 9812 10436
rect 9876 10372 9877 10436
rect 9811 10371 9877 10372
rect 9627 10300 9693 10301
rect 9627 10236 9628 10300
rect 9692 10236 9693 10300
rect 9627 10235 9693 10236
rect 9259 10028 9325 10029
rect 9259 9964 9260 10028
rect 9324 9964 9325 10028
rect 9259 9963 9325 9964
rect 10363 9756 10429 9757
rect 10363 9692 10364 9756
rect 10428 9692 10429 9756
rect 10363 9691 10429 9692
rect 8707 5948 8773 5949
rect 8707 5884 8708 5948
rect 8772 5884 8773 5948
rect 8707 5883 8773 5884
rect 8526 5750 8954 5810
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8195 4928
rect 7874 3840 8195 4864
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8195 3840
rect 7874 2752 8195 3776
rect 8894 3501 8954 5750
rect 9443 5540 9509 5541
rect 9443 5476 9444 5540
rect 9508 5476 9509 5540
rect 9443 5475 9509 5476
rect 8891 3500 8957 3501
rect 8891 3436 8892 3500
rect 8956 3436 8957 3500
rect 8891 3435 8957 3436
rect 9446 2821 9506 5475
rect 10366 3093 10426 9691
rect 10550 8397 10610 16763
rect 11340 16352 11660 17376
rect 14805 20160 15125 20720
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 19072 15125 20096
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 17984 15125 19008
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 16896 15125 17920
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 11835 16556 11901 16557
rect 11835 16492 11836 16556
rect 11900 16492 11901 16556
rect 11835 16491 11901 16492
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11099 13836 11165 13837
rect 11099 13772 11100 13836
rect 11164 13772 11165 13836
rect 11099 13771 11165 13772
rect 10915 13428 10981 13429
rect 10915 13364 10916 13428
rect 10980 13364 10981 13428
rect 10915 13363 10981 13364
rect 10547 8396 10613 8397
rect 10547 8332 10548 8396
rect 10612 8332 10613 8396
rect 10547 8331 10613 8332
rect 10918 8261 10978 13363
rect 11102 12477 11162 13771
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11099 12476 11165 12477
rect 11099 12412 11100 12476
rect 11164 12412 11165 12476
rect 11099 12411 11165 12412
rect 11102 10437 11162 12411
rect 11340 12000 11660 13024
rect 11838 12341 11898 16491
rect 14805 15808 15125 16832
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 12571 15332 12637 15333
rect 12571 15268 12572 15332
rect 12636 15268 12637 15332
rect 12571 15267 12637 15268
rect 11835 12340 11901 12341
rect 11835 12276 11836 12340
rect 11900 12276 11901 12340
rect 11835 12275 11901 12276
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 12019 11932 12085 11933
rect 12019 11868 12020 11932
rect 12084 11868 12085 11932
rect 12019 11867 12085 11868
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11099 10436 11165 10437
rect 11099 10372 11100 10436
rect 11164 10372 11165 10436
rect 11099 10371 11165 10372
rect 11340 9824 11660 10848
rect 11835 10300 11901 10301
rect 11835 10236 11836 10300
rect 11900 10236 11901 10300
rect 11835 10235 11901 10236
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11099 8804 11165 8805
rect 11099 8740 11100 8804
rect 11164 8740 11165 8804
rect 11099 8739 11165 8740
rect 10915 8260 10981 8261
rect 10915 8196 10916 8260
rect 10980 8196 10981 8260
rect 10915 8195 10981 8196
rect 11102 7173 11162 8739
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11099 7172 11165 7173
rect 11099 7108 11100 7172
rect 11164 7108 11165 7172
rect 11099 7107 11165 7108
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11838 5133 11898 10235
rect 12022 6493 12082 11867
rect 12574 11117 12634 15267
rect 14805 14720 15125 15744
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 13632 15125 14656
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 12544 15125 13568
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 11456 15125 12480
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 12571 11116 12637 11117
rect 12571 11052 12572 11116
rect 12636 11052 12637 11116
rect 12571 11051 12637 11052
rect 12574 9349 12634 11051
rect 14805 10368 15125 11392
rect 18270 20704 18591 20720
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18591 20704
rect 18270 19616 18591 20640
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18591 19616
rect 18270 18528 18591 19552
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18591 18528
rect 18270 17440 18591 18464
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18591 17440
rect 18270 16352 18591 17376
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18591 16352
rect 18270 15264 18591 16288
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18591 15264
rect 18270 14176 18591 15200
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18591 14176
rect 18270 13088 18591 14112
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18591 13088
rect 18270 12000 18591 13024
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18591 12000
rect 17907 11116 17973 11117
rect 17907 11052 17908 11116
rect 17972 11052 17973 11116
rect 17907 11051 17973 11052
rect 17910 10845 17970 11051
rect 18270 10912 18591 11936
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18591 10912
rect 17907 10844 17973 10845
rect 17907 10780 17908 10844
rect 17972 10780 17973 10844
rect 17907 10779 17973 10780
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 12571 9348 12637 9349
rect 12571 9284 12572 9348
rect 12636 9284 12637 9348
rect 12571 9283 12637 9284
rect 14805 9280 15125 10304
rect 17907 10300 17973 10301
rect 17907 10236 17908 10300
rect 17972 10236 17973 10300
rect 17907 10235 17973 10236
rect 17910 10029 17970 10235
rect 17907 10028 17973 10029
rect 17907 9964 17908 10028
rect 17972 9964 17973 10028
rect 17907 9963 17973 9964
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14043 9212 14109 9213
rect 14043 9148 14044 9212
rect 14108 9148 14109 9212
rect 14043 9147 14109 9148
rect 13123 8668 13189 8669
rect 13123 8604 13124 8668
rect 13188 8604 13189 8668
rect 13123 8603 13189 8604
rect 13126 8397 13186 8603
rect 13123 8396 13189 8397
rect 13123 8332 13124 8396
rect 13188 8332 13189 8396
rect 13123 8331 13189 8332
rect 12019 6492 12085 6493
rect 12019 6428 12020 6492
rect 12084 6428 12085 6492
rect 12019 6427 12085 6428
rect 11835 5132 11901 5133
rect 11835 5068 11836 5132
rect 11900 5068 11901 5132
rect 11835 5067 11901 5068
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 14046 4181 14106 9147
rect 14805 8192 15125 9216
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 7104 15125 8128
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 6016 15125 7040
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 4928 15125 5952
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14043 4180 14109 4181
rect 14043 4116 14044 4180
rect 14108 4116 14109 4180
rect 14043 4115 14109 4116
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 10363 3092 10429 3093
rect 10363 3028 10364 3092
rect 10428 3028 10429 3092
rect 10363 3027 10429 3028
rect 9443 2820 9509 2821
rect 9443 2756 9444 2820
rect 9508 2756 9509 2820
rect 9443 2755 9509 2756
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8195 2752
rect 7874 2128 8195 2688
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 14805 3840 15125 4864
rect 18270 9824 18591 10848
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18591 9824
rect 18270 8736 18591 9760
rect 19195 9212 19261 9213
rect 19195 9148 19196 9212
rect 19260 9148 19261 9212
rect 19195 9147 19261 9148
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18591 8736
rect 18270 7648 18591 8672
rect 18827 8668 18893 8669
rect 18827 8604 18828 8668
rect 18892 8604 18893 8668
rect 18827 8603 18893 8604
rect 18830 8397 18890 8603
rect 18827 8396 18893 8397
rect 18827 8332 18828 8396
rect 18892 8332 18893 8396
rect 18827 8331 18893 8332
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18591 7648
rect 18270 6560 18591 7584
rect 19198 6629 19258 9147
rect 19195 6628 19261 6629
rect 19195 6564 19196 6628
rect 19260 6564 19261 6628
rect 19195 6563 19261 6564
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18591 6560
rect 18270 5472 18591 6496
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18591 5472
rect 17907 4588 17973 4589
rect 17907 4524 17908 4588
rect 17972 4524 17973 4588
rect 17907 4523 17973 4524
rect 17910 4181 17970 4523
rect 18270 4384 18591 5408
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18591 4384
rect 17907 4180 17973 4181
rect 17907 4116 17908 4180
rect 17972 4116 17973 4180
rect 17907 4115 17973 4116
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 2752 15125 3776
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2128 15125 2688
rect 18270 3296 18591 4320
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18591 3296
rect 18270 2208 18591 3232
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18591 2208
rect 18270 2128 18591 2144
use sky130_fd_sc_hd__fill_2  FILLER_1_11 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1380 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2484 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A1 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608910539
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2484 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3036 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 3128 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_4__A0
timestamp 1608910539
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_4__A1
timestamp 1608910539
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1608910539
transform 1 0 3312 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _051_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3312 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32
timestamp 1608910539
transform 1 0 4048 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608910539
transform 1 0 4140 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_4_
timestamp 1608910539
transform 1 0 4140 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 4324 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_1_51
timestamp 1608910539
transform 1 0 5796 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A0
timestamp 1608910539
transform 1 0 5796 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608910539
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608910539
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1608910539
transform 1 0 4968 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1608910539
transform 1 0 5980 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_2_
timestamp 1608910539
transform 1 0 5888 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63
timestamp 1608910539
transform 1 0 6900 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_4__A0
timestamp 1608910539
transform 1 0 6992 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_4__A1
timestamp 1608910539
transform 1 0 7176 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 8464 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_5_
timestamp 1608910539
transform 1 0 8188 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_4_
timestamp 1608910539
transform 1 0 7360 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 6992 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90
timestamp 1608910539
transform 1 0 9384 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 9200 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 9016 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608910539
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 10580 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1608910539
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1608910539
transform 1 0 9016 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9844 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_1_111
timestamp 1608910539
transform 1 0 11316 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1608910539
transform 1 0 11316 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1608910539
transform 1 0 11408 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A0
timestamp 1608910539
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1608910539
transform 1 0 11500 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _096_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 11592 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608910539
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608910539
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1608910539
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 12420 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_1_145
timestamp 1608910539
transform 1 0 14444 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 13892 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1608910539
transform 1 0 14168 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1608910539
transform 1 0 13800 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1608910539
transform 1 0 13432 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_150
timestamp 1608910539
transform 1 0 14904 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 14536 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1608910539
transform 1 0 14996 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1608910539
transform 1 0 14536 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1608910539
transform 1 0 15088 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608910539
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 15364 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1608910539
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_164
timestamp 1608910539
transform 1 0 16192 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1608910539
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 15916 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1608910539
transform 1 0 15824 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_173
timestamp 1608910539
transform 1 0 17020 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 16836 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1608910539
transform 1 0 17112 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1608910539
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1608910539
transform 1 0 16836 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1608910539
transform 1 0 16468 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1608910539
transform 1 0 16468 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_184
timestamp 1608910539
transform 1 0 18032 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_185
timestamp 1608910539
transform 1 0 18124 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1608910539
transform 1 0 17572 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1608910539
transform 1 0 17756 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 17940 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608910539
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608910539
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1608910539
transform 1 0 18124 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1608910539
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1608910539
transform 1 0 19228 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1608910539
transform 1 0 19044 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1608910539
transform 1 0 18952 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1608910539
transform 1 0 18676 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_207
timestamp 1608910539
transform 1 0 20148 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 19780 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 19412 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1608910539
transform 1 0 19964 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1608910539
transform 1 0 19596 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1608910539
transform 1 0 20148 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1608910539
transform 1 0 19780 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1608910539
transform 1 0 21068 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_222
timestamp 1608910539
transform 1 0 21528 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_218 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 21160 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1608910539
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1608910539
transform 1 0 20884 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608910539
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608910539
transform -1 0 21896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608910539
transform -1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1608910539
transform 1 0 20516 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_11
timestamp 1608910539
transform 1 0 2116 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1608910539
transform 1 0 1380 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608910539
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1608910539
transform 1 0 2300 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608910539
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1608910539
transform 1 0 3128 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4048 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_48
timestamp 1608910539
transform 1 0 5520 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 5704 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_1_
timestamp 1608910539
transform 1 0 5888 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 6716 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 8556 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_5__A0
timestamp 1608910539
transform 1 0 8372 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_5__A1
timestamp 1608910539
transform 1 0 8188 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8740 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608910539
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9660 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_111
timestamp 1608910539
transform 1 0 11316 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 11132 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 11500 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1608910539
transform 1 0 13800 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1608910539
transform 1 0 12972 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608910539
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1608910539
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1608910539
transform 1 0 16100 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1608910539
transform 1 0 14628 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1608910539
transform 1 0 18124 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 16652 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1608910539
transform 1 0 18952 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1608910539
transform 1 0 19780 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_215
timestamp 1608910539
transform 1 0 20884 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_210
timestamp 1608910539
transform 1 0 20424 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608910539
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608910539
transform -1 0 21896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1608910539
transform 1 0 1380 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608910539
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1608910539
transform 1 0 1932 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 2760 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_34
timestamp 1608910539
transform 1 0 4232 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_62
timestamp 1608910539
transform 1 0 6808 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_60
timestamp 1608910539
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608910539
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1608910539
transform 1 0 5796 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1608910539
transform 1 0 4968 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_81
timestamp 1608910539
transform 1 0 8556 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1608910539
transform 1 0 8648 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1608910539
transform 1 0 6900 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_3_104
timestamp 1608910539
transform 1 0 10672 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1608910539
transform 1 0 9844 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_110
timestamp 1608910539
transform 1 0 11224 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1608910539
transform 1 0 12604 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608910539
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1608910539
transform 1 0 11316 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 12788 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1608910539
transform 1 0 13800 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12972 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_147
timestamp 1608910539
transform 1 0 14628 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_4__A0
timestamp 1608910539
transform 1 0 15916 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_4_
timestamp 1608910539
transform 1 0 15088 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 16100 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1608910539
transform 1 0 14720 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1608910539
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A0
timestamp 1608910539
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608910539
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 18032 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1608910539
transform 1 0 19504 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_3_211
timestamp 1608910539
transform 1 0 20516 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 20332 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608910539
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_19
timestamp 1608910539
transform 1 0 2852 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 2944 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608910539
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 1380 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_4_39
timestamp 1608910539
transform 1 0 4692 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_35
timestamp 1608910539
transform 1 0 4324 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 4508 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608910539
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1608910539
transform 1 0 3128 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1608910539
transform 1 0 4784 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1608910539
transform 1 0 4048 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 5612 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l5_in_0_
timestamp 1608910539
transform 1 0 7084 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1608910539
transform 1 0 7912 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8740 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_104
timestamp 1608910539
transform 1 0 10672 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608910539
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1608910539
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_125
timestamp 1608910539
transform 1 0 12604 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_120
timestamp 1608910539
transform 1 0 12144 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_4__A1
timestamp 1608910539
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A0
timestamp 1608910539
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 10948 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 11960 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1608910539
transform 1 0 11132 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1608910539
transform 1 0 14168 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12696 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_4__A1
timestamp 1608910539
transform 1 0 15272 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608910539
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 15456 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_174
timestamp 1608910539
transform 1 0 17112 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1608910539
transform 1 0 16928 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 17480 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1608910539
transform 1 0 17664 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_4_207
timestamp 1608910539
transform 1 0 20148 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1608910539
transform 1 0 19320 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1608910539
transform 1 0 18492 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_215
timestamp 1608910539
transform 1 0 20884 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_213
timestamp 1608910539
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608910539
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608910539
transform -1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1608910539
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608910539
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 1748 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1608910539
transform 1 0 4692 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 3220 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_5_62
timestamp 1608910539
transform 1 0 6808 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608910539
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1608910539
transform 1 0 5520 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_77
timestamp 1608910539
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_67
timestamp 1608910539
transform 1 0 7268 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 6900 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 7084 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_3_
timestamp 1608910539
transform 1 0 7360 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1608910539
transform 1 0 8280 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1608910539
transform 1 0 10580 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 9108 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_5_121
timestamp 1608910539
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608910539
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_4_
timestamp 1608910539
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1608910539
transform 1 0 11408 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_132
timestamp 1608910539
transform 1 0 13248 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_4_
timestamp 1608910539
transform 1 0 14168 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1608910539
transform 1 0 13340 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_151
timestamp 1608910539
transform 1 0 14996 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 15088 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_5_184
timestamp 1608910539
transform 1 0 18032 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_177
timestamp 1608910539
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608910539
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1608910539
transform 1 0 16560 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 18124 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1608910539
transform 1 0 19596 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_222
timestamp 1608910539
transform 1 0 21528 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_210
timestamp 1608910539
transform 1 0 20424 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608910539
transform -1 0 21896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_9
timestamp 1608910539
transform 1 0 1932 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1608910539
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1608910539
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608910539
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608910539
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1656 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_12
timestamp 1608910539
transform 1 0 2208 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_4__A1
timestamp 1608910539
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1608910539
transform 1 0 2300 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1608910539
transform 1 0 2024 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_7_31
timestamp 1608910539
transform 1 0 3956 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_21
timestamp 1608910539
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_32
timestamp 1608910539
transform 1 0 4048 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608910539
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1608910539
transform 1 0 3128 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_3_
timestamp 1608910539
transform 1 0 3128 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1608910539
transform 1 0 4692 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4140 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_6_51
timestamp 1608910539
transform 1 0 5796 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6072 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 5704 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 5612 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608910539
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1608910539
transform 1 0 6256 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1608910539
transform 1 0 5888 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1608910539
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_7_80
timestamp 1608910539
transform 1 0 8464 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__A0
timestamp 1608910539
transform 1 0 7084 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__A1
timestamp 1608910539
transform 1 0 7268 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_4_
timestamp 1608910539
transform 1 0 8556 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_7_
timestamp 1608910539
transform 1 0 7636 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_6_
timestamp 1608910539
transform 1 0 7728 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1608910539
transform 1 0 8556 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1608910539
transform 1 0 7452 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_103
timestamp 1608910539
transform 1 0 10580 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 10672 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 9384 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_4__A0
timestamp 1608910539
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608910539
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1608910539
transform 1 0 9568 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9660 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 10856 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1608910539
transform 1 0 11040 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1608910539
transform 1 0 11132 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_7_119
timestamp 1608910539
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_123
timestamp 1608910539
transform 1 0 12420 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_118
timestamp 1608910539
transform 1 0 11960 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 11868 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 12236 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_4__A0
timestamp 1608910539
transform 1 0 12052 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608910539
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1608910539
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12512 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_134
timestamp 1608910539
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_4__A0
timestamp 1608910539
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_4__A1
timestamp 1608910539
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 13984 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 14168 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1608910539
transform 1 0 14352 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 14168 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_7_158
timestamp 1608910539
transform 1 0 15640 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_156
timestamp 1608910539
transform 1 0 15456 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1608910539
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__A0
timestamp 1608910539
transform 1 0 15548 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608910539
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 15732 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_3_
timestamp 1608910539
transform 1 0 15732 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 16560 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1608910539
transform 1 0 16560 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1608910539
transform 1 0 16744 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_7_184
timestamp 1608910539
transform 1 0 18032 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_180
timestamp 1608910539
transform 1 0 17664 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608910539
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1608910539
transform 1 0 18124 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1608910539
transform 1 0 17572 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1608910539
transform 1 0 17388 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_194
timestamp 1608910539
transform 1 0 18952 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_190
timestamp 1608910539
transform 1 0 18584 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 18400 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 20148 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 19228 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 18676 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1608910539
transform 1 0 21436 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_213
timestamp 1608910539
transform 1 0 20700 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_215
timestamp 1608910539
transform 1 0 20884 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1608910539
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608910539
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608910539
transform -1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608910539
transform -1 0 21896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1608910539
transform 1 0 1380 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_4__A0
timestamp 1608910539
transform 1 0 1472 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608910539
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1608910539
transform 1 0 1932 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_4_
timestamp 1608910539
transform 1 0 2760 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1608910539
transform 1 0 1656 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1608910539
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608910539
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4048 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 5520 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 8556 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A0
timestamp 1608910539
transform 1 0 8188 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 8004 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_7__A1
timestamp 1608910539
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1608910539
transform 1 0 6992 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_8_87
timestamp 1608910539
transform 1 0 9108 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8924 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_4__A1
timestamp 1608910539
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608910539
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_3_
timestamp 1608910539
transform 1 0 9844 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1608910539
transform 1 0 10672 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_111
timestamp 1608910539
transform 1 0 11316 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_107
timestamp 1608910539
transform 1 0 10948 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 11408 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 11592 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 14168 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1608910539
transform 1 0 13064 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1608910539
transform 1 0 13892 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_159
timestamp 1608910539
transform 1 0 15732 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_154
timestamp 1608910539
transform 1 0 15272 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 16008 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 15548 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 15364 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608910539
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1608910539
transform 1 0 16192 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 17848 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1608910539
transform 1 0 18032 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1608910539
transform 1 0 17020 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_2_
timestamp 1608910539
transform 1 0 18860 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_7_
timestamp 1608910539
transform 1 0 19688 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_219
timestamp 1608910539
transform 1 0 21252 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1608910539
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_4__A0
timestamp 1608910539
transform 1 0 21068 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_4__A1
timestamp 1608910539
transform 1 0 20884 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_7__A1
timestamp 1608910539
transform 1 0 20516 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608910539
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608910539
transform -1 0 21896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1608910539
transform 1 0 1748 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1608910539
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608910539
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 1840 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_9_37
timestamp 1608910539
transform 1 0 4508 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_24
timestamp 1608910539
transform 1 0 3312 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1608910539
transform 1 0 3680 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_60
timestamp 1608910539
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608910539
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1608910539
transform 1 0 5796 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1608910539
transform 1 0 4968 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1608910539
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 7636 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 10304 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A0
timestamp 1608910539
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 10672 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1608910539
transform 1 0 9108 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_115
timestamp 1608910539
transform 1 0 11684 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_4__A0
timestamp 1608910539
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_4__A1
timestamp 1608910539
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608910539
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1608910539
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1608910539
transform 1 0 10856 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1608910539
transform 1 0 14076 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_4_
timestamp 1608910539
transform 1 0 13248 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_150
timestamp 1608910539
transform 1 0 14904 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 14996 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1608910539
transform 1 0 15180 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1608910539
transform 1 0 16008 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_175
timestamp 1608910539
transform 1 0 17204 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__A1
timestamp 1608910539
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__A0
timestamp 1608910539
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 16836 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608910539
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_6_
timestamp 1608910539
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_195
timestamp 1608910539
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_4_
timestamp 1608910539
transform 1 0 19504 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1608910539
transform 1 0 19228 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_222
timestamp 1608910539
transform 1 0 21528 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 21344 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 21160 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608910539
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1608910539
transform 1 0 20332 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_5
timestamp 1608910539
transform 1 0 1564 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_7__A1
timestamp 1608910539
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608910539
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 1656 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_10_38
timestamp 1608910539
transform 1 0 4600 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_32
timestamp 1608910539
transform 1 0 4048 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 4692 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608910539
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1608910539
transform 1 0 3128 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1608910539
transform 1 0 6716 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_3_
timestamp 1608910539
transform 1 0 5060 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_2_
timestamp 1608910539
transform 1 0 5888 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_70
timestamp 1608910539
transform 1 0 7544 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 7636 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1608910539
transform 1 0 7912 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8740 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_93
timestamp 1608910539
transform 1 0 9660 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 9936 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 9752 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608910539
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1608910539
transform 1 0 10120 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 12420 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 10948 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12696 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1608910539
transform 1 0 14352 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1608910539
transform 1 0 13524 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_163
timestamp 1608910539
transform 1 0 16100 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608910539
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16192 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_2_
timestamp 1608910539
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_173
timestamp 1608910539
transform 1 0 17020 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1608910539
transform 1 0 17112 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 17940 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_203
timestamp 1608910539
transform 1 0 19780 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 19596 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_5__A1
timestamp 1608910539
transform 1 0 19412 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1608910539
transform 1 0 19964 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_219
timestamp 1608910539
transform 1 0 21252 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A0
timestamp 1608910539
transform 1 0 21068 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 20884 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 21436 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608910539
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608910539
transform -1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_18
timestamp 1608910539
transform 1 0 2760 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608910539
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1380 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1608910539
transform 1 0 1932 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 2852 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_39
timestamp 1608910539
transform 1 0 4692 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_35
timestamp 1608910539
transform 1 0 4324 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 4784 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1608910539
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608910539
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1608910539
transform 1 0 6256 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_79
timestamp 1608910539
transform 1 0 8372 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_67
timestamp 1608910539
transform 1 0 7268 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 7084 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1608910539
transform 1 0 7360 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 8464 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1608910539
transform 1 0 9936 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_105
timestamp 1608910539
transform 1 0 10764 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608910539
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1608910539
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10856 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_132
timestamp 1608910539
transform 1 0 13248 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 13524 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 13340 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 13708 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 15180 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608910539
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_5_
timestamp 1608910539
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_3_
timestamp 1608910539
transform 1 0 16652 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1608910539
transform 1 0 17480 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1608910539
transform 1 0 18860 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1608910539
transform 1 0 19688 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_222
timestamp 1608910539
transform 1 0 21528 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 21344 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608910539
transform -1 0 21896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1608910539
transform 1 0 20516 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_4__A1
timestamp 1608910539
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608910539
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_7_
timestamp 1608910539
transform 1 0 1564 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_4_
timestamp 1608910539
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_12_28
timestamp 1608910539
transform 1 0 3680 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_4__A0
timestamp 1608910539
transform 1 0 3496 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608910539
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4048 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1608910539
transform 1 0 3220 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 5520 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 5704 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_12_73
timestamp 1608910539
transform 1 0 7820 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 7636 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 7452 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 7176 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1608910539
transform 1 0 7912 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1608910539
transform 1 0 8740 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608910539
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1608910539
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_115
timestamp 1608910539
transform 1 0 11684 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1608910539
transform 1 0 10856 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_145
timestamp 1608910539
transform 1 0 14444 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_140
timestamp 1608910539
transform 1 0 13984 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_127
timestamp 1608910539
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 14260 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 14076 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 12972 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1608910539
transform 1 0 13156 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_157
timestamp 1608910539
transform 1 0 15548 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1608910539
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 14536 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 14720 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 14904 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608910539
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 15640 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1608910539
transform 1 0 17112 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_3_
timestamp 1608910539
transform 1 0 17940 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 18768 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_12_215
timestamp 1608910539
transform 1 0 20884 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_210
timestamp 1608910539
transform 1 0 20424 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608910539
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608910539
transform -1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_9
timestamp 1608910539
transform 1 0 1932 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3
timestamp 1608910539
transform 1 0 1380 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_5__A0
timestamp 1608910539
transform 1 0 2852 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_5__A1
timestamp 1608910539
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608910539
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608910539
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_3_
timestamp 1608910539
transform 1 0 1564 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_2_
timestamp 1608910539
transform 1 0 2024 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_5_
timestamp 1608910539
transform 1 0 2392 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_14_25
timestamp 1608910539
transform 1 0 3404 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_6__A0
timestamp 1608910539
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_6__A1
timestamp 1608910539
transform 1 0 3036 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_6_
timestamp 1608910539
transform 1 0 3220 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_32
timestamp 1608910539
transform 1 0 4048 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 4140 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608910539
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1608910539
transform 1 0 4324 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1608910539
transform 1 0 4232 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_44
timestamp 1608910539
transform 1 0 5152 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 6072 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608910539
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l4_in_0_
timestamp 1608910539
transform 1 0 5244 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_1_
timestamp 1608910539
transform 1 0 5060 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1608910539
transform 1 0 6256 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1608910539
transform 1 0 5888 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_13_80
timestamp 1608910539
transform 1 0 8464 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7084 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1608910539
transform 1 0 7912 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1608910539
transform 1 0 8740 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 6992 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 8740 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_13_102
timestamp 1608910539
transform 1 0 10488 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608910539
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 9660 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1608910539
transform 1 0 10212 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_109
timestamp 1608910539
transform 1 0 11132 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_123
timestamp 1608910539
transform 1 0 12420 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 11224 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608910539
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l4_in_0_
timestamp 1608910539
transform 1 0 11408 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1608910539
transform 1 0 12512 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10856 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 12236 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 14076 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 14444 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 13892 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 13708 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 14168 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1608910539
transform 1 0 13340 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1608910539
transform 1 0 14260 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1608910539
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 14628 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608910539
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_2_
timestamp 1608910539
transform 1 0 14812 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1608910539
transform 1 0 16100 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1608910539
transform 1 0 15640 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1608910539
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_176
timestamp 1608910539
transform 1 0 17296 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 17112 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 16928 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1608910539
transform 1 0 16468 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_13_184
timestamp 1608910539
transform 1 0 18032 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1608910539
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 17480 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_5__A0
timestamp 1608910539
transform 1 0 17664 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608910539
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_1_
timestamp 1608910539
transform 1 0 18124 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 17388 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 19044 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 18860 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 19228 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1608910539
transform 1 0 18952 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_14_215
timestamp 1608910539
transform 1 0 20884 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1608910539
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_219
timestamp 1608910539
transform 1 0 21252 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608910539
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608910539
transform -1 0 21896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608910539
transform -1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1608910539
transform 1 0 20424 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1608910539
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608910539
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_1_
timestamp 1608910539
transform 1 0 1472 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 2300 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_29
timestamp 1608910539
transform 1 0 3772 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1608910539
transform 1 0 4692 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1608910539
transform 1 0 3864 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 5520 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608910539
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_1_
timestamp 1608910539
transform 1 0 5704 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 6808 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1608910539
transform 1 0 8280 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1608910539
transform 1 0 9108 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9936 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_123
timestamp 1608910539
transform 1 0 12420 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1608910539
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608910539
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1608910539
transform 1 0 11408 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 12512 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1608910539
transform 1 0 13984 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_151
timestamp 1608910539
transform 1 0 14996 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1608910539
transform 1 0 15088 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 15916 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_182
timestamp 1608910539
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_177
timestamp 1608910539
transform 1 0 17388 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 17480 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 17664 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608910539
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1608910539
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 19136 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l5_in_0_
timestamp 1608910539
transform 1 0 19320 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 20148 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1608910539
transform 1 0 18860 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_219
timestamp 1608910539
transform 1 0 21252 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608910539
transform -1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 20700 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608910539
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 1748 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1608910539
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_32
timestamp 1608910539
transform 1 0 4048 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_23
timestamp 1608910539
transform 1 0 3220 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A0
timestamp 1608910539
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608910539
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1608910539
transform 1 0 4140 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_44
timestamp 1608910539
transform 1 0 5152 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 4968 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_3_
timestamp 1608910539
transform 1 0 5244 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_2_
timestamp 1608910539
transform 1 0 6072 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 7728 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 8740 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1608910539
transform 1 0 7912 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1608910539
transform 1 0 6900 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_95
timestamp 1608910539
transform 1 0 9844 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 10396 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608910539
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1608910539
transform 1 0 12236 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 13340 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 13064 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_3_
timestamp 1608910539
transform 1 0 14352 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_2_
timestamp 1608910539
transform 1 0 13524 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608910539
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16100 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_1_
timestamp 1608910539
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_181
timestamp 1608910539
transform 1 0 17756 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1608910539
transform 1 0 16928 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1608910539
transform 1 0 17848 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_16_200
timestamp 1608910539
transform 1 0 19504 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1608910539
transform 1 0 18676 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_219
timestamp 1608910539
transform 1 0 21252 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1608910539
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608910539
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608910539
transform -1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1608910539
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1608910539
transform 1 0 1380 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608910539
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1608910539
transform 1 0 1472 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1608910539
transform 1 0 2944 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_24
timestamp 1608910539
transform 1 0 3312 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1608910539
transform 1 0 4232 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1608910539
transform 1 0 3404 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_62
timestamp 1608910539
transform 1 0 6808 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 5060 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1608910539
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 5244 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6900 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1608910539
transform 1 0 7084 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1608910539
transform 1 0 7912 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1608910539
transform 1 0 8740 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 9752 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 9568 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10304 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1608910539
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_118
timestamp 1608910539
transform 1 0 11960 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 12052 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1608910539
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 13432 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_17_152
timestamp 1608910539
transform 1 0 15088 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 14904 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1608910539
transform 1 0 15364 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 16192 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_184
timestamp 1608910539
transform 1 0 18032 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_180
timestamp 1608910539
transform 1 0 17664 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1608910539
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1608910539
transform 1 0 18124 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_17_198
timestamp 1608910539
transform 1 0 19320 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 19136 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 18952 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_222
timestamp 1608910539
transform 1 0 21528 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_210
timestamp 1608910539
transform 1 0 20424 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608910539
transform -1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1608910539
transform 1 0 21160 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1608910539
transform 1 0 20792 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_17
timestamp 1608910539
transform 1 0 2668 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1608910539
transform 1 0 1380 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608910539
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l5_in_0_
timestamp 1608910539
transform 1 0 1840 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1608910539
transform 1 0 2760 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1608910539
transform 1 0 1472 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1608910539
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 4324 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1608910539
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1608910539
transform 1 0 4508 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1608910539
transform 1 0 4048 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_48
timestamp 1608910539
transform 1 0 5520 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 5612 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 5336 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 5796 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_18_70
timestamp 1608910539
transform 1 0 7544 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 7636 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 7268 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 8004 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_18_93
timestamp 1608910539
transform 1 0 9660 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1608910539
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9752 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 9936 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1608910539
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1608910539
transform 1 0 10120 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_18_125
timestamp 1608910539
transform 1 0 12604 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_3_
timestamp 1608910539
transform 1 0 11776 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10948 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_18_145
timestamp 1608910539
transform 1 0 14444 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12696 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1608910539
transform 1 0 14168 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1608910539
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 14720 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 14904 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1608910539
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15272 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 17112 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 16744 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 16928 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 17296 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_203
timestamp 1608910539
transform 1 0 19780 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 19596 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19964 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1608910539
transform 1 0 18768 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_215
timestamp 1608910539
transform 1 0 20884 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_211
timestamp 1608910539
transform 1 0 20516 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1608910539
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608910539
transform -1 0 21896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1608910539
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1608910539
transform 1 0 1748 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1608910539
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608910539
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608910539
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1656 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__059__A
timestamp 1608910539
transform 1 0 2944 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1608910539
transform 1 0 2576 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1608910539
transform 1 0 2208 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 1840 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_19_38
timestamp 1608910539
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_24
timestamp 1608910539
transform 1 0 3312 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1608910539
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1608910539
transform 1 0 3128 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1608910539
transform 1 0 4784 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1608910539
transform 1 0 3772 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 4048 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_20_51
timestamp 1608910539
transform 1 0 5796 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_49
timestamp 1608910539
transform 1 0 5612 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 5704 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 5888 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 5520 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1608910539
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_2_
timestamp 1608910539
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1608910539
transform 1 0 6072 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l4_in_0_
timestamp 1608910539
transform 1 0 5888 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_19_71
timestamp 1608910539
transform 1 0 7636 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1608910539
transform 1 0 8372 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1608910539
transform 1 0 7728 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8556 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 6900 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1608910539
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1608910539
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1608910539
transform 1 0 9568 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_2_
timestamp 1608910539
transform 1 0 10672 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 10396 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1608910539
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_1_
timestamp 1608910539
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 11500 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1608910539
transform 1 0 11868 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_129
timestamp 1608910539
transform 1 0 12972 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 14352 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 14076 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1608910539
transform 1 0 13524 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1608910539
transform 1 0 14352 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l4_in_0_
timestamp 1608910539
transform 1 0 13248 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_19_159
timestamp 1608910539
transform 1 0 15732 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 14536 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 14720 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1608910539
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_3_
timestamp 1608910539
transform 1 0 16100 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1608910539
transform 1 0 14904 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1608910539
transform 1 0 16008 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1608910539
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_172
timestamp 1608910539
transform 1 0 16928 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_173
timestamp 1608910539
transform 1 0 17020 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 16836 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1608910539
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1608910539
transform 1 0 17020 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1608910539
transform 1 0 17848 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1608910539
transform 1 0 17112 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 18032 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_20_200
timestamp 1608910539
transform 1 0 19504 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_197
timestamp 1608910539
transform 1 0 19228 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_191
timestamp 1608910539
transform 1 0 18676 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 19320 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1608910539
transform 1 0 19504 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_212
timestamp 1608910539
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_213
timestamp 1608910539
transform 1 0 20700 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_209
timestamp 1608910539
transform 1 0 20332 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_218
timestamp 1608910539
transform 1 0 21160 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1608910539
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1608910539
transform 1 0 20792 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1608910539
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1608910539
transform 1 0 21436 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_222
timestamp 1608910539
transform 1 0 21528 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1608910539
transform 1 0 21252 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608910539
transform -1 0 21896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608910539
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_15
timestamp 1608910539
transform 1 0 2484 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A
timestamp 1608910539
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608910539
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1932 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 2576 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1608910539
transform 1 0 1564 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_32
timestamp 1608910539
transform 1 0 4048 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 4416 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1608910539
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1608910539
transform 1 0 5888 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1608910539
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 8464 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 8648 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1608910539
transform 1 0 7636 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1608910539
transform 1 0 10488 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1608910539
transform 1 0 8832 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1608910539
transform 1 0 9660 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_125
timestamp 1608910539
transform 1 0 12604 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1608910539
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_115
timestamp 1608910539
transform 1 0 11684 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 11500 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 11316 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1608910539
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l4_in_0_
timestamp 1608910539
transform 1 0 12696 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 13524 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_2_
timestamp 1608910539
transform 1 0 15824 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1608910539
transform 1 0 14996 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_21_176
timestamp 1608910539
transform 1 0 17296 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 17112 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 16928 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1608910539
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_2_
timestamp 1608910539
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1608910539
transform 1 0 16652 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_202
timestamp 1608910539
transform 1 0 19688 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_1_
timestamp 1608910539
transform 1 0 18860 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  Test_en_N_FTB01
timestamp 1608910539
transform 1 0 20240 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_222
timestamp 1608910539
transform 1 0 21528 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1608910539
transform 1 0 21344 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_N_FTB01_A
timestamp 1608910539
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608910539
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1608910539
transform 1 0 20792 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1608910539
transform 1 0 1380 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_7__A1
timestamp 1608910539
transform 1 0 1472 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__A0
timestamp 1608910539
transform 1 0 2576 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608910539
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_7_
timestamp 1608910539
transform 1 0 2760 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2024 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1608910539
transform 1 0 1656 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__A0
timestamp 1608910539
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1608910539
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1608910539
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1608910539
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_45
timestamp 1608910539
transform 1 0 5244 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 6532 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 6348 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__A1
timestamp 1608910539
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1608910539
transform 1 0 6716 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1608910539
transform 1 0 5520 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7544 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_22_93
timestamp 1608910539
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_90
timestamp 1608910539
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 9752 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1608910539
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1608910539
transform 1 0 10212 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1608910539
transform 1 0 9936 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 12052 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 11868 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 12236 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1608910539
transform 1 0 11040 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1608910539
transform 1 0 12512 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_22_135
timestamp 1608910539
transform 1 0 13524 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 13340 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 13616 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_22_152
timestamp 1608910539
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1608910539
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 15272 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_22_170
timestamp 1608910539
transform 1 0 16744 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 17480 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_22_203
timestamp 1608910539
transform 1 0 19780 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19872 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_3_
timestamp 1608910539
transform 1 0 18952 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1608910539
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1608910539
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608910539
transform -1 0 21896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1608910539
transform 1 0 21252 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1608910539
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__A1
timestamp 1608910539
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608910539
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_3_
timestamp 1608910539
transform 1 0 1932 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_6_
timestamp 1608910539
transform 1 0 2760 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1608910539
transform 1 0 1564 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_30
timestamp 1608910539
transform 1 0 3864 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_4_
timestamp 1608910539
transform 1 0 3956 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4784 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1608910539
transform 1 0 3588 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_58
timestamp 1608910539
transform 1 0 6440 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__A1
timestamp 1608910539
transform 1 0 6256 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1608910539
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_79
timestamp 1608910539
transform 1 0 8372 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_64
timestamp 1608910539
transform 1 0 6992 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__A0
timestamp 1608910539
transform 1 0 7084 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 8096 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_3_
timestamp 1608910539
transform 1 0 7268 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 8464 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_23_96
timestamp 1608910539
transform 1 0 9936 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1608910539
transform 1 0 10028 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_108
timestamp 1608910539
transform 1 0 11040 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 10856 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 11316 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1608910539
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_2_
timestamp 1608910539
transform 1 0 11500 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12420 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_23_142
timestamp 1608910539
transform 1 0 14168 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1608910539
transform 1 0 13892 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_163
timestamp 1608910539
transform 1 0 16100 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_148
timestamp 1608910539
transform 1 0 14720 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 15916 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 15640 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_1_
timestamp 1608910539
transform 1 0 14812 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 16284 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_181
timestamp 1608910539
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1608910539
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 18032 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_23_203
timestamp 1608910539
transform 1 0 19780 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19872 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1608910539
transform 1 0 19504 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_220
timestamp 1608910539
transform 1 0 21344 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_210
timestamp 1608910539
transform 1 0 20424 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1608910539
transform 1 0 21160 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608910539
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1608910539
transform 1 0 20792 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1608910539
transform 1 0 1380 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1608910539
transform 1 0 1472 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1608910539
transform 1 0 1656 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608910539
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1840 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 2392 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_24_32
timestamp 1608910539
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_30
timestamp 1608910539
transform 1 0 3864 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1608910539
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_5_
timestamp 1608910539
transform 1 0 4416 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1608910539
transform 1 0 6072 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 5244 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_24_82
timestamp 1608910539
transform 1 0 8648 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_78
timestamp 1608910539
transform 1 0 8280 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_75
timestamp 1608910539
transform 1 0 8004 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 8096 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8740 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1608910539
transform 1 0 6900 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1608910539
transform 1 0 7728 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1608910539
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 9660 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_24_109
timestamp 1608910539
transform 1 0 11132 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 11224 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_1_
timestamp 1608910539
transform 1 0 11408 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1608910539
transform 1 0 12236 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_3_
timestamp 1608910539
transform 1 0 13892 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1608910539
transform 1 0 13064 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_24_150
timestamp 1608910539
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 14720 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1608910539
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_3_
timestamp 1608910539
transform 1 0 16100 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1608910539
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_24_180
timestamp 1608910539
transform 1 0 17664 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_176
timestamp 1608910539
transform 1 0 17296 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 17112 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 16928 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l4_in_0_
timestamp 1608910539
transform 1 0 17756 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_24_202
timestamp 1608910539
transform 1 0 19688 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1608910539
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1608910539
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1608910539
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1608910539
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608910539
transform -1 0 21896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1608910539
transform 1 0 21252 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1608910539
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608910539
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_1_
timestamp 1608910539
transform 1 0 2852 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1608910539
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1608910539
transform 1 0 2484 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1608910539
transform 1 0 2116 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1608910539
transform 1 0 1748 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 4692 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 4876 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1608910539
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_2_
timestamp 1608910539
transform 1 0 3680 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__A0
timestamp 1608910539
transform 1 0 5060 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1608910539
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 6808 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 5244 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1608910539
transform 1 0 8280 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_25_91
timestamp 1608910539
transform 1 0 9476 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_87
timestamp 1608910539
transform 1 0 9108 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9568 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp 1608910539
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 12052 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 11868 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1608910539
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1608910539
transform 1 0 11040 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 12420 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 14076 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 13892 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 14260 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_159
timestamp 1608910539
transform 1 0 15732 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15916 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1608910539
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_180
timestamp 1608910539
transform 1 0 17664 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1608910539
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1608910539
transform 1 0 17388 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_204
timestamp 1608910539
transform 1 0 19872 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_196
timestamp 1608910539
transform 1 0 19136 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1608910539
transform 1 0 20056 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1608910539
transform 1 0 20240 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_222
timestamp 1608910539
transform 1 0 21528 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608910539
transform -1 0 21896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1608910539
transform 1 0 20424 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1608910539
transform 1 0 21160 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1608910539
transform 1 0 20792 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_3
timestamp 1608910539
transform 1 0 1380 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_3
timestamp 1608910539
transform 1 0 1380 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1608910539
transform 1 0 1656 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608910539
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608910539
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1608910539
transform 1 0 1840 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1608910539
transform 1 0 2668 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 1840 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1608910539
transform 1 0 1472 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_32
timestamp 1608910539
transform 1 0 4048 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_30
timestamp 1608910539
transform 1 0 3864 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A
timestamp 1608910539
transform 1 0 3680 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1608910539
transform 1 0 3496 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1608910539
transform 1 0 3312 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1608910539
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1608910539
transform 1 0 4140 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4140 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A0
timestamp 1608910539
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1608910539
transform 1 0 5152 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 5612 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__A0
timestamp 1608910539
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1608910539
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1608910539
transform 1 0 6440 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_62
timestamp 1608910539
transform 1 0 6808 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__A1
timestamp 1608910539
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7728 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_4_
timestamp 1608910539
transform 1 0 6900 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1608910539
transform 1 0 8740 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 7268 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_27_85
timestamp 1608910539
transform 1 0 8924 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 9476 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 9660 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 10488 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1608910539
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1608910539
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_3_
timestamp 1608910539
transform 1 0 10672 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_2_
timestamp 1608910539
transform 1 0 9844 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_121
timestamp 1608910539
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_115
timestamp 1608910539
transform 1 0 11684 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 11040 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1608910539
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12052 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1608910539
transform 1 0 11224 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 12420 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l4_in_0_
timestamp 1608910539
transform 1 0 13708 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1608910539
transform 1 0 12880 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 13892 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_26_150
timestamp 1608910539
transform 1 0 14904 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_146
timestamp 1608910539
transform 1 0 14536 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1608910539
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1608910539
transform 1 0 16192 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1608910539
transform 1 0 15364 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 15272 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1608910539
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 1608910539
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_173
timestamp 1608910539
transform 1 0 17020 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_179
timestamp 1608910539
transform 1 0 17572 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1608910539
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16744 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_27_196
timestamp 1608910539
transform 1 0 19136 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_203
timestamp 1608910539
transform 1 0 19780 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_191
timestamp 1608910539
transform 1 0 18676 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19872 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_210
timestamp 1608910539
transform 1 0 20424 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_211
timestamp 1608910539
transform 1 0 20516 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_S_FTB01_A
timestamp 1608910539
transform 1 0 20516 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1608910539
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_S_FTB01
timestamp 1608910539
transform 1 0 20700 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1608910539
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_3_S_FTB01_A
timestamp 1608910539
transform 1 0 21436 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1608910539
transform 1 0 21252 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1608910539
transform 1 0 21252 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608910539
transform -1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608910539
transform -1 0 21896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1608910539
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1608910539
transform 1 0 2300 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1748 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1608910539
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1608910539
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l5_in_0_
timestamp 1608910539
transform 1 0 4876 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1608910539
transform 1 0 3128 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1608910539
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_28_50
timestamp 1608910539
transform 1 0 5704 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 6256 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1608910539
transform 1 0 6440 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_28_70
timestamp 1608910539
transform 1 0 7544 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_67
timestamp 1608910539
transform 1 0 7268 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 7360 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A0
timestamp 1608910539
transform 1 0 7636 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 8648 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1608910539
transform 1 0 7820 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_28_93
timestamp 1608910539
transform 1 0 9660 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_84
timestamp 1608910539
transform 1 0 8832 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 9752 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1608910539
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9936 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_28_125
timestamp 1608910539
transform 1 0 12604 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 12420 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_1_
timestamp 1608910539
transform 1 0 11592 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1608910539
transform 1 0 10764 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 13340 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 13524 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1608910539
transform 1 0 13708 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_28_150
timestamp 1608910539
transform 1 0 14904 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_146
timestamp 1608910539
transform 1 0 14536 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1608910539
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 16100 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1608910539
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_28_181
timestamp 1608910539
transform 1 0 17756 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_169
timestamp 1608910539
transform 1 0 16652 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_201
timestamp 1608910539
transform 1 0 19596 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_193
timestamp 1608910539
transform 1 0 18860 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1608910539
transform 1 0 19688 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_S_FTB01
timestamp 1608910539
transform 1 0 20240 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1608910539
transform 1 0 19872 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_2_S_FTB01_A
timestamp 1608910539
transform 1 0 21436 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1608910539
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1608910539
transform -1 0 21896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  clk_2_S_FTB01
timestamp 1608910539
transform 1 0 20884 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1608910539
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1608910539
transform 1 0 2852 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1608910539
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1608910539
transform 1 0 2484 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1608910539
transform 1 0 2116 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1608910539
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 4876 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 4692 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1608910539
transform 1 0 3036 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1608910539
transform 1 0 3864 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_29_51
timestamp 1608910539
transform 1 0 5796 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_45
timestamp 1608910539
transform 1 0 5244 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 5060 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1608910539
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1608910539
transform 1 0 5888 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1608910539
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_79
timestamp 1608910539
transform 1 0 8372 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_65
timestamp 1608910539
transform 1 0 7084 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8188 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1608910539
transform 1 0 7360 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 8648 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 10120 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_29_121
timestamp 1608910539
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_117
timestamp 1608910539
transform 1 0 11868 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1608910539
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12420 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1608910539
transform 1 0 11592 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_145
timestamp 1608910539
transform 1 0 14444 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 13892 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_165
timestamp 1608910539
transform 1 0 16284 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_157
timestamp 1608910539
transform 1 0 15548 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_184
timestamp 1608910539
transform 1 0 18032 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1608910539
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1608910539
transform 1 0 18308 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1608910539
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _132_
timestamp 1608910539
transform 1 0 16468 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_206
timestamp 1608910539
transform 1 0 20056 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_197
timestamp 1608910539
transform 1 0 19228 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_193
timestamp 1608910539
transform 1 0 18860 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_E_FTB01_A
timestamp 1608910539
transform 1 0 20148 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_W_FTB01_A
timestamp 1608910539
transform 1 0 19872 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1608910539
transform 1 0 19320 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1608910539
transform 1 0 19504 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1608910539
transform 1 0 18492 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_3_S_FTB01_A
timestamp 1608910539
transform 1 0 20332 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1608910539
transform 1 0 20516 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1608910539
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  clk_3_S_FTB01
timestamp 1608910539
transform 1 0 20700 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1608910539
transform 1 0 21252 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_13
timestamp 1608910539
transform 1 0 2300 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1608910539
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 2668 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1608910539
transform 1 0 2116 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1608910539
transform 1 0 2852 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1608910539
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1608910539
transform 1 0 1748 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_32
timestamp 1608910539
transform 1 0 4048 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_23
timestamp 1608910539
transform 1 0 3220 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 3036 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 4140 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1608910539
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1608910539
transform 1 0 4324 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_30_44
timestamp 1608910539
transform 1 0 5152 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 5244 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1608910539
transform 1 0 5428 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1608910539
transform 1 0 6256 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_30_65
timestamp 1608910539
transform 1 0 7084 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8004 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1608910539
transform 1 0 7176 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8188 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_30_93
timestamp 1608910539
transform 1 0 9660 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_86
timestamp 1608910539
transform 1 0 9016 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1608910539
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1608910539
transform 1 0 9752 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 10580 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_30_119
timestamp 1608910539
transform 1 0 12052 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_142
timestamp 1608910539
transform 1 0 14168 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_137
timestamp 1608910539
transform 1 0 13708 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_133
timestamp 1608910539
transform 1 0 13340 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_129
timestamp 1608910539
transform 1 0 12972 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A
timestamp 1608910539
transform 1 0 14352 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1608910539
transform 1 0 13984 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1608910539
transform 1 0 13524 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A
timestamp 1608910539
transform 1 0 13156 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1608910539
transform 1 0 12788 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_165
timestamp 1608910539
transform 1 0 16284 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_160
timestamp 1608910539
transform 1 0 15824 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_154
timestamp 1608910539
transform 1 0 15272 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_152
timestamp 1608910539
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_146
timestamp 1608910539
transform 1 0 14536 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_1_W_FTB01_A
timestamp 1608910539
transform 1 0 16100 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__A
timestamp 1608910539
transform 1 0 15916 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1608910539
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_174
timestamp 1608910539
transform 1 0 17112 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_171
timestamp 1608910539
transform 1 0 16836 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_3_W_FTB01_A
timestamp 1608910539
transform 1 0 17848 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__A
timestamp 1608910539
transform 1 0 16928 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_W_FTB01
timestamp 1608910539
transform 1 0 18032 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_207
timestamp 1608910539
transform 1 0 20148 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_204
timestamp 1608910539
transform 1 0 19872 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_3_E_FTB01_A
timestamp 1608910539
transform 1 0 19964 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_3_W_FTB01_A
timestamp 1608910539
transform 1 0 19688 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_W_FTB01
timestamp 1608910539
transform 1 0 19136 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_E_FTB01
timestamp 1608910539
transform 1 0 20240 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_3_W_FTB01
timestamp 1608910539
transform 1 0 18584 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_3_N_FTB01_A
timestamp 1608910539
transform 1 0 21436 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1608910539
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1608910539
transform -1 0 21896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  clk_3_N_FTB01
timestamp 1608910539
transform 1 0 20884 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_13
timestamp 1608910539
transform 1 0 2300 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1608910539
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1608910539
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1608910539
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1608910539
transform 1 0 1748 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_21
timestamp 1608910539
transform 1 0 3036 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 3220 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 3772 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_31_62
timestamp 1608910539
transform 1 0 6808 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1608910539
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 5244 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8372 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 6900 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_31_100
timestamp 1608910539
transform 1 0 10304 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 9752 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1608910539
transform 1 0 10396 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 9200 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_121
timestamp 1608910539
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 12052 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1608910539
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 12420 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l4_in_0_
timestamp 1608910539
transform 1 0 11224 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_31_141
timestamp 1608910539
transform 1 0 14076 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1608910539
transform 1 0 14168 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1608910539
transform 1 0 13708 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1608910539
transform 1 0 13340 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1608910539
transform 1 0 12972 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_156
timestamp 1608910539
transform 1 0 15456 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__A
timestamp 1608910539
transform 1 0 15272 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  prog_clk_1_W_FTB01
timestamp 1608910539
transform 1 0 15548 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _130_
timestamp 1608910539
transform 1 0 16100 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _127_
timestamp 1608910539
transform 1 0 14904 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _126_
timestamp 1608910539
transform 1 0 14536 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_178
timestamp 1608910539
transform 1 0 17480 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_173
timestamp 1608910539
transform 1 0 17020 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A
timestamp 1608910539
transform 1 0 18032 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__A
timestamp 1608910539
transform 1 0 16836 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1608910539
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  clk_1_W_FTB01
timestamp 1608910539
transform 1 0 18216 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _134_
timestamp 1608910539
transform 1 0 17572 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _133_
timestamp 1608910539
transform 1 0 17112 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _131_
timestamp 1608910539
transform 1 0 16468 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_192
timestamp 1608910539
transform 1 0 18768 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_1_W_FTB01_A
timestamp 1608910539
transform 1 0 19964 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 18860 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  clk_3_E_FTB01
timestamp 1608910539
transform 1 0 20148 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1608910539
transform 1 0 21436 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_2_E_FTB01_A
timestamp 1608910539
transform 1 0 21252 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1608910539
transform -1 0 21896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  clk_2_E_FTB01
timestamp 1608910539
transform 1 0 20700 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1608910539
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1608910539
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1608910539
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1608910539
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1608910539
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4048 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_32_48
timestamp 1608910539
transform 1 0 5520 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 5796 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 7268 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 7452 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8648 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8464 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1608910539
transform 1 0 7636 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_32_98
timestamp 1608910539
transform 1 0 10120 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_93
timestamp 1608910539
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_84
timestamp 1608910539
transform 1 0 8832 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1608910539
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 10304 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1608910539
transform 1 0 9752 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_122
timestamp 1608910539
transform 1 0 12328 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_110
timestamp 1608910539
transform 1 0 11224 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1608910539
transform 1 0 12144 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1608910539
transform 1 0 11408 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1608910539
transform 1 0 11776 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1608910539
transform 1 0 10856 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_134
timestamp 1608910539
transform 1 0 13432 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1608910539
transform 1 0 13064 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_160
timestamp 1608910539
transform 1 0 15824 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_150
timestamp 1608910539
transform 1 0 14904 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A
timestamp 1608910539
transform 1 0 15640 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1608910539
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _129_
timestamp 1608910539
transform 1 0 15272 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _128_
timestamp 1608910539
transform 1 0 14536 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_186
timestamp 1608910539
transform 1 0 18216 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_178
timestamp 1608910539
transform 1 0 17480 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1608910539
transform 1 0 16928 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _135_
timestamp 1608910539
transform 1 0 17112 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_201
timestamp 1608910539
transform 1 0 19596 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_194
timestamp 1608910539
transform 1 0 18952 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_E_FTB01
timestamp 1608910539
transform 1 0 19688 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_1_E_FTB01
timestamp 1608910539
transform 1 0 20240 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_2_W_FTB01
timestamp 1608910539
transform 1 0 18400 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_1_E_FTB01
timestamp 1608910539
transform 1 0 19044 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_2_N_FTB01_A
timestamp 1608910539
transform 1 0 21436 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1608910539
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1608910539
transform -1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  clk_2_N_FTB01
timestamp 1608910539
transform 1 0 20884 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1608910539
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1608910539
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1608910539
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_32
timestamp 1608910539
transform 1 0 4048 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_27
timestamp 1608910539
transform 1 0 3588 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1608910539
transform 1 0 3956 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1608910539
transform 1 0 4600 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_54
timestamp 1608910539
transform 1 0 6072 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_42
timestamp 1608910539
transform 1 0 4968 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1608910539
transform 1 0 6808 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_72
timestamp 1608910539
transform 1 0 7728 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1608910539
transform 1 0 6900 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_33_94
timestamp 1608910539
transform 1 0 9752 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_92
timestamp 1608910539
transform 1 0 9568 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_84
timestamp 1608910539
transform 1 0 8832 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1608910539
transform 1 0 9660 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1608910539
transform 1 0 12604 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_118
timestamp 1608910539
transform 1 0 11960 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_106
timestamp 1608910539
transform 1 0 10856 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1608910539
transform 1 0 12512 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_137
timestamp 1608910539
transform 1 0 13708 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_156
timestamp 1608910539
transform 1 0 15456 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_149
timestamp 1608910539
transform 1 0 14812 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1608910539
transform 1 0 15364 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_187
timestamp 1608910539
transform 1 0 18308 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_180
timestamp 1608910539
transform 1 0 17664 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_168
timestamp 1608910539
transform 1 0 16560 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1608910539
transform 1 0 18216 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_197
timestamp 1608910539
transform 1 0 19228 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_3_E_FTB01_A
timestamp 1608910539
transform 1 0 19596 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_3_N_FTB01_A
timestamp 1608910539
transform 1 0 19780 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_2_W_FTB01_A
timestamp 1608910539
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_1_E_FTB01_A
timestamp 1608910539
transform 1 0 18860 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_N_FTB01
timestamp 1608910539
transform 1 0 19964 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_222
timestamp 1608910539
transform 1 0 21528 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_N_FTB01_A
timestamp 1608910539
transform 1 0 21344 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_1_E_FTB01_A
timestamp 1608910539
transform 1 0 21160 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1608910539
transform 1 0 21068 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1608910539
transform -1 0 21896 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_N_FTB01
timestamp 1608910539
transform 1 0 20516 0 1 20128
box -38 -48 590 592
<< labels >>
rlabel metal2 s 18602 22200 18658 23000 6 Test_en_N_out
port 0 nsew signal tristate
rlabel metal2 s 21086 0 21142 800 6 Test_en_S_in
port 1 nsew signal input
rlabel metal2 s 202 0 258 800 6 bottom_left_grid_pin_42_
port 2 nsew signal input
rlabel metal2 s 570 0 626 800 6 bottom_left_grid_pin_43_
port 3 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 bottom_left_grid_pin_44_
port 4 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 bottom_left_grid_pin_45_
port 5 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 bottom_left_grid_pin_46_
port 6 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 bottom_left_grid_pin_47_
port 7 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 bottom_left_grid_pin_48_
port 8 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 bottom_left_grid_pin_49_
port 9 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 ccff_head
port 10 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 ccff_tail
port 11 nsew signal tristate
rlabel metal3 s 0 3544 800 3664 6 chanx_left_in[0]
port 12 nsew signal input
rlabel metal3 s 0 7760 800 7880 6 chanx_left_in[10]
port 13 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 chanx_left_in[11]
port 14 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 chanx_left_in[12]
port 15 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[13]
port 16 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[14]
port 17 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 chanx_left_in[15]
port 18 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[16]
port 19 nsew signal input
rlabel metal3 s 0 10752 800 10872 6 chanx_left_in[17]
port 20 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 chanx_left_in[18]
port 21 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 chanx_left_in[19]
port 22 nsew signal input
rlabel metal3 s 0 3952 800 4072 6 chanx_left_in[1]
port 23 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 chanx_left_in[2]
port 24 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 chanx_left_in[3]
port 25 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 chanx_left_in[4]
port 26 nsew signal input
rlabel metal3 s 0 5584 800 5704 6 chanx_left_in[5]
port 27 nsew signal input
rlabel metal3 s 0 5992 800 6112 6 chanx_left_in[6]
port 28 nsew signal input
rlabel metal3 s 0 6400 800 6520 6 chanx_left_in[7]
port 29 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 chanx_left_in[8]
port 30 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 chanx_left_in[9]
port 31 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 chanx_left_out[0]
port 32 nsew signal tristate
rlabel metal3 s 0 16192 800 16312 6 chanx_left_out[10]
port 33 nsew signal tristate
rlabel metal3 s 0 16736 800 16856 6 chanx_left_out[11]
port 34 nsew signal tristate
rlabel metal3 s 0 17144 800 17264 6 chanx_left_out[12]
port 35 nsew signal tristate
rlabel metal3 s 0 17552 800 17672 6 chanx_left_out[13]
port 36 nsew signal tristate
rlabel metal3 s 0 17960 800 18080 6 chanx_left_out[14]
port 37 nsew signal tristate
rlabel metal3 s 0 18368 800 18488 6 chanx_left_out[15]
port 38 nsew signal tristate
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[16]
port 39 nsew signal tristate
rlabel metal3 s 0 19184 800 19304 6 chanx_left_out[17]
port 40 nsew signal tristate
rlabel metal3 s 0 19592 800 19712 6 chanx_left_out[18]
port 41 nsew signal tristate
rlabel metal3 s 0 20136 800 20256 6 chanx_left_out[19]
port 42 nsew signal tristate
rlabel metal3 s 0 12384 800 12504 6 chanx_left_out[1]
port 43 nsew signal tristate
rlabel metal3 s 0 12792 800 12912 6 chanx_left_out[2]
port 44 nsew signal tristate
rlabel metal3 s 0 13336 800 13456 6 chanx_left_out[3]
port 45 nsew signal tristate
rlabel metal3 s 0 13744 800 13864 6 chanx_left_out[4]
port 46 nsew signal tristate
rlabel metal3 s 0 14152 800 14272 6 chanx_left_out[5]
port 47 nsew signal tristate
rlabel metal3 s 0 14560 800 14680 6 chanx_left_out[6]
port 48 nsew signal tristate
rlabel metal3 s 0 14968 800 15088 6 chanx_left_out[7]
port 49 nsew signal tristate
rlabel metal3 s 0 15376 800 15496 6 chanx_left_out[8]
port 50 nsew signal tristate
rlabel metal3 s 0 15784 800 15904 6 chanx_left_out[9]
port 51 nsew signal tristate
rlabel metal3 s 22200 3544 23000 3664 6 chanx_right_in[0]
port 52 nsew signal input
rlabel metal3 s 22200 7760 23000 7880 6 chanx_right_in[10]
port 53 nsew signal input
rlabel metal3 s 22200 8168 23000 8288 6 chanx_right_in[11]
port 54 nsew signal input
rlabel metal3 s 22200 8576 23000 8696 6 chanx_right_in[12]
port 55 nsew signal input
rlabel metal3 s 22200 8984 23000 9104 6 chanx_right_in[13]
port 56 nsew signal input
rlabel metal3 s 22200 9392 23000 9512 6 chanx_right_in[14]
port 57 nsew signal input
rlabel metal3 s 22200 9800 23000 9920 6 chanx_right_in[15]
port 58 nsew signal input
rlabel metal3 s 22200 10344 23000 10464 6 chanx_right_in[16]
port 59 nsew signal input
rlabel metal3 s 22200 10752 23000 10872 6 chanx_right_in[17]
port 60 nsew signal input
rlabel metal3 s 22200 11160 23000 11280 6 chanx_right_in[18]
port 61 nsew signal input
rlabel metal3 s 22200 11568 23000 11688 6 chanx_right_in[19]
port 62 nsew signal input
rlabel metal3 s 22200 3952 23000 4072 6 chanx_right_in[1]
port 63 nsew signal input
rlabel metal3 s 22200 4360 23000 4480 6 chanx_right_in[2]
port 64 nsew signal input
rlabel metal3 s 22200 4768 23000 4888 6 chanx_right_in[3]
port 65 nsew signal input
rlabel metal3 s 22200 5176 23000 5296 6 chanx_right_in[4]
port 66 nsew signal input
rlabel metal3 s 22200 5584 23000 5704 6 chanx_right_in[5]
port 67 nsew signal input
rlabel metal3 s 22200 5992 23000 6112 6 chanx_right_in[6]
port 68 nsew signal input
rlabel metal3 s 22200 6400 23000 6520 6 chanx_right_in[7]
port 69 nsew signal input
rlabel metal3 s 22200 6944 23000 7064 6 chanx_right_in[8]
port 70 nsew signal input
rlabel metal3 s 22200 7352 23000 7472 6 chanx_right_in[9]
port 71 nsew signal input
rlabel metal3 s 22200 11976 23000 12096 6 chanx_right_out[0]
port 72 nsew signal tristate
rlabel metal3 s 22200 16192 23000 16312 6 chanx_right_out[10]
port 73 nsew signal tristate
rlabel metal3 s 22200 16736 23000 16856 6 chanx_right_out[11]
port 74 nsew signal tristate
rlabel metal3 s 22200 17144 23000 17264 6 chanx_right_out[12]
port 75 nsew signal tristate
rlabel metal3 s 22200 17552 23000 17672 6 chanx_right_out[13]
port 76 nsew signal tristate
rlabel metal3 s 22200 17960 23000 18080 6 chanx_right_out[14]
port 77 nsew signal tristate
rlabel metal3 s 22200 18368 23000 18488 6 chanx_right_out[15]
port 78 nsew signal tristate
rlabel metal3 s 22200 18776 23000 18896 6 chanx_right_out[16]
port 79 nsew signal tristate
rlabel metal3 s 22200 19184 23000 19304 6 chanx_right_out[17]
port 80 nsew signal tristate
rlabel metal3 s 22200 19592 23000 19712 6 chanx_right_out[18]
port 81 nsew signal tristate
rlabel metal3 s 22200 20136 23000 20256 6 chanx_right_out[19]
port 82 nsew signal tristate
rlabel metal3 s 22200 12384 23000 12504 6 chanx_right_out[1]
port 83 nsew signal tristate
rlabel metal3 s 22200 12792 23000 12912 6 chanx_right_out[2]
port 84 nsew signal tristate
rlabel metal3 s 22200 13336 23000 13456 6 chanx_right_out[3]
port 85 nsew signal tristate
rlabel metal3 s 22200 13744 23000 13864 6 chanx_right_out[4]
port 86 nsew signal tristate
rlabel metal3 s 22200 14152 23000 14272 6 chanx_right_out[5]
port 87 nsew signal tristate
rlabel metal3 s 22200 14560 23000 14680 6 chanx_right_out[6]
port 88 nsew signal tristate
rlabel metal3 s 22200 14968 23000 15088 6 chanx_right_out[7]
port 89 nsew signal tristate
rlabel metal3 s 22200 15376 23000 15496 6 chanx_right_out[8]
port 90 nsew signal tristate
rlabel metal3 s 22200 15784 23000 15904 6 chanx_right_out[9]
port 91 nsew signal tristate
rlabel metal2 s 4342 0 4398 800 6 chany_bottom_in[0]
port 92 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 chany_bottom_in[10]
port 93 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 chany_bottom_in[11]
port 94 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 chany_bottom_in[12]
port 95 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 chany_bottom_in[13]
port 96 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 chany_bottom_in[14]
port 97 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 chany_bottom_in[15]
port 98 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 chany_bottom_in[16]
port 99 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 chany_bottom_in[17]
port 100 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 chany_bottom_in[18]
port 101 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 chany_bottom_in[19]
port 102 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 chany_bottom_in[1]
port 103 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 chany_bottom_in[2]
port 104 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 chany_bottom_in[3]
port 105 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 chany_bottom_in[4]
port 106 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 chany_bottom_in[5]
port 107 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 chany_bottom_in[6]
port 108 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 chany_bottom_in[7]
port 109 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 chany_bottom_in[8]
port 110 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 chany_bottom_in[9]
port 111 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 chany_bottom_out[0]
port 112 nsew signal tristate
rlabel metal2 s 16854 0 16910 800 6 chany_bottom_out[10]
port 113 nsew signal tristate
rlabel metal2 s 17314 0 17370 800 6 chany_bottom_out[11]
port 114 nsew signal tristate
rlabel metal2 s 17682 0 17738 800 6 chany_bottom_out[12]
port 115 nsew signal tristate
rlabel metal2 s 18142 0 18198 800 6 chany_bottom_out[13]
port 116 nsew signal tristate
rlabel metal2 s 18602 0 18658 800 6 chany_bottom_out[14]
port 117 nsew signal tristate
rlabel metal2 s 18970 0 19026 800 6 chany_bottom_out[15]
port 118 nsew signal tristate
rlabel metal2 s 19430 0 19486 800 6 chany_bottom_out[16]
port 119 nsew signal tristate
rlabel metal2 s 19798 0 19854 800 6 chany_bottom_out[17]
port 120 nsew signal tristate
rlabel metal2 s 20258 0 20314 800 6 chany_bottom_out[18]
port 121 nsew signal tristate
rlabel metal2 s 20626 0 20682 800 6 chany_bottom_out[19]
port 122 nsew signal tristate
rlabel metal2 s 13082 0 13138 800 6 chany_bottom_out[1]
port 123 nsew signal tristate
rlabel metal2 s 13542 0 13598 800 6 chany_bottom_out[2]
port 124 nsew signal tristate
rlabel metal2 s 14002 0 14058 800 6 chany_bottom_out[3]
port 125 nsew signal tristate
rlabel metal2 s 14370 0 14426 800 6 chany_bottom_out[4]
port 126 nsew signal tristate
rlabel metal2 s 14830 0 14886 800 6 chany_bottom_out[5]
port 127 nsew signal tristate
rlabel metal2 s 15198 0 15254 800 6 chany_bottom_out[6]
port 128 nsew signal tristate
rlabel metal2 s 15658 0 15714 800 6 chany_bottom_out[7]
port 129 nsew signal tristate
rlabel metal2 s 16026 0 16082 800 6 chany_bottom_out[8]
port 130 nsew signal tristate
rlabel metal2 s 16486 0 16542 800 6 chany_bottom_out[9]
port 131 nsew signal tristate
rlabel metal2 s 3238 22200 3294 23000 6 chany_top_in[0]
port 132 nsew signal input
rlabel metal2 s 7102 22200 7158 23000 6 chany_top_in[10]
port 133 nsew signal input
rlabel metal2 s 7470 22200 7526 23000 6 chany_top_in[11]
port 134 nsew signal input
rlabel metal2 s 7838 22200 7894 23000 6 chany_top_in[12]
port 135 nsew signal input
rlabel metal2 s 8206 22200 8262 23000 6 chany_top_in[13]
port 136 nsew signal input
rlabel metal2 s 8574 22200 8630 23000 6 chany_top_in[14]
port 137 nsew signal input
rlabel metal2 s 8942 22200 8998 23000 6 chany_top_in[15]
port 138 nsew signal input
rlabel metal2 s 9402 22200 9458 23000 6 chany_top_in[16]
port 139 nsew signal input
rlabel metal2 s 9770 22200 9826 23000 6 chany_top_in[17]
port 140 nsew signal input
rlabel metal2 s 10138 22200 10194 23000 6 chany_top_in[18]
port 141 nsew signal input
rlabel metal2 s 10506 22200 10562 23000 6 chany_top_in[19]
port 142 nsew signal input
rlabel metal2 s 3606 22200 3662 23000 6 chany_top_in[1]
port 143 nsew signal input
rlabel metal2 s 3974 22200 4030 23000 6 chany_top_in[2]
port 144 nsew signal input
rlabel metal2 s 4342 22200 4398 23000 6 chany_top_in[3]
port 145 nsew signal input
rlabel metal2 s 4802 22200 4858 23000 6 chany_top_in[4]
port 146 nsew signal input
rlabel metal2 s 5170 22200 5226 23000 6 chany_top_in[5]
port 147 nsew signal input
rlabel metal2 s 5538 22200 5594 23000 6 chany_top_in[6]
port 148 nsew signal input
rlabel metal2 s 5906 22200 5962 23000 6 chany_top_in[7]
port 149 nsew signal input
rlabel metal2 s 6274 22200 6330 23000 6 chany_top_in[8]
port 150 nsew signal input
rlabel metal2 s 6642 22200 6698 23000 6 chany_top_in[9]
port 151 nsew signal input
rlabel metal2 s 10874 22200 10930 23000 6 chany_top_out[0]
port 152 nsew signal tristate
rlabel metal2 s 14738 22200 14794 23000 6 chany_top_out[10]
port 153 nsew signal tristate
rlabel metal2 s 15106 22200 15162 23000 6 chany_top_out[11]
port 154 nsew signal tristate
rlabel metal2 s 15474 22200 15530 23000 6 chany_top_out[12]
port 155 nsew signal tristate
rlabel metal2 s 15842 22200 15898 23000 6 chany_top_out[13]
port 156 nsew signal tristate
rlabel metal2 s 16302 22200 16358 23000 6 chany_top_out[14]
port 157 nsew signal tristate
rlabel metal2 s 16670 22200 16726 23000 6 chany_top_out[15]
port 158 nsew signal tristate
rlabel metal2 s 17038 22200 17094 23000 6 chany_top_out[16]
port 159 nsew signal tristate
rlabel metal2 s 17406 22200 17462 23000 6 chany_top_out[17]
port 160 nsew signal tristate
rlabel metal2 s 17774 22200 17830 23000 6 chany_top_out[18]
port 161 nsew signal tristate
rlabel metal2 s 18142 22200 18198 23000 6 chany_top_out[19]
port 162 nsew signal tristate
rlabel metal2 s 11242 22200 11298 23000 6 chany_top_out[1]
port 163 nsew signal tristate
rlabel metal2 s 11702 22200 11758 23000 6 chany_top_out[2]
port 164 nsew signal tristate
rlabel metal2 s 12070 22200 12126 23000 6 chany_top_out[3]
port 165 nsew signal tristate
rlabel metal2 s 12438 22200 12494 23000 6 chany_top_out[4]
port 166 nsew signal tristate
rlabel metal2 s 12806 22200 12862 23000 6 chany_top_out[5]
port 167 nsew signal tristate
rlabel metal2 s 13174 22200 13230 23000 6 chany_top_out[6]
port 168 nsew signal tristate
rlabel metal2 s 13542 22200 13598 23000 6 chany_top_out[7]
port 169 nsew signal tristate
rlabel metal2 s 14002 22200 14058 23000 6 chany_top_out[8]
port 170 nsew signal tristate
rlabel metal2 s 14370 22200 14426 23000 6 chany_top_out[9]
port 171 nsew signal tristate
rlabel metal3 s 22200 20544 23000 20664 6 clk_1_E_out
port 172 nsew signal tristate
rlabel metal2 s 18970 22200 19026 23000 6 clk_1_N_in
port 173 nsew signal input
rlabel metal3 s 0 20544 800 20664 6 clk_1_W_out
port 174 nsew signal tristate
rlabel metal3 s 22200 20952 23000 21072 6 clk_2_E_out
port 175 nsew signal tristate
rlabel metal2 s 19338 22200 19394 23000 6 clk_2_N_in
port 176 nsew signal input
rlabel metal2 s 21638 22200 21694 23000 6 clk_2_N_out
port 177 nsew signal tristate
rlabel metal2 s 21454 0 21510 800 6 clk_2_S_out
port 178 nsew signal tristate
rlabel metal3 s 0 20952 800 21072 6 clk_2_W_out
port 179 nsew signal tristate
rlabel metal3 s 22200 21360 23000 21480 6 clk_3_E_out
port 180 nsew signal tristate
rlabel metal2 s 19706 22200 19762 23000 6 clk_3_N_in
port 181 nsew signal input
rlabel metal2 s 22006 22200 22062 23000 6 clk_3_N_out
port 182 nsew signal tristate
rlabel metal2 s 21914 0 21970 800 6 clk_3_S_out
port 183 nsew signal tristate
rlabel metal3 s 0 21360 800 21480 6 clk_3_W_out
port 184 nsew signal tristate
rlabel metal3 s 0 144 800 264 6 left_bottom_grid_pin_34_
port 185 nsew signal input
rlabel metal3 s 0 552 800 672 6 left_bottom_grid_pin_35_
port 186 nsew signal input
rlabel metal3 s 0 960 800 1080 6 left_bottom_grid_pin_36_
port 187 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 left_bottom_grid_pin_37_
port 188 nsew signal input
rlabel metal3 s 0 1776 800 1896 6 left_bottom_grid_pin_38_
port 189 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 left_bottom_grid_pin_39_
port 190 nsew signal input
rlabel metal3 s 0 2592 800 2712 6 left_bottom_grid_pin_40_
port 191 nsew signal input
rlabel metal3 s 0 3000 800 3120 6 left_bottom_grid_pin_41_
port 192 nsew signal input
rlabel metal2 s 20074 22200 20130 23000 6 prog_clk_0_N_in
port 193 nsew signal input
rlabel metal3 s 22200 21768 23000 21888 6 prog_clk_1_E_out
port 194 nsew signal tristate
rlabel metal2 s 20442 22200 20498 23000 6 prog_clk_1_N_in
port 195 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 prog_clk_1_W_out
port 196 nsew signal tristate
rlabel metal3 s 22200 22176 23000 22296 6 prog_clk_2_E_out
port 197 nsew signal tristate
rlabel metal2 s 20902 22200 20958 23000 6 prog_clk_2_N_in
port 198 nsew signal input
rlabel metal2 s 22374 22200 22430 23000 6 prog_clk_2_N_out
port 199 nsew signal tristate
rlabel metal2 s 22282 0 22338 800 6 prog_clk_2_S_out
port 200 nsew signal tristate
rlabel metal3 s 0 22176 800 22296 6 prog_clk_2_W_out
port 201 nsew signal tristate
rlabel metal3 s 22200 22584 23000 22704 6 prog_clk_3_E_out
port 202 nsew signal tristate
rlabel metal2 s 21270 22200 21326 23000 6 prog_clk_3_N_in
port 203 nsew signal input
rlabel metal2 s 22742 22200 22798 23000 6 prog_clk_3_N_out
port 204 nsew signal tristate
rlabel metal2 s 22742 0 22798 800 6 prog_clk_3_S_out
port 205 nsew signal tristate
rlabel metal3 s 0 22584 800 22704 6 prog_clk_3_W_out
port 206 nsew signal tristate
rlabel metal3 s 22200 144 23000 264 6 right_bottom_grid_pin_34_
port 207 nsew signal input
rlabel metal3 s 22200 552 23000 672 6 right_bottom_grid_pin_35_
port 208 nsew signal input
rlabel metal3 s 22200 960 23000 1080 6 right_bottom_grid_pin_36_
port 209 nsew signal input
rlabel metal3 s 22200 1368 23000 1488 6 right_bottom_grid_pin_37_
port 210 nsew signal input
rlabel metal3 s 22200 1776 23000 1896 6 right_bottom_grid_pin_38_
port 211 nsew signal input
rlabel metal3 s 22200 2184 23000 2304 6 right_bottom_grid_pin_39_
port 212 nsew signal input
rlabel metal3 s 22200 2592 23000 2712 6 right_bottom_grid_pin_40_
port 213 nsew signal input
rlabel metal3 s 22200 3000 23000 3120 6 right_bottom_grid_pin_41_
port 214 nsew signal input
rlabel metal2 s 202 22200 258 23000 6 top_left_grid_pin_42_
port 215 nsew signal input
rlabel metal2 s 570 22200 626 23000 6 top_left_grid_pin_43_
port 216 nsew signal input
rlabel metal2 s 938 22200 994 23000 6 top_left_grid_pin_44_
port 217 nsew signal input
rlabel metal2 s 1306 22200 1362 23000 6 top_left_grid_pin_45_
port 218 nsew signal input
rlabel metal2 s 1674 22200 1730 23000 6 top_left_grid_pin_46_
port 219 nsew signal input
rlabel metal2 s 2042 22200 2098 23000 6 top_left_grid_pin_47_
port 220 nsew signal input
rlabel metal2 s 2502 22200 2558 23000 6 top_left_grid_pin_48_
port 221 nsew signal input
rlabel metal2 s 2870 22200 2926 23000 6 top_left_grid_pin_49_
port 222 nsew signal input
rlabel metal4 s 18271 2128 18591 20720 6 VPWR
port 223 nsew power bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VPWR
port 224 nsew power bidirectional
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 225 nsew power bidirectional
rlabel metal4 s 14805 2128 15125 20720 6 VGND
port 226 nsew ground bidirectional
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 227 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
