VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_io_right
  CLASS BLOCK ;
  FOREIGN grid_io_right ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 2.400 8.800 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 2.400 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 4.800 140.000 5.400 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 2.400 25.800 ;
    END
  END address[3]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 2.400 ;
    END
  END enable
  PIN gfpga_pad_GPIO_PAD[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 15.000 140.000 15.600 ;
    END
  END gfpga_pad_GPIO_PAD[0]
  PIN gfpga_pad_GPIO_PAD[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 137.600 23.370 140.000 ;
    END
  END gfpga_pad_GPIO_PAD[1]
  PIN gfpga_pad_GPIO_PAD[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 25.880 140.000 26.480 ;
    END
  END gfpga_pad_GPIO_PAD[2]
  PIN gfpga_pad_GPIO_PAD[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 2.400 43.480 ;
    END
  END gfpga_pad_GPIO_PAD[3]
  PIN gfpga_pad_GPIO_PAD[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 36.760 140.000 37.360 ;
    END
  END gfpga_pad_GPIO_PAD[4]
  PIN gfpga_pad_GPIO_PAD[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 47.640 140.000 48.240 ;
    END
  END gfpga_pad_GPIO_PAD[5]
  PIN gfpga_pad_GPIO_PAD[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 58.520 140.000 59.120 ;
    END
  END gfpga_pad_GPIO_PAD[6]
  PIN gfpga_pad_GPIO_PAD[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 2.400 ;
    END
  END gfpga_pad_GPIO_PAD[7]
  PIN left_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 2.400 ;
    END
  END left_width_0_height_0__pin_0_
  PIN left_width_0_height_0__pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 2.400 ;
    END
  END left_width_0_height_0__pin_10_
  PIN left_width_0_height_0__pin_11_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 2.400 131.200 ;
    END
  END left_width_0_height_0__pin_11_
  PIN left_width_0_height_0__pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 123.120 140.000 123.720 ;
    END
  END left_width_0_height_0__pin_12_
  PIN left_width_0_height_0__pin_13_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 134.000 140.000 134.600 ;
    END
  END left_width_0_height_0__pin_13_
  PIN left_width_0_height_0__pin_14_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 137.600 69.830 140.000 ;
    END
  END left_width_0_height_0__pin_14_
  PIN left_width_0_height_0__pin_15_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.010 137.600 116.290 140.000 ;
    END
  END left_width_0_height_0__pin_15_
  PIN left_width_0_height_0__pin_1_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 69.400 140.000 70.000 ;
    END
  END left_width_0_height_0__pin_1_
  PIN left_width_0_height_0__pin_2_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 2.400 61.160 ;
    END
  END left_width_0_height_0__pin_2_
  PIN left_width_0_height_0__pin_3_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 2.400 78.840 ;
    END
  END left_width_0_height_0__pin_3_
  PIN left_width_0_height_0__pin_4_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 2.400 95.840 ;
    END
  END left_width_0_height_0__pin_4_
  PIN left_width_0_height_0__pin_5_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 2.400 113.520 ;
    END
  END left_width_0_height_0__pin_5_
  PIN left_width_0_height_0__pin_6_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 79.600 140.000 80.200 ;
    END
  END left_width_0_height_0__pin_6_
  PIN left_width_0_height_0__pin_7_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 90.480 140.000 91.080 ;
    END
  END left_width_0_height_0__pin_7_
  PIN left_width_0_height_0__pin_8_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 101.360 140.000 101.960 ;
    END
  END left_width_0_height_0__pin_8_
  PIN left_width_0_height_0__pin_9_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 112.240 140.000 112.840 ;
    END
  END left_width_0_height_0__pin_9_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 0.530 10.640 134.320 128.080 ;
      LAYER met2 ;
        RECT 0.550 2.680 138.370 128.080 ;
        RECT 0.550 0.155 11.310 2.680 ;
        RECT 12.150 0.155 34.310 2.680 ;
        RECT 35.150 0.155 57.770 2.680 ;
        RECT 58.610 0.155 81.230 2.680 ;
        RECT 82.070 0.155 104.230 2.680 ;
        RECT 105.070 0.155 127.690 2.680 ;
        RECT 128.530 0.155 138.370 2.680 ;
      LAYER met3 ;
        RECT 28.050 124.120 138.395 128.005 ;
        RECT 28.050 122.720 137.200 124.120 ;
        RECT 28.050 113.240 138.395 122.720 ;
        RECT 28.050 111.840 137.200 113.240 ;
        RECT 28.050 102.360 138.395 111.840 ;
        RECT 28.050 100.960 137.200 102.360 ;
        RECT 28.050 91.480 138.395 100.960 ;
        RECT 28.050 90.080 137.200 91.480 ;
        RECT 28.050 80.600 138.395 90.080 ;
        RECT 28.050 79.200 137.200 80.600 ;
        RECT 28.050 70.400 138.395 79.200 ;
        RECT 28.050 69.000 137.200 70.400 ;
        RECT 28.050 59.520 138.395 69.000 ;
        RECT 28.050 58.120 137.200 59.520 ;
        RECT 28.050 48.640 138.395 58.120 ;
        RECT 28.050 47.240 137.200 48.640 ;
        RECT 28.050 37.760 138.395 47.240 ;
        RECT 28.050 36.360 137.200 37.760 ;
        RECT 28.050 26.880 138.395 36.360 ;
        RECT 28.050 25.480 137.200 26.880 ;
        RECT 28.050 16.000 138.395 25.480 ;
        RECT 28.050 14.600 137.200 16.000 ;
        RECT 28.050 5.800 138.395 14.600 ;
        RECT 28.050 4.400 137.200 5.800 ;
        RECT 28.050 0.175 138.395 4.400 ;
      LAYER met4 ;
        RECT 30.055 10.640 50.985 128.080 ;
        RECT 53.385 10.640 122.985 128.080 ;
  END
END grid_io_right
END LIBRARY

